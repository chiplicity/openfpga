magic
tech sky130A
magscale 1 2
timestamp 1604668940
<< locali >>
rect 14013 25143 14047 25245
rect 949 22627 983 24837
rect 19257 24735 19291 24905
rect 3249 23035 3283 23137
rect 3341 22967 3375 23273
rect 6377 21335 6411 21437
rect 6653 21335 6687 21641
rect 3249 19771 3283 19941
rect 3525 19363 3559 19465
rect 10517 18751 10551 18921
rect 6377 18071 6411 18377
rect 18153 17595 18187 17765
rect 23305 16099 23339 16201
rect 21649 14875 21683 14977
rect 6929 13787 6963 13889
rect 4905 12767 4939 12937
rect 8125 12699 8159 12869
rect 5365 12223 5399 12325
rect 9413 11543 9447 11849
rect 12081 10455 12115 10625
rect 12081 9367 12115 9605
rect 19257 9367 19291 9605
rect 22201 7803 22235 7905
rect 13093 7327 13127 7497
rect 21189 7259 21223 7429
rect 7481 6171 7515 6273
rect 3249 4607 3283 4777
rect 21833 4471 21867 4709
rect 4629 3995 4663 4165
rect 14841 2839 14875 3009
rect 24869 2295 24903 2397
<< viali >>
rect 2697 25449 2731 25483
rect 10977 25449 11011 25483
rect 14473 25449 14507 25483
rect 21373 25449 21407 25483
rect 13001 25381 13035 25415
rect 18981 25381 19015 25415
rect 1409 25313 1443 25347
rect 2513 25313 2547 25347
rect 4077 25313 4111 25347
rect 7849 25313 7883 25347
rect 9597 25313 9631 25347
rect 9873 25313 9907 25347
rect 10885 25313 10919 25347
rect 11345 25313 11379 25347
rect 12081 25313 12115 25347
rect 14289 25313 14323 25347
rect 16865 25313 16899 25347
rect 19993 25313 20027 25347
rect 21189 25313 21223 25347
rect 5181 25245 5215 25279
rect 7941 25245 7975 25279
rect 8125 25245 8159 25279
rect 11437 25245 11471 25279
rect 11529 25245 11563 25279
rect 13093 25245 13127 25279
rect 13277 25245 13311 25279
rect 14013 25245 14047 25279
rect 16129 25245 16163 25279
rect 16957 25245 16991 25279
rect 17049 25245 17083 25279
rect 17693 25245 17727 25279
rect 19073 25245 19107 25279
rect 19165 25245 19199 25279
rect 2421 25177 2455 25211
rect 4721 25177 4755 25211
rect 7297 25177 7331 25211
rect 8861 25177 8895 25211
rect 10057 25177 10091 25211
rect 10517 25177 10551 25211
rect 12633 25177 12667 25211
rect 1593 25109 1627 25143
rect 2053 25109 2087 25143
rect 3157 25109 3191 25143
rect 3709 25109 3743 25143
rect 4261 25109 4295 25143
rect 4997 25109 5031 25143
rect 5641 25109 5675 25143
rect 6745 25109 6779 25143
rect 7481 25109 7515 25143
rect 8585 25109 8619 25143
rect 12357 25109 12391 25143
rect 14013 25109 14047 25143
rect 14197 25109 14231 25143
rect 14841 25109 14875 25143
rect 15853 25109 15887 25143
rect 16497 25109 16531 25143
rect 18153 25109 18187 25143
rect 18613 25109 18647 25143
rect 19717 25109 19751 25143
rect 4629 24905 4663 24939
rect 6653 24905 6687 24939
rect 19257 24905 19291 24939
rect 949 24837 983 24871
rect 3801 24837 3835 24871
rect 15117 24837 15151 24871
rect 3065 24769 3099 24803
rect 3433 24769 3467 24803
rect 4169 24769 4203 24803
rect 5181 24769 5215 24803
rect 8769 24769 8803 24803
rect 10333 24769 10367 24803
rect 12173 24769 12207 24803
rect 13093 24769 13127 24803
rect 14749 24769 14783 24803
rect 16313 24769 16347 24803
rect 17877 24769 17911 24803
rect 18613 24769 18647 24803
rect 20177 24769 20211 24803
rect 1409 24701 1443 24735
rect 2329 24701 2363 24735
rect 2513 24701 2547 24735
rect 3617 24701 3651 24735
rect 4997 24701 5031 24735
rect 7113 24701 7147 24735
rect 8677 24701 8711 24735
rect 9689 24701 9723 24735
rect 10241 24701 10275 24735
rect 11897 24701 11931 24735
rect 16129 24701 16163 24735
rect 17141 24701 17175 24735
rect 18429 24701 18463 24735
rect 19073 24701 19107 24735
rect 19257 24701 19291 24735
rect 19533 24701 19567 24735
rect 21649 24701 21683 24735
rect 22201 24701 22235 24735
rect 23949 24701 23983 24735
rect 24501 24701 24535 24735
rect 5641 24633 5675 24667
rect 9321 24633 9355 24667
rect 10149 24633 10183 24667
rect 11345 24633 11379 24667
rect 12909 24633 12943 24667
rect 14013 24633 14047 24667
rect 15577 24633 15611 24667
rect 19993 24633 20027 24667
rect 1593 24565 1627 24599
rect 2053 24565 2087 24599
rect 2697 24565 2731 24599
rect 4445 24565 4479 24599
rect 5089 24565 5123 24599
rect 6009 24565 6043 24599
rect 7297 24565 7331 24599
rect 7757 24565 7791 24599
rect 8125 24565 8159 24599
rect 8217 24565 8251 24599
rect 8585 24565 8619 24599
rect 9781 24565 9815 24599
rect 11069 24565 11103 24599
rect 12541 24565 12575 24599
rect 13001 24565 13035 24599
rect 13645 24565 13679 24599
rect 14105 24565 14139 24599
rect 14473 24565 14507 24599
rect 14565 24565 14599 24599
rect 15761 24565 15795 24599
rect 16221 24565 16255 24599
rect 16865 24565 16899 24599
rect 18061 24565 18095 24599
rect 18521 24565 18555 24599
rect 19625 24565 19659 24599
rect 20085 24565 20119 24599
rect 20637 24565 20671 24599
rect 21189 24565 21223 24599
rect 21833 24565 21867 24599
rect 24133 24565 24167 24599
rect 2145 24361 2179 24395
rect 4537 24361 4571 24395
rect 12725 24361 12759 24395
rect 13461 24361 13495 24395
rect 15485 24361 15519 24395
rect 18613 24361 18647 24395
rect 19533 24361 19567 24395
rect 19901 24361 19935 24395
rect 21373 24361 21407 24395
rect 21925 24361 21959 24395
rect 22661 24361 22695 24395
rect 24685 24361 24719 24395
rect 2053 24293 2087 24327
rect 10762 24293 10796 24327
rect 15117 24293 15151 24327
rect 16957 24293 16991 24327
rect 18521 24293 18555 24327
rect 4905 24225 4939 24259
rect 6920 24225 6954 24259
rect 13369 24225 13403 24259
rect 15301 24225 15335 24259
rect 19165 24225 19199 24259
rect 19717 24225 19751 24259
rect 21281 24225 21315 24259
rect 22477 24225 22511 24259
rect 24501 24225 24535 24259
rect 2329 24157 2363 24191
rect 2789 24157 2823 24191
rect 4997 24157 5031 24191
rect 5089 24157 5123 24191
rect 5917 24157 5951 24191
rect 6653 24157 6687 24191
rect 10517 24157 10551 24191
rect 13645 24157 13679 24191
rect 17049 24157 17083 24191
rect 17233 24157 17267 24191
rect 18705 24157 18739 24191
rect 21465 24157 21499 24191
rect 3525 24089 3559 24123
rect 14749 24089 14783 24123
rect 16497 24089 16531 24123
rect 17693 24089 17727 24123
rect 18061 24089 18095 24123
rect 20545 24089 20579 24123
rect 20913 24089 20947 24123
rect 1685 24021 1719 24055
rect 3157 24021 3191 24055
rect 3893 24021 3927 24055
rect 4445 24021 4479 24055
rect 5641 24021 5675 24055
rect 6561 24021 6595 24055
rect 8033 24021 8067 24055
rect 8677 24021 8711 24055
rect 9505 24021 9539 24055
rect 9965 24021 9999 24055
rect 10425 24021 10459 24055
rect 11897 24021 11931 24055
rect 13001 24021 13035 24055
rect 14197 24021 14231 24055
rect 15853 24021 15887 24055
rect 16589 24021 16623 24055
rect 18153 24021 18187 24055
rect 3617 23817 3651 23851
rect 6193 23817 6227 23851
rect 6561 23817 6595 23851
rect 8033 23817 8067 23851
rect 10149 23817 10183 23851
rect 12265 23817 12299 23851
rect 14381 23817 14415 23851
rect 20545 23817 20579 23851
rect 21557 23817 21591 23851
rect 22293 23817 22327 23851
rect 24777 23817 24811 23851
rect 5181 23749 5215 23783
rect 15209 23749 15243 23783
rect 2145 23681 2179 23715
rect 2329 23681 2363 23715
rect 4077 23681 4111 23715
rect 4261 23681 4295 23715
rect 4721 23681 4755 23715
rect 5641 23681 5675 23715
rect 5825 23681 5859 23715
rect 7481 23681 7515 23715
rect 8217 23681 8251 23715
rect 11253 23681 11287 23715
rect 11437 23681 11471 23715
rect 21097 23681 21131 23715
rect 25145 23681 25179 23715
rect 3525 23613 3559 23647
rect 6837 23613 6871 23647
rect 10609 23613 10643 23647
rect 12449 23613 12483 23647
rect 14749 23613 14783 23647
rect 15301 23613 15335 23647
rect 15557 23613 15591 23647
rect 17785 23613 17819 23647
rect 18061 23613 18095 23647
rect 22109 23613 22143 23647
rect 24593 23613 24627 23647
rect 2053 23545 2087 23579
rect 5089 23545 5123 23579
rect 5549 23545 5583 23579
rect 8484 23545 8518 23579
rect 11897 23545 11931 23579
rect 12694 23545 12728 23579
rect 18306 23545 18340 23579
rect 20085 23545 20119 23579
rect 20913 23545 20947 23579
rect 1685 23477 1719 23511
rect 2789 23477 2823 23511
rect 3157 23477 3191 23511
rect 3985 23477 4019 23511
rect 7021 23477 7055 23511
rect 9597 23477 9631 23511
rect 10793 23477 10827 23511
rect 11161 23477 11195 23511
rect 13829 23477 13863 23511
rect 16681 23477 16715 23511
rect 17509 23477 17543 23511
rect 19441 23477 19475 23511
rect 20361 23477 20395 23511
rect 21005 23477 21039 23511
rect 21925 23477 21959 23511
rect 22661 23477 22695 23511
rect 24501 23477 24535 23511
rect 1593 23273 1627 23307
rect 2421 23273 2455 23307
rect 2789 23273 2823 23307
rect 3341 23273 3375 23307
rect 4537 23273 4571 23307
rect 7205 23273 7239 23307
rect 7849 23273 7883 23307
rect 9137 23273 9171 23307
rect 10057 23273 10091 23307
rect 10149 23273 10183 23307
rect 11253 23273 11287 23307
rect 12817 23273 12851 23307
rect 13185 23273 13219 23307
rect 15853 23273 15887 23307
rect 18797 23273 18831 23307
rect 19349 23273 19383 23307
rect 20269 23273 20303 23307
rect 20637 23273 20671 23307
rect 22017 23273 22051 23307
rect 22937 23273 22971 23307
rect 24777 23273 24811 23307
rect 1401 23137 1435 23171
rect 3249 23137 3283 23171
rect 2329 23069 2363 23103
rect 2881 23069 2915 23103
rect 3065 23069 3099 23103
rect 3249 23001 3283 23035
rect 10885 23205 10919 23239
rect 11713 23205 11747 23239
rect 13921 23205 13955 23239
rect 16764 23205 16798 23239
rect 23489 23205 23523 23239
rect 4905 23137 4939 23171
rect 5172 23137 5206 23171
rect 8401 23137 8435 23171
rect 9505 23137 9539 23171
rect 11621 23137 11655 23171
rect 13277 23137 13311 23171
rect 14749 23137 14783 23171
rect 15301 23137 15335 23171
rect 19441 23137 19475 23171
rect 21281 23137 21315 23171
rect 22845 23137 22879 23171
rect 24593 23137 24627 23171
rect 8493 23069 8527 23103
rect 8585 23069 8619 23103
rect 10333 23069 10367 23103
rect 11805 23069 11839 23103
rect 13461 23069 13495 23103
rect 16497 23069 16531 23103
rect 19533 23069 19567 23103
rect 21373 23069 21407 23103
rect 21465 23069 21499 23103
rect 23029 23069 23063 23103
rect 3525 23001 3559 23035
rect 8033 23001 8067 23035
rect 9689 23001 9723 23035
rect 15485 23001 15519 23035
rect 1961 22933 1995 22967
rect 3341 22933 3375 22967
rect 3893 22933 3927 22967
rect 6285 22933 6319 22967
rect 6929 22933 6963 22967
rect 12449 22933 12483 22967
rect 14473 22933 14507 22967
rect 16313 22933 16347 22967
rect 17877 22933 17911 22967
rect 18429 22933 18463 22967
rect 18981 22933 19015 22967
rect 20913 22933 20947 22967
rect 22293 22933 22327 22967
rect 22477 22933 22511 22967
rect 2697 22729 2731 22763
rect 3709 22729 3743 22763
rect 6837 22729 6871 22763
rect 8401 22729 8435 22763
rect 10701 22729 10735 22763
rect 11437 22729 11471 22763
rect 12173 22729 12207 22763
rect 12449 22729 12483 22763
rect 13461 22729 13495 22763
rect 15761 22729 15795 22763
rect 17049 22729 17083 22763
rect 18705 22729 18739 22763
rect 22845 22729 22879 22763
rect 23857 22729 23891 22763
rect 1593 22661 1627 22695
rect 11069 22661 11103 22695
rect 20913 22661 20947 22695
rect 21189 22661 21223 22695
rect 949 22593 983 22627
rect 1961 22593 1995 22627
rect 2605 22593 2639 22627
rect 3341 22593 3375 22627
rect 6285 22593 6319 22627
rect 7481 22593 7515 22627
rect 8585 22593 8619 22627
rect 13001 22593 13035 22627
rect 18429 22593 18463 22627
rect 21925 22593 21959 22627
rect 22569 22593 22603 22627
rect 24593 22593 24627 22627
rect 1409 22525 1443 22559
rect 3157 22525 3191 22559
rect 4169 22525 4203 22559
rect 4261 22525 4295 22559
rect 11253 22525 11287 22559
rect 12817 22525 12851 22559
rect 14197 22525 14231 22559
rect 14381 22525 14415 22559
rect 14637 22525 14671 22559
rect 16865 22525 16899 22559
rect 17417 22525 17451 22559
rect 18889 22525 18923 22559
rect 19156 22525 19190 22559
rect 21833 22525 21867 22559
rect 23673 22525 23707 22559
rect 24225 22525 24259 22559
rect 24777 22525 24811 22559
rect 4506 22457 4540 22491
rect 6653 22457 6687 22491
rect 7297 22457 7331 22491
rect 8125 22457 8159 22491
rect 8852 22457 8886 22491
rect 12909 22457 12943 22491
rect 13829 22457 13863 22491
rect 25237 22457 25271 22491
rect 3065 22389 3099 22423
rect 5641 22389 5675 22423
rect 7205 22389 7239 22423
rect 9965 22389 9999 22423
rect 11805 22389 11839 22423
rect 16497 22389 16531 22423
rect 17785 22389 17819 22423
rect 20269 22389 20303 22423
rect 21373 22389 21407 22423
rect 21741 22389 21775 22423
rect 23213 22389 23247 22423
rect 24961 22389 24995 22423
rect 1961 22185 1995 22219
rect 5733 22185 5767 22219
rect 6469 22185 6503 22219
rect 9413 22185 9447 22219
rect 10333 22185 10367 22219
rect 12357 22185 12391 22219
rect 12909 22185 12943 22219
rect 13461 22185 13495 22219
rect 17785 22185 17819 22219
rect 19073 22185 19107 22219
rect 20729 22185 20763 22219
rect 22845 22185 22879 22219
rect 23213 22185 23247 22219
rect 4629 22117 4663 22151
rect 6837 22117 6871 22151
rect 8401 22117 8435 22151
rect 13829 22117 13863 22151
rect 13921 22117 13955 22151
rect 24409 22117 24443 22151
rect 1869 22049 1903 22083
rect 2329 22049 2363 22083
rect 4721 22049 4755 22083
rect 6377 22049 6411 22083
rect 9137 22049 9171 22083
rect 9689 22049 9723 22083
rect 11244 22049 11278 22083
rect 14473 22049 14507 22083
rect 15568 22049 15602 22083
rect 17233 22049 17267 22083
rect 18153 22049 18187 22083
rect 19349 22049 19383 22083
rect 21649 22049 21683 22083
rect 22753 22049 22787 22083
rect 23949 22049 23983 22083
rect 25421 22049 25455 22083
rect 2421 21981 2455 22015
rect 2605 21981 2639 22015
rect 4813 21981 4847 22015
rect 6929 21981 6963 22015
rect 7113 21981 7147 22015
rect 8493 21981 8527 22015
rect 8585 21981 8619 22015
rect 10977 21981 11011 22015
rect 14013 21981 14047 22015
rect 15301 21981 15335 22015
rect 18245 21981 18279 22015
rect 18337 21981 18371 22015
rect 21741 21981 21775 22015
rect 21833 21981 21867 22015
rect 23305 21981 23339 22015
rect 23397 21981 23431 22015
rect 3065 21913 3099 21947
rect 5365 21913 5399 21947
rect 8033 21913 8067 21947
rect 9873 21913 9907 21947
rect 16681 21913 16715 21947
rect 17693 21913 17727 21947
rect 19533 21913 19567 21947
rect 20361 21913 20395 21947
rect 21281 21913 21315 21947
rect 3617 21845 3651 21879
rect 4261 21845 4295 21879
rect 7665 21845 7699 21879
rect 10701 21845 10735 21879
rect 13369 21845 13403 21879
rect 14841 21845 14875 21879
rect 19993 21845 20027 21879
rect 21097 21845 21131 21879
rect 22293 21845 22327 21879
rect 25605 21845 25639 21879
rect 1777 21641 1811 21675
rect 1961 21641 1995 21675
rect 3525 21641 3559 21675
rect 5089 21641 5123 21675
rect 6653 21641 6687 21675
rect 7573 21641 7607 21675
rect 9045 21641 9079 21675
rect 11529 21641 11563 21675
rect 12725 21641 12759 21675
rect 16313 21641 16347 21675
rect 16405 21641 16439 21675
rect 17509 21641 17543 21675
rect 17877 21641 17911 21675
rect 21465 21641 21499 21675
rect 23213 21641 23247 21675
rect 25421 21641 25455 21675
rect 3341 21573 3375 21607
rect 4905 21573 4939 21607
rect 2421 21505 2455 21539
rect 2605 21505 2639 21539
rect 3985 21505 4019 21539
rect 4077 21505 4111 21539
rect 5641 21505 5675 21539
rect 2329 21437 2363 21471
rect 2973 21437 3007 21471
rect 5457 21437 5491 21471
rect 6377 21437 6411 21471
rect 6193 21369 6227 21403
rect 10149 21573 10183 21607
rect 26157 21573 26191 21607
rect 10609 21505 10643 21539
rect 10793 21505 10827 21539
rect 16957 21505 16991 21539
rect 18797 21505 18831 21539
rect 18981 21505 19015 21539
rect 20545 21505 20579 21539
rect 22109 21505 22143 21539
rect 22293 21505 22327 21539
rect 24133 21505 24167 21539
rect 24225 21505 24259 21539
rect 7021 21437 7055 21471
rect 7665 21437 7699 21471
rect 11161 21437 11195 21471
rect 13277 21437 13311 21471
rect 15301 21437 15335 21471
rect 16773 21437 16807 21471
rect 18705 21437 18739 21471
rect 20361 21437 20395 21471
rect 24041 21437 24075 21471
rect 25237 21437 25271 21471
rect 25789 21437 25823 21471
rect 7932 21369 7966 21403
rect 9781 21369 9815 21403
rect 13544 21369 13578 21403
rect 16865 21369 16899 21403
rect 19717 21369 19751 21403
rect 20269 21369 20303 21403
rect 21097 21369 21131 21403
rect 24685 21369 24719 21403
rect 3893 21301 3927 21335
rect 4629 21301 4663 21335
rect 5549 21301 5583 21335
rect 6377 21301 6411 21335
rect 6561 21301 6595 21335
rect 6653 21301 6687 21335
rect 10517 21301 10551 21335
rect 11897 21301 11931 21335
rect 13185 21301 13219 21335
rect 14657 21301 14691 21335
rect 15669 21301 15703 21335
rect 18337 21301 18371 21335
rect 19349 21301 19383 21335
rect 19901 21301 19935 21335
rect 21649 21301 21683 21335
rect 22017 21301 22051 21335
rect 22937 21301 22971 21335
rect 23673 21301 23707 21335
rect 1961 21097 1995 21131
rect 2329 21097 2363 21131
rect 4077 21097 4111 21131
rect 4537 21097 4571 21131
rect 7573 21097 7607 21131
rect 9045 21097 9079 21131
rect 11069 21097 11103 21131
rect 12173 21097 12207 21131
rect 13553 21097 13587 21131
rect 14289 21097 14323 21131
rect 15301 21097 15335 21131
rect 16865 21097 16899 21131
rect 16957 21097 16991 21131
rect 18061 21097 18095 21131
rect 18981 21097 19015 21131
rect 19625 21097 19659 21131
rect 20361 21097 20395 21131
rect 20729 21097 20763 21131
rect 21741 21097 21775 21131
rect 24225 21097 24259 21131
rect 24777 21097 24811 21131
rect 1777 21029 1811 21063
rect 6101 21029 6135 21063
rect 9934 21029 9968 21063
rect 13829 21029 13863 21063
rect 17325 21029 17359 21063
rect 18429 21029 18463 21063
rect 19993 21029 20027 21063
rect 22192 21029 22226 21063
rect 23949 21029 23983 21063
rect 4445 20961 4479 20995
rect 6009 20961 6043 20995
rect 7113 20961 7147 20995
rect 8309 20961 8343 20995
rect 12081 20961 12115 20995
rect 12541 20961 12575 20995
rect 12633 20961 12667 20995
rect 14105 20961 14139 20995
rect 15669 20961 15703 20995
rect 16497 20961 16531 20995
rect 17417 20961 17451 20995
rect 18889 20961 18923 20995
rect 2421 20893 2455 20927
rect 2605 20893 2639 20927
rect 3249 20893 3283 20927
rect 4629 20893 4663 20927
rect 5089 20893 5123 20927
rect 6193 20893 6227 20927
rect 7665 20893 7699 20927
rect 7757 20893 7791 20927
rect 9689 20893 9723 20927
rect 11621 20893 11655 20927
rect 12725 20893 12759 20927
rect 15761 20893 15795 20927
rect 15945 20893 15979 20927
rect 17509 20893 17543 20927
rect 19073 20893 19107 20927
rect 20913 20893 20947 20927
rect 21925 20893 21959 20927
rect 24869 20893 24903 20927
rect 25053 20893 25087 20927
rect 5457 20825 5491 20859
rect 5641 20825 5675 20859
rect 6653 20825 6687 20859
rect 8677 20825 8711 20859
rect 3617 20757 3651 20791
rect 7205 20757 7239 20791
rect 9413 20757 9447 20791
rect 14657 20757 14691 20791
rect 15025 20757 15059 20791
rect 18521 20757 18555 20791
rect 23305 20757 23339 20791
rect 24409 20757 24443 20791
rect 1777 20553 1811 20587
rect 1961 20553 1995 20587
rect 3065 20553 3099 20587
rect 6193 20553 6227 20587
rect 6469 20553 6503 20587
rect 7389 20553 7423 20587
rect 10333 20553 10367 20587
rect 12449 20553 12483 20587
rect 13461 20553 13495 20587
rect 16221 20553 16255 20587
rect 16405 20553 16439 20587
rect 17509 20553 17543 20587
rect 18981 20553 19015 20587
rect 21189 20553 21223 20587
rect 23489 20553 23523 20587
rect 25421 20553 25455 20587
rect 26249 20553 26283 20587
rect 3341 20485 3375 20519
rect 10241 20485 10275 20519
rect 13921 20485 13955 20519
rect 18245 20485 18279 20519
rect 23673 20485 23707 20519
rect 2421 20417 2455 20451
rect 2605 20417 2639 20451
rect 6837 20417 6871 20451
rect 10885 20417 10919 20451
rect 11345 20417 11379 20451
rect 11805 20417 11839 20451
rect 13001 20417 13035 20451
rect 14565 20417 14599 20451
rect 16957 20417 16991 20451
rect 22293 20417 22327 20451
rect 24133 20417 24167 20451
rect 24317 20417 24351 20451
rect 24685 20417 24719 20451
rect 3801 20349 3835 20383
rect 4068 20349 4102 20383
rect 5733 20349 5767 20383
rect 7849 20349 7883 20383
rect 8105 20349 8139 20383
rect 10793 20349 10827 20383
rect 12909 20349 12943 20383
rect 15669 20349 15703 20383
rect 16773 20349 16807 20383
rect 18061 20349 18095 20383
rect 18613 20349 18647 20383
rect 19165 20349 19199 20383
rect 21557 20349 21591 20383
rect 22017 20349 22051 20383
rect 22109 20349 22143 20383
rect 25237 20349 25271 20383
rect 25789 20349 25823 20383
rect 14473 20281 14507 20315
rect 16865 20281 16899 20315
rect 17785 20281 17819 20315
rect 19432 20281 19466 20315
rect 23121 20281 23155 20315
rect 24041 20281 24075 20315
rect 2329 20213 2363 20247
rect 5181 20213 5215 20247
rect 7665 20213 7699 20247
rect 9229 20213 9263 20247
rect 9873 20213 9907 20247
rect 10701 20213 10735 20247
rect 12173 20213 12207 20247
rect 12817 20213 12851 20247
rect 14013 20213 14047 20247
rect 14381 20213 14415 20247
rect 15301 20213 15335 20247
rect 20545 20213 20579 20247
rect 21649 20213 21683 20247
rect 22661 20213 22695 20247
rect 25053 20213 25087 20247
rect 1961 20009 1995 20043
rect 5089 20009 5123 20043
rect 6929 20009 6963 20043
rect 7849 20009 7883 20043
rect 8033 20009 8067 20043
rect 9689 20009 9723 20043
rect 11161 20009 11195 20043
rect 12541 20009 12575 20043
rect 14105 20009 14139 20043
rect 15117 20009 15151 20043
rect 15761 20009 15795 20043
rect 16497 20009 16531 20043
rect 19073 20009 19107 20043
rect 19625 20009 19659 20043
rect 20269 20009 20303 20043
rect 22845 20009 22879 20043
rect 2881 19941 2915 19975
rect 3249 19941 3283 19975
rect 3525 19941 3559 19975
rect 4721 19941 4755 19975
rect 5794 19941 5828 19975
rect 8401 19941 8435 19975
rect 12081 19941 12115 19975
rect 12992 19941 13026 19975
rect 23642 19941 23676 19975
rect 2789 19873 2823 19907
rect 1409 19805 1443 19839
rect 3065 19805 3099 19839
rect 4077 19873 4111 19907
rect 11069 19873 11103 19907
rect 12725 19873 12759 19907
rect 15669 19873 15703 19907
rect 17417 19873 17451 19907
rect 17509 19873 17543 19907
rect 18981 19873 19015 19907
rect 20913 19873 20947 19907
rect 21180 19873 21214 19907
rect 5549 19805 5583 19839
rect 7573 19805 7607 19839
rect 8493 19805 8527 19839
rect 8585 19805 8619 19839
rect 11345 19805 11379 19839
rect 11713 19805 11747 19839
rect 15853 19805 15887 19839
rect 17601 19805 17635 19839
rect 19257 19805 19291 19839
rect 23397 19805 23431 19839
rect 3249 19737 3283 19771
rect 10701 19737 10735 19771
rect 14657 19737 14691 19771
rect 18153 19737 18187 19771
rect 18521 19737 18555 19771
rect 22293 19737 22327 19771
rect 2421 19669 2455 19703
rect 3801 19669 3835 19703
rect 4261 19669 4295 19703
rect 5457 19669 5491 19703
rect 9137 19669 9171 19703
rect 9505 19669 9539 19703
rect 10333 19669 10367 19703
rect 15301 19669 15335 19703
rect 16957 19669 16991 19703
rect 17049 19669 17083 19703
rect 18613 19669 18647 19703
rect 20729 19669 20763 19703
rect 23305 19669 23339 19703
rect 24777 19669 24811 19703
rect 3525 19465 3559 19499
rect 4077 19465 4111 19499
rect 6561 19465 6595 19499
rect 9413 19465 9447 19499
rect 11897 19465 11931 19499
rect 14565 19465 14599 19499
rect 14933 19465 14967 19499
rect 16865 19465 16899 19499
rect 21557 19465 21591 19499
rect 24685 19465 24719 19499
rect 10793 19397 10827 19431
rect 12173 19397 12207 19431
rect 21189 19397 21223 19431
rect 3341 19329 3375 19363
rect 3525 19329 3559 19363
rect 7849 19329 7883 19363
rect 8033 19329 8067 19363
rect 11345 19329 11379 19363
rect 12817 19329 12851 19363
rect 13737 19329 13771 19363
rect 15669 19329 15703 19363
rect 19257 19329 19291 19363
rect 20729 19329 20763 19363
rect 22569 19329 22603 19363
rect 23397 19329 23431 19363
rect 24225 19329 24259 19363
rect 1409 19261 1443 19295
rect 2053 19261 2087 19295
rect 3065 19261 3099 19295
rect 4261 19261 4295 19295
rect 4528 19261 4562 19295
rect 6837 19261 6871 19295
rect 11253 19261 11287 19295
rect 13645 19261 13679 19295
rect 14289 19261 14323 19295
rect 15577 19261 15611 19295
rect 16957 19261 16991 19295
rect 19625 19261 19659 19295
rect 22477 19261 22511 19295
rect 24133 19261 24167 19295
rect 25237 19261 25271 19295
rect 25789 19261 25823 19295
rect 2605 19193 2639 19227
rect 3801 19193 3835 19227
rect 8278 19193 8312 19227
rect 10333 19193 10367 19227
rect 15485 19193 15519 19227
rect 17417 19193 17451 19227
rect 20085 19193 20119 19227
rect 20545 19193 20579 19227
rect 24041 19193 24075 19227
rect 25053 19193 25087 19227
rect 1593 19125 1627 19159
rect 2697 19125 2731 19159
rect 3157 19125 3191 19159
rect 5641 19125 5675 19159
rect 6285 19125 6319 19159
rect 7021 19125 7055 19159
rect 7481 19125 7515 19159
rect 10701 19125 10735 19159
rect 11161 19125 11195 19159
rect 13185 19125 13219 19159
rect 13553 19125 13587 19159
rect 15117 19125 15151 19159
rect 16129 19125 16163 19159
rect 17141 19125 17175 19159
rect 17785 19125 17819 19159
rect 18429 19125 18463 19159
rect 18613 19125 18647 19159
rect 18981 19125 19015 19159
rect 19073 19125 19107 19159
rect 20177 19125 20211 19159
rect 20637 19125 20671 19159
rect 22017 19125 22051 19159
rect 22385 19125 22419 19159
rect 23029 19125 23063 19159
rect 23673 19125 23707 19159
rect 25421 19125 25455 19159
rect 1593 18921 1627 18955
rect 1961 18921 1995 18955
rect 2881 18921 2915 18955
rect 3525 18921 3559 18955
rect 3893 18921 3927 18955
rect 4629 18921 4663 18955
rect 6745 18921 6779 18955
rect 8033 18921 8067 18955
rect 8493 18921 8527 18955
rect 9505 18921 9539 18955
rect 9873 18921 9907 18955
rect 10517 18921 10551 18955
rect 12173 18921 12207 18955
rect 12725 18921 12759 18955
rect 13277 18921 13311 18955
rect 15117 18921 15151 18955
rect 16129 18921 16163 18955
rect 17693 18921 17727 18955
rect 19257 18921 19291 18955
rect 19809 18921 19843 18955
rect 20177 18921 20211 18955
rect 20729 18921 20763 18955
rect 21465 18921 21499 18955
rect 22109 18921 22143 18955
rect 23949 18921 23983 18955
rect 25237 18921 25271 18955
rect 5632 18853 5666 18887
rect 7481 18853 7515 18887
rect 9045 18853 9079 18887
rect 1409 18785 1443 18819
rect 2789 18785 2823 18819
rect 4077 18785 4111 18819
rect 5365 18785 5399 18819
rect 8401 18785 8435 18819
rect 9689 18785 9723 18819
rect 11060 18853 11094 18887
rect 22814 18853 22848 18887
rect 10793 18785 10827 18819
rect 13737 18785 13771 18819
rect 15301 18785 15335 18819
rect 16313 18785 16347 18819
rect 16580 18785 16614 18819
rect 19165 18785 19199 18819
rect 21373 18785 21407 18819
rect 22569 18785 22603 18819
rect 24501 18785 24535 18819
rect 25053 18785 25087 18819
rect 2329 18717 2363 18751
rect 3065 18717 3099 18751
rect 5181 18717 5215 18751
rect 8585 18717 8619 18751
rect 10241 18717 10275 18751
rect 10517 18717 10551 18751
rect 10609 18717 10643 18751
rect 13829 18717 13863 18751
rect 14013 18717 14047 18751
rect 18337 18717 18371 18751
rect 19349 18717 19383 18751
rect 21557 18717 21591 18751
rect 15485 18649 15519 18683
rect 21005 18649 21039 18683
rect 2421 18581 2455 18615
rect 4261 18581 4295 18615
rect 7941 18581 7975 18615
rect 13369 18581 13403 18615
rect 14381 18581 14415 18615
rect 15853 18581 15887 18615
rect 18613 18581 18647 18615
rect 18797 18581 18831 18615
rect 22385 18581 22419 18615
rect 1777 18377 1811 18411
rect 3617 18377 3651 18411
rect 4537 18377 4571 18411
rect 5089 18377 5123 18411
rect 6377 18377 6411 18411
rect 8953 18377 8987 18411
rect 9229 18377 9263 18411
rect 10793 18377 10827 18411
rect 11805 18377 11839 18411
rect 13093 18377 13127 18411
rect 13553 18377 13587 18411
rect 14565 18377 14599 18411
rect 17417 18377 17451 18411
rect 17877 18377 17911 18411
rect 18613 18377 18647 18411
rect 20453 18377 20487 18411
rect 21005 18377 21039 18411
rect 21373 18377 21407 18411
rect 23673 18377 23707 18411
rect 24685 18377 24719 18411
rect 25053 18377 25087 18411
rect 25421 18377 25455 18411
rect 2145 18309 2179 18343
rect 4261 18309 4295 18343
rect 2237 18241 2271 18275
rect 5733 18241 5767 18275
rect 2504 18173 2538 18207
rect 5549 18105 5583 18139
rect 7113 18309 7147 18343
rect 12173 18309 12207 18343
rect 16497 18309 16531 18343
rect 23489 18309 23523 18343
rect 6653 18241 6687 18275
rect 8033 18241 8067 18275
rect 8217 18241 8251 18275
rect 8585 18241 8619 18275
rect 9689 18241 9723 18275
rect 9781 18241 9815 18275
rect 11345 18241 11379 18275
rect 12541 18241 12575 18275
rect 14197 18241 14231 18275
rect 22201 18241 22235 18275
rect 23121 18241 23155 18275
rect 24133 18241 24167 18275
rect 24225 18241 24259 18275
rect 7481 18173 7515 18207
rect 7941 18173 7975 18207
rect 9597 18173 9631 18207
rect 10333 18173 10367 18207
rect 13921 18173 13955 18207
rect 15117 18173 15151 18207
rect 15384 18173 15418 18207
rect 18061 18173 18095 18207
rect 18889 18173 18923 18207
rect 19073 18173 19107 18207
rect 19329 18173 19363 18207
rect 21925 18173 21959 18207
rect 24041 18173 24075 18207
rect 25237 18173 25271 18207
rect 25789 18173 25823 18207
rect 11161 18105 11195 18139
rect 14013 18105 14047 18139
rect 5181 18037 5215 18071
rect 5641 18037 5675 18071
rect 6285 18037 6319 18071
rect 6377 18037 6411 18071
rect 7573 18037 7607 18071
rect 10701 18037 10735 18071
rect 11253 18037 11287 18071
rect 13369 18037 13403 18071
rect 14933 18037 14967 18071
rect 17049 18037 17083 18071
rect 18245 18037 18279 18071
rect 21557 18037 21591 18071
rect 22017 18037 22051 18071
rect 22661 18037 22695 18071
rect 3893 17833 3927 17867
rect 4905 17833 4939 17867
rect 6285 17833 6319 17867
rect 7941 17833 7975 17867
rect 8493 17833 8527 17867
rect 9689 17833 9723 17867
rect 10885 17833 10919 17867
rect 14933 17833 14967 17867
rect 17601 17833 17635 17867
rect 17969 17833 18003 17867
rect 19717 17833 19751 17867
rect 20269 17833 20303 17867
rect 20729 17833 20763 17867
rect 22569 17833 22603 17867
rect 25421 17833 25455 17867
rect 1768 17765 1802 17799
rect 3433 17765 3467 17799
rect 11621 17765 11655 17799
rect 13921 17765 13955 17799
rect 14565 17765 14599 17799
rect 15568 17765 15602 17799
rect 18153 17765 18187 17799
rect 21281 17765 21315 17799
rect 25053 17765 25087 17799
rect 1501 17697 1535 17731
rect 4813 17697 4847 17731
rect 5273 17697 5307 17731
rect 6837 17697 6871 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 11713 17697 11747 17731
rect 12265 17697 12299 17731
rect 13185 17697 13219 17731
rect 5365 17629 5399 17663
rect 5457 17629 5491 17663
rect 6929 17629 6963 17663
rect 7021 17629 7055 17663
rect 8677 17629 8711 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 11805 17629 11839 17663
rect 13277 17629 13311 17663
rect 13461 17629 13495 17663
rect 15301 17629 15335 17663
rect 18593 17697 18627 17731
rect 23009 17697 23043 17731
rect 25237 17697 25271 17731
rect 18337 17629 18371 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 22753 17629 22787 17663
rect 4445 17561 4479 17595
rect 5917 17561 5951 17595
rect 9229 17561 9263 17595
rect 14197 17561 14231 17595
rect 18153 17561 18187 17595
rect 24685 17561 24719 17595
rect 2881 17493 2915 17527
rect 6469 17493 6503 17527
rect 7481 17493 7515 17527
rect 8033 17493 8067 17527
rect 11253 17493 11287 17527
rect 12633 17493 12667 17527
rect 12817 17493 12851 17527
rect 16681 17493 16715 17527
rect 17325 17493 17359 17527
rect 20913 17493 20947 17527
rect 21925 17493 21959 17527
rect 24133 17493 24167 17527
rect 1685 17289 1719 17323
rect 2053 17289 2087 17323
rect 4261 17289 4295 17323
rect 5181 17289 5215 17323
rect 8769 17289 8803 17323
rect 9413 17289 9447 17323
rect 12173 17289 12207 17323
rect 16221 17289 16255 17323
rect 17509 17289 17543 17323
rect 17877 17289 17911 17323
rect 20453 17289 20487 17323
rect 23489 17289 23523 17323
rect 25421 17289 25455 17323
rect 4629 17221 4663 17255
rect 9689 17221 9723 17255
rect 15301 17221 15335 17255
rect 18521 17221 18555 17255
rect 18889 17221 18923 17255
rect 21465 17221 21499 17255
rect 2145 17153 2179 17187
rect 5733 17153 5767 17187
rect 12449 17153 12483 17187
rect 15393 17153 15427 17187
rect 16865 17153 16899 17187
rect 17049 17153 17083 17187
rect 19073 17153 19107 17187
rect 22109 17153 22143 17187
rect 24133 17153 24167 17187
rect 24225 17153 24259 17187
rect 5089 17085 5123 17119
rect 5641 17085 5675 17119
rect 6837 17085 6871 17119
rect 9873 17085 9907 17119
rect 16773 17085 16807 17119
rect 19340 17085 19374 17119
rect 21925 17085 21959 17119
rect 24685 17085 24719 17119
rect 25237 17085 25271 17119
rect 25789 17085 25823 17119
rect 2412 17017 2446 17051
rect 5549 17017 5583 17051
rect 7082 17017 7116 17051
rect 10118 17017 10152 17051
rect 11805 17017 11839 17051
rect 12694 17017 12728 17051
rect 14381 17017 14415 17051
rect 22017 17017 22051 17051
rect 23029 17017 23063 17051
rect 24041 17017 24075 17051
rect 3525 16949 3559 16983
rect 6561 16949 6595 16983
rect 8217 16949 8251 16983
rect 11253 16949 11287 16983
rect 13829 16949 13863 16983
rect 14933 16949 14967 16983
rect 15853 16949 15887 16983
rect 16405 16949 16439 16983
rect 18061 16949 18095 16983
rect 21005 16949 21039 16983
rect 21557 16949 21591 16983
rect 22753 16949 22787 16983
rect 23673 16949 23707 16983
rect 25145 16949 25179 16983
rect 1593 16745 1627 16779
rect 3525 16745 3559 16779
rect 3801 16745 3835 16779
rect 6377 16745 6411 16779
rect 7941 16745 7975 16779
rect 8493 16745 8527 16779
rect 9413 16745 9447 16779
rect 9965 16745 9999 16779
rect 11713 16745 11747 16779
rect 12817 16745 12851 16779
rect 14197 16745 14231 16779
rect 14565 16745 14599 16779
rect 17141 16745 17175 16779
rect 18705 16745 18739 16779
rect 19717 16745 19751 16779
rect 20269 16745 20303 16779
rect 20637 16745 20671 16779
rect 20913 16745 20947 16779
rect 22661 16745 22695 16779
rect 24685 16745 24719 16779
rect 25421 16745 25455 16779
rect 2145 16677 2179 16711
rect 2881 16677 2915 16711
rect 4322 16677 4356 16711
rect 6806 16677 6840 16711
rect 10578 16677 10612 16711
rect 13185 16677 13219 16711
rect 14933 16677 14967 16711
rect 15669 16677 15703 16711
rect 18797 16677 18831 16711
rect 19441 16677 19475 16711
rect 21373 16677 21407 16711
rect 22998 16677 23032 16711
rect 25053 16677 25087 16711
rect 1409 16609 1443 16643
rect 2789 16609 2823 16643
rect 4077 16609 4111 16643
rect 6101 16609 6135 16643
rect 9045 16609 9079 16643
rect 10333 16609 10367 16643
rect 13829 16609 13863 16643
rect 15761 16609 15795 16643
rect 17233 16609 17267 16643
rect 21281 16609 21315 16643
rect 25237 16609 25271 16643
rect 2973 16541 3007 16575
rect 6561 16541 6595 16575
rect 13277 16541 13311 16575
rect 13461 16541 13495 16575
rect 17417 16541 17451 16575
rect 18981 16541 19015 16575
rect 21465 16541 21499 16575
rect 22753 16541 22787 16575
rect 16497 16473 16531 16507
rect 21925 16473 21959 16507
rect 2421 16405 2455 16439
rect 5457 16405 5491 16439
rect 12541 16405 12575 16439
rect 16773 16405 16807 16439
rect 18061 16405 18095 16439
rect 18337 16405 18371 16439
rect 24133 16405 24167 16439
rect 3065 16201 3099 16235
rect 5089 16201 5123 16235
rect 6193 16201 6227 16235
rect 8125 16201 8159 16235
rect 10793 16201 10827 16235
rect 12541 16201 12575 16235
rect 13645 16201 13679 16235
rect 15945 16201 15979 16235
rect 16405 16201 16439 16235
rect 17877 16201 17911 16235
rect 19073 16201 19107 16235
rect 19625 16201 19659 16235
rect 20729 16201 20763 16235
rect 22385 16201 22419 16235
rect 22753 16201 22787 16235
rect 23305 16201 23339 16235
rect 23397 16201 23431 16235
rect 23673 16201 23707 16235
rect 24685 16201 24719 16235
rect 25421 16201 25455 16235
rect 5181 16133 5215 16167
rect 12173 16133 12207 16167
rect 17417 16133 17451 16167
rect 21189 16133 21223 16167
rect 26157 16133 26191 16167
rect 2697 16065 2731 16099
rect 4077 16065 4111 16099
rect 4169 16065 4203 16099
rect 5825 16065 5859 16099
rect 8677 16065 8711 16099
rect 8861 16065 8895 16099
rect 10333 16065 10367 16099
rect 11161 16065 11195 16099
rect 11897 16065 11931 16099
rect 13001 16065 13035 16099
rect 13185 16065 13219 16099
rect 14749 16065 14783 16099
rect 15485 16065 15519 16099
rect 17049 16065 17083 16099
rect 18521 16065 18555 16099
rect 18705 16065 18739 16099
rect 20085 16065 20119 16099
rect 20269 16065 20303 16099
rect 21833 16065 21867 16099
rect 23305 16065 23339 16099
rect 24225 16065 24259 16099
rect 1961 15997 1995 16031
rect 6837 15997 6871 16031
rect 7481 15997 7515 16031
rect 8585 15997 8619 16031
rect 9689 15997 9723 16031
rect 10241 15997 10275 16031
rect 18429 15997 18463 16031
rect 19993 15997 20027 16031
rect 21557 15997 21591 16031
rect 24133 15997 24167 16031
rect 25237 15997 25271 16031
rect 25789 15997 25823 16031
rect 2513 15929 2547 15963
rect 5641 15929 5675 15963
rect 9321 15929 9355 15963
rect 10149 15929 10183 15963
rect 11345 15929 11379 15963
rect 12909 15929 12943 15963
rect 14013 15929 14047 15963
rect 15301 15929 15335 15963
rect 2053 15861 2087 15895
rect 2421 15861 2455 15895
rect 3433 15861 3467 15895
rect 3617 15861 3651 15895
rect 3985 15861 4019 15895
rect 4629 15861 4663 15895
rect 5549 15861 5583 15895
rect 6561 15861 6595 15895
rect 7021 15861 7055 15895
rect 8217 15861 8251 15895
rect 9781 15861 9815 15895
rect 14289 15861 14323 15895
rect 14841 15861 14875 15895
rect 15209 15861 15243 15895
rect 16313 15861 16347 15895
rect 16773 15861 16807 15895
rect 16865 15861 16899 15895
rect 18061 15861 18095 15895
rect 19533 15861 19567 15895
rect 21005 15861 21039 15895
rect 21649 15861 21683 15895
rect 24041 15861 24075 15895
rect 25053 15861 25087 15895
rect 3709 15657 3743 15691
rect 6285 15657 6319 15691
rect 7205 15657 7239 15691
rect 7941 15657 7975 15691
rect 8493 15657 8527 15691
rect 9413 15657 9447 15691
rect 9689 15657 9723 15691
rect 10149 15657 10183 15691
rect 13829 15657 13863 15691
rect 14381 15657 14415 15691
rect 14749 15657 14783 15691
rect 15577 15657 15611 15691
rect 17141 15657 17175 15691
rect 17693 15657 17727 15691
rect 18705 15657 18739 15691
rect 19993 15657 20027 15691
rect 21097 15657 21131 15691
rect 24501 15657 24535 15691
rect 25513 15657 25547 15691
rect 2789 15589 2823 15623
rect 4813 15589 4847 15623
rect 5172 15589 5206 15623
rect 7573 15589 7607 15623
rect 11130 15589 11164 15623
rect 12909 15589 12943 15623
rect 13737 15589 13771 15623
rect 19257 15589 19291 15623
rect 19717 15589 19751 15623
rect 21833 15589 21867 15623
rect 24317 15589 24351 15623
rect 1409 15521 1443 15555
rect 2881 15521 2915 15555
rect 4905 15521 4939 15555
rect 8401 15521 8435 15555
rect 10885 15521 10919 15555
rect 15761 15521 15795 15555
rect 16028 15521 16062 15555
rect 18613 15521 18647 15555
rect 19809 15521 19843 15555
rect 20913 15521 20947 15555
rect 22017 15521 22051 15555
rect 22284 15521 22318 15555
rect 24869 15521 24903 15555
rect 3065 15453 3099 15487
rect 4353 15453 4387 15487
rect 8585 15453 8619 15487
rect 14013 15453 14047 15487
rect 18797 15453 18831 15487
rect 20729 15453 20763 15487
rect 24961 15453 24995 15487
rect 25053 15453 25087 15487
rect 1593 15385 1627 15419
rect 8033 15385 8067 15419
rect 13277 15385 13311 15419
rect 18245 15385 18279 15419
rect 21557 15385 21591 15419
rect 2145 15317 2179 15351
rect 2421 15317 2455 15351
rect 9045 15317 9079 15351
rect 10517 15317 10551 15351
rect 12265 15317 12299 15351
rect 13369 15317 13403 15351
rect 18061 15317 18095 15351
rect 20361 15317 20395 15351
rect 23397 15317 23431 15351
rect 24041 15317 24075 15351
rect 7113 15113 7147 15147
rect 8217 15113 8251 15147
rect 8585 15113 8619 15147
rect 10885 15113 10919 15147
rect 13553 15113 13587 15147
rect 14289 15113 14323 15147
rect 17417 15113 17451 15147
rect 17877 15113 17911 15147
rect 20821 15113 20855 15147
rect 22937 15113 22971 15147
rect 23489 15113 23523 15147
rect 25421 15113 25455 15147
rect 26157 15113 26191 15147
rect 1593 15045 1627 15079
rect 3709 15045 3743 15079
rect 14565 15045 14599 15079
rect 21833 15045 21867 15079
rect 25053 15045 25087 15079
rect 3065 14977 3099 15011
rect 3249 14977 3283 15011
rect 7665 14977 7699 15011
rect 11713 14977 11747 15011
rect 12265 14977 12299 15011
rect 13093 14977 13127 15011
rect 13921 14977 13955 15011
rect 21373 14977 21407 15011
rect 21649 14977 21683 15011
rect 22569 14977 22603 15011
rect 24225 14977 24259 15011
rect 1409 14909 1443 14943
rect 2973 14909 3007 14943
rect 4169 14909 4203 14943
rect 4436 14909 4470 14943
rect 7573 14909 7607 14943
rect 8677 14909 8711 14943
rect 14105 14909 14139 14943
rect 15393 14909 15427 14943
rect 15485 14909 15519 14943
rect 18337 14909 18371 14943
rect 19349 14909 19383 14943
rect 19441 14909 19475 14943
rect 22385 14909 22419 14943
rect 24685 14909 24719 14943
rect 25237 14909 25271 14943
rect 25789 14909 25823 14943
rect 2513 14841 2547 14875
rect 4077 14841 4111 14875
rect 6653 14841 6687 14875
rect 7481 14841 7515 14875
rect 8922 14841 8956 14875
rect 12909 14841 12943 14875
rect 15025 14841 15059 14875
rect 15752 14841 15786 14875
rect 18889 14841 18923 14875
rect 19708 14841 19742 14875
rect 21649 14841 21683 14875
rect 24041 14841 24075 14875
rect 2053 14773 2087 14807
rect 2605 14773 2639 14807
rect 5549 14773 5583 14807
rect 6193 14773 6227 14807
rect 10057 14773 10091 14807
rect 11161 14773 11195 14807
rect 12541 14773 12575 14807
rect 13001 14773 13035 14807
rect 16865 14773 16899 14807
rect 18521 14773 18555 14807
rect 21925 14773 21959 14807
rect 22293 14773 22327 14807
rect 23673 14773 23707 14807
rect 24133 14773 24167 14807
rect 1961 14569 1995 14603
rect 2421 14569 2455 14603
rect 3801 14569 3835 14603
rect 6285 14569 6319 14603
rect 7481 14569 7515 14603
rect 7849 14569 7883 14603
rect 11069 14569 11103 14603
rect 11345 14569 11379 14603
rect 13553 14569 13587 14603
rect 14105 14569 14139 14603
rect 14841 14569 14875 14603
rect 16313 14569 16347 14603
rect 18797 14569 18831 14603
rect 21097 14569 21131 14603
rect 21925 14569 21959 14603
rect 23397 14569 23431 14603
rect 24961 14569 24995 14603
rect 2881 14501 2915 14535
rect 3525 14501 3559 14535
rect 4620 14501 4654 14535
rect 12440 14501 12474 14535
rect 14565 14501 14599 14535
rect 16764 14501 16798 14535
rect 20729 14501 20763 14535
rect 1409 14433 1443 14467
rect 2789 14433 2823 14467
rect 4353 14433 4387 14467
rect 6837 14433 6871 14467
rect 8401 14433 8435 14467
rect 10333 14433 10367 14467
rect 11713 14433 11747 14467
rect 16497 14433 16531 14467
rect 19349 14433 19383 14467
rect 20085 14433 20119 14467
rect 20913 14433 20947 14467
rect 22017 14433 22051 14467
rect 22284 14433 22318 14467
rect 23949 14433 23983 14467
rect 24869 14433 24903 14467
rect 2973 14365 3007 14399
rect 8493 14365 8527 14399
rect 8585 14365 8619 14399
rect 10425 14365 10459 14399
rect 10609 14365 10643 14399
rect 12173 14365 12207 14399
rect 15301 14365 15335 14399
rect 19441 14365 19475 14399
rect 19533 14365 19567 14399
rect 25053 14365 25087 14399
rect 7021 14297 7055 14331
rect 8033 14297 8067 14331
rect 15853 14297 15887 14331
rect 18981 14297 19015 14331
rect 21465 14297 21499 14331
rect 24317 14297 24351 14331
rect 1593 14229 1627 14263
rect 2329 14229 2363 14263
rect 5733 14229 5767 14263
rect 6653 14229 6687 14263
rect 9045 14229 9079 14263
rect 9505 14229 9539 14263
rect 9965 14229 9999 14263
rect 17877 14229 17911 14263
rect 18521 14229 18555 14263
rect 24501 14229 24535 14263
rect 25513 14229 25547 14263
rect 3433 14025 3467 14059
rect 9229 14025 9263 14059
rect 9781 14025 9815 14059
rect 11253 14025 11287 14059
rect 12173 14025 12207 14059
rect 12449 14025 12483 14059
rect 13461 14025 13495 14059
rect 15761 14025 15795 14059
rect 16865 14025 16899 14059
rect 17325 14025 17359 14059
rect 19073 14025 19107 14059
rect 20729 14025 20763 14059
rect 21281 14025 21315 14059
rect 21833 14025 21867 14059
rect 22845 14025 22879 14059
rect 23397 14025 23431 14059
rect 24685 14025 24719 14059
rect 25053 14025 25087 14059
rect 25421 14025 25455 14059
rect 1593 13957 1627 13991
rect 3341 13957 3375 13991
rect 4997 13957 5031 13991
rect 8585 13957 8619 13991
rect 23673 13957 23707 13991
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 3893 13889 3927 13923
rect 3985 13889 4019 13923
rect 5641 13889 5675 13923
rect 6009 13889 6043 13923
rect 6929 13889 6963 13923
rect 7205 13889 7239 13923
rect 11897 13889 11931 13923
rect 13093 13889 13127 13923
rect 14565 13889 14599 13923
rect 15393 13889 15427 13923
rect 16405 13889 16439 13923
rect 19349 13889 19383 13923
rect 21741 13889 21775 13923
rect 22385 13889 22419 13923
rect 24225 13889 24259 13923
rect 2053 13821 2087 13855
rect 4905 13821 4939 13855
rect 5457 13821 5491 13855
rect 7461 13821 7495 13855
rect 9873 13821 9907 13855
rect 12909 13821 12943 13855
rect 14473 13821 14507 13855
rect 16221 13821 16255 13855
rect 16313 13821 16347 13855
rect 17785 13821 17819 13855
rect 22201 13821 22235 13855
rect 24133 13821 24167 13855
rect 25237 13821 25271 13855
rect 25789 13821 25823 13855
rect 26249 13821 26283 13855
rect 4537 13753 4571 13787
rect 5365 13753 5399 13787
rect 6929 13753 6963 13787
rect 7021 13753 7055 13787
rect 10118 13753 10152 13787
rect 12817 13753 12851 13787
rect 14381 13753 14415 13787
rect 19594 13753 19628 13787
rect 22293 13753 22327 13787
rect 1961 13685 1995 13719
rect 3801 13685 3835 13719
rect 6561 13685 6595 13719
rect 13921 13685 13955 13719
rect 14013 13685 14047 13719
rect 15853 13685 15887 13719
rect 18337 13685 18371 13719
rect 24041 13685 24075 13719
rect 1685 13481 1719 13515
rect 2329 13481 2363 13515
rect 3249 13481 3283 13515
rect 4721 13481 4755 13515
rect 4905 13481 4939 13515
rect 7849 13481 7883 13515
rect 8769 13481 8803 13515
rect 9505 13481 9539 13515
rect 11621 13481 11655 13515
rect 13921 13481 13955 13515
rect 14565 13481 14599 13515
rect 15853 13481 15887 13515
rect 16405 13481 16439 13515
rect 17325 13481 17359 13515
rect 17877 13481 17911 13515
rect 18245 13481 18279 13515
rect 20913 13481 20947 13515
rect 21281 13481 21315 13515
rect 21373 13481 21407 13515
rect 22569 13481 22603 13515
rect 24593 13481 24627 13515
rect 2973 13413 3007 13447
rect 5365 13413 5399 13447
rect 6714 13413 6748 13447
rect 12541 13413 12575 13447
rect 20361 13413 20395 13447
rect 23029 13413 23063 13447
rect 23673 13413 23707 13447
rect 2237 13345 2271 13379
rect 5273 13345 5307 13379
rect 10057 13345 10091 13379
rect 10701 13345 10735 13379
rect 11069 13345 11103 13379
rect 13185 13345 13219 13379
rect 16313 13345 16347 13379
rect 18593 13345 18627 13379
rect 22385 13345 22419 13379
rect 22937 13345 22971 13379
rect 24501 13345 24535 13379
rect 2513 13277 2547 13311
rect 5457 13277 5491 13311
rect 6469 13277 6503 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 11713 13277 11747 13311
rect 11805 13277 11839 13311
rect 13277 13277 13311 13311
rect 13461 13277 13495 13311
rect 16497 13277 16531 13311
rect 18337 13277 18371 13311
rect 21465 13277 21499 13311
rect 23121 13277 23155 13311
rect 24685 13277 24719 13311
rect 25145 13277 25179 13311
rect 1869 13209 1903 13243
rect 3617 13209 3651 13243
rect 4445 13209 4479 13243
rect 8493 13209 8527 13243
rect 11253 13209 11287 13243
rect 14197 13209 14231 13243
rect 15945 13209 15979 13243
rect 6009 13141 6043 13175
rect 6285 13141 6319 13175
rect 9689 13141 9723 13175
rect 12817 13141 12851 13175
rect 14933 13141 14967 13175
rect 17049 13141 17083 13175
rect 19717 13141 19751 13175
rect 20729 13141 20763 13175
rect 22109 13141 22143 13175
rect 24133 13141 24167 13175
rect 25513 13141 25547 13175
rect 25881 13141 25915 13175
rect 26249 13141 26283 13175
rect 1869 12937 1903 12971
rect 2053 12937 2087 12971
rect 3065 12937 3099 12971
rect 3617 12937 3651 12971
rect 4905 12937 4939 12971
rect 4997 12937 5031 12971
rect 8401 12937 8435 12971
rect 9965 12937 9999 12971
rect 11345 12937 11379 12971
rect 12909 12937 12943 12971
rect 14105 12937 14139 12971
rect 15577 12937 15611 12971
rect 16037 12937 16071 12971
rect 20913 12937 20947 12971
rect 21741 12937 21775 12971
rect 22845 12937 22879 12971
rect 23489 12937 23523 12971
rect 23673 12937 23707 12971
rect 24685 12937 24719 12971
rect 25421 12937 25455 12971
rect 26249 12937 26283 12971
rect 4721 12869 4755 12903
rect 2513 12801 2547 12835
rect 2697 12801 2731 12835
rect 4077 12801 4111 12835
rect 4169 12801 4203 12835
rect 8125 12869 8159 12903
rect 9413 12869 9447 12903
rect 13001 12869 13035 12903
rect 14381 12869 14415 12903
rect 5825 12801 5859 12835
rect 7389 12801 7423 12835
rect 3525 12733 3559 12767
rect 4905 12733 4939 12767
rect 7205 12733 7239 12767
rect 7849 12733 7883 12767
rect 8953 12801 8987 12835
rect 10609 12801 10643 12835
rect 11621 12801 11655 12835
rect 13645 12801 13679 12835
rect 15117 12801 15151 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 17877 12801 17911 12835
rect 21649 12801 21683 12835
rect 22385 12801 22419 12835
rect 24225 12801 24259 12835
rect 14933 12733 14967 12767
rect 16773 12733 16807 12767
rect 17417 12733 17451 12767
rect 18705 12733 18739 12767
rect 25053 12733 25087 12767
rect 25237 12733 25271 12767
rect 25789 12733 25823 12767
rect 5641 12665 5675 12699
rect 8125 12665 8159 12699
rect 8309 12665 8343 12699
rect 8769 12665 8803 12699
rect 10425 12665 10459 12699
rect 12173 12665 12207 12699
rect 18972 12665 19006 12699
rect 22201 12665 22235 12699
rect 24041 12665 24075 12699
rect 2421 12597 2455 12631
rect 3985 12597 4019 12631
rect 5181 12597 5215 12631
rect 5549 12597 5583 12631
rect 6561 12597 6595 12631
rect 6837 12597 6871 12631
rect 7297 12597 7331 12631
rect 8861 12597 8895 12631
rect 9781 12597 9815 12631
rect 10333 12597 10367 12631
rect 13369 12597 13403 12631
rect 13461 12597 13495 12631
rect 14565 12597 14599 12631
rect 15025 12597 15059 12631
rect 16405 12597 16439 12631
rect 18337 12597 18371 12631
rect 20085 12597 20119 12631
rect 22109 12597 22143 12631
rect 24133 12597 24167 12631
rect 1593 12393 1627 12427
rect 2881 12393 2915 12427
rect 4261 12393 4295 12427
rect 6837 12393 6871 12427
rect 8769 12393 8803 12427
rect 9505 12393 9539 12427
rect 9965 12393 9999 12427
rect 14657 12393 14691 12427
rect 16037 12393 16071 12427
rect 16681 12393 16715 12427
rect 18429 12393 18463 12427
rect 20361 12393 20395 12427
rect 21557 12393 21591 12427
rect 22661 12393 22695 12427
rect 23029 12393 23063 12427
rect 23121 12393 23155 12427
rect 24501 12393 24535 12427
rect 24685 12393 24719 12427
rect 2053 12325 2087 12359
rect 5365 12325 5399 12359
rect 14197 12325 14231 12359
rect 17601 12325 17635 12359
rect 19993 12325 20027 12359
rect 21465 12325 21499 12359
rect 26065 12325 26099 12359
rect 1409 12257 1443 12291
rect 2789 12257 2823 12291
rect 4077 12257 4111 12291
rect 4629 12257 4663 12291
rect 5917 12257 5951 12291
rect 7481 12257 7515 12291
rect 7573 12257 7607 12291
rect 10692 12257 10726 12291
rect 13553 12257 13587 12291
rect 16589 12257 16623 12291
rect 17233 12257 17267 12291
rect 19257 12257 19291 12291
rect 21925 12257 21959 12291
rect 23489 12257 23523 12291
rect 25053 12257 25087 12291
rect 25145 12257 25179 12291
rect 3065 12189 3099 12223
rect 3525 12189 3559 12223
rect 5365 12189 5399 12223
rect 6009 12189 6043 12223
rect 6193 12189 6227 12223
rect 7665 12189 7699 12223
rect 8401 12189 8435 12223
rect 10425 12189 10459 12223
rect 13093 12189 13127 12223
rect 13645 12189 13679 12223
rect 13737 12189 13771 12223
rect 16865 12189 16899 12223
rect 17877 12189 17911 12223
rect 19349 12189 19383 12223
rect 19441 12189 19475 12223
rect 20729 12189 20763 12223
rect 22017 12189 22051 12223
rect 22201 12189 22235 12223
rect 23581 12189 23615 12223
rect 23673 12189 23707 12223
rect 24225 12189 24259 12223
rect 25237 12189 25271 12223
rect 3801 12121 3835 12155
rect 12725 12121 12759 12155
rect 2421 12053 2455 12087
rect 5273 12053 5307 12087
rect 5549 12053 5583 12087
rect 7113 12053 7147 12087
rect 11805 12053 11839 12087
rect 13185 12053 13219 12087
rect 14933 12053 14967 12087
rect 15577 12053 15611 12087
rect 16221 12053 16255 12087
rect 18705 12053 18739 12087
rect 18889 12053 18923 12087
rect 25697 12053 25731 12087
rect 1593 11849 1627 11883
rect 2881 11849 2915 11883
rect 5641 11849 5675 11883
rect 6285 11849 6319 11883
rect 8769 11849 8803 11883
rect 9413 11849 9447 11883
rect 9689 11849 9723 11883
rect 14749 11849 14783 11883
rect 20085 11849 20119 11883
rect 20821 11849 20855 11883
rect 21649 11849 21683 11883
rect 22753 11849 22787 11883
rect 25421 11849 25455 11883
rect 26249 11849 26283 11883
rect 2237 11713 2271 11747
rect 2421 11713 2455 11747
rect 2145 11645 2179 11679
rect 3249 11645 3283 11679
rect 3341 11645 3375 11679
rect 6653 11645 6687 11679
rect 6837 11645 6871 11679
rect 3608 11577 3642 11611
rect 7104 11577 7138 11611
rect 19441 11781 19475 11815
rect 23673 11781 23707 11815
rect 25789 11781 25823 11815
rect 9781 11713 9815 11747
rect 12449 11713 12483 11747
rect 22293 11713 22327 11747
rect 23029 11713 23063 11747
rect 24317 11713 24351 11747
rect 15393 11645 15427 11679
rect 15485 11645 15519 11679
rect 17785 11645 17819 11679
rect 18061 11645 18095 11679
rect 20637 11645 20671 11679
rect 25053 11645 25087 11679
rect 25237 11645 25271 11679
rect 10026 11577 10060 11611
rect 12694 11577 12728 11611
rect 14381 11577 14415 11611
rect 15730 11577 15764 11611
rect 18306 11577 18340 11611
rect 20361 11577 20395 11611
rect 21465 11577 21499 11611
rect 22017 11577 22051 11611
rect 1777 11509 1811 11543
rect 4721 11509 4755 11543
rect 8217 11509 8251 11543
rect 9229 11509 9263 11543
rect 9413 11509 9447 11543
rect 11161 11509 11195 11543
rect 11713 11509 11747 11543
rect 12265 11509 12299 11543
rect 13829 11509 13863 11543
rect 16865 11509 16899 11543
rect 17417 11509 17451 11543
rect 21097 11509 21131 11543
rect 22109 11509 22143 11543
rect 23489 11509 23523 11543
rect 24041 11509 24075 11543
rect 24133 11509 24167 11543
rect 24777 11509 24811 11543
rect 1961 11305 1995 11339
rect 2329 11305 2363 11339
rect 2789 11305 2823 11339
rect 2881 11305 2915 11339
rect 3525 11305 3559 11339
rect 4353 11305 4387 11339
rect 6469 11305 6503 11339
rect 6929 11305 6963 11339
rect 7297 11305 7331 11339
rect 7757 11305 7791 11339
rect 8309 11305 8343 11339
rect 10241 11305 10275 11339
rect 11529 11305 11563 11339
rect 11897 11305 11931 11339
rect 14105 11305 14139 11339
rect 15485 11305 15519 11339
rect 15761 11305 15795 11339
rect 16313 11305 16347 11339
rect 17969 11305 18003 11339
rect 18521 11305 18555 11339
rect 19533 11305 19567 11339
rect 20913 11305 20947 11339
rect 21281 11305 21315 11339
rect 21925 11305 21959 11339
rect 22477 11305 22511 11339
rect 22937 11305 22971 11339
rect 24041 11305 24075 11339
rect 24409 11305 24443 11339
rect 24501 11305 24535 11339
rect 25145 11305 25179 11339
rect 25789 11305 25823 11339
rect 12992 11237 13026 11271
rect 14657 11237 14691 11271
rect 21373 11237 21407 11271
rect 25421 11237 25455 11271
rect 1409 11169 1443 11203
rect 4537 11169 4571 11203
rect 4793 11169 4827 11203
rect 8217 11169 8251 11203
rect 10885 11169 10919 11203
rect 12725 11169 12759 11203
rect 15301 11169 15335 11203
rect 16856 11169 16890 11203
rect 19441 11169 19475 11203
rect 22385 11169 22419 11203
rect 22845 11169 22879 11203
rect 3065 11101 3099 11135
rect 8401 11101 8435 11135
rect 10977 11101 11011 11135
rect 11161 11101 11195 11135
rect 12449 11101 12483 11135
rect 16589 11101 16623 11135
rect 19625 11101 19659 11135
rect 21465 11101 21499 11135
rect 23121 11101 23155 11135
rect 24593 11101 24627 11135
rect 1593 11033 1627 11067
rect 2421 11033 2455 11067
rect 5917 11033 5951 11067
rect 7849 11033 7883 11067
rect 10517 11033 10551 11067
rect 15025 11033 15059 11067
rect 18889 11033 18923 11067
rect 19073 11033 19107 11067
rect 3893 10965 3927 10999
rect 9229 10965 9263 10999
rect 9965 10965 9999 10999
rect 20085 10965 20119 10999
rect 20729 10965 20763 10999
rect 23765 10965 23799 10999
rect 26157 10965 26191 10999
rect 1593 10761 1627 10795
rect 4997 10761 5031 10795
rect 5181 10761 5215 10795
rect 6193 10761 6227 10795
rect 6561 10761 6595 10795
rect 9137 10761 9171 10795
rect 12449 10761 12483 10795
rect 16681 10761 16715 10795
rect 20729 10761 20763 10795
rect 22201 10761 22235 10795
rect 22661 10761 22695 10795
rect 23305 10761 23339 10795
rect 24409 10761 24443 10795
rect 25513 10761 25547 10795
rect 4629 10693 4663 10727
rect 7297 10693 7331 10727
rect 15669 10693 15703 10727
rect 19625 10693 19659 10727
rect 24777 10693 24811 10727
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 7849 10625 7883 10659
rect 9689 10625 9723 10659
rect 10241 10625 10275 10659
rect 10609 10625 10643 10659
rect 11253 10625 11287 10659
rect 12081 10625 12115 10659
rect 13093 10625 13127 10659
rect 13553 10625 13587 10659
rect 18521 10625 18555 10659
rect 18705 10625 18739 10659
rect 19533 10625 19567 10659
rect 20269 10625 20303 10659
rect 21741 10625 21775 10659
rect 25881 10625 25915 10659
rect 1409 10557 1443 10591
rect 2605 10557 2639 10591
rect 2697 10557 2731 10591
rect 5549 10557 5583 10591
rect 7205 10557 7239 10591
rect 7757 10557 7791 10591
rect 8953 10557 8987 10591
rect 9597 10557 9631 10591
rect 11161 10557 11195 10591
rect 2964 10489 2998 10523
rect 7665 10489 7699 10523
rect 8401 10489 8435 10523
rect 12909 10557 12943 10591
rect 14197 10557 14231 10591
rect 14289 10557 14323 10591
rect 14545 10557 14579 10591
rect 16773 10557 16807 10591
rect 17509 10557 17543 10591
rect 19993 10557 20027 10591
rect 21557 10557 21591 10591
rect 24593 10557 24627 10591
rect 25145 10557 25179 10591
rect 12817 10489 12851 10523
rect 17785 10489 17819 10523
rect 18429 10489 18463 10523
rect 21097 10489 21131 10523
rect 21649 10489 21683 10523
rect 24041 10489 24075 10523
rect 2053 10421 2087 10455
rect 4077 10421 4111 10455
rect 9505 10421 9539 10455
rect 10701 10421 10735 10455
rect 11069 10421 11103 10455
rect 11897 10421 11931 10455
rect 12081 10421 12115 10455
rect 12173 10421 12207 10455
rect 16221 10421 16255 10455
rect 18061 10421 18095 10455
rect 19073 10421 19107 10455
rect 20085 10421 20119 10455
rect 21189 10421 21223 10455
rect 22937 10421 22971 10455
rect 26341 10421 26375 10455
rect 2329 10217 2363 10251
rect 4077 10217 4111 10251
rect 4445 10217 4479 10251
rect 4537 10217 4571 10251
rect 5181 10217 5215 10251
rect 5641 10217 5675 10251
rect 5917 10217 5951 10251
rect 7757 10217 7791 10251
rect 8125 10217 8159 10251
rect 8769 10217 8803 10251
rect 9873 10217 9907 10251
rect 10149 10217 10183 10251
rect 11345 10217 11379 10251
rect 12449 10217 12483 10251
rect 13829 10217 13863 10251
rect 14657 10217 14691 10251
rect 15485 10217 15519 10251
rect 16957 10217 16991 10251
rect 17509 10217 17543 10251
rect 17969 10217 18003 10251
rect 18521 10217 18555 10251
rect 18889 10217 18923 10251
rect 19441 10217 19475 10251
rect 21925 10217 21959 10251
rect 22293 10217 22327 10251
rect 23029 10217 23063 10251
rect 23489 10217 23523 10251
rect 23765 10217 23799 10251
rect 24501 10217 24535 10251
rect 25513 10217 25547 10251
rect 25881 10217 25915 10251
rect 26341 10217 26375 10251
rect 2789 10149 2823 10183
rect 7389 10149 7423 10183
rect 10701 10149 10735 10183
rect 17325 10149 17359 10183
rect 24041 10149 24075 10183
rect 2881 10081 2915 10115
rect 6561 10081 6595 10115
rect 9689 10081 9723 10115
rect 11253 10081 11287 10115
rect 11897 10081 11931 10115
rect 12817 10081 12851 10115
rect 14197 10081 14231 10115
rect 16313 10081 16347 10115
rect 17877 10081 17911 10115
rect 21281 10081 21315 10115
rect 21373 10081 21407 10115
rect 22569 10081 22603 10115
rect 23581 10081 23615 10115
rect 24593 10081 24627 10115
rect 25145 10081 25179 10115
rect 2973 10013 3007 10047
rect 4629 10013 4663 10047
rect 6653 10013 6687 10047
rect 6745 10013 6779 10047
rect 8217 10013 8251 10047
rect 8401 10013 8435 10047
rect 11437 10013 11471 10047
rect 12357 10013 12391 10047
rect 12909 10013 12943 10047
rect 13093 10013 13127 10047
rect 16405 10013 16439 10047
rect 16589 10013 16623 10047
rect 18061 10013 18095 10047
rect 19533 10013 19567 10047
rect 19717 10013 19751 10047
rect 21557 10013 21591 10047
rect 2421 9945 2455 9979
rect 6193 9945 6227 9979
rect 10885 9945 10919 9979
rect 15025 9945 15059 9979
rect 15945 9945 15979 9979
rect 22753 9945 22787 9979
rect 24777 9945 24811 9979
rect 1961 9877 1995 9911
rect 3525 9877 3559 9911
rect 3801 9877 3835 9911
rect 9137 9877 9171 9911
rect 13461 9877 13495 9911
rect 19073 9877 19107 9911
rect 20085 9877 20119 9911
rect 20729 9877 20763 9911
rect 20913 9877 20947 9911
rect 5917 9673 5951 9707
rect 8217 9673 8251 9707
rect 11069 9673 11103 9707
rect 11345 9673 11379 9707
rect 12449 9673 12483 9707
rect 15209 9673 15243 9707
rect 18061 9673 18095 9707
rect 20913 9673 20947 9707
rect 22661 9673 22695 9707
rect 22937 9673 22971 9707
rect 23857 9673 23891 9707
rect 24409 9673 24443 9707
rect 7113 9605 7147 9639
rect 12081 9605 12115 9639
rect 13829 9605 13863 9639
rect 16681 9605 16715 9639
rect 19073 9605 19107 9639
rect 19257 9605 19291 9639
rect 19441 9605 19475 9639
rect 21189 9605 21223 9639
rect 24777 9605 24811 9639
rect 25881 9605 25915 9639
rect 26341 9605 26375 9639
rect 1685 9537 1719 9571
rect 2421 9537 2455 9571
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 7665 9537 7699 9571
rect 8493 9537 8527 9571
rect 11897 9537 11931 9571
rect 6285 9469 6319 9503
rect 7481 9469 7515 9503
rect 9045 9469 9079 9503
rect 2237 9401 2271 9435
rect 2789 9401 2823 9435
rect 3608 9401 3642 9435
rect 5273 9401 5307 9435
rect 9312 9401 9346 9435
rect 13001 9537 13035 9571
rect 13461 9537 13495 9571
rect 14841 9537 14875 9571
rect 15853 9537 15887 9571
rect 16405 9537 16439 9571
rect 18613 9537 18647 9571
rect 14013 9469 14047 9503
rect 16865 9469 16899 9503
rect 12909 9401 12943 9435
rect 17877 9401 17911 9435
rect 20269 9537 20303 9571
rect 21649 9537 21683 9571
rect 21833 9537 21867 9571
rect 22201 9537 22235 9571
rect 25145 9537 25179 9571
rect 19993 9469 20027 9503
rect 21557 9469 21591 9503
rect 24593 9469 24627 9503
rect 25513 9469 25547 9503
rect 1777 9333 1811 9367
rect 2145 9333 2179 9367
rect 4721 9333 4755 9367
rect 6561 9333 6595 9367
rect 7573 9333 7607 9367
rect 8861 9333 8895 9367
rect 10425 9333 10459 9367
rect 12081 9333 12115 9367
rect 12173 9333 12207 9367
rect 12817 9333 12851 9367
rect 15301 9333 15335 9367
rect 15669 9333 15703 9367
rect 15761 9333 15795 9367
rect 17417 9333 17451 9367
rect 18429 9333 18463 9367
rect 18521 9333 18555 9367
rect 19257 9333 19291 9367
rect 19625 9333 19659 9367
rect 20085 9333 20119 9367
rect 23305 9333 23339 9367
rect 2237 9129 2271 9163
rect 2421 9129 2455 9163
rect 4353 9129 4387 9163
rect 4629 9129 4663 9163
rect 5365 9129 5399 9163
rect 8401 9129 8435 9163
rect 9137 9129 9171 9163
rect 13645 9129 13679 9163
rect 14565 9129 14599 9163
rect 15117 9129 15151 9163
rect 20729 9129 20763 9163
rect 20913 9129 20947 9163
rect 21373 9129 21407 9163
rect 21925 9129 21959 9163
rect 23305 9129 23339 9163
rect 24409 9129 24443 9163
rect 24777 9129 24811 9163
rect 25881 9129 25915 9163
rect 2789 9061 2823 9095
rect 5273 9061 5307 9095
rect 9413 9061 9447 9095
rect 10946 9061 10980 9095
rect 13553 9061 13587 9095
rect 14197 9061 14231 9095
rect 15546 9061 15580 9095
rect 21281 9061 21315 9095
rect 24041 9061 24075 9095
rect 2881 8993 2915 9027
rect 6469 8993 6503 9027
rect 6736 8993 6770 9027
rect 10701 8993 10735 9027
rect 18153 8993 18187 9027
rect 19717 8993 19751 9027
rect 22477 8993 22511 9027
rect 23581 8993 23615 9027
rect 24593 8993 24627 9027
rect 25145 8993 25179 9027
rect 1409 8925 1443 8959
rect 2973 8925 3007 8959
rect 3433 8925 3467 8959
rect 5549 8925 5583 8959
rect 9689 8925 9723 8959
rect 12633 8925 12667 8959
rect 13737 8925 13771 8959
rect 15301 8925 15335 8959
rect 17325 8925 17359 8959
rect 18245 8925 18279 8959
rect 18337 8925 18371 8959
rect 19441 8925 19475 8959
rect 20269 8925 20303 8959
rect 21465 8925 21499 8959
rect 22937 8925 22971 8959
rect 6009 8857 6043 8891
rect 13185 8857 13219 8891
rect 17693 8857 17727 8891
rect 22661 8857 22695 8891
rect 23765 8857 23799 8891
rect 1869 8789 1903 8823
rect 3893 8789 3927 8823
rect 4905 8789 4939 8823
rect 6285 8789 6319 8823
rect 7849 8789 7883 8823
rect 10333 8789 10367 8823
rect 12081 8789 12115 8823
rect 13093 8789 13127 8823
rect 16681 8789 16715 8823
rect 17785 8789 17819 8823
rect 19073 8789 19107 8823
rect 19901 8789 19935 8823
rect 22293 8789 22327 8823
rect 25605 8789 25639 8823
rect 26249 8789 26283 8823
rect 1593 8585 1627 8619
rect 2881 8585 2915 8619
rect 4261 8585 4295 8619
rect 7205 8585 7239 8619
rect 9045 8585 9079 8619
rect 9689 8585 9723 8619
rect 10241 8585 10275 8619
rect 11253 8585 11287 8619
rect 12173 8585 12207 8619
rect 12817 8585 12851 8619
rect 14657 8585 14691 8619
rect 15761 8585 15795 8619
rect 20085 8585 20119 8619
rect 20545 8585 20579 8619
rect 21557 8585 21591 8619
rect 24501 8585 24535 8619
rect 25513 8585 25547 8619
rect 25973 8585 26007 8619
rect 26341 8585 26375 8619
rect 2513 8517 2547 8551
rect 4445 8517 4479 8551
rect 13093 8517 13127 8551
rect 16773 8517 16807 8551
rect 17785 8517 17819 8551
rect 19441 8517 19475 8551
rect 20361 8517 20395 8551
rect 22293 8517 22327 8551
rect 24869 8517 24903 8551
rect 3341 8449 3375 8483
rect 3525 8449 3559 8483
rect 4997 8449 5031 8483
rect 5457 8449 5491 8483
rect 7481 8449 7515 8483
rect 7665 8449 7699 8483
rect 10793 8449 10827 8483
rect 16313 8449 16347 8483
rect 18061 8449 18095 8483
rect 21005 8449 21039 8483
rect 21097 8449 21131 8483
rect 23489 8449 23523 8483
rect 1409 8381 1443 8415
rect 4813 8381 4847 8415
rect 4905 8381 4939 8415
rect 6469 8381 6503 8415
rect 10609 8381 10643 8415
rect 13277 8381 13311 8415
rect 16129 8381 16163 8415
rect 20913 8381 20947 8415
rect 21925 8381 21959 8415
rect 22109 8381 22143 8415
rect 22661 8381 22695 8415
rect 23029 8381 23063 8415
rect 23673 8381 23707 8415
rect 24133 8381 24167 8415
rect 24685 8381 24719 8415
rect 2145 8313 2179 8347
rect 3985 8313 4019 8347
rect 7910 8313 7944 8347
rect 10701 8313 10735 8347
rect 11621 8313 11655 8347
rect 13544 8313 13578 8347
rect 15209 8313 15243 8347
rect 15577 8313 15611 8347
rect 16221 8313 16255 8347
rect 17509 8313 17543 8347
rect 18328 8313 18362 8347
rect 25145 8313 25179 8347
rect 3249 8245 3283 8279
rect 6193 8245 6227 8279
rect 10149 8245 10183 8279
rect 23857 8245 23891 8279
rect 2237 8041 2271 8075
rect 2421 8041 2455 8075
rect 2789 8041 2823 8075
rect 3433 8041 3467 8075
rect 4261 8041 4295 8075
rect 4721 8041 4755 8075
rect 9505 8041 9539 8075
rect 9781 8041 9815 8075
rect 10149 8041 10183 8075
rect 10241 8041 10275 8075
rect 11621 8041 11655 8075
rect 13829 8041 13863 8075
rect 14197 8041 14231 8075
rect 15117 8041 15151 8075
rect 16681 8041 16715 8075
rect 17785 8041 17819 8075
rect 19165 8041 19199 8075
rect 20269 8041 20303 8075
rect 22937 8041 22971 8075
rect 2881 7973 2915 8007
rect 4997 7973 5031 8007
rect 5540 7973 5574 8007
rect 7757 7973 7791 8007
rect 10793 7973 10827 8007
rect 12142 7973 12176 8007
rect 4077 7905 4111 7939
rect 5273 7905 5307 7939
rect 8401 7905 8435 7939
rect 11897 7905 11931 7939
rect 15301 7905 15335 7939
rect 15568 7905 15602 7939
rect 17601 7905 17635 7939
rect 18153 7905 18187 7939
rect 18245 7905 18279 7939
rect 19349 7905 19383 7939
rect 19901 7905 19935 7939
rect 21281 7905 21315 7939
rect 22201 7905 22235 7939
rect 22385 7905 22419 7939
rect 22845 7905 22879 7939
rect 24041 7905 24075 7939
rect 25145 7905 25179 7939
rect 1409 7837 1443 7871
rect 2973 7837 3007 7871
rect 8493 7837 8527 7871
rect 8585 7837 8619 7871
rect 10333 7837 10367 7871
rect 18337 7837 18371 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 23029 7837 23063 7871
rect 24593 7837 24627 7871
rect 7389 7769 7423 7803
rect 9137 7769 9171 7803
rect 18797 7769 18831 7803
rect 20913 7769 20947 7803
rect 22201 7769 22235 7803
rect 24225 7769 24259 7803
rect 1869 7701 1903 7735
rect 3801 7701 3835 7735
rect 6653 7701 6687 7735
rect 8033 7701 8067 7735
rect 11253 7701 11287 7735
rect 13277 7701 13311 7735
rect 14657 7701 14691 7735
rect 17233 7701 17267 7735
rect 19533 7701 19567 7735
rect 20729 7701 20763 7735
rect 21925 7701 21959 7735
rect 22477 7701 22511 7735
rect 23489 7701 23523 7735
rect 23949 7701 23983 7735
rect 24961 7701 24995 7735
rect 25329 7701 25363 7735
rect 25697 7701 25731 7735
rect 26065 7701 26099 7735
rect 1593 7497 1627 7531
rect 3157 7497 3191 7531
rect 4629 7497 4663 7531
rect 6193 7497 6227 7531
rect 7665 7497 7699 7531
rect 8677 7497 8711 7531
rect 10333 7497 10367 7531
rect 11897 7497 11931 7531
rect 13093 7497 13127 7531
rect 13277 7497 13311 7531
rect 15393 7497 15427 7531
rect 15853 7497 15887 7531
rect 17141 7497 17175 7531
rect 18153 7497 18187 7531
rect 19441 7497 19475 7531
rect 19717 7497 19751 7531
rect 21281 7497 21315 7531
rect 22845 7497 22879 7531
rect 23213 7497 23247 7531
rect 24685 7497 24719 7531
rect 25329 7497 25363 7531
rect 25789 7497 25823 7531
rect 26065 7497 26099 7531
rect 7205 7429 7239 7463
rect 10609 7429 10643 7463
rect 2053 7361 2087 7395
rect 2237 7361 2271 7395
rect 3065 7361 3099 7395
rect 3801 7361 3835 7395
rect 5273 7361 5307 7395
rect 8217 7361 8251 7395
rect 9873 7361 9907 7395
rect 11437 7361 11471 7395
rect 12909 7361 12943 7395
rect 21189 7429 21223 7463
rect 24225 7429 24259 7463
rect 15761 7361 15795 7395
rect 16405 7361 16439 7395
rect 18705 7361 18739 7395
rect 20269 7361 20303 7395
rect 3617 7293 3651 7327
rect 5089 7293 5123 7327
rect 9137 7293 9171 7327
rect 9689 7293 9723 7327
rect 11161 7293 11195 7327
rect 13093 7293 13127 7327
rect 13369 7293 13403 7327
rect 13636 7293 13670 7327
rect 17509 7293 17543 7327
rect 18521 7293 18555 7327
rect 20085 7293 20119 7327
rect 21833 7361 21867 7395
rect 23673 7293 23707 7327
rect 24777 7293 24811 7327
rect 26433 7293 26467 7327
rect 1961 7225 1995 7259
rect 3525 7225 3559 7259
rect 4261 7225 4295 7259
rect 5733 7225 5767 7259
rect 6653 7225 6687 7259
rect 8033 7225 8067 7259
rect 11253 7225 11287 7259
rect 20177 7225 20211 7259
rect 21189 7225 21223 7259
rect 21649 7225 21683 7259
rect 2605 7157 2639 7191
rect 4721 7157 4755 7191
rect 5181 7157 5215 7191
rect 7481 7157 7515 7191
rect 8125 7157 8159 7191
rect 9229 7157 9263 7191
rect 9597 7157 9631 7191
rect 10793 7157 10827 7191
rect 14749 7157 14783 7191
rect 16221 7157 16255 7191
rect 16313 7157 16347 7191
rect 17877 7157 17911 7191
rect 18613 7157 18647 7191
rect 21005 7157 21039 7191
rect 21741 7157 21775 7191
rect 22569 7157 22603 7191
rect 23857 7157 23891 7191
rect 24961 7157 24995 7191
rect 2421 6953 2455 6987
rect 2789 6953 2823 6987
rect 4445 6953 4479 6987
rect 6469 6953 6503 6987
rect 9229 6953 9263 6987
rect 9965 6953 9999 6987
rect 12265 6953 12299 6987
rect 18613 6953 18647 6987
rect 19625 6953 19659 6987
rect 21281 6953 21315 6987
rect 22845 6953 22879 6987
rect 24777 6953 24811 6987
rect 1685 6885 1719 6919
rect 8401 6885 8435 6919
rect 13185 6885 13219 6919
rect 2881 6817 2915 6851
rect 4537 6817 4571 6851
rect 5825 6817 5859 6851
rect 7757 6817 7791 6851
rect 10600 6817 10634 6851
rect 15025 6817 15059 6851
rect 15577 6817 15611 6851
rect 16681 6817 16715 6851
rect 16937 6817 16971 6851
rect 19533 6817 19567 6851
rect 21373 6817 21407 6851
rect 22385 6817 22419 6851
rect 22937 6817 22971 6851
rect 23673 6817 23707 6851
rect 24041 6817 24075 6851
rect 25145 6817 25179 6851
rect 2973 6749 3007 6783
rect 4629 6749 4663 6783
rect 6561 6749 6595 6783
rect 6653 6749 6687 6783
rect 8493 6749 8527 6783
rect 8677 6749 8711 6783
rect 10333 6749 10367 6783
rect 13277 6749 13311 6783
rect 13369 6749 13403 6783
rect 13921 6749 13955 6783
rect 18981 6749 19015 6783
rect 19717 6749 19751 6783
rect 21465 6749 21499 6783
rect 23121 6749 23155 6783
rect 3801 6681 3835 6715
rect 5549 6681 5583 6715
rect 6101 6681 6135 6715
rect 7389 6681 7423 6715
rect 12817 6681 12851 6715
rect 14381 6681 14415 6715
rect 20913 6681 20947 6715
rect 22477 6681 22511 6715
rect 2329 6613 2363 6647
rect 3433 6613 3467 6647
rect 4077 6613 4111 6647
rect 5181 6613 5215 6647
rect 8033 6613 8067 6647
rect 11713 6613 11747 6647
rect 12725 6613 12759 6647
rect 14749 6613 14783 6647
rect 15761 6613 15795 6647
rect 16129 6613 16163 6647
rect 16589 6613 16623 6647
rect 18061 6613 18095 6647
rect 19165 6613 19199 6647
rect 20177 6613 20211 6647
rect 20729 6613 20763 6647
rect 22017 6613 22051 6647
rect 24225 6613 24259 6647
rect 25329 6613 25363 6647
rect 25697 6613 25731 6647
rect 26065 6613 26099 6647
rect 2053 6409 2087 6443
rect 2237 6409 2271 6443
rect 3249 6409 3283 6443
rect 6101 6409 6135 6443
rect 6561 6409 6595 6443
rect 7297 6409 7331 6443
rect 10425 6409 10459 6443
rect 11621 6409 11655 6443
rect 16405 6409 16439 6443
rect 18061 6409 18095 6443
rect 21005 6409 21039 6443
rect 21189 6409 21223 6443
rect 24685 6409 24719 6443
rect 25145 6409 25179 6443
rect 25789 6409 25823 6443
rect 1777 6341 1811 6375
rect 5825 6341 5859 6375
rect 10057 6341 10091 6375
rect 19073 6341 19107 6375
rect 2789 6273 2823 6307
rect 7481 6273 7515 6307
rect 7757 6273 7791 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11989 6273 12023 6307
rect 16313 6273 16347 6307
rect 17049 6273 17083 6307
rect 18705 6273 18739 6307
rect 20177 6273 20211 6307
rect 21741 6273 21775 6307
rect 24225 6273 24259 6307
rect 2605 6205 2639 6239
rect 3801 6205 3835 6239
rect 10885 6205 10919 6239
rect 13001 6205 13035 6239
rect 13268 6205 13302 6239
rect 16865 6205 16899 6239
rect 21557 6205 21591 6239
rect 23029 6205 23063 6239
rect 25237 6205 25271 6239
rect 4046 6137 4080 6171
rect 7481 6137 7515 6171
rect 7573 6137 7607 6171
rect 8024 6137 8058 6171
rect 15761 6137 15795 6171
rect 16773 6137 16807 6171
rect 17785 6137 17819 6171
rect 18429 6137 18463 6171
rect 19441 6137 19475 6171
rect 20085 6137 20119 6171
rect 22293 6137 22327 6171
rect 22661 6137 22695 6171
rect 23489 6137 23523 6171
rect 24041 6137 24075 6171
rect 24133 6137 24167 6171
rect 2697 6069 2731 6103
rect 3617 6069 3651 6103
rect 5181 6069 5215 6103
rect 9137 6069 9171 6103
rect 10517 6069 10551 6103
rect 12817 6069 12851 6103
rect 14381 6069 14415 6103
rect 14933 6069 14967 6103
rect 15393 6069 15427 6103
rect 17417 6069 17451 6103
rect 18521 6069 18555 6103
rect 19625 6069 19659 6103
rect 19993 6069 20027 6103
rect 21649 6069 21683 6103
rect 23673 6069 23707 6103
rect 25421 6069 25455 6103
rect 26249 6069 26283 6103
rect 2421 5865 2455 5899
rect 2789 5865 2823 5899
rect 5181 5865 5215 5899
rect 5273 5865 5307 5899
rect 6285 5865 6319 5899
rect 6745 5865 6779 5899
rect 8217 5865 8251 5899
rect 8769 5865 8803 5899
rect 12633 5865 12667 5899
rect 14105 5865 14139 5899
rect 15301 5865 15335 5899
rect 15761 5865 15795 5899
rect 16405 5865 16439 5899
rect 16773 5865 16807 5899
rect 19349 5865 19383 5899
rect 21373 5865 21407 5899
rect 22293 5865 22327 5899
rect 22937 5865 22971 5899
rect 24409 5865 24443 5899
rect 25421 5865 25455 5899
rect 9505 5797 9539 5831
rect 17202 5797 17236 5831
rect 18889 5797 18923 5831
rect 22845 5797 22879 5831
rect 24501 5797 24535 5831
rect 25053 5797 25087 5831
rect 25789 5797 25823 5831
rect 2329 5729 2363 5763
rect 5641 5729 5675 5763
rect 7104 5729 7138 5763
rect 9945 5729 9979 5763
rect 12981 5729 13015 5763
rect 15669 5729 15703 5763
rect 19441 5729 19475 5763
rect 21281 5729 21315 5763
rect 2881 5661 2915 5695
rect 3065 5661 3099 5695
rect 3801 5661 3835 5695
rect 4261 5661 4295 5695
rect 5733 5661 5767 5695
rect 5917 5661 5951 5695
rect 6837 5661 6871 5695
rect 9689 5661 9723 5695
rect 12173 5661 12207 5695
rect 12725 5661 12759 5695
rect 15117 5661 15151 5695
rect 15853 5661 15887 5695
rect 16957 5661 16991 5695
rect 21465 5661 21499 5695
rect 23029 5661 23063 5695
rect 24685 5661 24719 5695
rect 4813 5593 4847 5627
rect 18337 5593 18371 5627
rect 20913 5593 20947 5627
rect 22477 5593 22511 5627
rect 24041 5593 24075 5627
rect 1961 5525 1995 5559
rect 3433 5525 3467 5559
rect 11069 5525 11103 5559
rect 11713 5525 11747 5559
rect 14749 5525 14783 5559
rect 19625 5525 19659 5559
rect 19993 5525 20027 5559
rect 20729 5525 20763 5559
rect 21925 5525 21959 5559
rect 23673 5525 23707 5559
rect 26249 5525 26283 5559
rect 5181 5321 5215 5355
rect 6285 5321 6319 5355
rect 7297 5321 7331 5355
rect 10425 5321 10459 5355
rect 12265 5321 12299 5355
rect 13829 5321 13863 5355
rect 14933 5321 14967 5355
rect 15301 5321 15335 5355
rect 17785 5321 17819 5355
rect 19625 5321 19659 5355
rect 22937 5321 22971 5355
rect 23673 5321 23707 5355
rect 24685 5321 24719 5355
rect 25881 5321 25915 5355
rect 13921 5253 13955 5287
rect 22569 5253 22603 5287
rect 26249 5253 26283 5287
rect 1777 5185 1811 5219
rect 2605 5185 2639 5219
rect 5089 5185 5123 5219
rect 5825 5185 5859 5219
rect 8309 5185 8343 5219
rect 8769 5185 8803 5219
rect 10977 5185 11011 5219
rect 11437 5185 11471 5219
rect 14565 5185 14599 5219
rect 18613 5185 18647 5219
rect 20177 5185 20211 5219
rect 20637 5185 20671 5219
rect 21741 5185 21775 5219
rect 24225 5185 24259 5219
rect 4721 5117 4755 5151
rect 5641 5117 5675 5151
rect 9137 5117 9171 5151
rect 9321 5117 9355 5151
rect 10333 5117 10367 5151
rect 12817 5117 12851 5151
rect 14289 5117 14323 5151
rect 15485 5117 15519 5151
rect 17417 5117 17451 5151
rect 19533 5117 19567 5151
rect 20085 5117 20119 5151
rect 21557 5117 21591 5151
rect 24041 5117 24075 5151
rect 25237 5117 25271 5151
rect 2145 5049 2179 5083
rect 2872 5049 2906 5083
rect 5549 5049 5583 5083
rect 7665 5049 7699 5083
rect 8125 5049 8159 5083
rect 9965 5049 9999 5083
rect 10885 5049 10919 5083
rect 13461 5049 13495 5083
rect 15752 5049 15786 5083
rect 21649 5049 21683 5083
rect 2421 4981 2455 5015
rect 3985 4981 4019 5015
rect 6561 4981 6595 5015
rect 7757 4981 7791 5015
rect 8217 4981 8251 5015
rect 10793 4981 10827 5015
rect 11897 4981 11931 5015
rect 12633 4981 12667 5015
rect 13001 4981 13035 5015
rect 14381 4981 14415 5015
rect 16865 4981 16899 5015
rect 18061 4981 18095 5015
rect 18429 4981 18463 5015
rect 18521 4981 18555 5015
rect 19073 4981 19107 5015
rect 19993 4981 20027 5015
rect 21005 4981 21039 5015
rect 21189 4981 21223 5015
rect 23489 4981 23523 5015
rect 24133 4981 24167 5015
rect 25053 4981 25087 5015
rect 25421 4981 25455 5015
rect 1961 4777 1995 4811
rect 2421 4777 2455 4811
rect 2881 4777 2915 4811
rect 3249 4777 3283 4811
rect 3525 4777 3559 4811
rect 8585 4777 8619 4811
rect 10241 4777 10275 4811
rect 11805 4777 11839 4811
rect 14105 4777 14139 4811
rect 15025 4777 15059 4811
rect 15669 4777 15703 4811
rect 16865 4777 16899 4811
rect 18153 4777 18187 4811
rect 18429 4777 18463 4811
rect 18797 4777 18831 4811
rect 18889 4777 18923 4811
rect 19625 4777 19659 4811
rect 20085 4777 20119 4811
rect 20361 4777 20395 4811
rect 22385 4777 22419 4811
rect 23765 4777 23799 4811
rect 24133 4777 24167 4811
rect 1409 4641 1443 4675
rect 2789 4641 2823 4675
rect 4322 4709 4356 4743
rect 9965 4709 9999 4743
rect 14749 4709 14783 4743
rect 15761 4709 15795 4743
rect 21833 4709 21867 4743
rect 21925 4709 21959 4743
rect 6469 4641 6503 4675
rect 6828 4641 6862 4675
rect 10609 4641 10643 4675
rect 12173 4641 12207 4675
rect 12265 4641 12299 4675
rect 14013 4641 14047 4675
rect 16773 4641 16807 4675
rect 17233 4641 17267 4675
rect 21281 4641 21315 4675
rect 3065 4573 3099 4607
rect 3249 4573 3283 4607
rect 4077 4573 4111 4607
rect 6561 4573 6595 4607
rect 10701 4573 10735 4607
rect 10793 4573 10827 4607
rect 12357 4573 12391 4607
rect 13185 4573 13219 4607
rect 14289 4573 14323 4607
rect 15945 4573 15979 4607
rect 17325 4573 17359 4607
rect 17509 4573 17543 4607
rect 18981 4573 19015 4607
rect 21373 4573 21407 4607
rect 21557 4573 21591 4607
rect 1593 4505 1627 4539
rect 5457 4505 5491 4539
rect 12909 4505 12943 4539
rect 22845 4641 22879 4675
rect 22937 4641 22971 4675
rect 24501 4641 24535 4675
rect 23029 4573 23063 4607
rect 25421 4573 25455 4607
rect 25789 4573 25823 4607
rect 2329 4437 2363 4471
rect 3801 4437 3835 4471
rect 6101 4437 6135 4471
rect 7941 4437 7975 4471
rect 8953 4437 8987 4471
rect 9321 4437 9355 4471
rect 11253 4437 11287 4471
rect 11713 4437 11747 4471
rect 13645 4437 13679 4471
rect 15301 4437 15335 4471
rect 16313 4437 16347 4471
rect 20913 4437 20947 4471
rect 21833 4437 21867 4471
rect 22477 4437 22511 4471
rect 24685 4437 24719 4471
rect 25053 4437 25087 4471
rect 26249 4437 26283 4471
rect 3341 4233 3375 4267
rect 4353 4233 4387 4267
rect 10701 4233 10735 4267
rect 11253 4233 11287 4267
rect 19073 4233 19107 4267
rect 24685 4233 24719 4267
rect 4629 4165 4663 4199
rect 4905 4165 4939 4199
rect 14197 4165 14231 4199
rect 15853 4165 15887 4199
rect 2421 4097 2455 4131
rect 3893 4097 3927 4131
rect 2237 4029 2271 4063
rect 3249 4029 3283 4063
rect 3801 4029 3835 4063
rect 5457 4097 5491 4131
rect 9781 4097 9815 4131
rect 9873 4097 9907 4131
rect 12265 4097 12299 4131
rect 13369 4097 13403 4131
rect 14749 4097 14783 4131
rect 14933 4097 14967 4131
rect 16589 4097 16623 4131
rect 17877 4097 17911 4131
rect 18613 4097 18647 4131
rect 20085 4097 20119 4131
rect 20269 4097 20303 4131
rect 21741 4097 21775 4131
rect 22201 4097 22235 4131
rect 24225 4097 24259 4131
rect 5273 4029 5307 4063
rect 6837 4029 6871 4063
rect 9229 4029 9263 4063
rect 9689 4029 9723 4063
rect 11345 4029 11379 4063
rect 13093 4029 13127 4063
rect 14657 4029 14691 4063
rect 15485 4029 15519 4063
rect 16313 4029 16347 4063
rect 18429 4029 18463 4063
rect 19441 4029 19475 4063
rect 21649 4029 21683 4063
rect 22937 4029 22971 4063
rect 24133 4029 24167 4063
rect 25237 4029 25271 4063
rect 25789 4029 25823 4063
rect 1685 3961 1719 3995
rect 2145 3961 2179 3995
rect 4629 3961 4663 3995
rect 4813 3961 4847 3995
rect 5365 3961 5399 3995
rect 7104 3961 7138 3995
rect 19993 3961 20027 3995
rect 21557 3961 21591 3995
rect 26249 3961 26283 3995
rect 1777 3893 1811 3927
rect 2789 3893 2823 3927
rect 3709 3893 3743 3927
rect 6193 3893 6227 3927
rect 6561 3893 6595 3927
rect 8217 3893 8251 3927
rect 8861 3893 8895 3927
rect 9321 3893 9355 3927
rect 10333 3893 10367 3927
rect 11897 3893 11931 3927
rect 12725 3893 12759 3927
rect 13185 3893 13219 3927
rect 13829 3893 13863 3927
rect 14289 3893 14323 3927
rect 15945 3893 15979 3927
rect 16405 3893 16439 3927
rect 16957 3893 16991 3927
rect 17325 3893 17359 3927
rect 18061 3893 18095 3927
rect 18521 3893 18555 3927
rect 19625 3893 19659 3927
rect 20729 3893 20763 3927
rect 21005 3893 21039 3927
rect 21189 3893 21223 3927
rect 22661 3893 22695 3927
rect 23489 3893 23523 3927
rect 23673 3893 23707 3927
rect 24041 3893 24075 3927
rect 25053 3893 25087 3927
rect 25421 3893 25455 3927
rect 1593 3689 1627 3723
rect 1961 3689 1995 3723
rect 2329 3689 2363 3723
rect 2421 3689 2455 3723
rect 2881 3689 2915 3723
rect 4077 3689 4111 3723
rect 5089 3689 5123 3723
rect 7205 3689 7239 3723
rect 9689 3689 9723 3723
rect 10057 3689 10091 3723
rect 10793 3689 10827 3723
rect 12265 3689 12299 3723
rect 12817 3689 12851 3723
rect 13553 3689 13587 3723
rect 14013 3689 14047 3723
rect 16037 3689 16071 3723
rect 16129 3689 16163 3723
rect 16957 3689 16991 3723
rect 17601 3689 17635 3723
rect 18797 3689 18831 3723
rect 20913 3689 20947 3723
rect 22293 3689 22327 3723
rect 22477 3689 22511 3723
rect 24501 3689 24535 3723
rect 2789 3621 2823 3655
rect 4445 3621 4479 3655
rect 5733 3621 5767 3655
rect 11621 3621 11655 3655
rect 14105 3621 14139 3655
rect 18521 3621 18555 3655
rect 19257 3621 19291 3655
rect 19809 3621 19843 3655
rect 20637 3621 20671 3655
rect 25421 3621 25455 3655
rect 26249 3621 26283 3655
rect 1409 3553 1443 3587
rect 4537 3553 4571 3587
rect 5825 3553 5859 3587
rect 6092 3553 6126 3587
rect 9505 3553 9539 3587
rect 11161 3553 11195 3587
rect 14749 3553 14783 3587
rect 19165 3553 19199 3587
rect 21281 3553 21315 3587
rect 22845 3553 22879 3587
rect 22937 3553 22971 3587
rect 24409 3553 24443 3587
rect 3065 3485 3099 3519
rect 3525 3485 3559 3519
rect 3893 3485 3927 3519
rect 4721 3485 4755 3519
rect 8585 3485 8619 3519
rect 10149 3485 10183 3519
rect 10333 3485 10367 3519
rect 11713 3485 11747 3519
rect 11805 3485 11839 3519
rect 14289 3485 14323 3519
rect 15117 3485 15151 3519
rect 15577 3485 15611 3519
rect 16313 3485 16347 3519
rect 17693 3485 17727 3519
rect 17785 3485 17819 3519
rect 19349 3485 19383 3519
rect 21373 3485 21407 3519
rect 21465 3485 21499 3519
rect 21925 3485 21959 3519
rect 23029 3485 23063 3519
rect 23857 3485 23891 3519
rect 24593 3485 24627 3519
rect 7849 3417 7883 3451
rect 9045 3417 9079 3451
rect 13185 3417 13219 3451
rect 15669 3417 15703 3451
rect 25789 3417 25823 3451
rect 8493 3349 8527 3383
rect 11253 3349 11287 3383
rect 13645 3349 13679 3383
rect 17233 3349 17267 3383
rect 20177 3349 20211 3383
rect 23489 3349 23523 3383
rect 24041 3349 24075 3383
rect 25053 3349 25087 3383
rect 1869 3145 1903 3179
rect 3525 3145 3559 3179
rect 6837 3145 6871 3179
rect 9781 3145 9815 3179
rect 10701 3145 10735 3179
rect 13829 3145 13863 3179
rect 16497 3145 16531 3179
rect 17509 3145 17543 3179
rect 18061 3145 18095 3179
rect 19073 3145 19107 3179
rect 19625 3145 19659 3179
rect 22201 3145 22235 3179
rect 23489 3145 23523 3179
rect 25053 3145 25087 3179
rect 4537 3077 4571 3111
rect 4997 3077 5031 3111
rect 5089 3077 5123 3111
rect 6561 3077 6595 3111
rect 10333 3077 10367 3111
rect 11437 3077 11471 3111
rect 17049 3077 17083 3111
rect 19533 3077 19567 3111
rect 20729 3077 20763 3111
rect 21189 3077 21223 3111
rect 22937 3077 22971 3111
rect 24777 3077 24811 3111
rect 2513 3009 2547 3043
rect 3065 3009 3099 3043
rect 4077 3009 4111 3043
rect 5641 3009 5675 3043
rect 7389 3009 7423 3043
rect 14841 3009 14875 3043
rect 17877 3009 17911 3043
rect 18613 3009 18647 3043
rect 20269 3009 20303 3043
rect 21741 3009 21775 3043
rect 24133 3009 24167 3043
rect 24225 3009 24259 3043
rect 2421 2941 2455 2975
rect 5457 2941 5491 2975
rect 5549 2941 5583 2975
rect 7205 2941 7239 2975
rect 7849 2941 7883 2975
rect 8401 2941 8435 2975
rect 8668 2941 8702 2975
rect 11253 2941 11287 2975
rect 12449 2941 12483 2975
rect 2329 2873 2363 2907
rect 3433 2873 3467 2907
rect 7297 2873 7331 2907
rect 11897 2873 11931 2907
rect 12716 2873 12750 2907
rect 15117 2941 15151 2975
rect 15384 2941 15418 2975
rect 18429 2941 18463 2975
rect 18521 2941 18555 2975
rect 19993 2941 20027 2975
rect 20085 2941 20119 2975
rect 25237 2941 25271 2975
rect 25789 2941 25823 2975
rect 22569 2873 22603 2907
rect 24041 2873 24075 2907
rect 1961 2805 1995 2839
rect 3893 2805 3927 2839
rect 3985 2805 4019 2839
rect 6101 2805 6135 2839
rect 8217 2805 8251 2839
rect 11161 2805 11195 2839
rect 12173 2805 12207 2839
rect 14657 2805 14691 2839
rect 14841 2805 14875 2839
rect 15025 2805 15059 2839
rect 21097 2805 21131 2839
rect 21557 2805 21591 2839
rect 21649 2805 21683 2839
rect 23673 2805 23707 2839
rect 25421 2805 25455 2839
rect 26249 2805 26283 2839
rect 2421 2601 2455 2635
rect 2789 2601 2823 2635
rect 5733 2601 5767 2635
rect 6653 2601 6687 2635
rect 8309 2601 8343 2635
rect 12449 2601 12483 2635
rect 14289 2601 14323 2635
rect 16865 2601 16899 2635
rect 18061 2601 18095 2635
rect 18797 2601 18831 2635
rect 21189 2601 21223 2635
rect 23305 2601 23339 2635
rect 23673 2601 23707 2635
rect 24041 2601 24075 2635
rect 25421 2601 25455 2635
rect 25789 2601 25823 2635
rect 2881 2533 2915 2567
rect 3617 2533 3651 2567
rect 7196 2533 7230 2567
rect 8861 2533 8895 2567
rect 9505 2533 9539 2567
rect 10048 2533 10082 2567
rect 12081 2533 12115 2567
rect 13176 2533 13210 2567
rect 14933 2533 14967 2567
rect 15752 2533 15786 2567
rect 19717 2533 19751 2567
rect 22201 2533 22235 2567
rect 24409 2533 24443 2567
rect 26433 2533 26467 2567
rect 1409 2465 1443 2499
rect 4353 2465 4387 2499
rect 4620 2465 4654 2499
rect 6285 2465 6319 2499
rect 6929 2465 6963 2499
rect 9781 2465 9815 2499
rect 12909 2465 12943 2499
rect 15301 2465 15335 2499
rect 15485 2465 15519 2499
rect 18705 2465 18739 2499
rect 19901 2465 19935 2499
rect 21557 2465 21591 2499
rect 21649 2465 21683 2499
rect 22753 2465 22787 2499
rect 25605 2465 25639 2499
rect 2329 2397 2363 2431
rect 3065 2397 3099 2431
rect 18889 2397 18923 2431
rect 21833 2397 21867 2431
rect 22569 2397 22603 2431
rect 24501 2397 24535 2431
rect 24685 2397 24719 2431
rect 24869 2397 24903 2431
rect 20545 2329 20579 2363
rect 26065 2329 26099 2363
rect 1593 2261 1627 2295
rect 1961 2261 1995 2295
rect 11161 2261 11195 2295
rect 17693 2261 17727 2295
rect 18337 2261 18371 2295
rect 20085 2261 20119 2295
rect 20913 2261 20947 2295
rect 22937 2261 22971 2295
rect 24869 2261 24903 2295
rect 25053 2261 25087 2295
<< metal1 >>
rect 18230 26664 18236 26716
rect 18288 26704 18294 26716
rect 24762 26704 24768 26716
rect 18288 26676 24768 26704
rect 18288 26664 18294 26676
rect 24762 26664 24768 26676
rect 24820 26664 24826 26716
rect 22002 26392 22008 26444
rect 22060 26432 22066 26444
rect 24762 26432 24768 26444
rect 22060 26404 24768 26432
rect 22060 26392 22066 26404
rect 24762 26392 24768 26404
rect 24820 26392 24826 26444
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 16574 26228 16580 26240
rect 10100 26200 16580 26228
rect 10100 26188 10106 26200
rect 16574 26188 16580 26200
rect 16632 26188 16638 26240
rect 6362 26120 6368 26172
rect 6420 26160 6426 26172
rect 17402 26160 17408 26172
rect 6420 26132 17408 26160
rect 6420 26120 6426 26132
rect 17402 26120 17408 26132
rect 17460 26120 17466 26172
rect 9122 26052 9128 26104
rect 9180 26092 9186 26104
rect 23474 26092 23480 26104
rect 9180 26064 23480 26092
rect 9180 26052 9186 26064
rect 23474 26052 23480 26064
rect 23532 26052 23538 26104
rect 11238 25984 11244 26036
rect 11296 26024 11302 26036
rect 20346 26024 20352 26036
rect 11296 25996 20352 26024
rect 11296 25984 11302 25996
rect 20346 25984 20352 25996
rect 20404 25984 20410 26036
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 9490 25956 9496 25968
rect 6972 25928 9496 25956
rect 6972 25916 6978 25928
rect 9490 25916 9496 25928
rect 9548 25916 9554 25968
rect 12158 25916 12164 25968
rect 12216 25956 12222 25968
rect 19426 25956 19432 25968
rect 12216 25928 19432 25956
rect 12216 25916 12222 25928
rect 19426 25916 19432 25928
rect 19484 25916 19490 25968
rect 1762 25848 1768 25900
rect 1820 25888 1826 25900
rect 11974 25888 11980 25900
rect 1820 25860 11980 25888
rect 1820 25848 1826 25860
rect 11974 25848 11980 25860
rect 12032 25848 12038 25900
rect 13446 25848 13452 25900
rect 13504 25888 13510 25900
rect 18966 25888 18972 25900
rect 13504 25860 18972 25888
rect 13504 25848 13510 25860
rect 18966 25848 18972 25860
rect 19024 25848 19030 25900
rect 6086 25780 6092 25832
rect 6144 25820 6150 25832
rect 9490 25820 9496 25832
rect 6144 25792 9496 25820
rect 6144 25780 6150 25792
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 10962 25780 10968 25832
rect 11020 25820 11026 25832
rect 21358 25820 21364 25832
rect 11020 25792 21364 25820
rect 11020 25780 11026 25792
rect 21358 25780 21364 25792
rect 21416 25780 21422 25832
rect 10778 25712 10784 25764
rect 10836 25752 10842 25764
rect 19334 25752 19340 25764
rect 10836 25724 19340 25752
rect 10836 25712 10842 25724
rect 19334 25712 19340 25724
rect 19392 25712 19398 25764
rect 4890 25644 4896 25696
rect 4948 25684 4954 25696
rect 13998 25684 14004 25696
rect 4948 25656 14004 25684
rect 4948 25644 4954 25656
rect 13998 25644 14004 25656
rect 14056 25644 14062 25696
rect 15470 25644 15476 25696
rect 15528 25684 15534 25696
rect 24670 25684 24676 25696
rect 15528 25656 24676 25684
rect 15528 25644 15534 25656
rect 24670 25644 24676 25656
rect 24728 25644 24734 25696
rect 1104 25594 26864 25616
rect 1104 25542 10315 25594
rect 10367 25542 10379 25594
rect 10431 25542 10443 25594
rect 10495 25542 10507 25594
rect 10559 25542 19648 25594
rect 19700 25542 19712 25594
rect 19764 25542 19776 25594
rect 19828 25542 19840 25594
rect 19892 25542 26864 25594
rect 1104 25520 26864 25542
rect 2685 25483 2743 25489
rect 2685 25449 2697 25483
rect 2731 25480 2743 25483
rect 3234 25480 3240 25492
rect 2731 25452 3240 25480
rect 2731 25449 2743 25452
rect 2685 25443 2743 25449
rect 3234 25440 3240 25452
rect 3292 25440 3298 25492
rect 7834 25440 7840 25492
rect 7892 25480 7898 25492
rect 10962 25480 10968 25492
rect 7892 25452 10456 25480
rect 10923 25452 10968 25480
rect 7892 25440 7898 25452
rect 6270 25372 6276 25424
rect 6328 25412 6334 25424
rect 6328 25384 8248 25412
rect 6328 25372 6334 25384
rect 1397 25347 1455 25353
rect 1397 25313 1409 25347
rect 1443 25344 1455 25347
rect 2130 25344 2136 25356
rect 1443 25316 2136 25344
rect 1443 25313 1455 25316
rect 1397 25307 1455 25313
rect 2130 25304 2136 25316
rect 2188 25304 2194 25356
rect 2501 25347 2559 25353
rect 2501 25313 2513 25347
rect 2547 25344 2559 25347
rect 3418 25344 3424 25356
rect 2547 25316 3424 25344
rect 2547 25313 2559 25316
rect 2501 25307 2559 25313
rect 3418 25304 3424 25316
rect 3476 25304 3482 25356
rect 4065 25347 4123 25353
rect 4065 25313 4077 25347
rect 4111 25344 4123 25347
rect 4154 25344 4160 25356
rect 4111 25316 4160 25344
rect 4111 25313 4123 25316
rect 4065 25307 4123 25313
rect 4154 25304 4160 25316
rect 4212 25304 4218 25356
rect 7837 25347 7895 25353
rect 7837 25313 7849 25347
rect 7883 25313 7895 25347
rect 7837 25307 7895 25313
rect 5166 25276 5172 25288
rect 5127 25248 5172 25276
rect 5166 25236 5172 25248
rect 5224 25236 5230 25288
rect 2409 25211 2467 25217
rect 2409 25177 2421 25211
rect 2455 25208 2467 25211
rect 3050 25208 3056 25220
rect 2455 25180 3056 25208
rect 2455 25177 2467 25180
rect 2409 25171 2467 25177
rect 3050 25168 3056 25180
rect 3108 25168 3114 25220
rect 4709 25211 4767 25217
rect 4709 25177 4721 25211
rect 4755 25208 4767 25211
rect 5074 25208 5080 25220
rect 4755 25180 5080 25208
rect 4755 25177 4767 25180
rect 4709 25171 4767 25177
rect 5074 25168 5080 25180
rect 5132 25168 5138 25220
rect 5258 25168 5264 25220
rect 5316 25208 5322 25220
rect 7285 25211 7343 25217
rect 7285 25208 7297 25211
rect 5316 25180 7297 25208
rect 5316 25168 5322 25180
rect 7285 25177 7297 25180
rect 7331 25208 7343 25211
rect 7852 25208 7880 25307
rect 7929 25279 7987 25285
rect 7929 25245 7941 25279
rect 7975 25245 7987 25279
rect 8110 25276 8116 25288
rect 8071 25248 8116 25276
rect 7929 25239 7987 25245
rect 7331 25180 7880 25208
rect 7944 25208 7972 25239
rect 8110 25236 8116 25248
rect 8168 25236 8174 25288
rect 8220 25276 8248 25384
rect 9585 25347 9643 25353
rect 9585 25313 9597 25347
rect 9631 25344 9643 25347
rect 9858 25344 9864 25356
rect 9631 25316 9864 25344
rect 9631 25313 9643 25316
rect 9585 25307 9643 25313
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10428 25344 10456 25452
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 11054 25440 11060 25492
rect 11112 25480 11118 25492
rect 14461 25483 14519 25489
rect 11112 25452 14412 25480
rect 11112 25440 11118 25452
rect 12434 25372 12440 25424
rect 12492 25412 12498 25424
rect 12989 25415 13047 25421
rect 12989 25412 13001 25415
rect 12492 25384 13001 25412
rect 12492 25372 12498 25384
rect 12989 25381 13001 25384
rect 13035 25381 13047 25415
rect 14384 25412 14412 25452
rect 14461 25449 14473 25483
rect 14507 25480 14519 25483
rect 18322 25480 18328 25492
rect 14507 25452 18328 25480
rect 14507 25449 14519 25452
rect 14461 25443 14519 25449
rect 18322 25440 18328 25452
rect 18380 25440 18386 25492
rect 21361 25483 21419 25489
rect 21361 25449 21373 25483
rect 21407 25480 21419 25483
rect 22370 25480 22376 25492
rect 21407 25452 22376 25480
rect 21407 25449 21419 25452
rect 21361 25443 21419 25449
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 14384 25384 16712 25412
rect 12989 25375 13047 25381
rect 10873 25347 10931 25353
rect 10873 25344 10885 25347
rect 10428 25316 10885 25344
rect 10873 25313 10885 25316
rect 10919 25344 10931 25347
rect 11238 25344 11244 25356
rect 10919 25316 11244 25344
rect 10919 25313 10931 25316
rect 10873 25307 10931 25313
rect 11238 25304 11244 25316
rect 11296 25344 11302 25356
rect 11333 25347 11391 25353
rect 11333 25344 11345 25347
rect 11296 25316 11345 25344
rect 11296 25304 11302 25316
rect 11333 25313 11345 25316
rect 11379 25313 11391 25347
rect 11333 25307 11391 25313
rect 12069 25347 12127 25353
rect 12069 25313 12081 25347
rect 12115 25344 12127 25347
rect 14277 25347 14335 25353
rect 12115 25316 13308 25344
rect 12115 25313 12127 25316
rect 12069 25307 12127 25313
rect 10962 25276 10968 25288
rect 8220 25248 10968 25276
rect 10962 25236 10968 25248
rect 11020 25236 11026 25288
rect 11054 25236 11060 25288
rect 11112 25276 11118 25288
rect 11425 25279 11483 25285
rect 11425 25276 11437 25279
rect 11112 25248 11437 25276
rect 11112 25236 11118 25248
rect 11425 25245 11437 25248
rect 11471 25245 11483 25279
rect 11425 25239 11483 25245
rect 11517 25279 11575 25285
rect 11517 25245 11529 25279
rect 11563 25245 11575 25279
rect 13078 25276 13084 25288
rect 13039 25248 13084 25276
rect 11517 25239 11575 25245
rect 8018 25208 8024 25220
rect 7944 25180 8024 25208
rect 7331 25177 7343 25180
rect 7285 25171 7343 25177
rect 8018 25168 8024 25180
rect 8076 25168 8082 25220
rect 8294 25168 8300 25220
rect 8352 25208 8358 25220
rect 8849 25211 8907 25217
rect 8849 25208 8861 25211
rect 8352 25180 8861 25208
rect 8352 25168 8358 25180
rect 8849 25177 8861 25180
rect 8895 25177 8907 25211
rect 10042 25208 10048 25220
rect 10003 25180 10048 25208
rect 8849 25171 8907 25177
rect 10042 25168 10048 25180
rect 10100 25168 10106 25220
rect 10505 25211 10563 25217
rect 10505 25177 10517 25211
rect 10551 25208 10563 25211
rect 11532 25208 11560 25239
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13280 25285 13308 25316
rect 14277 25313 14289 25347
rect 14323 25344 14335 25347
rect 15286 25344 15292 25356
rect 14323 25316 15292 25344
rect 14323 25313 14335 25316
rect 14277 25307 14335 25313
rect 15286 25304 15292 25316
rect 15344 25304 15350 25356
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 14001 25279 14059 25285
rect 14001 25276 14013 25279
rect 13311 25248 14013 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 14001 25245 14013 25248
rect 14047 25245 14059 25279
rect 14001 25239 14059 25245
rect 15378 25236 15384 25288
rect 15436 25276 15442 25288
rect 16117 25279 16175 25285
rect 16117 25276 16129 25279
rect 15436 25248 16129 25276
rect 15436 25236 15442 25248
rect 16117 25245 16129 25248
rect 16163 25245 16175 25279
rect 16117 25239 16175 25245
rect 11790 25208 11796 25220
rect 10551 25180 11796 25208
rect 10551 25177 10563 25180
rect 10505 25171 10563 25177
rect 11790 25168 11796 25180
rect 11848 25168 11854 25220
rect 12621 25211 12679 25217
rect 12621 25177 12633 25211
rect 12667 25208 12679 25211
rect 16684 25208 16712 25384
rect 17862 25372 17868 25424
rect 17920 25412 17926 25424
rect 18969 25415 19027 25421
rect 18969 25412 18981 25415
rect 17920 25384 18981 25412
rect 17920 25372 17926 25384
rect 18969 25381 18981 25384
rect 19015 25412 19027 25415
rect 24854 25412 24860 25424
rect 19015 25384 24860 25412
rect 19015 25381 19027 25384
rect 18969 25375 19027 25381
rect 24854 25372 24860 25384
rect 24912 25372 24918 25424
rect 16853 25347 16911 25353
rect 16853 25313 16865 25347
rect 16899 25344 16911 25347
rect 17126 25344 17132 25356
rect 16899 25316 17132 25344
rect 16899 25313 16911 25316
rect 16853 25307 16911 25313
rect 17126 25304 17132 25316
rect 17184 25304 17190 25356
rect 19981 25347 20039 25353
rect 19981 25344 19993 25347
rect 19168 25316 19993 25344
rect 19168 25288 19196 25316
rect 19981 25313 19993 25316
rect 20027 25313 20039 25347
rect 19981 25307 20039 25313
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 21177 25347 21235 25353
rect 21177 25344 21189 25347
rect 21140 25316 21189 25344
rect 21140 25304 21146 25316
rect 21177 25313 21189 25316
rect 21223 25313 21235 25347
rect 21177 25307 21235 25313
rect 16942 25276 16948 25288
rect 16903 25248 16948 25276
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17037 25279 17095 25285
rect 17037 25245 17049 25279
rect 17083 25276 17095 25279
rect 17218 25276 17224 25288
rect 17083 25248 17224 25276
rect 17083 25245 17095 25248
rect 17037 25239 17095 25245
rect 17218 25236 17224 25248
rect 17276 25276 17282 25288
rect 17681 25279 17739 25285
rect 17681 25276 17693 25279
rect 17276 25248 17693 25276
rect 17276 25236 17282 25248
rect 17681 25245 17693 25248
rect 17727 25245 17739 25279
rect 19058 25276 19064 25288
rect 19019 25248 19064 25276
rect 17681 25239 17739 25245
rect 19058 25236 19064 25248
rect 19116 25236 19122 25288
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19208 25248 19253 25276
rect 19208 25236 19214 25248
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 22830 25276 22836 25288
rect 19392 25248 22836 25276
rect 19392 25236 19398 25248
rect 22830 25236 22836 25248
rect 22888 25236 22894 25288
rect 25774 25208 25780 25220
rect 12667 25180 16160 25208
rect 16684 25180 25780 25208
rect 12667 25177 12679 25180
rect 12621 25171 12679 25177
rect 16132 25152 16160 25180
rect 25774 25168 25780 25180
rect 25832 25168 25838 25220
rect 1394 25100 1400 25152
rect 1452 25140 1458 25152
rect 1581 25143 1639 25149
rect 1581 25140 1593 25143
rect 1452 25112 1593 25140
rect 1452 25100 1458 25112
rect 1581 25109 1593 25112
rect 1627 25109 1639 25143
rect 2038 25140 2044 25152
rect 1999 25112 2044 25140
rect 1581 25103 1639 25109
rect 2038 25100 2044 25112
rect 2096 25100 2102 25152
rect 3145 25143 3203 25149
rect 3145 25109 3157 25143
rect 3191 25140 3203 25143
rect 3510 25140 3516 25152
rect 3191 25112 3516 25140
rect 3191 25109 3203 25112
rect 3145 25103 3203 25109
rect 3510 25100 3516 25112
rect 3568 25100 3574 25152
rect 3694 25140 3700 25152
rect 3655 25112 3700 25140
rect 3694 25100 3700 25112
rect 3752 25100 3758 25152
rect 3970 25100 3976 25152
rect 4028 25140 4034 25152
rect 4249 25143 4307 25149
rect 4249 25140 4261 25143
rect 4028 25112 4261 25140
rect 4028 25100 4034 25112
rect 4249 25109 4261 25112
rect 4295 25109 4307 25143
rect 4982 25140 4988 25152
rect 4943 25112 4988 25140
rect 4249 25103 4307 25109
rect 4982 25100 4988 25112
rect 5040 25100 5046 25152
rect 5350 25100 5356 25152
rect 5408 25140 5414 25152
rect 5629 25143 5687 25149
rect 5629 25140 5641 25143
rect 5408 25112 5641 25140
rect 5408 25100 5414 25112
rect 5629 25109 5641 25112
rect 5675 25109 5687 25143
rect 5629 25103 5687 25109
rect 6733 25143 6791 25149
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 7098 25140 7104 25152
rect 6779 25112 7104 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 7098 25100 7104 25112
rect 7156 25100 7162 25152
rect 7469 25143 7527 25149
rect 7469 25109 7481 25143
rect 7515 25140 7527 25143
rect 7926 25140 7932 25152
rect 7515 25112 7932 25140
rect 7515 25109 7527 25112
rect 7469 25103 7527 25109
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 8573 25143 8631 25149
rect 8573 25109 8585 25143
rect 8619 25140 8631 25143
rect 8938 25140 8944 25152
rect 8619 25112 8944 25140
rect 8619 25109 8631 25112
rect 8573 25103 8631 25109
rect 8938 25100 8944 25112
rect 8996 25100 9002 25152
rect 12250 25100 12256 25152
rect 12308 25140 12314 25152
rect 12345 25143 12403 25149
rect 12345 25140 12357 25143
rect 12308 25112 12357 25140
rect 12308 25100 12314 25112
rect 12345 25109 12357 25112
rect 12391 25109 12403 25143
rect 12345 25103 12403 25109
rect 14001 25143 14059 25149
rect 14001 25109 14013 25143
rect 14047 25140 14059 25143
rect 14185 25143 14243 25149
rect 14185 25140 14197 25143
rect 14047 25112 14197 25140
rect 14047 25109 14059 25112
rect 14001 25103 14059 25109
rect 14185 25109 14197 25112
rect 14231 25140 14243 25143
rect 14366 25140 14372 25152
rect 14231 25112 14372 25140
rect 14231 25109 14243 25112
rect 14185 25103 14243 25109
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 14734 25100 14740 25152
rect 14792 25140 14798 25152
rect 14829 25143 14887 25149
rect 14829 25140 14841 25143
rect 14792 25112 14841 25140
rect 14792 25100 14798 25112
rect 14829 25109 14841 25112
rect 14875 25109 14887 25143
rect 15838 25140 15844 25152
rect 15799 25112 15844 25140
rect 14829 25103 14887 25109
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 16114 25100 16120 25152
rect 16172 25100 16178 25152
rect 16485 25143 16543 25149
rect 16485 25109 16497 25143
rect 16531 25140 16543 25143
rect 16758 25140 16764 25152
rect 16531 25112 16764 25140
rect 16531 25109 16543 25112
rect 16485 25103 16543 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 18141 25143 18199 25149
rect 18141 25109 18153 25143
rect 18187 25140 18199 25143
rect 18230 25140 18236 25152
rect 18187 25112 18236 25140
rect 18187 25109 18199 25112
rect 18141 25103 18199 25109
rect 18230 25100 18236 25112
rect 18288 25100 18294 25152
rect 18598 25140 18604 25152
rect 18559 25112 18604 25140
rect 18598 25100 18604 25112
rect 18656 25100 18662 25152
rect 19702 25140 19708 25152
rect 19663 25112 19708 25140
rect 19702 25100 19708 25112
rect 19760 25100 19766 25152
rect 1104 25050 26864 25072
rect 1104 24998 5648 25050
rect 5700 24998 5712 25050
rect 5764 24998 5776 25050
rect 5828 24998 5840 25050
rect 5892 24998 14982 25050
rect 15034 24998 15046 25050
rect 15098 24998 15110 25050
rect 15162 24998 15174 25050
rect 15226 24998 24315 25050
rect 24367 24998 24379 25050
rect 24431 24998 24443 25050
rect 24495 24998 24507 25050
rect 24559 24998 26864 25050
rect 1104 24976 26864 24998
rect 3050 24896 3056 24948
rect 3108 24936 3114 24948
rect 4617 24939 4675 24945
rect 4617 24936 4629 24939
rect 3108 24908 4629 24936
rect 3108 24896 3114 24908
rect 4617 24905 4629 24908
rect 4663 24905 4675 24939
rect 6638 24936 6644 24948
rect 6551 24908 6644 24936
rect 4617 24899 4675 24905
rect 6638 24896 6644 24908
rect 6696 24936 6702 24948
rect 8018 24936 8024 24948
rect 6696 24908 8024 24936
rect 6696 24896 6702 24908
rect 8018 24896 8024 24908
rect 8076 24896 8082 24948
rect 12066 24936 12072 24948
rect 9600 24908 12072 24936
rect 937 24871 995 24877
rect 937 24837 949 24871
rect 983 24868 995 24871
rect 1762 24868 1768 24880
rect 983 24840 1768 24868
rect 983 24837 995 24840
rect 937 24831 995 24837
rect 1762 24828 1768 24840
rect 1820 24828 1826 24880
rect 3789 24871 3847 24877
rect 3789 24868 3801 24871
rect 3436 24840 3801 24868
rect 3436 24812 3464 24840
rect 3789 24837 3801 24840
rect 3835 24837 3847 24871
rect 3789 24831 3847 24837
rect 4430 24828 4436 24880
rect 4488 24868 4494 24880
rect 4488 24840 5212 24868
rect 4488 24828 4494 24840
rect 3053 24803 3111 24809
rect 3053 24800 3065 24803
rect 2608 24772 3065 24800
rect 1397 24735 1455 24741
rect 1397 24701 1409 24735
rect 1443 24732 1455 24735
rect 1578 24732 1584 24744
rect 1443 24704 1584 24732
rect 1443 24701 1455 24704
rect 1397 24695 1455 24701
rect 1578 24692 1584 24704
rect 1636 24732 1642 24744
rect 2317 24735 2375 24741
rect 2317 24732 2329 24735
rect 1636 24704 2329 24732
rect 1636 24692 1642 24704
rect 2317 24701 2329 24704
rect 2363 24701 2375 24735
rect 2498 24732 2504 24744
rect 2411 24704 2504 24732
rect 2317 24695 2375 24701
rect 2498 24692 2504 24704
rect 2556 24732 2562 24744
rect 2608 24732 2636 24772
rect 3053 24769 3065 24772
rect 3099 24769 3111 24803
rect 3418 24800 3424 24812
rect 3379 24772 3424 24800
rect 3053 24763 3111 24769
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 4154 24800 4160 24812
rect 4067 24772 4160 24800
rect 4154 24760 4160 24772
rect 4212 24800 4218 24812
rect 4890 24800 4896 24812
rect 4212 24772 4896 24800
rect 4212 24760 4218 24772
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 5184 24809 5212 24840
rect 8110 24828 8116 24880
rect 8168 24868 8174 24880
rect 8168 24840 8800 24868
rect 8168 24828 8174 24840
rect 8772 24809 8800 24840
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24769 5227 24803
rect 5169 24763 5227 24769
rect 8757 24803 8815 24809
rect 8757 24769 8769 24803
rect 8803 24769 8815 24803
rect 8757 24763 8815 24769
rect 2556 24704 2636 24732
rect 2556 24692 2562 24704
rect 2774 24692 2780 24744
rect 2832 24732 2838 24744
rect 3605 24735 3663 24741
rect 3605 24732 3617 24735
rect 2832 24704 3617 24732
rect 2832 24692 2838 24704
rect 3605 24701 3617 24704
rect 3651 24701 3663 24735
rect 4982 24732 4988 24744
rect 4943 24704 4988 24732
rect 3605 24695 3663 24701
rect 2958 24664 2964 24676
rect 1596 24636 2964 24664
rect 1596 24605 1624 24636
rect 2958 24624 2964 24636
rect 3016 24624 3022 24676
rect 3620 24664 3648 24695
rect 4982 24692 4988 24704
rect 5040 24692 5046 24744
rect 7098 24732 7104 24744
rect 7011 24704 7104 24732
rect 7098 24692 7104 24704
rect 7156 24732 7162 24744
rect 8386 24732 8392 24744
rect 7156 24704 8392 24732
rect 7156 24692 7162 24704
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 8665 24735 8723 24741
rect 8665 24701 8677 24735
rect 8711 24732 8723 24735
rect 8938 24732 8944 24744
rect 8711 24704 8944 24732
rect 8711 24701 8723 24704
rect 8665 24695 8723 24701
rect 8938 24692 8944 24704
rect 8996 24732 9002 24744
rect 9600 24732 9628 24908
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 19058 24896 19064 24948
rect 19116 24936 19122 24948
rect 19245 24939 19303 24945
rect 19245 24936 19257 24939
rect 19116 24908 19257 24936
rect 19116 24896 19122 24908
rect 19245 24905 19257 24908
rect 19291 24936 19303 24939
rect 24762 24936 24768 24948
rect 19291 24908 24768 24936
rect 19291 24905 19303 24908
rect 19245 24899 19303 24905
rect 24762 24896 24768 24908
rect 24820 24896 24826 24948
rect 9858 24828 9864 24880
rect 9916 24868 9922 24880
rect 15010 24868 15016 24880
rect 9916 24840 15016 24868
rect 9916 24828 9922 24840
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 15105 24871 15163 24877
rect 15105 24837 15117 24871
rect 15151 24868 15163 24871
rect 15286 24868 15292 24880
rect 15151 24840 15292 24868
rect 15151 24837 15163 24840
rect 15105 24831 15163 24837
rect 15286 24828 15292 24840
rect 15344 24868 15350 24880
rect 16390 24868 16396 24880
rect 15344 24840 16396 24868
rect 15344 24828 15350 24840
rect 16390 24828 16396 24840
rect 16448 24828 16454 24880
rect 19702 24868 19708 24880
rect 16868 24840 19708 24868
rect 9950 24760 9956 24812
rect 10008 24800 10014 24812
rect 10321 24803 10379 24809
rect 10321 24800 10333 24803
rect 10008 24772 10333 24800
rect 10008 24760 10014 24772
rect 10321 24769 10333 24772
rect 10367 24769 10379 24803
rect 10321 24763 10379 24769
rect 11974 24760 11980 24812
rect 12032 24800 12038 24812
rect 12161 24803 12219 24809
rect 12161 24800 12173 24803
rect 12032 24772 12173 24800
rect 12032 24760 12038 24772
rect 12161 24769 12173 24772
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12250 24760 12256 24812
rect 12308 24800 12314 24812
rect 12618 24800 12624 24812
rect 12308 24772 12624 24800
rect 12308 24760 12314 24772
rect 12618 24760 12624 24772
rect 12676 24800 12682 24812
rect 13081 24803 13139 24809
rect 13081 24800 13093 24803
rect 12676 24772 13093 24800
rect 12676 24760 12682 24772
rect 13081 24769 13093 24772
rect 13127 24800 13139 24803
rect 13630 24800 13636 24812
rect 13127 24772 13636 24800
rect 13127 24769 13139 24772
rect 13081 24763 13139 24769
rect 13630 24760 13636 24772
rect 13688 24760 13694 24812
rect 14366 24760 14372 24812
rect 14424 24800 14430 24812
rect 14737 24803 14795 24809
rect 14737 24800 14749 24803
rect 14424 24772 14749 24800
rect 14424 24760 14430 24772
rect 14737 24769 14749 24772
rect 14783 24800 14795 24803
rect 15746 24800 15752 24812
rect 14783 24772 15752 24800
rect 14783 24769 14795 24772
rect 14737 24763 14795 24769
rect 15746 24760 15752 24772
rect 15804 24800 15810 24812
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 15804 24772 16313 24800
rect 15804 24760 15810 24772
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 8996 24704 9628 24732
rect 9677 24735 9735 24741
rect 8996 24692 9002 24704
rect 9677 24701 9689 24735
rect 9723 24732 9735 24735
rect 9858 24732 9864 24744
rect 9723 24704 9864 24732
rect 9723 24701 9735 24704
rect 9677 24695 9735 24701
rect 9858 24692 9864 24704
rect 9916 24732 9922 24744
rect 10229 24735 10287 24741
rect 10229 24732 10241 24735
rect 9916 24704 10241 24732
rect 9916 24692 9922 24704
rect 10229 24701 10241 24704
rect 10275 24701 10287 24735
rect 10229 24695 10287 24701
rect 11885 24735 11943 24741
rect 11885 24701 11897 24735
rect 11931 24732 11943 24735
rect 12342 24732 12348 24744
rect 11931 24704 12348 24732
rect 11931 24701 11943 24704
rect 11885 24695 11943 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12526 24692 12532 24744
rect 12584 24732 12590 24744
rect 12584 24704 15608 24732
rect 12584 24692 12590 24704
rect 5629 24667 5687 24673
rect 5629 24664 5641 24667
rect 3620 24636 5641 24664
rect 5629 24633 5641 24636
rect 5675 24633 5687 24667
rect 5629 24627 5687 24633
rect 7834 24624 7840 24676
rect 7892 24664 7898 24676
rect 9309 24667 9367 24673
rect 7892 24636 8248 24664
rect 7892 24624 7898 24636
rect 1581 24599 1639 24605
rect 1581 24565 1593 24599
rect 1627 24565 1639 24599
rect 1581 24559 1639 24565
rect 2041 24599 2099 24605
rect 2041 24565 2053 24599
rect 2087 24596 2099 24599
rect 2130 24596 2136 24608
rect 2087 24568 2136 24596
rect 2087 24565 2099 24568
rect 2041 24559 2099 24565
rect 2130 24556 2136 24568
rect 2188 24556 2194 24608
rect 2682 24596 2688 24608
rect 2643 24568 2688 24596
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 4430 24596 4436 24608
rect 4391 24568 4436 24596
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 5074 24596 5080 24608
rect 5035 24568 5080 24596
rect 5074 24556 5080 24568
rect 5132 24556 5138 24608
rect 5994 24596 6000 24608
rect 5955 24568 6000 24596
rect 5994 24556 6000 24568
rect 6052 24556 6058 24608
rect 7282 24596 7288 24608
rect 7243 24568 7288 24596
rect 7282 24556 7288 24568
rect 7340 24556 7346 24608
rect 7745 24599 7803 24605
rect 7745 24565 7757 24599
rect 7791 24596 7803 24599
rect 8110 24596 8116 24608
rect 7791 24568 8116 24596
rect 7791 24565 7803 24568
rect 7745 24559 7803 24565
rect 8110 24556 8116 24568
rect 8168 24556 8174 24608
rect 8220 24605 8248 24636
rect 9309 24633 9321 24667
rect 9355 24664 9367 24667
rect 10137 24667 10195 24673
rect 10137 24664 10149 24667
rect 9355 24636 10149 24664
rect 9355 24633 9367 24636
rect 9309 24627 9367 24633
rect 10137 24633 10149 24636
rect 10183 24664 10195 24667
rect 11333 24667 11391 24673
rect 11333 24664 11345 24667
rect 10183 24636 11345 24664
rect 10183 24633 10195 24636
rect 10137 24627 10195 24633
rect 11333 24633 11345 24636
rect 11379 24633 11391 24667
rect 11333 24627 11391 24633
rect 11974 24624 11980 24676
rect 12032 24664 12038 24676
rect 12897 24667 12955 24673
rect 12897 24664 12909 24667
rect 12032 24636 12909 24664
rect 12032 24624 12038 24636
rect 12897 24633 12909 24636
rect 12943 24664 12955 24667
rect 13170 24664 13176 24676
rect 12943 24636 13176 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 13170 24624 13176 24636
rect 13228 24624 13234 24676
rect 13998 24664 14004 24676
rect 13911 24636 14004 24664
rect 13998 24624 14004 24636
rect 14056 24664 14062 24676
rect 15580 24673 15608 24704
rect 15838 24692 15844 24744
rect 15896 24732 15902 24744
rect 16117 24735 16175 24741
rect 16117 24732 16129 24735
rect 15896 24704 16129 24732
rect 15896 24692 15902 24704
rect 16117 24701 16129 24704
rect 16163 24732 16175 24735
rect 16868 24732 16896 24840
rect 19702 24828 19708 24840
rect 19760 24828 19766 24880
rect 20990 24828 20996 24880
rect 21048 24868 21054 24880
rect 24210 24868 24216 24880
rect 21048 24840 24216 24868
rect 21048 24828 21054 24840
rect 24210 24828 24216 24840
rect 24268 24828 24274 24880
rect 17862 24800 17868 24812
rect 17823 24772 17868 24800
rect 17862 24760 17868 24772
rect 17920 24760 17926 24812
rect 18601 24803 18659 24809
rect 18601 24800 18613 24803
rect 17972 24772 18613 24800
rect 17126 24732 17132 24744
rect 16163 24704 16896 24732
rect 17087 24704 17132 24732
rect 16163 24701 16175 24704
rect 16117 24695 16175 24701
rect 17126 24692 17132 24704
rect 17184 24692 17190 24744
rect 17218 24692 17224 24744
rect 17276 24732 17282 24744
rect 17972 24732 18000 24772
rect 18601 24769 18613 24772
rect 18647 24800 18659 24803
rect 19150 24800 19156 24812
rect 18647 24772 19156 24800
rect 18647 24769 18659 24772
rect 18601 24763 18659 24769
rect 19150 24760 19156 24772
rect 19208 24800 19214 24812
rect 20165 24803 20223 24809
rect 20165 24800 20177 24803
rect 19208 24772 20177 24800
rect 19208 24760 19214 24772
rect 20165 24769 20177 24772
rect 20211 24800 20223 24803
rect 20438 24800 20444 24812
rect 20211 24772 20444 24800
rect 20211 24769 20223 24772
rect 20165 24763 20223 24769
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 17276 24704 18000 24732
rect 17276 24692 17282 24704
rect 18046 24692 18052 24744
rect 18104 24732 18110 24744
rect 18417 24735 18475 24741
rect 18417 24732 18429 24735
rect 18104 24704 18429 24732
rect 18104 24692 18110 24704
rect 18417 24701 18429 24704
rect 18463 24701 18475 24735
rect 18417 24695 18475 24701
rect 18506 24692 18512 24744
rect 18564 24732 18570 24744
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18564 24704 19073 24732
rect 18564 24692 18570 24704
rect 19061 24701 19073 24704
rect 19107 24732 19119 24735
rect 19245 24735 19303 24741
rect 19245 24732 19257 24735
rect 19107 24704 19257 24732
rect 19107 24701 19119 24704
rect 19061 24695 19119 24701
rect 19245 24701 19257 24704
rect 19291 24701 19303 24735
rect 19245 24695 19303 24701
rect 19521 24735 19579 24741
rect 19521 24701 19533 24735
rect 19567 24732 19579 24735
rect 19567 24704 20484 24732
rect 19567 24701 19579 24704
rect 19521 24695 19579 24701
rect 15565 24667 15623 24673
rect 14056 24636 14596 24664
rect 14056 24624 14062 24636
rect 8205 24599 8263 24605
rect 8205 24565 8217 24599
rect 8251 24565 8263 24599
rect 8205 24559 8263 24565
rect 8294 24556 8300 24608
rect 8352 24596 8358 24608
rect 8573 24599 8631 24605
rect 8573 24596 8585 24599
rect 8352 24568 8585 24596
rect 8352 24556 8358 24568
rect 8573 24565 8585 24568
rect 8619 24565 8631 24599
rect 9766 24596 9772 24608
rect 9727 24568 9772 24596
rect 8573 24559 8631 24565
rect 9766 24556 9772 24568
rect 9824 24556 9830 24608
rect 11054 24596 11060 24608
rect 11015 24568 11060 24596
rect 11054 24556 11060 24568
rect 11112 24556 11118 24608
rect 12529 24599 12587 24605
rect 12529 24565 12541 24599
rect 12575 24596 12587 24599
rect 12710 24596 12716 24608
rect 12575 24568 12716 24596
rect 12575 24565 12587 24568
rect 12529 24559 12587 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 12989 24599 13047 24605
rect 12989 24565 13001 24599
rect 13035 24596 13047 24599
rect 13633 24599 13691 24605
rect 13633 24596 13645 24599
rect 13035 24568 13645 24596
rect 13035 24565 13047 24568
rect 12989 24559 13047 24565
rect 13633 24565 13645 24568
rect 13679 24596 13691 24599
rect 13722 24596 13728 24608
rect 13679 24568 13728 24596
rect 13679 24565 13691 24568
rect 13633 24559 13691 24565
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14458 24596 14464 24608
rect 14419 24568 14464 24596
rect 14458 24556 14464 24568
rect 14516 24556 14522 24608
rect 14568 24605 14596 24636
rect 15565 24633 15577 24667
rect 15611 24664 15623 24667
rect 17310 24664 17316 24676
rect 15611 24636 15884 24664
rect 15611 24633 15623 24636
rect 15565 24627 15623 24633
rect 14553 24599 14611 24605
rect 14553 24565 14565 24599
rect 14599 24596 14611 24599
rect 14642 24596 14648 24608
rect 14599 24568 14648 24596
rect 14599 24565 14611 24568
rect 14553 24559 14611 24565
rect 14642 24556 14648 24568
rect 14700 24556 14706 24608
rect 15654 24556 15660 24608
rect 15712 24596 15718 24608
rect 15749 24599 15807 24605
rect 15749 24596 15761 24599
rect 15712 24568 15761 24596
rect 15712 24556 15718 24568
rect 15749 24565 15761 24568
rect 15795 24565 15807 24599
rect 15856 24596 15884 24636
rect 16592 24636 17316 24664
rect 16209 24599 16267 24605
rect 16209 24596 16221 24599
rect 15856 24568 16221 24596
rect 15749 24559 15807 24565
rect 16209 24565 16221 24568
rect 16255 24596 16267 24599
rect 16592 24596 16620 24636
rect 17310 24624 17316 24636
rect 17368 24624 17374 24676
rect 19702 24624 19708 24676
rect 19760 24664 19766 24676
rect 19981 24667 20039 24673
rect 19981 24664 19993 24667
rect 19760 24636 19993 24664
rect 19760 24624 19766 24636
rect 19981 24633 19993 24636
rect 20027 24664 20039 24667
rect 20162 24664 20168 24676
rect 20027 24636 20168 24664
rect 20027 24633 20039 24636
rect 19981 24627 20039 24633
rect 20162 24624 20168 24636
rect 20220 24624 20226 24676
rect 20456 24664 20484 24704
rect 21174 24692 21180 24744
rect 21232 24732 21238 24744
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21232 24704 21649 24732
rect 21232 24692 21238 24704
rect 21637 24701 21649 24704
rect 21683 24732 21695 24735
rect 22189 24735 22247 24741
rect 22189 24732 22201 24735
rect 21683 24704 22201 24732
rect 21683 24701 21695 24704
rect 21637 24695 21695 24701
rect 22189 24701 22201 24704
rect 22235 24701 22247 24735
rect 23934 24732 23940 24744
rect 23895 24704 23940 24732
rect 22189 24695 22247 24701
rect 23934 24692 23940 24704
rect 23992 24732 23998 24744
rect 24489 24735 24547 24741
rect 24489 24732 24501 24735
rect 23992 24704 24501 24732
rect 23992 24692 23998 24704
rect 24489 24701 24501 24704
rect 24535 24701 24547 24735
rect 24489 24695 24547 24701
rect 27246 24664 27252 24676
rect 20456 24636 27252 24664
rect 16850 24596 16856 24608
rect 16255 24568 16620 24596
rect 16811 24568 16856 24596
rect 16255 24565 16267 24568
rect 16209 24559 16267 24565
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 17862 24556 17868 24608
rect 17920 24596 17926 24608
rect 18049 24599 18107 24605
rect 18049 24596 18061 24599
rect 17920 24568 18061 24596
rect 17920 24556 17926 24568
rect 18049 24565 18061 24568
rect 18095 24565 18107 24599
rect 18049 24559 18107 24565
rect 18230 24556 18236 24608
rect 18288 24596 18294 24608
rect 18509 24599 18567 24605
rect 18509 24596 18521 24599
rect 18288 24568 18521 24596
rect 18288 24556 18294 24568
rect 18509 24565 18521 24568
rect 18555 24565 18567 24599
rect 18509 24559 18567 24565
rect 19518 24556 19524 24608
rect 19576 24596 19582 24608
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19576 24568 19625 24596
rect 19576 24556 19582 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 19613 24559 19671 24565
rect 20073 24599 20131 24605
rect 20073 24565 20085 24599
rect 20119 24596 20131 24599
rect 20254 24596 20260 24608
rect 20119 24568 20260 24596
rect 20119 24565 20131 24568
rect 20073 24559 20131 24565
rect 20254 24556 20260 24568
rect 20312 24596 20318 24608
rect 20456 24596 20484 24636
rect 27246 24624 27252 24636
rect 27304 24624 27310 24676
rect 20622 24596 20628 24608
rect 20312 24568 20484 24596
rect 20583 24568 20628 24596
rect 20312 24556 20318 24568
rect 20622 24556 20628 24568
rect 20680 24556 20686 24608
rect 21082 24556 21088 24608
rect 21140 24596 21146 24608
rect 21177 24599 21235 24605
rect 21177 24596 21189 24599
rect 21140 24568 21189 24596
rect 21140 24556 21146 24568
rect 21177 24565 21189 24568
rect 21223 24565 21235 24599
rect 21818 24596 21824 24608
rect 21779 24568 21824 24596
rect 21177 24559 21235 24565
rect 21818 24556 21824 24568
rect 21876 24556 21882 24608
rect 24121 24599 24179 24605
rect 24121 24565 24133 24599
rect 24167 24596 24179 24599
rect 24210 24596 24216 24608
rect 24167 24568 24216 24596
rect 24167 24565 24179 24568
rect 24121 24559 24179 24565
rect 24210 24556 24216 24568
rect 24268 24556 24274 24608
rect 1104 24506 26864 24528
rect 1104 24454 10315 24506
rect 10367 24454 10379 24506
rect 10431 24454 10443 24506
rect 10495 24454 10507 24506
rect 10559 24454 19648 24506
rect 19700 24454 19712 24506
rect 19764 24454 19776 24506
rect 19828 24454 19840 24506
rect 19892 24454 26864 24506
rect 1104 24432 26864 24454
rect 2133 24395 2191 24401
rect 2133 24361 2145 24395
rect 2179 24392 2191 24395
rect 2406 24392 2412 24404
rect 2179 24364 2412 24392
rect 2179 24361 2191 24364
rect 2133 24355 2191 24361
rect 2406 24352 2412 24364
rect 2464 24352 2470 24404
rect 4525 24395 4583 24401
rect 4525 24361 4537 24395
rect 4571 24392 4583 24395
rect 4982 24392 4988 24404
rect 4571 24364 4988 24392
rect 4571 24361 4583 24364
rect 4525 24355 4583 24361
rect 4982 24352 4988 24364
rect 5040 24352 5046 24404
rect 9674 24352 9680 24404
rect 9732 24392 9738 24404
rect 12713 24395 12771 24401
rect 9732 24364 10916 24392
rect 9732 24352 9738 24364
rect 1946 24284 1952 24336
rect 2004 24324 2010 24336
rect 2041 24327 2099 24333
rect 2041 24324 2053 24327
rect 2004 24296 2053 24324
rect 2004 24284 2010 24296
rect 2041 24293 2053 24296
rect 2087 24324 2099 24327
rect 5350 24324 5356 24336
rect 2087 24296 5356 24324
rect 2087 24293 2099 24296
rect 2041 24287 2099 24293
rect 5350 24284 5356 24296
rect 5408 24284 5414 24336
rect 9950 24284 9956 24336
rect 10008 24324 10014 24336
rect 10750 24327 10808 24333
rect 10750 24324 10762 24327
rect 10008 24296 10762 24324
rect 10008 24284 10014 24296
rect 10750 24293 10762 24296
rect 10796 24293 10808 24327
rect 10888 24324 10916 24364
rect 12713 24361 12725 24395
rect 12759 24392 12771 24395
rect 13078 24392 13084 24404
rect 12759 24364 13084 24392
rect 12759 24361 12771 24364
rect 12713 24355 12771 24361
rect 13078 24352 13084 24364
rect 13136 24352 13142 24404
rect 13446 24392 13452 24404
rect 13407 24364 13452 24392
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 15470 24392 15476 24404
rect 15431 24364 15476 24392
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 18598 24392 18604 24404
rect 18559 24364 18604 24392
rect 18598 24352 18604 24364
rect 18656 24392 18662 24404
rect 19521 24395 19579 24401
rect 19521 24392 19533 24395
rect 18656 24364 19533 24392
rect 18656 24352 18662 24364
rect 19521 24361 19533 24364
rect 19567 24361 19579 24395
rect 19521 24355 19579 24361
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19978 24392 19984 24404
rect 19935 24364 19984 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 21358 24392 21364 24404
rect 21319 24364 21364 24392
rect 21358 24352 21364 24364
rect 21416 24392 21422 24404
rect 21913 24395 21971 24401
rect 21913 24392 21925 24395
rect 21416 24364 21925 24392
rect 21416 24352 21422 24364
rect 21913 24361 21925 24364
rect 21959 24361 21971 24395
rect 21913 24355 21971 24361
rect 22649 24395 22707 24401
rect 22649 24361 22661 24395
rect 22695 24392 22707 24395
rect 24118 24392 24124 24404
rect 22695 24364 24124 24392
rect 22695 24361 22707 24364
rect 22649 24355 22707 24361
rect 24118 24352 24124 24364
rect 24176 24352 24182 24404
rect 24670 24392 24676 24404
rect 24631 24364 24676 24392
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 11330 24324 11336 24336
rect 10888 24296 11336 24324
rect 10750 24287 10808 24293
rect 11330 24284 11336 24296
rect 11388 24324 11394 24336
rect 14458 24324 14464 24336
rect 11388 24296 14464 24324
rect 11388 24284 11394 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 15102 24324 15108 24336
rect 15063 24296 15108 24324
rect 15102 24284 15108 24296
rect 15160 24284 15166 24336
rect 15194 24284 15200 24336
rect 15252 24324 15258 24336
rect 16206 24324 16212 24336
rect 15252 24296 16212 24324
rect 15252 24284 15258 24296
rect 16206 24284 16212 24296
rect 16264 24284 16270 24336
rect 16942 24324 16948 24336
rect 16903 24296 16948 24324
rect 16942 24284 16948 24296
rect 17000 24284 17006 24336
rect 18509 24327 18567 24333
rect 18509 24293 18521 24327
rect 18555 24324 18567 24327
rect 20622 24324 20628 24336
rect 18555 24296 20628 24324
rect 18555 24293 18567 24296
rect 18509 24287 18567 24293
rect 20622 24284 20628 24296
rect 20680 24284 20686 24336
rect 4893 24259 4951 24265
rect 4893 24225 4905 24259
rect 4939 24256 4951 24259
rect 5166 24256 5172 24268
rect 4939 24228 5172 24256
rect 4939 24225 4951 24228
rect 4893 24219 4951 24225
rect 5166 24216 5172 24228
rect 5224 24256 5230 24268
rect 6178 24256 6184 24268
rect 5224 24228 6184 24256
rect 5224 24216 5230 24228
rect 6178 24216 6184 24228
rect 6236 24216 6242 24268
rect 6908 24259 6966 24265
rect 6908 24225 6920 24259
rect 6954 24256 6966 24259
rect 7190 24256 7196 24268
rect 6954 24228 7196 24256
rect 6954 24225 6966 24228
rect 6908 24219 6966 24225
rect 7190 24216 7196 24228
rect 7248 24216 7254 24268
rect 13354 24256 13360 24268
rect 13267 24228 13360 24256
rect 13354 24216 13360 24228
rect 13412 24256 13418 24268
rect 13906 24256 13912 24268
rect 13412 24228 13912 24256
rect 13412 24216 13418 24228
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 14366 24216 14372 24268
rect 14424 24256 14430 24268
rect 14826 24256 14832 24268
rect 14424 24228 14832 24256
rect 14424 24216 14430 24228
rect 14826 24216 14832 24228
rect 14884 24216 14890 24268
rect 15286 24256 15292 24268
rect 15247 24228 15292 24256
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 19150 24256 19156 24268
rect 16960 24228 19012 24256
rect 19111 24228 19156 24256
rect 2317 24191 2375 24197
rect 2317 24157 2329 24191
rect 2363 24188 2375 24191
rect 2498 24188 2504 24200
rect 2363 24160 2504 24188
rect 2363 24157 2375 24160
rect 2317 24151 2375 24157
rect 2498 24148 2504 24160
rect 2556 24188 2562 24200
rect 2777 24191 2835 24197
rect 2777 24188 2789 24191
rect 2556 24160 2789 24188
rect 2556 24148 2562 24160
rect 2777 24157 2789 24160
rect 2823 24188 2835 24191
rect 3326 24188 3332 24200
rect 2823 24160 3332 24188
rect 2823 24157 2835 24160
rect 2777 24151 2835 24157
rect 3326 24148 3332 24160
rect 3384 24148 3390 24200
rect 3418 24148 3424 24200
rect 3476 24188 3482 24200
rect 3476 24160 4200 24188
rect 3476 24148 3482 24160
rect 3513 24123 3571 24129
rect 3513 24089 3525 24123
rect 3559 24120 3571 24123
rect 4062 24120 4068 24132
rect 3559 24092 4068 24120
rect 3559 24089 3571 24092
rect 3513 24083 3571 24089
rect 4062 24080 4068 24092
rect 4120 24080 4126 24132
rect 4172 24120 4200 24160
rect 4246 24148 4252 24200
rect 4304 24188 4310 24200
rect 4985 24191 5043 24197
rect 4985 24188 4997 24191
rect 4304 24160 4997 24188
rect 4304 24148 4310 24160
rect 4985 24157 4997 24160
rect 5031 24157 5043 24191
rect 4985 24151 5043 24157
rect 5077 24191 5135 24197
rect 5077 24157 5089 24191
rect 5123 24157 5135 24191
rect 5902 24188 5908 24200
rect 5863 24160 5908 24188
rect 5077 24151 5135 24157
rect 4172 24092 4476 24120
rect 1673 24055 1731 24061
rect 1673 24021 1685 24055
rect 1719 24052 1731 24055
rect 1762 24052 1768 24064
rect 1719 24024 1768 24052
rect 1719 24021 1731 24024
rect 1673 24015 1731 24021
rect 1762 24012 1768 24024
rect 1820 24012 1826 24064
rect 3142 24052 3148 24064
rect 3103 24024 3148 24052
rect 3142 24012 3148 24024
rect 3200 24012 3206 24064
rect 3881 24055 3939 24061
rect 3881 24021 3893 24055
rect 3927 24052 3939 24055
rect 4154 24052 4160 24064
rect 3927 24024 4160 24052
rect 3927 24021 3939 24024
rect 3881 24015 3939 24021
rect 4154 24012 4160 24024
rect 4212 24012 4218 24064
rect 4448 24061 4476 24092
rect 4433 24055 4491 24061
rect 4433 24021 4445 24055
rect 4479 24052 4491 24055
rect 5092 24052 5120 24151
rect 5902 24148 5908 24160
rect 5960 24148 5966 24200
rect 6546 24148 6552 24200
rect 6604 24188 6610 24200
rect 6641 24191 6699 24197
rect 6641 24188 6653 24191
rect 6604 24160 6653 24188
rect 6604 24148 6610 24160
rect 6641 24157 6653 24160
rect 6687 24157 6699 24191
rect 10502 24188 10508 24200
rect 10463 24160 10508 24188
rect 6641 24151 6699 24157
rect 10502 24148 10508 24160
rect 10560 24148 10566 24200
rect 11514 24148 11520 24200
rect 11572 24188 11578 24200
rect 12250 24188 12256 24200
rect 11572 24160 12256 24188
rect 11572 24148 11578 24160
rect 12250 24148 12256 24160
rect 12308 24188 12314 24200
rect 13446 24188 13452 24200
rect 12308 24160 13452 24188
rect 12308 24148 12314 24160
rect 13446 24148 13452 24160
rect 13504 24148 13510 24200
rect 13630 24188 13636 24200
rect 13591 24160 13636 24188
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 16960 24188 16988 24228
rect 14660 24160 16988 24188
rect 17037 24191 17095 24197
rect 13262 24080 13268 24132
rect 13320 24120 13326 24132
rect 14660 24120 14688 24160
rect 17037 24157 17049 24191
rect 17083 24157 17095 24191
rect 17037 24151 17095 24157
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24188 17279 24191
rect 17494 24188 17500 24200
rect 17267 24160 17500 24188
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 13320 24092 14688 24120
rect 14737 24123 14795 24129
rect 13320 24080 13326 24092
rect 14737 24089 14749 24123
rect 14783 24120 14795 24123
rect 14826 24120 14832 24132
rect 14783 24092 14832 24120
rect 14783 24089 14795 24092
rect 14737 24083 14795 24089
rect 14826 24080 14832 24092
rect 14884 24080 14890 24132
rect 16485 24123 16543 24129
rect 16485 24089 16497 24123
rect 16531 24120 16543 24123
rect 16942 24120 16948 24132
rect 16531 24092 16948 24120
rect 16531 24089 16543 24092
rect 16485 24083 16543 24089
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 17052 24120 17080 24151
rect 17494 24148 17500 24160
rect 17552 24188 17558 24200
rect 18693 24191 18751 24197
rect 18693 24188 18705 24191
rect 17552 24160 18705 24188
rect 17552 24148 17558 24160
rect 18693 24157 18705 24160
rect 18739 24157 18751 24191
rect 18984 24188 19012 24228
rect 19150 24216 19156 24228
rect 19208 24216 19214 24268
rect 19702 24256 19708 24268
rect 19663 24228 19708 24256
rect 19702 24216 19708 24228
rect 19760 24216 19766 24268
rect 21269 24259 21327 24265
rect 21269 24256 21281 24259
rect 19904 24228 21281 24256
rect 19904 24188 19932 24228
rect 21269 24225 21281 24228
rect 21315 24256 21327 24259
rect 21542 24256 21548 24268
rect 21315 24228 21548 24256
rect 21315 24225 21327 24228
rect 21269 24219 21327 24225
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 22465 24259 22523 24265
rect 22465 24225 22477 24259
rect 22511 24256 22523 24259
rect 22646 24256 22652 24268
rect 22511 24228 22652 24256
rect 22511 24225 22523 24228
rect 22465 24219 22523 24225
rect 22646 24216 22652 24228
rect 22704 24216 22710 24268
rect 24489 24259 24547 24265
rect 24489 24225 24501 24259
rect 24535 24256 24547 24259
rect 24670 24256 24676 24268
rect 24535 24228 24676 24256
rect 24535 24225 24547 24228
rect 24489 24219 24547 24225
rect 24670 24216 24676 24228
rect 24728 24216 24734 24268
rect 18984 24160 19932 24188
rect 18693 24151 18751 24157
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20346 24188 20352 24200
rect 20220 24160 20352 24188
rect 20220 24148 20226 24160
rect 20346 24148 20352 24160
rect 20404 24148 20410 24200
rect 21453 24191 21511 24197
rect 21453 24188 21465 24191
rect 20548 24160 21465 24188
rect 17678 24120 17684 24132
rect 17052 24092 17684 24120
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 18046 24120 18052 24132
rect 18007 24092 18052 24120
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 19978 24120 19984 24132
rect 19392 24092 19984 24120
rect 19392 24080 19398 24092
rect 19978 24080 19984 24092
rect 20036 24080 20042 24132
rect 20438 24080 20444 24132
rect 20496 24120 20502 24132
rect 20548 24129 20576 24160
rect 21453 24157 21465 24160
rect 21499 24157 21511 24191
rect 21453 24151 21511 24157
rect 20533 24123 20591 24129
rect 20533 24120 20545 24123
rect 20496 24092 20545 24120
rect 20496 24080 20502 24092
rect 20533 24089 20545 24092
rect 20579 24089 20591 24123
rect 20898 24120 20904 24132
rect 20859 24092 20904 24120
rect 20533 24083 20591 24089
rect 20898 24080 20904 24092
rect 20956 24080 20962 24132
rect 5629 24055 5687 24061
rect 5629 24052 5641 24055
rect 4479 24024 5641 24052
rect 4479 24021 4491 24024
rect 4433 24015 4491 24021
rect 5629 24021 5641 24024
rect 5675 24052 5687 24055
rect 5994 24052 6000 24064
rect 5675 24024 6000 24052
rect 5675 24021 5687 24024
rect 5629 24015 5687 24021
rect 5994 24012 6000 24024
rect 6052 24012 6058 24064
rect 6549 24055 6607 24061
rect 6549 24021 6561 24055
rect 6595 24052 6607 24055
rect 7282 24052 7288 24064
rect 6595 24024 7288 24052
rect 6595 24021 6607 24024
rect 6549 24015 6607 24021
rect 7282 24012 7288 24024
rect 7340 24012 7346 24064
rect 7558 24012 7564 24064
rect 7616 24052 7622 24064
rect 8021 24055 8079 24061
rect 8021 24052 8033 24055
rect 7616 24024 8033 24052
rect 7616 24012 7622 24024
rect 8021 24021 8033 24024
rect 8067 24021 8079 24055
rect 8021 24015 8079 24021
rect 8665 24055 8723 24061
rect 8665 24021 8677 24055
rect 8711 24052 8723 24055
rect 9306 24052 9312 24064
rect 8711 24024 9312 24052
rect 8711 24021 8723 24024
rect 8665 24015 8723 24021
rect 9306 24012 9312 24024
rect 9364 24012 9370 24064
rect 9490 24052 9496 24064
rect 9451 24024 9496 24052
rect 9490 24012 9496 24024
rect 9548 24012 9554 24064
rect 9950 24052 9956 24064
rect 9911 24024 9956 24052
rect 9950 24012 9956 24024
rect 10008 24012 10014 24064
rect 10413 24055 10471 24061
rect 10413 24021 10425 24055
rect 10459 24052 10471 24055
rect 11238 24052 11244 24064
rect 10459 24024 11244 24052
rect 10459 24021 10471 24024
rect 10413 24015 10471 24021
rect 11238 24012 11244 24024
rect 11296 24012 11302 24064
rect 11422 24012 11428 24064
rect 11480 24052 11486 24064
rect 11885 24055 11943 24061
rect 11885 24052 11897 24055
rect 11480 24024 11897 24052
rect 11480 24012 11486 24024
rect 11885 24021 11897 24024
rect 11931 24021 11943 24055
rect 12986 24052 12992 24064
rect 12947 24024 12992 24052
rect 11885 24015 11943 24021
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 14185 24055 14243 24061
rect 14185 24021 14197 24055
rect 14231 24052 14243 24055
rect 14458 24052 14464 24064
rect 14231 24024 14464 24052
rect 14231 24021 14243 24024
rect 14185 24015 14243 24021
rect 14458 24012 14464 24024
rect 14516 24012 14522 24064
rect 15746 24012 15752 24064
rect 15804 24052 15810 24064
rect 15841 24055 15899 24061
rect 15841 24052 15853 24055
rect 15804 24024 15853 24052
rect 15804 24012 15810 24024
rect 15841 24021 15853 24024
rect 15887 24021 15899 24055
rect 16574 24052 16580 24064
rect 16535 24024 16580 24052
rect 15841 24015 15899 24021
rect 16574 24012 16580 24024
rect 16632 24012 16638 24064
rect 16960 24052 16988 24080
rect 17218 24052 17224 24064
rect 16960 24024 17224 24052
rect 17218 24012 17224 24024
rect 17276 24012 17282 24064
rect 18138 24052 18144 24064
rect 18099 24024 18144 24052
rect 18138 24012 18144 24024
rect 18196 24012 18202 24064
rect 1104 23962 26864 23984
rect 1104 23910 5648 23962
rect 5700 23910 5712 23962
rect 5764 23910 5776 23962
rect 5828 23910 5840 23962
rect 5892 23910 14982 23962
rect 15034 23910 15046 23962
rect 15098 23910 15110 23962
rect 15162 23910 15174 23962
rect 15226 23910 24315 23962
rect 24367 23910 24379 23962
rect 24431 23910 24443 23962
rect 24495 23910 24507 23962
rect 24559 23910 26864 23962
rect 1104 23888 26864 23910
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 3605 23851 3663 23857
rect 3605 23848 3617 23851
rect 3568 23820 3617 23848
rect 3568 23808 3574 23820
rect 3605 23817 3617 23820
rect 3651 23817 3663 23851
rect 6178 23848 6184 23860
rect 6139 23820 6184 23848
rect 3605 23811 3663 23817
rect 6178 23808 6184 23820
rect 6236 23808 6242 23860
rect 6546 23848 6552 23860
rect 6507 23820 6552 23848
rect 6546 23808 6552 23820
rect 6604 23848 6610 23860
rect 8021 23851 8079 23857
rect 8021 23848 8033 23851
rect 6604 23820 8033 23848
rect 6604 23808 6610 23820
rect 8021 23817 8033 23820
rect 8067 23817 8079 23851
rect 8021 23811 8079 23817
rect 5169 23783 5227 23789
rect 5169 23780 5181 23783
rect 4080 23752 5181 23780
rect 2038 23672 2044 23724
rect 2096 23712 2102 23724
rect 2133 23715 2191 23721
rect 2133 23712 2145 23715
rect 2096 23684 2145 23712
rect 2096 23672 2102 23684
rect 2133 23681 2145 23684
rect 2179 23681 2191 23715
rect 2133 23675 2191 23681
rect 2317 23715 2375 23721
rect 2317 23681 2329 23715
rect 2363 23712 2375 23715
rect 2498 23712 2504 23724
rect 2363 23684 2504 23712
rect 2363 23681 2375 23684
rect 2317 23675 2375 23681
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 3142 23672 3148 23724
rect 3200 23712 3206 23724
rect 4080 23721 4108 23752
rect 5169 23749 5181 23752
rect 5215 23749 5227 23783
rect 5169 23743 5227 23749
rect 4065 23715 4123 23721
rect 4065 23712 4077 23715
rect 3200 23684 4077 23712
rect 3200 23672 3206 23684
rect 4065 23681 4077 23684
rect 4111 23681 4123 23715
rect 4065 23675 4123 23681
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23712 4307 23715
rect 4430 23712 4436 23724
rect 4295 23684 4436 23712
rect 4295 23681 4307 23684
rect 4249 23675 4307 23681
rect 3513 23647 3571 23653
rect 3513 23613 3525 23647
rect 3559 23644 3571 23647
rect 4264 23644 4292 23675
rect 4430 23672 4436 23684
rect 4488 23672 4494 23724
rect 4709 23715 4767 23721
rect 4709 23681 4721 23715
rect 4755 23712 4767 23715
rect 5534 23712 5540 23724
rect 4755 23684 5540 23712
rect 4755 23681 4767 23684
rect 4709 23675 4767 23681
rect 5534 23672 5540 23684
rect 5592 23712 5598 23724
rect 5629 23715 5687 23721
rect 5629 23712 5641 23715
rect 5592 23684 5641 23712
rect 5592 23672 5598 23684
rect 5629 23681 5641 23684
rect 5675 23681 5687 23715
rect 5629 23675 5687 23681
rect 5813 23715 5871 23721
rect 5813 23681 5825 23715
rect 5859 23712 5871 23715
rect 5994 23712 6000 23724
rect 5859 23684 6000 23712
rect 5859 23681 5871 23684
rect 5813 23675 5871 23681
rect 5994 23672 6000 23684
rect 6052 23672 6058 23724
rect 7466 23712 7472 23724
rect 7427 23684 7472 23712
rect 7466 23672 7472 23684
rect 7524 23672 7530 23724
rect 8036 23712 8064 23811
rect 9950 23808 9956 23860
rect 10008 23848 10014 23860
rect 10137 23851 10195 23857
rect 10137 23848 10149 23851
rect 10008 23820 10149 23848
rect 10008 23808 10014 23820
rect 10137 23817 10149 23820
rect 10183 23817 10195 23851
rect 12250 23848 12256 23860
rect 12211 23820 12256 23848
rect 10137 23811 10195 23817
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12452 23820 13584 23848
rect 10962 23740 10968 23792
rect 11020 23780 11026 23792
rect 11020 23752 11468 23780
rect 11020 23740 11026 23752
rect 11440 23724 11468 23752
rect 11790 23740 11796 23792
rect 11848 23780 11854 23792
rect 12452 23780 12480 23820
rect 11848 23752 12480 23780
rect 11848 23740 11854 23752
rect 8205 23715 8263 23721
rect 8205 23712 8217 23715
rect 8036 23684 8217 23712
rect 8205 23681 8217 23684
rect 8251 23681 8263 23715
rect 11238 23712 11244 23724
rect 11199 23684 11244 23712
rect 8205 23675 8263 23681
rect 3559 23616 4292 23644
rect 6825 23647 6883 23653
rect 3559 23613 3571 23616
rect 3513 23607 3571 23613
rect 6825 23613 6837 23647
rect 6871 23644 6883 23647
rect 7484 23644 7512 23672
rect 6871 23616 7512 23644
rect 8220 23644 8248 23675
rect 11238 23672 11244 23684
rect 11296 23672 11302 23724
rect 11422 23712 11428 23724
rect 11383 23684 11428 23712
rect 11422 23672 11428 23684
rect 11480 23672 11486 23724
rect 13556 23712 13584 23820
rect 13630 23808 13636 23860
rect 13688 23848 13694 23860
rect 13998 23848 14004 23860
rect 13688 23820 14004 23848
rect 13688 23808 13694 23820
rect 13998 23808 14004 23820
rect 14056 23848 14062 23860
rect 14369 23851 14427 23857
rect 14369 23848 14381 23851
rect 14056 23820 14381 23848
rect 14056 23808 14062 23820
rect 14369 23817 14381 23820
rect 14415 23817 14427 23851
rect 14369 23811 14427 23817
rect 14458 23808 14464 23860
rect 14516 23848 14522 23860
rect 20254 23848 20260 23860
rect 14516 23820 20260 23848
rect 14516 23808 14522 23820
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 20533 23851 20591 23857
rect 20533 23817 20545 23851
rect 20579 23848 20591 23851
rect 20622 23848 20628 23860
rect 20579 23820 20628 23848
rect 20579 23817 20591 23820
rect 20533 23811 20591 23817
rect 20622 23808 20628 23820
rect 20680 23808 20686 23860
rect 21542 23848 21548 23860
rect 21503 23820 21548 23848
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 21910 23808 21916 23860
rect 21968 23848 21974 23860
rect 22281 23851 22339 23857
rect 22281 23848 22293 23851
rect 21968 23820 22293 23848
rect 21968 23808 21974 23820
rect 22281 23817 22293 23820
rect 22327 23817 22339 23851
rect 24762 23848 24768 23860
rect 24723 23820 24768 23848
rect 22281 23811 22339 23817
rect 24762 23808 24768 23820
rect 24820 23808 24826 23860
rect 15194 23780 15200 23792
rect 15155 23752 15200 23780
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 16298 23740 16304 23792
rect 16356 23780 16362 23792
rect 16482 23780 16488 23792
rect 16356 23752 16488 23780
rect 16356 23740 16362 23752
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 13556 23684 15424 23712
rect 8294 23644 8300 23656
rect 8220 23616 8300 23644
rect 6871 23613 6883 23616
rect 6825 23607 6883 23613
rect 8294 23604 8300 23616
rect 8352 23604 8358 23656
rect 10502 23604 10508 23656
rect 10560 23644 10566 23656
rect 10597 23647 10655 23653
rect 10597 23644 10609 23647
rect 10560 23616 10609 23644
rect 10560 23604 10566 23616
rect 10597 23613 10609 23616
rect 10643 23644 10655 23647
rect 10778 23644 10784 23656
rect 10643 23616 10784 23644
rect 10643 23613 10655 23616
rect 10597 23607 10655 23613
rect 10778 23604 10784 23616
rect 10836 23604 10842 23656
rect 11256 23644 11284 23672
rect 12342 23644 12348 23656
rect 11256 23616 12348 23644
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12437 23647 12495 23653
rect 12437 23613 12449 23647
rect 12483 23644 12495 23647
rect 12526 23644 12532 23656
rect 12483 23616 12532 23644
rect 12483 23613 12495 23616
rect 12437 23607 12495 23613
rect 12526 23604 12532 23616
rect 12584 23644 12590 23656
rect 14737 23647 14795 23653
rect 14737 23644 14749 23647
rect 12584 23616 14749 23644
rect 12584 23604 12590 23616
rect 14737 23613 14749 23616
rect 14783 23644 14795 23647
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 14783 23616 15301 23644
rect 14783 23613 14795 23616
rect 14737 23607 14795 23613
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15396 23644 15424 23684
rect 20438 23672 20444 23724
rect 20496 23712 20502 23724
rect 21085 23715 21143 23721
rect 21085 23712 21097 23715
rect 20496 23684 21097 23712
rect 20496 23672 20502 23684
rect 21085 23681 21097 23684
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 24302 23672 24308 23724
rect 24360 23712 24366 23724
rect 24670 23712 24676 23724
rect 24360 23684 24676 23712
rect 24360 23672 24366 23684
rect 24670 23672 24676 23684
rect 24728 23712 24734 23724
rect 25133 23715 25191 23721
rect 25133 23712 25145 23715
rect 24728 23684 25145 23712
rect 24728 23672 24734 23684
rect 25133 23681 25145 23684
rect 25179 23681 25191 23715
rect 25133 23675 25191 23681
rect 15562 23653 15568 23656
rect 15545 23647 15568 23653
rect 15545 23644 15557 23647
rect 15396 23616 15557 23644
rect 15289 23607 15347 23613
rect 15545 23613 15557 23616
rect 15620 23644 15626 23656
rect 15620 23616 15693 23644
rect 15545 23607 15568 23613
rect 15562 23604 15568 23607
rect 15620 23604 15626 23616
rect 16482 23604 16488 23656
rect 16540 23644 16546 23656
rect 17773 23647 17831 23653
rect 17773 23644 17785 23647
rect 16540 23616 17785 23644
rect 16540 23604 16546 23616
rect 17773 23613 17785 23616
rect 17819 23644 17831 23647
rect 18049 23647 18107 23653
rect 18049 23644 18061 23647
rect 17819 23616 18061 23644
rect 17819 23613 17831 23616
rect 17773 23607 17831 23613
rect 18049 23613 18061 23616
rect 18095 23644 18107 23647
rect 18690 23644 18696 23656
rect 18095 23616 18696 23644
rect 18095 23613 18107 23616
rect 18049 23607 18107 23613
rect 18690 23604 18696 23616
rect 18748 23604 18754 23656
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23613 22155 23647
rect 24581 23647 24639 23653
rect 24581 23644 24593 23647
rect 22097 23607 22155 23613
rect 24504 23616 24593 23644
rect 2041 23579 2099 23585
rect 2041 23545 2053 23579
rect 2087 23576 2099 23579
rect 2222 23576 2228 23588
rect 2087 23548 2228 23576
rect 2087 23545 2099 23548
rect 2041 23539 2099 23545
rect 2222 23536 2228 23548
rect 2280 23536 2286 23588
rect 5077 23579 5135 23585
rect 5077 23545 5089 23579
rect 5123 23576 5135 23579
rect 5537 23579 5595 23585
rect 5537 23576 5549 23579
rect 5123 23548 5549 23576
rect 5123 23545 5135 23548
rect 5077 23539 5135 23545
rect 5537 23545 5549 23548
rect 5583 23576 5595 23579
rect 6086 23576 6092 23588
rect 5583 23548 6092 23576
rect 5583 23545 5595 23548
rect 5537 23539 5595 23545
rect 6086 23536 6092 23548
rect 6144 23536 6150 23588
rect 8472 23579 8530 23585
rect 8472 23545 8484 23579
rect 8518 23576 8530 23579
rect 9306 23576 9312 23588
rect 8518 23548 9312 23576
rect 8518 23545 8530 23548
rect 8472 23539 8530 23545
rect 9306 23536 9312 23548
rect 9364 23536 9370 23588
rect 11885 23579 11943 23585
rect 11885 23545 11897 23579
rect 11931 23576 11943 23579
rect 12618 23576 12624 23588
rect 11931 23548 12624 23576
rect 11931 23545 11943 23548
rect 11885 23539 11943 23545
rect 12618 23536 12624 23548
rect 12676 23585 12682 23588
rect 12676 23579 12740 23585
rect 12676 23545 12694 23579
rect 12728 23545 12740 23579
rect 18294 23579 18352 23585
rect 18294 23576 18306 23579
rect 12676 23539 12740 23545
rect 17512 23548 18306 23576
rect 12676 23536 12682 23539
rect 17512 23520 17540 23548
rect 18294 23545 18306 23548
rect 18340 23545 18352 23579
rect 18294 23539 18352 23545
rect 18598 23536 18604 23588
rect 18656 23576 18662 23588
rect 18656 23548 19656 23576
rect 18656 23536 18662 23548
rect 1486 23468 1492 23520
rect 1544 23508 1550 23520
rect 1673 23511 1731 23517
rect 1673 23508 1685 23511
rect 1544 23480 1685 23508
rect 1544 23468 1550 23480
rect 1673 23477 1685 23480
rect 1719 23477 1731 23511
rect 1673 23471 1731 23477
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 3145 23511 3203 23517
rect 2832 23480 2877 23508
rect 2832 23468 2838 23480
rect 3145 23477 3157 23511
rect 3191 23508 3203 23511
rect 3326 23508 3332 23520
rect 3191 23480 3332 23508
rect 3191 23477 3203 23480
rect 3145 23471 3203 23477
rect 3326 23468 3332 23480
rect 3384 23468 3390 23520
rect 3694 23468 3700 23520
rect 3752 23508 3758 23520
rect 3973 23511 4031 23517
rect 3973 23508 3985 23511
rect 3752 23480 3985 23508
rect 3752 23468 3758 23480
rect 3973 23477 3985 23480
rect 4019 23477 4031 23511
rect 7006 23508 7012 23520
rect 6967 23480 7012 23508
rect 3973 23471 4031 23477
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 8570 23468 8576 23520
rect 8628 23508 8634 23520
rect 9585 23511 9643 23517
rect 9585 23508 9597 23511
rect 8628 23480 9597 23508
rect 8628 23468 8634 23480
rect 9585 23477 9597 23480
rect 9631 23477 9643 23511
rect 9585 23471 9643 23477
rect 9674 23468 9680 23520
rect 9732 23508 9738 23520
rect 10781 23511 10839 23517
rect 10781 23508 10793 23511
rect 9732 23480 10793 23508
rect 9732 23468 9738 23480
rect 10781 23477 10793 23480
rect 10827 23477 10839 23511
rect 11146 23508 11152 23520
rect 11107 23480 11152 23508
rect 10781 23471 10839 23477
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 13814 23508 13820 23520
rect 13775 23480 13820 23508
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 16669 23511 16727 23517
rect 16669 23477 16681 23511
rect 16715 23508 16727 23511
rect 16942 23508 16948 23520
rect 16715 23480 16948 23508
rect 16715 23477 16727 23480
rect 16669 23471 16727 23477
rect 16942 23468 16948 23480
rect 17000 23468 17006 23520
rect 17494 23508 17500 23520
rect 17455 23480 17500 23508
rect 17494 23468 17500 23480
rect 17552 23468 17558 23520
rect 19429 23511 19487 23517
rect 19429 23477 19441 23511
rect 19475 23508 19487 23511
rect 19518 23508 19524 23520
rect 19475 23480 19524 23508
rect 19475 23477 19487 23480
rect 19429 23471 19487 23477
rect 19518 23468 19524 23480
rect 19576 23468 19582 23520
rect 19628 23508 19656 23548
rect 19702 23536 19708 23588
rect 19760 23576 19766 23588
rect 20073 23579 20131 23585
rect 20073 23576 20085 23579
rect 19760 23548 20085 23576
rect 19760 23536 19766 23548
rect 20073 23545 20085 23548
rect 20119 23576 20131 23579
rect 20622 23576 20628 23588
rect 20119 23548 20628 23576
rect 20119 23545 20131 23548
rect 20073 23539 20131 23545
rect 20622 23536 20628 23548
rect 20680 23536 20686 23588
rect 20714 23536 20720 23588
rect 20772 23576 20778 23588
rect 20901 23579 20959 23585
rect 20901 23576 20913 23579
rect 20772 23548 20913 23576
rect 20772 23536 20778 23548
rect 20901 23545 20913 23548
rect 20947 23576 20959 23579
rect 22002 23576 22008 23588
rect 20947 23548 22008 23576
rect 20947 23545 20959 23548
rect 20901 23539 20959 23545
rect 22002 23536 22008 23548
rect 22060 23536 22066 23588
rect 20349 23511 20407 23517
rect 20349 23508 20361 23511
rect 19628 23480 20361 23508
rect 20349 23477 20361 23480
rect 20395 23508 20407 23511
rect 20990 23508 20996 23520
rect 20395 23480 20996 23508
rect 20395 23477 20407 23480
rect 20349 23471 20407 23477
rect 20990 23468 20996 23480
rect 21048 23468 21054 23520
rect 21910 23508 21916 23520
rect 21823 23480 21916 23508
rect 21910 23468 21916 23480
rect 21968 23508 21974 23520
rect 22112 23508 22140 23607
rect 24504 23520 24532 23616
rect 24581 23613 24593 23616
rect 24627 23613 24639 23647
rect 24581 23607 24639 23613
rect 22646 23508 22652 23520
rect 21968 23480 22140 23508
rect 22607 23480 22652 23508
rect 21968 23468 21974 23480
rect 22646 23468 22652 23480
rect 22704 23468 22710 23520
rect 24486 23508 24492 23520
rect 24447 23480 24492 23508
rect 24486 23468 24492 23480
rect 24544 23468 24550 23520
rect 1104 23418 26864 23440
rect 1104 23366 10315 23418
rect 10367 23366 10379 23418
rect 10431 23366 10443 23418
rect 10495 23366 10507 23418
rect 10559 23366 19648 23418
rect 19700 23366 19712 23418
rect 19764 23366 19776 23418
rect 19828 23366 19840 23418
rect 19892 23366 26864 23418
rect 1104 23344 26864 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 1670 23264 1676 23316
rect 1728 23304 1734 23316
rect 1946 23304 1952 23316
rect 1728 23276 1952 23304
rect 1728 23264 1734 23276
rect 1946 23264 1952 23276
rect 2004 23264 2010 23316
rect 2406 23304 2412 23316
rect 2367 23276 2412 23304
rect 2406 23264 2412 23276
rect 2464 23264 2470 23316
rect 2777 23307 2835 23313
rect 2777 23273 2789 23307
rect 2823 23304 2835 23307
rect 2866 23304 2872 23316
rect 2823 23276 2872 23304
rect 2823 23273 2835 23276
rect 2777 23267 2835 23273
rect 2866 23264 2872 23276
rect 2924 23264 2930 23316
rect 3326 23304 3332 23316
rect 3287 23276 3332 23304
rect 3326 23264 3332 23276
rect 3384 23264 3390 23316
rect 4246 23264 4252 23316
rect 4304 23304 4310 23316
rect 4522 23304 4528 23316
rect 4304 23276 4528 23304
rect 4304 23264 4310 23276
rect 4522 23264 4528 23276
rect 4580 23264 4586 23316
rect 7190 23304 7196 23316
rect 7151 23276 7196 23304
rect 7190 23264 7196 23276
rect 7248 23304 7254 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 7248 23276 7849 23304
rect 7248 23264 7254 23276
rect 7837 23273 7849 23276
rect 7883 23273 7895 23307
rect 7837 23267 7895 23273
rect 9125 23307 9183 23313
rect 9125 23273 9137 23307
rect 9171 23304 9183 23307
rect 9766 23304 9772 23316
rect 9171 23276 9772 23304
rect 9171 23273 9183 23276
rect 9125 23267 9183 23273
rect 3602 23236 3608 23248
rect 1412 23208 3608 23236
rect 1412 23177 1440 23208
rect 3602 23196 3608 23208
rect 3660 23196 3666 23248
rect 5442 23236 5448 23248
rect 4908 23208 5448 23236
rect 1389 23171 1447 23177
rect 1389 23137 1401 23171
rect 1435 23137 1447 23171
rect 1389 23131 1447 23137
rect 3237 23171 3295 23177
rect 3237 23137 3249 23171
rect 3283 23168 3295 23171
rect 3418 23168 3424 23180
rect 3283 23140 3424 23168
rect 3283 23137 3295 23140
rect 3237 23131 3295 23137
rect 3418 23128 3424 23140
rect 3476 23128 3482 23180
rect 4908 23177 4936 23208
rect 5442 23196 5448 23208
rect 5500 23196 5506 23248
rect 7852 23236 7880 23267
rect 9766 23264 9772 23276
rect 9824 23304 9830 23316
rect 10045 23307 10103 23313
rect 10045 23304 10057 23307
rect 9824 23276 10057 23304
rect 9824 23264 9830 23276
rect 10045 23273 10057 23276
rect 10091 23273 10103 23307
rect 10045 23267 10103 23273
rect 10134 23264 10140 23316
rect 10192 23304 10198 23316
rect 11241 23307 11299 23313
rect 11241 23304 11253 23307
rect 10192 23276 11253 23304
rect 10192 23264 10198 23276
rect 11241 23273 11253 23276
rect 11287 23273 11299 23307
rect 12802 23304 12808 23316
rect 12763 23276 12808 23304
rect 11241 23267 11299 23273
rect 12802 23264 12808 23276
rect 12860 23264 12866 23316
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 13173 23307 13231 23313
rect 13173 23304 13185 23307
rect 13136 23276 13185 23304
rect 13136 23264 13142 23276
rect 13173 23273 13185 23276
rect 13219 23273 13231 23307
rect 13173 23267 13231 23273
rect 15562 23264 15568 23316
rect 15620 23304 15626 23316
rect 15841 23307 15899 23313
rect 15841 23304 15853 23307
rect 15620 23276 15853 23304
rect 15620 23264 15626 23276
rect 15841 23273 15853 23276
rect 15887 23273 15899 23307
rect 15841 23267 15899 23273
rect 16666 23264 16672 23316
rect 16724 23264 16730 23316
rect 18138 23264 18144 23316
rect 18196 23304 18202 23316
rect 18785 23307 18843 23313
rect 18785 23304 18797 23307
rect 18196 23276 18797 23304
rect 18196 23264 18202 23276
rect 18785 23273 18797 23276
rect 18831 23304 18843 23307
rect 19337 23307 19395 23313
rect 19337 23304 19349 23307
rect 18831 23276 19349 23304
rect 18831 23273 18843 23276
rect 18785 23267 18843 23273
rect 19337 23273 19349 23276
rect 19383 23273 19395 23307
rect 19337 23267 19395 23273
rect 20257 23307 20315 23313
rect 20257 23273 20269 23307
rect 20303 23304 20315 23307
rect 20438 23304 20444 23316
rect 20303 23276 20444 23304
rect 20303 23273 20315 23276
rect 20257 23267 20315 23273
rect 20438 23264 20444 23276
rect 20496 23264 20502 23316
rect 20625 23307 20683 23313
rect 20625 23273 20637 23307
rect 20671 23304 20683 23307
rect 20714 23304 20720 23316
rect 20671 23276 20720 23304
rect 20671 23273 20683 23276
rect 20625 23267 20683 23273
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 22002 23304 22008 23316
rect 21963 23276 22008 23304
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 22830 23264 22836 23316
rect 22888 23304 22894 23316
rect 22925 23307 22983 23313
rect 22925 23304 22937 23307
rect 22888 23276 22937 23304
rect 22888 23264 22894 23276
rect 22925 23273 22937 23276
rect 22971 23273 22983 23307
rect 24762 23304 24768 23316
rect 24723 23276 24768 23304
rect 22925 23267 22983 23273
rect 24762 23264 24768 23276
rect 24820 23264 24826 23316
rect 8570 23236 8576 23248
rect 7852 23208 8576 23236
rect 8570 23196 8576 23208
rect 8628 23196 8634 23248
rect 10873 23239 10931 23245
rect 10873 23205 10885 23239
rect 10919 23236 10931 23239
rect 10962 23236 10968 23248
rect 10919 23208 10968 23236
rect 10919 23205 10931 23208
rect 10873 23199 10931 23205
rect 4893 23171 4951 23177
rect 4893 23137 4905 23171
rect 4939 23137 4951 23171
rect 4893 23131 4951 23137
rect 5160 23171 5218 23177
rect 5160 23137 5172 23171
rect 5206 23168 5218 23171
rect 5994 23168 6000 23180
rect 5206 23140 6000 23168
rect 5206 23137 5218 23140
rect 5160 23131 5218 23137
rect 5994 23128 6000 23140
rect 6052 23128 6058 23180
rect 8389 23171 8447 23177
rect 8389 23168 8401 23171
rect 8312 23140 8401 23168
rect 2317 23103 2375 23109
rect 2317 23069 2329 23103
rect 2363 23100 2375 23103
rect 2406 23100 2412 23112
rect 2363 23072 2412 23100
rect 2363 23069 2375 23072
rect 2317 23063 2375 23069
rect 2406 23060 2412 23072
rect 2464 23060 2470 23112
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 1949 22967 2007 22973
rect 1949 22933 1961 22967
rect 1995 22964 2007 22967
rect 2406 22964 2412 22976
rect 1995 22936 2412 22964
rect 1995 22933 2007 22936
rect 1949 22927 2007 22933
rect 2406 22924 2412 22936
rect 2464 22964 2470 22976
rect 2774 22964 2780 22976
rect 2464 22936 2780 22964
rect 2464 22924 2470 22936
rect 2774 22924 2780 22936
rect 2832 22924 2838 22976
rect 2884 22964 2912 23063
rect 3068 23032 3096 23063
rect 3237 23035 3295 23041
rect 3237 23032 3249 23035
rect 3068 23004 3249 23032
rect 3237 23001 3249 23004
rect 3283 23001 3295 23035
rect 3237 22995 3295 23001
rect 3513 23035 3571 23041
rect 3513 23001 3525 23035
rect 3559 23032 3571 23035
rect 3602 23032 3608 23044
rect 3559 23004 3608 23032
rect 3559 23001 3571 23004
rect 3513 22995 3571 23001
rect 3602 22992 3608 23004
rect 3660 22992 3666 23044
rect 8018 23032 8024 23044
rect 7979 23004 8024 23032
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 8312 23032 8340 23140
rect 8389 23137 8401 23140
rect 8435 23137 8447 23171
rect 8389 23131 8447 23137
rect 8478 23100 8484 23112
rect 8439 23072 8484 23100
rect 8478 23060 8484 23072
rect 8536 23060 8542 23112
rect 8588 23109 8616 23196
rect 9490 23168 9496 23180
rect 9451 23140 9496 23168
rect 9490 23128 9496 23140
rect 9548 23128 9554 23180
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 9306 23060 9312 23112
rect 9364 23100 9370 23112
rect 10321 23103 10379 23109
rect 10321 23100 10333 23103
rect 9364 23072 10333 23100
rect 9364 23060 9370 23072
rect 10321 23069 10333 23072
rect 10367 23100 10379 23103
rect 10888 23100 10916 23199
rect 10962 23196 10968 23208
rect 11020 23196 11026 23248
rect 11701 23239 11759 23245
rect 11701 23205 11713 23239
rect 11747 23236 11759 23239
rect 11790 23236 11796 23248
rect 11747 23208 11796 23236
rect 11747 23205 11759 23208
rect 11701 23199 11759 23205
rect 11790 23196 11796 23208
rect 11848 23196 11854 23248
rect 13906 23236 13912 23248
rect 13819 23208 13912 23236
rect 13906 23196 13912 23208
rect 13964 23236 13970 23248
rect 16684 23236 16712 23264
rect 13964 23208 16712 23236
rect 16752 23239 16810 23245
rect 13964 23196 13970 23208
rect 16752 23205 16764 23239
rect 16798 23236 16810 23239
rect 16942 23236 16948 23248
rect 16798 23208 16948 23236
rect 16798 23205 16810 23208
rect 16752 23199 16810 23205
rect 16942 23196 16948 23208
rect 17000 23196 17006 23248
rect 23474 23236 23480 23248
rect 23435 23208 23480 23236
rect 23474 23196 23480 23208
rect 23532 23196 23538 23248
rect 11054 23128 11060 23180
rect 11112 23168 11118 23180
rect 11609 23171 11667 23177
rect 11609 23168 11621 23171
rect 11112 23140 11621 23168
rect 11112 23128 11118 23140
rect 11609 23137 11621 23140
rect 11655 23137 11667 23171
rect 11609 23131 11667 23137
rect 13265 23171 13323 23177
rect 13265 23137 13277 23171
rect 13311 23168 13323 23171
rect 13538 23168 13544 23180
rect 13311 23140 13544 23168
rect 13311 23137 13323 23140
rect 13265 23131 13323 23137
rect 13538 23128 13544 23140
rect 13596 23168 13602 23180
rect 14737 23171 14795 23177
rect 14737 23168 14749 23171
rect 13596 23140 14749 23168
rect 13596 23128 13602 23140
rect 14737 23137 14749 23140
rect 14783 23137 14795 23171
rect 14737 23131 14795 23137
rect 15289 23171 15347 23177
rect 15289 23137 15301 23171
rect 15335 23168 15347 23171
rect 15378 23168 15384 23180
rect 15335 23140 15384 23168
rect 15335 23137 15347 23140
rect 15289 23131 15347 23137
rect 15378 23128 15384 23140
rect 15436 23128 15442 23180
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 19392 23140 19441 23168
rect 19392 23128 19398 23140
rect 19429 23137 19441 23140
rect 19475 23137 19487 23171
rect 19429 23131 19487 23137
rect 20162 23128 20168 23180
rect 20220 23168 20226 23180
rect 20438 23168 20444 23180
rect 20220 23140 20444 23168
rect 20220 23128 20226 23140
rect 20438 23128 20444 23140
rect 20496 23128 20502 23180
rect 21269 23171 21327 23177
rect 21269 23137 21281 23171
rect 21315 23168 21327 23171
rect 21634 23168 21640 23180
rect 21315 23140 21640 23168
rect 21315 23137 21327 23140
rect 21269 23131 21327 23137
rect 21634 23128 21640 23140
rect 21692 23128 21698 23180
rect 22830 23168 22836 23180
rect 22791 23140 22836 23168
rect 22830 23128 22836 23140
rect 22888 23128 22894 23180
rect 24581 23171 24639 23177
rect 24581 23137 24593 23171
rect 24627 23168 24639 23171
rect 24670 23168 24676 23180
rect 24627 23140 24676 23168
rect 24627 23137 24639 23140
rect 24581 23131 24639 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 10367 23072 10916 23100
rect 10367 23069 10379 23072
rect 10321 23063 10379 23069
rect 11146 23060 11152 23112
rect 11204 23100 11210 23112
rect 11793 23103 11851 23109
rect 11793 23100 11805 23103
rect 11204 23072 11805 23100
rect 11204 23060 11210 23072
rect 11793 23069 11805 23072
rect 11839 23100 11851 23103
rect 12158 23100 12164 23112
rect 11839 23072 12164 23100
rect 11839 23069 11851 23072
rect 11793 23063 11851 23069
rect 12158 23060 12164 23072
rect 12216 23100 12222 23112
rect 13449 23103 13507 23109
rect 13449 23100 13461 23103
rect 12216 23072 13461 23100
rect 12216 23060 12222 23072
rect 13449 23069 13461 23072
rect 13495 23100 13507 23103
rect 13722 23100 13728 23112
rect 13495 23072 13728 23100
rect 13495 23069 13507 23072
rect 13449 23063 13507 23069
rect 13722 23060 13728 23072
rect 13780 23060 13786 23112
rect 16482 23100 16488 23112
rect 16443 23072 16488 23100
rect 16482 23060 16488 23072
rect 16540 23060 16546 23112
rect 19518 23100 19524 23112
rect 19479 23072 19524 23100
rect 19518 23060 19524 23072
rect 19576 23060 19582 23112
rect 20898 23060 20904 23112
rect 20956 23100 20962 23112
rect 21361 23103 21419 23109
rect 21361 23100 21373 23103
rect 20956 23072 21373 23100
rect 20956 23060 20962 23072
rect 21361 23069 21373 23072
rect 21407 23069 21419 23103
rect 21361 23063 21419 23069
rect 21450 23060 21456 23112
rect 21508 23100 21514 23112
rect 23014 23100 23020 23112
rect 21508 23072 21553 23100
rect 22975 23072 23020 23100
rect 21508 23060 21514 23072
rect 23014 23060 23020 23072
rect 23072 23060 23078 23112
rect 9030 23032 9036 23044
rect 8312 23004 9036 23032
rect 9030 22992 9036 23004
rect 9088 23032 9094 23044
rect 9677 23035 9735 23041
rect 9677 23032 9689 23035
rect 9088 23004 9689 23032
rect 9088 22992 9094 23004
rect 9677 23001 9689 23004
rect 9723 23001 9735 23035
rect 9677 22995 9735 23001
rect 15473 23035 15531 23041
rect 15473 23001 15485 23035
rect 15519 23032 15531 23035
rect 15930 23032 15936 23044
rect 15519 23004 15936 23032
rect 15519 23001 15531 23004
rect 15473 22995 15531 23001
rect 15930 22992 15936 23004
rect 15988 22992 15994 23044
rect 19242 22992 19248 23044
rect 19300 23032 19306 23044
rect 21818 23032 21824 23044
rect 19300 23004 21824 23032
rect 19300 22992 19306 23004
rect 21818 22992 21824 23004
rect 21876 22992 21882 23044
rect 3050 22964 3056 22976
rect 2884 22936 3056 22964
rect 3050 22924 3056 22936
rect 3108 22924 3114 22976
rect 3329 22967 3387 22973
rect 3329 22933 3341 22967
rect 3375 22964 3387 22967
rect 3418 22964 3424 22976
rect 3375 22936 3424 22964
rect 3375 22933 3387 22936
rect 3329 22927 3387 22933
rect 3418 22924 3424 22936
rect 3476 22924 3482 22976
rect 3881 22967 3939 22973
rect 3881 22933 3893 22967
rect 3927 22964 3939 22967
rect 4430 22964 4436 22976
rect 3927 22936 4436 22964
rect 3927 22933 3939 22936
rect 3881 22927 3939 22933
rect 4430 22924 4436 22936
rect 4488 22964 4494 22976
rect 6273 22967 6331 22973
rect 6273 22964 6285 22967
rect 4488 22936 6285 22964
rect 4488 22924 4494 22936
rect 6273 22933 6285 22936
rect 6319 22933 6331 22967
rect 6273 22927 6331 22933
rect 6917 22967 6975 22973
rect 6917 22933 6929 22967
rect 6963 22964 6975 22967
rect 7190 22964 7196 22976
rect 6963 22936 7196 22964
rect 6963 22933 6975 22936
rect 6917 22927 6975 22933
rect 7190 22924 7196 22936
rect 7248 22924 7254 22976
rect 10778 22924 10784 22976
rect 10836 22964 10842 22976
rect 12437 22967 12495 22973
rect 12437 22964 12449 22967
rect 10836 22936 12449 22964
rect 10836 22924 10842 22936
rect 12437 22933 12449 22936
rect 12483 22964 12495 22967
rect 12526 22964 12532 22976
rect 12483 22936 12532 22964
rect 12483 22933 12495 22936
rect 12437 22927 12495 22933
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 14458 22964 14464 22976
rect 14419 22936 14464 22964
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 16298 22964 16304 22976
rect 16259 22936 16304 22964
rect 16298 22924 16304 22936
rect 16356 22964 16362 22976
rect 17494 22964 17500 22976
rect 16356 22936 17500 22964
rect 16356 22924 16362 22936
rect 17494 22924 17500 22936
rect 17552 22964 17558 22976
rect 17865 22967 17923 22973
rect 17865 22964 17877 22967
rect 17552 22936 17877 22964
rect 17552 22924 17558 22936
rect 17865 22933 17877 22936
rect 17911 22964 17923 22967
rect 18417 22967 18475 22973
rect 18417 22964 18429 22967
rect 17911 22936 18429 22964
rect 17911 22933 17923 22936
rect 17865 22927 17923 22933
rect 18417 22933 18429 22936
rect 18463 22933 18475 22967
rect 18417 22927 18475 22933
rect 18874 22924 18880 22976
rect 18932 22964 18938 22976
rect 18969 22967 19027 22973
rect 18969 22964 18981 22967
rect 18932 22936 18981 22964
rect 18932 22924 18938 22936
rect 18969 22933 18981 22936
rect 19015 22933 19027 22967
rect 18969 22927 19027 22933
rect 20714 22924 20720 22976
rect 20772 22964 20778 22976
rect 20901 22967 20959 22973
rect 20901 22964 20913 22967
rect 20772 22936 20913 22964
rect 20772 22924 20778 22936
rect 20901 22933 20913 22936
rect 20947 22933 20959 22967
rect 20901 22927 20959 22933
rect 22094 22924 22100 22976
rect 22152 22964 22158 22976
rect 22281 22967 22339 22973
rect 22281 22964 22293 22967
rect 22152 22936 22293 22964
rect 22152 22924 22158 22936
rect 22281 22933 22293 22936
rect 22327 22933 22339 22967
rect 22281 22927 22339 22933
rect 22465 22967 22523 22973
rect 22465 22933 22477 22967
rect 22511 22964 22523 22967
rect 23474 22964 23480 22976
rect 22511 22936 23480 22964
rect 22511 22933 22523 22936
rect 22465 22927 22523 22933
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 1104 22874 26864 22896
rect 1104 22822 5648 22874
rect 5700 22822 5712 22874
rect 5764 22822 5776 22874
rect 5828 22822 5840 22874
rect 5892 22822 14982 22874
rect 15034 22822 15046 22874
rect 15098 22822 15110 22874
rect 15162 22822 15174 22874
rect 15226 22822 24315 22874
rect 24367 22822 24379 22874
rect 24431 22822 24443 22874
rect 24495 22822 24507 22874
rect 24559 22822 26864 22874
rect 1104 22800 26864 22822
rect 1486 22720 1492 22772
rect 1544 22760 1550 22772
rect 1854 22760 1860 22772
rect 1544 22732 1860 22760
rect 1544 22720 1550 22732
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 2590 22720 2596 22772
rect 2648 22760 2654 22772
rect 2685 22763 2743 22769
rect 2685 22760 2697 22763
rect 2648 22732 2697 22760
rect 2648 22720 2654 22732
rect 2685 22729 2697 22732
rect 2731 22729 2743 22763
rect 2685 22723 2743 22729
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 3694 22760 3700 22772
rect 2924 22732 3700 22760
rect 2924 22720 2930 22732
rect 3694 22720 3700 22732
rect 3752 22720 3758 22772
rect 5534 22720 5540 22772
rect 5592 22760 5598 22772
rect 6825 22763 6883 22769
rect 6825 22760 6837 22763
rect 5592 22732 6837 22760
rect 5592 22720 5598 22732
rect 6825 22729 6837 22732
rect 6871 22729 6883 22763
rect 6825 22723 6883 22729
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8389 22763 8447 22769
rect 8389 22760 8401 22763
rect 8352 22732 8401 22760
rect 8352 22720 8358 22732
rect 8389 22729 8401 22732
rect 8435 22729 8447 22763
rect 8389 22723 8447 22729
rect 1581 22695 1639 22701
rect 1581 22661 1593 22695
rect 1627 22692 1639 22695
rect 2774 22692 2780 22704
rect 1627 22664 2780 22692
rect 1627 22661 1639 22664
rect 1581 22655 1639 22661
rect 2774 22652 2780 22664
rect 2832 22652 2838 22704
rect 937 22627 995 22633
rect 937 22593 949 22627
rect 983 22624 995 22627
rect 1949 22627 2007 22633
rect 1949 22624 1961 22627
rect 983 22596 1961 22624
rect 983 22593 995 22596
rect 937 22587 995 22593
rect 1412 22565 1440 22596
rect 1949 22593 1961 22596
rect 1995 22593 2007 22627
rect 1949 22587 2007 22593
rect 2593 22627 2651 22633
rect 2593 22593 2605 22627
rect 2639 22624 2651 22627
rect 3329 22627 3387 22633
rect 3329 22624 3341 22627
rect 2639 22596 3341 22624
rect 2639 22593 2651 22596
rect 2593 22587 2651 22593
rect 3329 22593 3341 22596
rect 3375 22624 3387 22627
rect 3375 22596 4108 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 1397 22559 1455 22565
rect 1397 22525 1409 22559
rect 1443 22556 1455 22559
rect 1443 22528 1477 22556
rect 1443 22525 1455 22528
rect 1397 22519 1455 22525
rect 1670 22516 1676 22568
rect 1728 22556 1734 22568
rect 2314 22556 2320 22568
rect 1728 22528 2320 22556
rect 1728 22516 1734 22528
rect 2314 22516 2320 22528
rect 2372 22516 2378 22568
rect 3145 22559 3203 22565
rect 3145 22525 3157 22559
rect 3191 22556 3203 22559
rect 3510 22556 3516 22568
rect 3191 22528 3516 22556
rect 3191 22525 3203 22528
rect 3145 22519 3203 22525
rect 3510 22516 3516 22528
rect 3568 22516 3574 22568
rect 1854 22448 1860 22500
rect 1912 22488 1918 22500
rect 2222 22488 2228 22500
rect 1912 22460 2228 22488
rect 1912 22448 1918 22460
rect 2222 22448 2228 22460
rect 2280 22448 2286 22500
rect 3053 22423 3111 22429
rect 3053 22389 3065 22423
rect 3099 22420 3111 22423
rect 3142 22420 3148 22432
rect 3099 22392 3148 22420
rect 3099 22389 3111 22392
rect 3053 22383 3111 22389
rect 3142 22380 3148 22392
rect 3200 22380 3206 22432
rect 4080 22420 4108 22596
rect 5994 22584 6000 22636
rect 6052 22624 6058 22636
rect 6273 22627 6331 22633
rect 6273 22624 6285 22627
rect 6052 22596 6285 22624
rect 6052 22584 6058 22596
rect 6273 22593 6285 22596
rect 6319 22624 6331 22627
rect 7469 22627 7527 22633
rect 7469 22624 7481 22627
rect 6319 22596 7481 22624
rect 6319 22593 6331 22596
rect 6273 22587 6331 22593
rect 7469 22593 7481 22596
rect 7515 22624 7527 22627
rect 7558 22624 7564 22636
rect 7515 22596 7564 22624
rect 7515 22593 7527 22596
rect 7469 22587 7527 22593
rect 7558 22584 7564 22596
rect 7616 22584 7622 22636
rect 8404 22624 8432 22723
rect 9950 22720 9956 22772
rect 10008 22760 10014 22772
rect 10689 22763 10747 22769
rect 10689 22760 10701 22763
rect 10008 22732 10701 22760
rect 10008 22720 10014 22732
rect 10689 22729 10701 22732
rect 10735 22760 10747 22763
rect 11146 22760 11152 22772
rect 10735 22732 11152 22760
rect 10735 22729 10747 22732
rect 10689 22723 10747 22729
rect 11146 22720 11152 22732
rect 11204 22720 11210 22772
rect 11422 22760 11428 22772
rect 11383 22732 11428 22760
rect 11422 22720 11428 22732
rect 11480 22720 11486 22772
rect 12158 22760 12164 22772
rect 12119 22732 12164 22760
rect 12158 22720 12164 22732
rect 12216 22720 12222 22772
rect 12434 22720 12440 22772
rect 12492 22760 12498 22772
rect 12492 22732 12537 22760
rect 12492 22720 12498 22732
rect 13078 22720 13084 22772
rect 13136 22760 13142 22772
rect 13449 22763 13507 22769
rect 13449 22760 13461 22763
rect 13136 22732 13461 22760
rect 13136 22720 13142 22732
rect 13449 22729 13461 22732
rect 13495 22729 13507 22763
rect 13449 22723 13507 22729
rect 15562 22720 15568 22772
rect 15620 22760 15626 22772
rect 15749 22763 15807 22769
rect 15749 22760 15761 22763
rect 15620 22732 15761 22760
rect 15620 22720 15626 22732
rect 15749 22729 15761 22732
rect 15795 22729 15807 22763
rect 17034 22760 17040 22772
rect 16995 22732 17040 22760
rect 15749 22723 15807 22729
rect 17034 22720 17040 22732
rect 17092 22720 17098 22772
rect 18690 22760 18696 22772
rect 18651 22732 18696 22760
rect 18690 22720 18696 22732
rect 18748 22720 18754 22772
rect 22830 22760 22836 22772
rect 18800 22732 22416 22760
rect 22791 22732 22836 22760
rect 11054 22692 11060 22704
rect 11015 22664 11060 22692
rect 11054 22652 11060 22664
rect 11112 22652 11118 22704
rect 11238 22652 11244 22704
rect 11296 22692 11302 22704
rect 13906 22692 13912 22704
rect 11296 22664 13912 22692
rect 11296 22652 11302 22664
rect 13906 22652 13912 22664
rect 13964 22652 13970 22704
rect 17218 22652 17224 22704
rect 17276 22692 17282 22704
rect 18800 22692 18828 22732
rect 20898 22692 20904 22704
rect 17276 22664 18828 22692
rect 20859 22664 20904 22692
rect 17276 22652 17282 22664
rect 20898 22652 20904 22664
rect 20956 22652 20962 22704
rect 20990 22652 20996 22704
rect 21048 22692 21054 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 21048 22664 21189 22692
rect 21048 22652 21054 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 21177 22655 21235 22661
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 8404 22596 8585 22624
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 12158 22584 12164 22636
rect 12216 22624 12222 22636
rect 12894 22624 12900 22636
rect 12216 22596 12900 22624
rect 12216 22584 12222 22596
rect 12894 22584 12900 22596
rect 12952 22624 12958 22636
rect 12989 22627 13047 22633
rect 12989 22624 13001 22627
rect 12952 22596 13001 22624
rect 12952 22584 12958 22596
rect 12989 22593 13001 22596
rect 13035 22593 13047 22627
rect 12989 22587 13047 22593
rect 15562 22584 15568 22636
rect 15620 22624 15626 22636
rect 15746 22624 15752 22636
rect 15620 22596 15752 22624
rect 15620 22584 15626 22596
rect 15746 22584 15752 22596
rect 15804 22584 15810 22636
rect 18322 22584 18328 22636
rect 18380 22624 18386 22636
rect 18417 22627 18475 22633
rect 18417 22624 18429 22627
rect 18380 22596 18429 22624
rect 18380 22584 18386 22596
rect 18417 22593 18429 22596
rect 18463 22624 18475 22627
rect 18463 22596 19012 22624
rect 18463 22593 18475 22596
rect 18417 22587 18475 22593
rect 4157 22559 4215 22565
rect 4157 22525 4169 22559
rect 4203 22556 4215 22559
rect 4249 22559 4307 22565
rect 4249 22556 4261 22559
rect 4203 22528 4261 22556
rect 4203 22525 4215 22528
rect 4157 22519 4215 22525
rect 4249 22525 4261 22528
rect 4295 22556 4307 22559
rect 5442 22556 5448 22568
rect 4295 22528 5448 22556
rect 4295 22525 4307 22528
rect 4249 22519 4307 22525
rect 5442 22516 5448 22528
rect 5500 22516 5506 22568
rect 11238 22556 11244 22568
rect 11199 22528 11244 22556
rect 11238 22516 11244 22528
rect 11296 22516 11302 22568
rect 12710 22516 12716 22568
rect 12768 22556 12774 22568
rect 12805 22559 12863 22565
rect 12805 22556 12817 22559
rect 12768 22528 12817 22556
rect 12768 22516 12774 22528
rect 12805 22525 12817 22528
rect 12851 22525 12863 22559
rect 12805 22519 12863 22525
rect 13354 22516 13360 22568
rect 13412 22556 13418 22568
rect 14185 22559 14243 22565
rect 14185 22556 14197 22559
rect 13412 22528 14197 22556
rect 13412 22516 13418 22528
rect 14185 22525 14197 22528
rect 14231 22556 14243 22559
rect 14369 22559 14427 22565
rect 14369 22556 14381 22559
rect 14231 22528 14381 22556
rect 14231 22525 14243 22528
rect 14185 22519 14243 22525
rect 14369 22525 14381 22528
rect 14415 22525 14427 22559
rect 14369 22519 14427 22525
rect 14458 22516 14464 22568
rect 14516 22556 14522 22568
rect 14642 22565 14648 22568
rect 14625 22559 14648 22565
rect 14625 22556 14637 22559
rect 14516 22528 14637 22556
rect 14516 22516 14522 22528
rect 14625 22525 14637 22528
rect 14700 22556 14706 22568
rect 16850 22556 16856 22568
rect 14700 22528 14773 22556
rect 16811 22528 16856 22556
rect 14625 22519 14648 22525
rect 14642 22516 14648 22519
rect 14700 22516 14706 22528
rect 16850 22516 16856 22528
rect 16908 22556 16914 22568
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 16908 22528 17417 22556
rect 16908 22516 16914 22528
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 18690 22516 18696 22568
rect 18748 22556 18754 22568
rect 18877 22559 18935 22565
rect 18877 22556 18889 22559
rect 18748 22528 18889 22556
rect 18748 22516 18754 22528
rect 18877 22525 18889 22528
rect 18923 22525 18935 22559
rect 18984 22556 19012 22596
rect 19150 22565 19156 22568
rect 19144 22556 19156 22565
rect 18984 22528 19156 22556
rect 18877 22519 18935 22525
rect 19144 22519 19156 22528
rect 19208 22556 19214 22568
rect 19518 22556 19524 22568
rect 19208 22528 19524 22556
rect 4430 22448 4436 22500
rect 4488 22497 4494 22500
rect 4488 22491 4552 22497
rect 4488 22457 4506 22491
rect 4540 22457 4552 22491
rect 4488 22451 4552 22457
rect 6641 22491 6699 22497
rect 6641 22457 6653 22491
rect 6687 22488 6699 22491
rect 6730 22488 6736 22500
rect 6687 22460 6736 22488
rect 6687 22457 6699 22460
rect 6641 22451 6699 22457
rect 4488 22448 4494 22451
rect 6730 22448 6736 22460
rect 6788 22488 6794 22500
rect 7285 22491 7343 22497
rect 7285 22488 7297 22491
rect 6788 22460 7297 22488
rect 6788 22448 6794 22460
rect 7285 22457 7297 22460
rect 7331 22457 7343 22491
rect 8110 22488 8116 22500
rect 8023 22460 8116 22488
rect 7285 22451 7343 22457
rect 8110 22448 8116 22460
rect 8168 22488 8174 22500
rect 8846 22497 8852 22500
rect 8840 22488 8852 22497
rect 8168 22460 8852 22488
rect 8168 22448 8174 22460
rect 8840 22451 8852 22460
rect 8846 22448 8852 22451
rect 8904 22448 8910 22500
rect 12897 22491 12955 22497
rect 12897 22457 12909 22491
rect 12943 22488 12955 22491
rect 12986 22488 12992 22500
rect 12943 22460 12992 22488
rect 12943 22457 12955 22460
rect 12897 22451 12955 22457
rect 12986 22448 12992 22460
rect 13044 22488 13050 22500
rect 13817 22491 13875 22497
rect 13817 22488 13829 22491
rect 13044 22460 13829 22488
rect 13044 22448 13050 22460
rect 13817 22457 13829 22460
rect 13863 22457 13875 22491
rect 18892 22488 18920 22519
rect 19150 22516 19156 22519
rect 19208 22516 19214 22528
rect 19518 22516 19524 22528
rect 19576 22516 19582 22568
rect 19978 22516 19984 22568
rect 20036 22556 20042 22568
rect 20898 22556 20904 22568
rect 20036 22528 20904 22556
rect 20036 22516 20042 22528
rect 20898 22516 20904 22528
rect 20956 22516 20962 22568
rect 19058 22488 19064 22500
rect 18892 22460 19064 22488
rect 13817 22451 13875 22457
rect 19058 22448 19064 22460
rect 19116 22448 19122 22500
rect 21192 22488 21220 22655
rect 21450 22584 21456 22636
rect 21508 22624 21514 22636
rect 21913 22627 21971 22633
rect 21913 22624 21925 22627
rect 21508 22596 21925 22624
rect 21508 22584 21514 22596
rect 21913 22593 21925 22596
rect 21959 22593 21971 22627
rect 21913 22587 21971 22593
rect 21726 22516 21732 22568
rect 21784 22556 21790 22568
rect 21821 22559 21879 22565
rect 21821 22556 21833 22559
rect 21784 22528 21833 22556
rect 21784 22516 21790 22528
rect 21821 22525 21833 22528
rect 21867 22556 21879 22559
rect 22002 22556 22008 22568
rect 21867 22528 22008 22556
rect 21867 22525 21879 22528
rect 21821 22519 21879 22525
rect 22002 22516 22008 22528
rect 22060 22516 22066 22568
rect 22388 22556 22416 22732
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 23845 22763 23903 22769
rect 23845 22729 23857 22763
rect 23891 22760 23903 22763
rect 24118 22760 24124 22772
rect 23891 22732 24124 22760
rect 23891 22729 23903 22732
rect 23845 22723 23903 22729
rect 24118 22720 24124 22732
rect 24176 22720 24182 22772
rect 22554 22624 22560 22636
rect 22467 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22624 22618 22636
rect 22738 22624 22744 22636
rect 22612 22596 22744 22624
rect 22612 22584 22618 22596
rect 22738 22584 22744 22596
rect 22796 22584 22802 22636
rect 23842 22624 23848 22636
rect 23492 22596 23848 22624
rect 23492 22556 23520 22596
rect 23842 22584 23848 22596
rect 23900 22624 23906 22636
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 23900 22596 24593 22624
rect 23900 22584 23906 22596
rect 24581 22593 24593 22596
rect 24627 22624 24639 22627
rect 24670 22624 24676 22636
rect 24627 22596 24676 22624
rect 24627 22593 24639 22596
rect 24581 22587 24639 22593
rect 24670 22584 24676 22596
rect 24728 22584 24734 22636
rect 23658 22556 23664 22568
rect 22388 22528 23520 22556
rect 23619 22528 23664 22556
rect 23658 22516 23664 22528
rect 23716 22556 23722 22568
rect 24213 22559 24271 22565
rect 24213 22556 24225 22559
rect 23716 22528 24225 22556
rect 23716 22516 23722 22528
rect 24213 22525 24225 22528
rect 24259 22525 24271 22559
rect 24213 22519 24271 22525
rect 24765 22559 24823 22565
rect 24765 22525 24777 22559
rect 24811 22525 24823 22559
rect 24765 22519 24823 22525
rect 21192 22460 21772 22488
rect 5629 22423 5687 22429
rect 5629 22420 5641 22423
rect 4080 22392 5641 22420
rect 5629 22389 5641 22392
rect 5675 22420 5687 22423
rect 5994 22420 6000 22432
rect 5675 22392 6000 22420
rect 5675 22389 5687 22392
rect 5629 22383 5687 22389
rect 5994 22380 6000 22392
rect 6052 22380 6058 22432
rect 7190 22420 7196 22432
rect 7151 22392 7196 22420
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 9950 22420 9956 22432
rect 9911 22392 9956 22420
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 11790 22420 11796 22432
rect 11751 22392 11796 22420
rect 11790 22380 11796 22392
rect 11848 22380 11854 22432
rect 11974 22380 11980 22432
rect 12032 22420 12038 22432
rect 13078 22420 13084 22432
rect 12032 22392 13084 22420
rect 12032 22380 12038 22392
rect 13078 22380 13084 22392
rect 13136 22380 13142 22432
rect 13262 22380 13268 22432
rect 13320 22420 13326 22432
rect 13446 22420 13452 22432
rect 13320 22392 13452 22420
rect 13320 22380 13326 22392
rect 13446 22380 13452 22392
rect 13504 22380 13510 22432
rect 15286 22380 15292 22432
rect 15344 22420 15350 22432
rect 16482 22420 16488 22432
rect 15344 22392 16488 22420
rect 15344 22380 15350 22392
rect 16482 22380 16488 22392
rect 16540 22380 16546 22432
rect 17770 22420 17776 22432
rect 17731 22392 17776 22420
rect 17770 22380 17776 22392
rect 17828 22380 17834 22432
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 20257 22423 20315 22429
rect 20257 22420 20269 22423
rect 19392 22392 20269 22420
rect 19392 22380 19398 22392
rect 20257 22389 20269 22392
rect 20303 22389 20315 22423
rect 21358 22420 21364 22432
rect 21319 22392 21364 22420
rect 20257 22383 20315 22389
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 21744 22429 21772 22460
rect 23750 22448 23756 22500
rect 23808 22488 23814 22500
rect 24780 22488 24808 22519
rect 25225 22491 25283 22497
rect 25225 22488 25237 22491
rect 23808 22460 25237 22488
rect 23808 22448 23814 22460
rect 25225 22457 25237 22460
rect 25271 22457 25283 22491
rect 25225 22451 25283 22457
rect 21729 22423 21787 22429
rect 21729 22389 21741 22423
rect 21775 22389 21787 22423
rect 21729 22383 21787 22389
rect 23014 22380 23020 22432
rect 23072 22420 23078 22432
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 23072 22392 23213 22420
rect 23072 22380 23078 22392
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 24946 22420 24952 22432
rect 24907 22392 24952 22420
rect 23201 22383 23259 22389
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 1104 22330 26864 22352
rect 1104 22278 10315 22330
rect 10367 22278 10379 22330
rect 10431 22278 10443 22330
rect 10495 22278 10507 22330
rect 10559 22278 19648 22330
rect 19700 22278 19712 22330
rect 19764 22278 19776 22330
rect 19828 22278 19840 22330
rect 19892 22278 26864 22330
rect 1104 22256 26864 22278
rect 1949 22219 2007 22225
rect 1949 22185 1961 22219
rect 1995 22216 2007 22219
rect 2038 22216 2044 22228
rect 1995 22188 2044 22216
rect 1995 22185 2007 22188
rect 1949 22179 2007 22185
rect 2038 22176 2044 22188
rect 2096 22176 2102 22228
rect 5721 22219 5779 22225
rect 5721 22185 5733 22219
rect 5767 22216 5779 22219
rect 5902 22216 5908 22228
rect 5767 22188 5908 22216
rect 5767 22185 5779 22188
rect 5721 22179 5779 22185
rect 5902 22176 5908 22188
rect 5960 22176 5966 22228
rect 6457 22219 6515 22225
rect 6457 22185 6469 22219
rect 6503 22216 6515 22219
rect 6638 22216 6644 22228
rect 6503 22188 6644 22216
rect 6503 22185 6515 22188
rect 6457 22179 6515 22185
rect 6638 22176 6644 22188
rect 6696 22176 6702 22228
rect 9306 22176 9312 22228
rect 9364 22216 9370 22228
rect 9401 22219 9459 22225
rect 9401 22216 9413 22219
rect 9364 22188 9413 22216
rect 9364 22176 9370 22188
rect 9401 22185 9413 22188
rect 9447 22185 9459 22219
rect 10134 22216 10140 22228
rect 9401 22179 9459 22185
rect 9692 22188 10140 22216
rect 2406 22108 2412 22160
rect 2464 22108 2470 22160
rect 4062 22108 4068 22160
rect 4120 22148 4126 22160
rect 4617 22151 4675 22157
rect 4617 22148 4629 22151
rect 4120 22120 4629 22148
rect 4120 22108 4126 22120
rect 4617 22117 4629 22120
rect 4663 22117 4675 22151
rect 4617 22111 4675 22117
rect 6825 22151 6883 22157
rect 6825 22117 6837 22151
rect 6871 22148 6883 22151
rect 7098 22148 7104 22160
rect 6871 22120 7104 22148
rect 6871 22117 6883 22120
rect 6825 22111 6883 22117
rect 7098 22108 7104 22120
rect 7156 22108 7162 22160
rect 8294 22108 8300 22160
rect 8352 22108 8358 22160
rect 8389 22151 8447 22157
rect 8389 22117 8401 22151
rect 8435 22148 8447 22151
rect 8570 22148 8576 22160
rect 8435 22120 8576 22148
rect 8435 22117 8447 22120
rect 8389 22111 8447 22117
rect 8570 22108 8576 22120
rect 8628 22108 8634 22160
rect 9692 22148 9720 22188
rect 10134 22176 10140 22188
rect 10192 22176 10198 22228
rect 10321 22219 10379 22225
rect 10321 22185 10333 22219
rect 10367 22216 10379 22219
rect 10686 22216 10692 22228
rect 10367 22188 10692 22216
rect 10367 22185 10379 22188
rect 10321 22179 10379 22185
rect 10686 22176 10692 22188
rect 10744 22216 10750 22228
rect 12250 22216 12256 22228
rect 10744 22188 12256 22216
rect 10744 22176 10750 22188
rect 12250 22176 12256 22188
rect 12308 22176 12314 22228
rect 12345 22219 12403 22225
rect 12345 22185 12357 22219
rect 12391 22216 12403 22219
rect 12434 22216 12440 22228
rect 12391 22188 12440 22216
rect 12391 22185 12403 22188
rect 12345 22179 12403 22185
rect 12434 22176 12440 22188
rect 12492 22216 12498 22228
rect 12618 22216 12624 22228
rect 12492 22188 12624 22216
rect 12492 22176 12498 22188
rect 12618 22176 12624 22188
rect 12676 22176 12682 22228
rect 12710 22176 12716 22228
rect 12768 22176 12774 22228
rect 12894 22216 12900 22228
rect 12855 22188 12900 22216
rect 12894 22176 12900 22188
rect 12952 22176 12958 22228
rect 13449 22219 13507 22225
rect 13449 22185 13461 22219
rect 13495 22216 13507 22219
rect 13538 22216 13544 22228
rect 13495 22188 13544 22216
rect 13495 22185 13507 22188
rect 13449 22179 13507 22185
rect 13538 22176 13544 22188
rect 13596 22176 13602 22228
rect 17770 22216 17776 22228
rect 13832 22188 17172 22216
rect 17731 22188 17776 22216
rect 9600 22120 9720 22148
rect 1857 22083 1915 22089
rect 1857 22049 1869 22083
rect 1903 22080 1915 22083
rect 2314 22080 2320 22092
rect 1903 22052 2320 22080
rect 1903 22049 1915 22052
rect 1857 22043 1915 22049
rect 2314 22040 2320 22052
rect 2372 22040 2378 22092
rect 2424 22080 2452 22108
rect 2424 22052 2636 22080
rect 2608 22024 2636 22052
rect 4080 22024 4108 22108
rect 4154 22040 4160 22092
rect 4212 22080 4218 22092
rect 4709 22083 4767 22089
rect 4709 22080 4721 22083
rect 4212 22052 4721 22080
rect 4212 22040 4218 22052
rect 4709 22049 4721 22052
rect 4755 22080 4767 22083
rect 5074 22080 5080 22092
rect 4755 22052 5080 22080
rect 4755 22049 4767 22052
rect 4709 22043 4767 22049
rect 5074 22040 5080 22052
rect 5132 22040 5138 22092
rect 6362 22080 6368 22092
rect 6323 22052 6368 22080
rect 6362 22040 6368 22052
rect 6420 22040 6426 22092
rect 6730 22040 6736 22092
rect 6788 22080 6794 22092
rect 7006 22080 7012 22092
rect 6788 22052 7012 22080
rect 6788 22040 6794 22052
rect 7006 22040 7012 22052
rect 7064 22040 7070 22092
rect 7558 22040 7564 22092
rect 7616 22080 7622 22092
rect 8312 22080 8340 22108
rect 7616 22052 8340 22080
rect 9125 22083 9183 22089
rect 7616 22040 7622 22052
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 9600 22080 9628 22120
rect 9950 22108 9956 22160
rect 10008 22148 10014 22160
rect 12728 22148 12756 22176
rect 13832 22160 13860 22188
rect 13814 22148 13820 22160
rect 10008 22120 11008 22148
rect 12728 22120 13676 22148
rect 13775 22120 13820 22148
rect 10008 22108 10014 22120
rect 9171 22052 9628 22080
rect 9677 22083 9735 22089
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 9677 22049 9689 22083
rect 9723 22080 9735 22083
rect 9766 22080 9772 22092
rect 9723 22052 9772 22080
rect 9723 22049 9735 22052
rect 9677 22043 9735 22049
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 9858 22040 9864 22092
rect 9916 22040 9922 22092
rect 10980 22080 11008 22120
rect 11232 22083 11290 22089
rect 11232 22080 11244 22083
rect 10980 22052 11244 22080
rect 11232 22049 11244 22052
rect 11278 22080 11290 22083
rect 11514 22080 11520 22092
rect 11278 22052 11520 22080
rect 11278 22049 11290 22052
rect 11232 22043 11290 22049
rect 11514 22040 11520 22052
rect 11572 22040 11578 22092
rect 13648 22080 13676 22120
rect 13814 22108 13820 22120
rect 13872 22108 13878 22160
rect 13909 22151 13967 22157
rect 13909 22117 13921 22151
rect 13955 22148 13967 22151
rect 14550 22148 14556 22160
rect 13955 22120 14556 22148
rect 13955 22117 13967 22120
rect 13909 22111 13967 22117
rect 14550 22108 14556 22120
rect 14608 22148 14614 22160
rect 15746 22148 15752 22160
rect 14608 22120 15752 22148
rect 14608 22108 14614 22120
rect 15746 22108 15752 22120
rect 15804 22108 15810 22160
rect 17144 22148 17172 22188
rect 17770 22176 17776 22188
rect 17828 22176 17834 22228
rect 19061 22219 19119 22225
rect 19061 22185 19073 22219
rect 19107 22216 19119 22219
rect 19150 22216 19156 22228
rect 19107 22188 19156 22216
rect 19107 22185 19119 22188
rect 19061 22179 19119 22185
rect 19150 22176 19156 22188
rect 19208 22176 19214 22228
rect 20717 22219 20775 22225
rect 20717 22185 20729 22219
rect 20763 22216 20775 22219
rect 21450 22216 21456 22228
rect 20763 22188 21456 22216
rect 20763 22185 20775 22188
rect 20717 22179 20775 22185
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 22833 22219 22891 22225
rect 22833 22216 22845 22219
rect 21652 22188 22845 22216
rect 19610 22148 19616 22160
rect 17144 22120 19616 22148
rect 19610 22108 19616 22120
rect 19668 22148 19674 22160
rect 20070 22148 20076 22160
rect 19668 22120 20076 22148
rect 19668 22108 19674 22120
rect 20070 22108 20076 22120
rect 20128 22108 20134 22160
rect 14461 22083 14519 22089
rect 14461 22080 14473 22083
rect 13648 22052 14473 22080
rect 14461 22049 14473 22052
rect 14507 22049 14519 22083
rect 14461 22043 14519 22049
rect 15556 22083 15614 22089
rect 15556 22049 15568 22083
rect 15602 22080 15614 22083
rect 15930 22080 15936 22092
rect 15602 22052 15936 22080
rect 15602 22049 15614 22052
rect 15556 22043 15614 22049
rect 15930 22040 15936 22052
rect 15988 22040 15994 22092
rect 16942 22040 16948 22092
rect 17000 22080 17006 22092
rect 17221 22083 17279 22089
rect 17221 22080 17233 22083
rect 17000 22052 17233 22080
rect 17000 22040 17006 22052
rect 17221 22049 17233 22052
rect 17267 22049 17279 22083
rect 18138 22080 18144 22092
rect 18099 22052 18144 22080
rect 17221 22043 17279 22049
rect 18138 22040 18144 22052
rect 18196 22040 18202 22092
rect 19337 22083 19395 22089
rect 19337 22049 19349 22083
rect 19383 22080 19395 22083
rect 19518 22080 19524 22092
rect 19383 22052 19524 22080
rect 19383 22049 19395 22052
rect 19337 22043 19395 22049
rect 19518 22040 19524 22052
rect 19576 22040 19582 22092
rect 20346 22040 20352 22092
rect 20404 22080 20410 22092
rect 21652 22089 21680 22188
rect 22833 22185 22845 22188
rect 22879 22185 22891 22219
rect 23198 22216 23204 22228
rect 23159 22188 23204 22216
rect 22833 22179 22891 22185
rect 23198 22176 23204 22188
rect 23256 22176 23262 22228
rect 24397 22151 24455 22157
rect 24397 22117 24409 22151
rect 24443 22148 24455 22151
rect 24670 22148 24676 22160
rect 24443 22120 24676 22148
rect 24443 22117 24455 22120
rect 24397 22111 24455 22117
rect 24670 22108 24676 22120
rect 24728 22108 24734 22160
rect 21637 22083 21695 22089
rect 21637 22080 21649 22083
rect 20404 22052 21649 22080
rect 20404 22040 20410 22052
rect 21637 22049 21649 22052
rect 21683 22049 21695 22083
rect 21637 22043 21695 22049
rect 22186 22040 22192 22092
rect 22244 22080 22250 22092
rect 22741 22083 22799 22089
rect 22741 22080 22753 22083
rect 22244 22052 22753 22080
rect 22244 22040 22250 22052
rect 22741 22049 22753 22052
rect 22787 22080 22799 22083
rect 23934 22080 23940 22092
rect 22787 22052 23428 22080
rect 23895 22052 23940 22080
rect 22787 22049 22799 22052
rect 22741 22043 22799 22049
rect 2406 22012 2412 22024
rect 2367 21984 2412 22012
rect 2406 21972 2412 21984
rect 2464 21972 2470 22024
rect 2590 21972 2596 22024
rect 2648 22012 2654 22024
rect 2648 21984 2741 22012
rect 2648 21972 2654 21984
rect 4062 21972 4068 22024
rect 4120 21972 4126 22024
rect 4614 21972 4620 22024
rect 4672 22012 4678 22024
rect 4801 22015 4859 22021
rect 4801 22012 4813 22015
rect 4672 21984 4813 22012
rect 4672 21972 4678 21984
rect 4801 21981 4813 21984
rect 4847 21981 4859 22015
rect 4801 21975 4859 21981
rect 6546 21972 6552 22024
rect 6604 22012 6610 22024
rect 6917 22015 6975 22021
rect 6917 22012 6929 22015
rect 6604 21984 6929 22012
rect 6604 21972 6610 21984
rect 6917 21981 6929 21984
rect 6963 21981 6975 22015
rect 6917 21975 6975 21981
rect 7101 22015 7159 22021
rect 7101 21981 7113 22015
rect 7147 22012 7159 22015
rect 8478 22012 8484 22024
rect 7147 21984 8340 22012
rect 8439 21984 8484 22012
rect 7147 21981 7159 21984
rect 7101 21975 7159 21981
rect 8312 21956 8340 21984
rect 8478 21972 8484 21984
rect 8536 21972 8542 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 3050 21944 3056 21956
rect 2963 21916 3056 21944
rect 3050 21904 3056 21916
rect 3108 21944 3114 21956
rect 5353 21947 5411 21953
rect 3108 21916 5203 21944
rect 3108 21904 3114 21916
rect 1210 21836 1216 21888
rect 1268 21876 1274 21888
rect 2314 21876 2320 21888
rect 1268 21848 2320 21876
rect 1268 21836 1274 21848
rect 2314 21836 2320 21848
rect 2372 21836 2378 21888
rect 3602 21876 3608 21888
rect 3563 21848 3608 21876
rect 3602 21836 3608 21848
rect 3660 21836 3666 21888
rect 3878 21836 3884 21888
rect 3936 21876 3942 21888
rect 4249 21879 4307 21885
rect 4249 21876 4261 21879
rect 3936 21848 4261 21876
rect 3936 21836 3942 21848
rect 4249 21845 4261 21848
rect 4295 21845 4307 21879
rect 5175 21876 5203 21916
rect 5353 21913 5365 21947
rect 5399 21944 5411 21947
rect 5442 21944 5448 21956
rect 5399 21916 5448 21944
rect 5399 21913 5411 21916
rect 5353 21907 5411 21913
rect 5442 21904 5448 21916
rect 5500 21944 5506 21956
rect 8021 21947 8079 21953
rect 5500 21916 7604 21944
rect 5500 21904 5506 21916
rect 7576 21888 7604 21916
rect 8021 21913 8033 21947
rect 8067 21944 8079 21947
rect 8202 21944 8208 21956
rect 8067 21916 8208 21944
rect 8067 21913 8079 21916
rect 8021 21907 8079 21913
rect 8202 21904 8208 21916
rect 8260 21904 8266 21956
rect 8294 21904 8300 21956
rect 8352 21944 8358 21956
rect 8588 21944 8616 21975
rect 9582 21972 9588 22024
rect 9640 22012 9646 22024
rect 9876 22012 9904 22040
rect 9640 21984 9904 22012
rect 9640 21972 9646 21984
rect 10778 21972 10784 22024
rect 10836 22012 10842 22024
rect 10962 22012 10968 22024
rect 10836 21984 10968 22012
rect 10836 21972 10842 21984
rect 10962 21972 10968 21984
rect 11020 21972 11026 22024
rect 13998 22012 14004 22024
rect 13959 21984 14004 22012
rect 13998 21972 14004 21984
rect 14056 21972 14062 22024
rect 15286 22012 15292 22024
rect 15247 21984 15292 22012
rect 15286 21972 15292 21984
rect 15344 21972 15350 22024
rect 17494 21972 17500 22024
rect 17552 22012 17558 22024
rect 18233 22015 18291 22021
rect 18233 22012 18245 22015
rect 17552 21984 18245 22012
rect 17552 21972 17558 21984
rect 18233 21981 18245 21984
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 20530 22012 20536 22024
rect 18380 21984 18425 22012
rect 19536 21984 20536 22012
rect 18380 21972 18386 21984
rect 8352 21916 8616 21944
rect 8352 21904 8358 21916
rect 9674 21904 9680 21956
rect 9732 21944 9738 21956
rect 9861 21947 9919 21953
rect 9861 21944 9873 21947
rect 9732 21916 9873 21944
rect 9732 21904 9738 21916
rect 9861 21913 9873 21916
rect 9907 21913 9919 21947
rect 16666 21944 16672 21956
rect 16627 21916 16672 21944
rect 9861 21907 9919 21913
rect 16666 21904 16672 21916
rect 16724 21904 16730 21956
rect 17681 21947 17739 21953
rect 17681 21913 17693 21947
rect 17727 21944 17739 21947
rect 18874 21944 18880 21956
rect 17727 21916 18880 21944
rect 17727 21913 17739 21916
rect 17681 21907 17739 21913
rect 18874 21904 18880 21916
rect 18932 21904 18938 21956
rect 19536 21953 19564 21984
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 21729 22015 21787 22021
rect 21729 22012 21741 22015
rect 20772 21984 21741 22012
rect 20772 21972 20778 21984
rect 21729 21981 21741 21984
rect 21775 21981 21787 22015
rect 21729 21975 21787 21981
rect 21818 21972 21824 22024
rect 21876 22012 21882 22024
rect 23290 22012 23296 22024
rect 21876 21984 21921 22012
rect 23251 21984 23296 22012
rect 21876 21972 21882 21984
rect 23290 21972 23296 21984
rect 23348 21972 23354 22024
rect 23400 22021 23428 22052
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 25314 22040 25320 22092
rect 25372 22080 25378 22092
rect 25409 22083 25467 22089
rect 25409 22080 25421 22083
rect 25372 22052 25421 22080
rect 25372 22040 25378 22052
rect 25409 22049 25421 22052
rect 25455 22049 25467 22083
rect 25409 22043 25467 22049
rect 23385 22015 23443 22021
rect 23385 21981 23397 22015
rect 23431 21981 23443 22015
rect 23385 21975 23443 21981
rect 19521 21947 19579 21953
rect 19521 21913 19533 21947
rect 19567 21913 19579 21947
rect 19521 21907 19579 21913
rect 20349 21947 20407 21953
rect 20349 21913 20361 21947
rect 20395 21944 20407 21947
rect 21266 21944 21272 21956
rect 20395 21916 21272 21944
rect 20395 21913 20407 21916
rect 20349 21907 20407 21913
rect 21266 21904 21272 21916
rect 21324 21904 21330 21956
rect 22462 21904 22468 21956
rect 22520 21944 22526 21956
rect 25774 21944 25780 21956
rect 22520 21916 25780 21944
rect 22520 21904 22526 21916
rect 25774 21904 25780 21916
rect 25832 21904 25838 21956
rect 6822 21876 6828 21888
rect 5175 21848 6828 21876
rect 4249 21839 4307 21845
rect 6822 21836 6828 21848
rect 6880 21836 6886 21888
rect 7558 21836 7564 21888
rect 7616 21876 7622 21888
rect 7653 21879 7711 21885
rect 7653 21876 7665 21879
rect 7616 21848 7665 21876
rect 7616 21836 7622 21848
rect 7653 21845 7665 21848
rect 7699 21845 7711 21879
rect 7653 21839 7711 21845
rect 9490 21836 9496 21888
rect 9548 21876 9554 21888
rect 10689 21879 10747 21885
rect 10689 21876 10701 21879
rect 9548 21848 10701 21876
rect 9548 21836 9554 21848
rect 10689 21845 10701 21848
rect 10735 21876 10747 21879
rect 10778 21876 10784 21888
rect 10735 21848 10784 21876
rect 10735 21845 10747 21848
rect 10689 21839 10747 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 13354 21876 13360 21888
rect 13315 21848 13360 21876
rect 13354 21836 13360 21848
rect 13412 21836 13418 21888
rect 14826 21876 14832 21888
rect 14787 21848 14832 21876
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 19981 21879 20039 21885
rect 19981 21845 19993 21879
rect 20027 21876 20039 21879
rect 20530 21876 20536 21888
rect 20027 21848 20536 21876
rect 20027 21845 20039 21848
rect 19981 21839 20039 21845
rect 20530 21836 20536 21848
rect 20588 21836 20594 21888
rect 21082 21876 21088 21888
rect 21043 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21876 21146 21888
rect 21634 21876 21640 21888
rect 21140 21848 21640 21876
rect 21140 21836 21146 21848
rect 21634 21836 21640 21848
rect 21692 21836 21698 21888
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 25593 21879 25651 21885
rect 25593 21845 25605 21879
rect 25639 21876 25651 21879
rect 26142 21876 26148 21888
rect 25639 21848 26148 21876
rect 25639 21845 25651 21848
rect 25593 21839 25651 21845
rect 26142 21836 26148 21848
rect 26200 21836 26206 21888
rect 1104 21786 26864 21808
rect 1104 21734 5648 21786
rect 5700 21734 5712 21786
rect 5764 21734 5776 21786
rect 5828 21734 5840 21786
rect 5892 21734 14982 21786
rect 15034 21734 15046 21786
rect 15098 21734 15110 21786
rect 15162 21734 15174 21786
rect 15226 21734 24315 21786
rect 24367 21734 24379 21786
rect 24431 21734 24443 21786
rect 24495 21734 24507 21786
rect 24559 21734 26864 21786
rect 1104 21712 26864 21734
rect 1302 21632 1308 21684
rect 1360 21672 1366 21684
rect 1765 21675 1823 21681
rect 1765 21672 1777 21675
rect 1360 21644 1777 21672
rect 1360 21632 1366 21644
rect 1765 21641 1777 21644
rect 1811 21641 1823 21675
rect 1765 21635 1823 21641
rect 1949 21675 2007 21681
rect 1949 21641 1961 21675
rect 1995 21672 2007 21675
rect 2498 21672 2504 21684
rect 1995 21644 2504 21672
rect 1995 21641 2007 21644
rect 1949 21635 2007 21641
rect 1780 21536 1808 21635
rect 2498 21632 2504 21644
rect 2556 21632 2562 21684
rect 3510 21672 3516 21684
rect 3471 21644 3516 21672
rect 3510 21632 3516 21644
rect 3568 21632 3574 21684
rect 5074 21672 5080 21684
rect 5035 21644 5080 21672
rect 5074 21632 5080 21644
rect 5132 21632 5138 21684
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 5408 21644 5580 21672
rect 5408 21632 5414 21644
rect 3329 21607 3387 21613
rect 3329 21604 3341 21607
rect 2424 21576 3341 21604
rect 2424 21545 2452 21576
rect 3329 21573 3341 21576
rect 3375 21604 3387 21607
rect 4893 21607 4951 21613
rect 4893 21604 4905 21607
rect 3375 21576 4905 21604
rect 3375 21573 3387 21576
rect 3329 21567 3387 21573
rect 2409 21539 2467 21545
rect 2409 21536 2421 21539
rect 1780 21508 2421 21536
rect 2409 21505 2421 21508
rect 2455 21505 2467 21539
rect 2590 21536 2596 21548
rect 2551 21508 2596 21536
rect 2409 21499 2467 21505
rect 2590 21496 2596 21508
rect 2648 21496 2654 21548
rect 3988 21545 4016 21576
rect 4893 21573 4905 21576
rect 4939 21604 4951 21607
rect 4939 21576 5488 21604
rect 4939 21573 4951 21576
rect 4893 21567 4951 21573
rect 3973 21539 4031 21545
rect 3973 21505 3985 21539
rect 4019 21505 4031 21539
rect 3973 21499 4031 21505
rect 4065 21539 4123 21545
rect 4065 21505 4077 21539
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 750 21428 756 21480
rect 808 21468 814 21480
rect 2317 21471 2375 21477
rect 2317 21468 2329 21471
rect 808 21440 2329 21468
rect 808 21428 814 21440
rect 2317 21437 2329 21440
rect 2363 21468 2375 21471
rect 2961 21471 3019 21477
rect 2961 21468 2973 21471
rect 2363 21440 2973 21468
rect 2363 21437 2375 21440
rect 2317 21431 2375 21437
rect 2961 21437 2973 21440
rect 3007 21468 3019 21471
rect 3510 21468 3516 21480
rect 3007 21440 3516 21468
rect 3007 21437 3019 21440
rect 2961 21431 3019 21437
rect 3510 21428 3516 21440
rect 3568 21428 3574 21480
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 4080 21468 4108 21499
rect 5460 21477 5488 21576
rect 5552 21536 5580 21644
rect 6546 21632 6552 21684
rect 6604 21672 6610 21684
rect 6641 21675 6699 21681
rect 6641 21672 6653 21675
rect 6604 21644 6653 21672
rect 6604 21632 6610 21644
rect 6641 21641 6653 21644
rect 6687 21641 6699 21675
rect 6641 21635 6699 21641
rect 7561 21675 7619 21681
rect 7561 21641 7573 21675
rect 7607 21672 7619 21675
rect 7650 21672 7656 21684
rect 7607 21644 7656 21672
rect 7607 21641 7619 21644
rect 7561 21635 7619 21641
rect 7650 21632 7656 21644
rect 7708 21632 7714 21684
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 9033 21675 9091 21681
rect 9033 21672 9045 21675
rect 8904 21644 9045 21672
rect 8904 21632 8910 21644
rect 9033 21641 9045 21644
rect 9079 21641 9091 21675
rect 11514 21672 11520 21684
rect 11475 21644 11520 21672
rect 9033 21635 9091 21641
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 12713 21675 12771 21681
rect 12713 21672 12725 21675
rect 12492 21644 12725 21672
rect 12492 21632 12498 21644
rect 12713 21641 12725 21644
rect 12759 21641 12771 21675
rect 12713 21635 12771 21641
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 14366 21672 14372 21684
rect 12952 21644 14372 21672
rect 12952 21632 12958 21644
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 16298 21672 16304 21684
rect 16259 21644 16304 21672
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16393 21675 16451 21681
rect 16393 21641 16405 21675
rect 16439 21672 16451 21675
rect 17494 21672 17500 21684
rect 16439 21644 17500 21672
rect 16439 21641 16451 21644
rect 16393 21635 16451 21641
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 17865 21675 17923 21681
rect 17865 21641 17877 21675
rect 17911 21672 17923 21675
rect 18322 21672 18328 21684
rect 17911 21644 18328 21672
rect 17911 21641 17923 21644
rect 17865 21635 17923 21641
rect 18322 21632 18328 21644
rect 18380 21632 18386 21684
rect 21450 21672 21456 21684
rect 21411 21644 21456 21672
rect 21450 21632 21456 21644
rect 21508 21632 21514 21684
rect 23198 21672 23204 21684
rect 23159 21644 23204 21672
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 25406 21672 25412 21684
rect 25367 21644 25412 21672
rect 25406 21632 25412 21644
rect 25464 21632 25470 21684
rect 10137 21607 10195 21613
rect 10137 21573 10149 21607
rect 10183 21604 10195 21607
rect 11054 21604 11060 21616
rect 10183 21576 11060 21604
rect 10183 21573 10195 21576
rect 10137 21567 10195 21573
rect 11054 21564 11060 21576
rect 11112 21564 11118 21616
rect 5629 21539 5687 21545
rect 5629 21536 5641 21539
rect 5552 21508 5641 21536
rect 5629 21505 5641 21508
rect 5675 21505 5687 21539
rect 5629 21499 5687 21505
rect 10597 21539 10655 21545
rect 10597 21505 10609 21539
rect 10643 21536 10655 21539
rect 10686 21536 10692 21548
rect 10643 21508 10692 21536
rect 10643 21505 10655 21508
rect 10597 21499 10655 21505
rect 10686 21496 10692 21508
rect 10744 21496 10750 21548
rect 10781 21539 10839 21545
rect 10781 21505 10793 21539
rect 10827 21536 10839 21539
rect 11882 21536 11888 21548
rect 10827 21508 11888 21536
rect 10827 21505 10839 21508
rect 10781 21499 10839 21505
rect 11882 21496 11888 21508
rect 11940 21496 11946 21548
rect 15378 21496 15384 21548
rect 15436 21536 15442 21548
rect 15838 21536 15844 21548
rect 15436 21508 15844 21536
rect 15436 21496 15442 21508
rect 15838 21496 15844 21508
rect 15896 21496 15902 21548
rect 16316 21536 16344 21632
rect 24854 21604 24860 21616
rect 24136 21576 24860 21604
rect 24136 21548 24164 21576
rect 24854 21564 24860 21576
rect 24912 21564 24918 21616
rect 25314 21564 25320 21616
rect 25372 21604 25378 21616
rect 26145 21607 26203 21613
rect 26145 21604 26157 21607
rect 25372 21576 26157 21604
rect 25372 21564 25378 21576
rect 26145 21573 26157 21576
rect 26191 21573 26203 21607
rect 26145 21567 26203 21573
rect 16945 21539 17003 21545
rect 16945 21536 16957 21539
rect 16316 21508 16957 21536
rect 16945 21505 16957 21508
rect 16991 21536 17003 21539
rect 17494 21536 17500 21548
rect 16991 21508 17500 21536
rect 16991 21505 17003 21508
rect 16945 21499 17003 21505
rect 17494 21496 17500 21508
rect 17552 21496 17558 21548
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21536 18843 21539
rect 18874 21536 18880 21548
rect 18831 21508 18880 21536
rect 18831 21505 18843 21508
rect 18785 21499 18843 21505
rect 18874 21496 18880 21508
rect 18932 21496 18938 21548
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 19242 21536 19248 21548
rect 19015 21508 19248 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 19242 21496 19248 21508
rect 19300 21496 19306 21548
rect 20530 21536 20536 21548
rect 20491 21508 20536 21536
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 21266 21496 21272 21548
rect 21324 21536 21330 21548
rect 22097 21539 22155 21545
rect 22097 21536 22109 21539
rect 21324 21508 22109 21536
rect 21324 21496 21330 21508
rect 22097 21505 22109 21508
rect 22143 21505 22155 21539
rect 22278 21536 22284 21548
rect 22239 21508 22284 21536
rect 22097 21499 22155 21505
rect 22278 21496 22284 21508
rect 22336 21496 22342 21548
rect 24118 21536 24124 21548
rect 24031 21508 24124 21536
rect 24118 21496 24124 21508
rect 24176 21496 24182 21548
rect 24213 21539 24271 21545
rect 24213 21505 24225 21539
rect 24259 21505 24271 21539
rect 24213 21499 24271 21505
rect 3660 21440 4108 21468
rect 3660 21428 3666 21440
rect 14 21360 20 21412
rect 72 21400 78 21412
rect 842 21400 848 21412
rect 72 21372 848 21400
rect 72 21360 78 21372
rect 842 21360 848 21372
rect 900 21360 906 21412
rect 4080 21400 4108 21440
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21437 5503 21471
rect 5445 21431 5503 21437
rect 6365 21471 6423 21477
rect 6365 21437 6377 21471
rect 6411 21468 6423 21471
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6411 21440 7021 21468
rect 6411 21437 6423 21440
rect 6365 21431 6423 21437
rect 7009 21437 7021 21440
rect 7055 21468 7067 21471
rect 7098 21468 7104 21480
rect 7055 21440 7104 21468
rect 7055 21437 7067 21440
rect 7009 21431 7067 21437
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7616 21440 7665 21468
rect 7616 21428 7622 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 10042 21428 10048 21480
rect 10100 21468 10106 21480
rect 10962 21468 10968 21480
rect 10100 21440 10968 21468
rect 10100 21428 10106 21440
rect 10962 21428 10968 21440
rect 11020 21468 11026 21480
rect 11149 21471 11207 21477
rect 11149 21468 11161 21471
rect 11020 21440 11161 21468
rect 11020 21428 11026 21440
rect 11149 21437 11161 21440
rect 11195 21468 11207 21471
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 11195 21440 13277 21468
rect 11195 21437 11207 21440
rect 11149 21431 11207 21437
rect 13265 21437 13277 21440
rect 13311 21468 13323 21471
rect 13354 21468 13360 21480
rect 13311 21440 13360 21468
rect 13311 21437 13323 21440
rect 13265 21431 13323 21437
rect 13354 21428 13360 21440
rect 13412 21468 13418 21480
rect 15286 21468 15292 21480
rect 13412 21440 15292 21468
rect 13412 21428 13418 21440
rect 15286 21428 15292 21440
rect 15344 21428 15350 21480
rect 16758 21468 16764 21480
rect 16719 21440 16764 21468
rect 16758 21428 16764 21440
rect 16816 21428 16822 21480
rect 17770 21428 17776 21480
rect 17828 21468 17834 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 17828 21440 18705 21468
rect 17828 21428 17834 21440
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 19610 21428 19616 21480
rect 19668 21468 19674 21480
rect 20070 21468 20076 21480
rect 19668 21440 20076 21468
rect 19668 21428 19674 21440
rect 20070 21428 20076 21440
rect 20128 21428 20134 21480
rect 20349 21471 20407 21477
rect 20349 21437 20361 21471
rect 20395 21468 20407 21471
rect 20622 21468 20628 21480
rect 20395 21440 20628 21468
rect 20395 21437 20407 21440
rect 20349 21431 20407 21437
rect 20622 21428 20628 21440
rect 20680 21428 20686 21480
rect 23934 21428 23940 21480
rect 23992 21468 23998 21480
rect 24029 21471 24087 21477
rect 24029 21468 24041 21471
rect 23992 21440 24041 21468
rect 23992 21428 23998 21440
rect 24029 21437 24041 21440
rect 24075 21437 24087 21471
rect 24029 21431 24087 21437
rect 6181 21403 6239 21409
rect 6181 21400 6193 21403
rect 4080 21372 6193 21400
rect 6181 21369 6193 21372
rect 6227 21400 6239 21403
rect 7920 21403 7978 21409
rect 7920 21400 7932 21403
rect 6227 21372 7932 21400
rect 6227 21369 6239 21372
rect 6181 21363 6239 21369
rect 7920 21369 7932 21372
rect 7966 21400 7978 21403
rect 8294 21400 8300 21412
rect 7966 21372 8300 21400
rect 7966 21369 7978 21372
rect 7920 21363 7978 21369
rect 8294 21360 8300 21372
rect 8352 21360 8358 21412
rect 9766 21400 9772 21412
rect 9679 21372 9772 21400
rect 9766 21360 9772 21372
rect 9824 21400 9830 21412
rect 13532 21403 13590 21409
rect 9824 21372 13216 21400
rect 9824 21360 9830 21372
rect 3602 21292 3608 21344
rect 3660 21332 3666 21344
rect 3881 21335 3939 21341
rect 3881 21332 3893 21335
rect 3660 21304 3893 21332
rect 3660 21292 3666 21304
rect 3881 21301 3893 21304
rect 3927 21301 3939 21335
rect 4614 21332 4620 21344
rect 4575 21304 4620 21332
rect 3881 21295 3939 21301
rect 4614 21292 4620 21304
rect 4672 21292 4678 21344
rect 5534 21292 5540 21344
rect 5592 21332 5598 21344
rect 6362 21332 6368 21344
rect 5592 21304 5637 21332
rect 6323 21304 6368 21332
rect 5592 21292 5598 21304
rect 6362 21292 6368 21304
rect 6420 21292 6426 21344
rect 6546 21332 6552 21344
rect 6507 21304 6552 21332
rect 6546 21292 6552 21304
rect 6604 21332 6610 21344
rect 6641 21335 6699 21341
rect 6641 21332 6653 21335
rect 6604 21304 6653 21332
rect 6604 21292 6610 21304
rect 6641 21301 6653 21304
rect 6687 21301 6699 21335
rect 6641 21295 6699 21301
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10778 21332 10784 21344
rect 10551 21304 10784 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 10778 21292 10784 21304
rect 10836 21332 10842 21344
rect 10962 21332 10968 21344
rect 10836 21304 10968 21332
rect 10836 21292 10842 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11882 21332 11888 21344
rect 11843 21304 11888 21332
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 13188 21341 13216 21372
rect 13532 21369 13544 21403
rect 13578 21400 13590 21403
rect 13630 21400 13636 21412
rect 13578 21372 13636 21400
rect 13578 21369 13590 21372
rect 13532 21363 13590 21369
rect 13630 21360 13636 21372
rect 13688 21360 13694 21412
rect 14182 21360 14188 21412
rect 14240 21400 14246 21412
rect 16298 21400 16304 21412
rect 14240 21372 16304 21400
rect 14240 21360 14246 21372
rect 16298 21360 16304 21372
rect 16356 21360 16362 21412
rect 16850 21400 16856 21412
rect 16763 21372 16856 21400
rect 16850 21360 16856 21372
rect 16908 21400 16914 21412
rect 17862 21400 17868 21412
rect 16908 21372 17868 21400
rect 16908 21360 16914 21372
rect 17862 21360 17868 21372
rect 17920 21360 17926 21412
rect 19702 21400 19708 21412
rect 19663 21372 19708 21400
rect 19702 21360 19708 21372
rect 19760 21400 19766 21412
rect 20257 21403 20315 21409
rect 20257 21400 20269 21403
rect 19760 21372 20269 21400
rect 19760 21360 19766 21372
rect 20257 21369 20269 21372
rect 20303 21369 20315 21403
rect 20257 21363 20315 21369
rect 21085 21403 21143 21409
rect 21085 21369 21097 21403
rect 21131 21400 21143 21403
rect 21818 21400 21824 21412
rect 21131 21372 21824 21400
rect 21131 21369 21143 21372
rect 21085 21363 21143 21369
rect 21818 21360 21824 21372
rect 21876 21360 21882 21412
rect 23014 21360 23020 21412
rect 23072 21400 23078 21412
rect 23198 21400 23204 21412
rect 23072 21372 23204 21400
rect 23072 21360 23078 21372
rect 23198 21360 23204 21372
rect 23256 21400 23262 21412
rect 24228 21400 24256 21499
rect 25130 21428 25136 21480
rect 25188 21468 25194 21480
rect 25225 21471 25283 21477
rect 25225 21468 25237 21471
rect 25188 21440 25237 21468
rect 25188 21428 25194 21440
rect 25225 21437 25237 21440
rect 25271 21468 25283 21471
rect 25777 21471 25835 21477
rect 25777 21468 25789 21471
rect 25271 21440 25789 21468
rect 25271 21437 25283 21440
rect 25225 21431 25283 21437
rect 25777 21437 25789 21440
rect 25823 21437 25835 21471
rect 25777 21431 25835 21437
rect 24673 21403 24731 21409
rect 24673 21400 24685 21403
rect 23256 21372 24685 21400
rect 23256 21360 23262 21372
rect 24673 21369 24685 21372
rect 24719 21369 24731 21403
rect 24673 21363 24731 21369
rect 13173 21335 13231 21341
rect 13173 21301 13185 21335
rect 13219 21332 13231 21335
rect 14458 21332 14464 21344
rect 13219 21304 14464 21332
rect 13219 21301 13231 21304
rect 13173 21295 13231 21301
rect 14458 21292 14464 21304
rect 14516 21292 14522 21344
rect 14645 21335 14703 21341
rect 14645 21301 14657 21335
rect 14691 21332 14703 21335
rect 15194 21332 15200 21344
rect 14691 21304 15200 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 15194 21292 15200 21304
rect 15252 21332 15258 21344
rect 15657 21335 15715 21341
rect 15657 21332 15669 21335
rect 15252 21304 15669 21332
rect 15252 21292 15258 21304
rect 15657 21301 15669 21304
rect 15703 21332 15715 21335
rect 15930 21332 15936 21344
rect 15703 21304 15936 21332
rect 15703 21301 15715 21304
rect 15657 21295 15715 21301
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 18325 21335 18383 21341
rect 18325 21301 18337 21335
rect 18371 21332 18383 21335
rect 18414 21332 18420 21344
rect 18371 21304 18420 21332
rect 18371 21301 18383 21304
rect 18325 21295 18383 21301
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 19337 21335 19395 21341
rect 19337 21332 19349 21335
rect 18840 21304 19349 21332
rect 18840 21292 18846 21304
rect 19337 21301 19349 21304
rect 19383 21332 19395 21335
rect 19518 21332 19524 21344
rect 19383 21304 19524 21332
rect 19383 21301 19395 21304
rect 19337 21295 19395 21301
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 19889 21335 19947 21341
rect 19889 21301 19901 21335
rect 19935 21332 19947 21335
rect 19978 21332 19984 21344
rect 19935 21304 19984 21332
rect 19935 21301 19947 21304
rect 19889 21295 19947 21301
rect 19978 21292 19984 21304
rect 20036 21292 20042 21344
rect 21634 21332 21640 21344
rect 21595 21304 21640 21332
rect 21634 21292 21640 21304
rect 21692 21292 21698 21344
rect 21910 21292 21916 21344
rect 21968 21332 21974 21344
rect 22005 21335 22063 21341
rect 22005 21332 22017 21335
rect 21968 21304 22017 21332
rect 21968 21292 21974 21304
rect 22005 21301 22017 21304
rect 22051 21301 22063 21335
rect 22005 21295 22063 21301
rect 22925 21335 22983 21341
rect 22925 21301 22937 21335
rect 22971 21332 22983 21335
rect 23382 21332 23388 21344
rect 22971 21304 23388 21332
rect 22971 21301 22983 21304
rect 22925 21295 22983 21301
rect 23382 21292 23388 21304
rect 23440 21292 23446 21344
rect 23658 21332 23664 21344
rect 23619 21304 23664 21332
rect 23658 21292 23664 21304
rect 23716 21292 23722 21344
rect 1104 21242 26864 21264
rect 1104 21190 10315 21242
rect 10367 21190 10379 21242
rect 10431 21190 10443 21242
rect 10495 21190 10507 21242
rect 10559 21190 19648 21242
rect 19700 21190 19712 21242
rect 19764 21190 19776 21242
rect 19828 21190 19840 21242
rect 19892 21190 26864 21242
rect 1104 21168 26864 21190
rect 1854 21088 1860 21140
rect 1912 21128 1918 21140
rect 1949 21131 2007 21137
rect 1949 21128 1961 21131
rect 1912 21100 1961 21128
rect 1912 21088 1918 21100
rect 1949 21097 1961 21100
rect 1995 21097 2007 21131
rect 2314 21128 2320 21140
rect 2275 21100 2320 21128
rect 1949 21091 2007 21097
rect 2314 21088 2320 21100
rect 2372 21128 2378 21140
rect 3142 21128 3148 21140
rect 2372 21100 3148 21128
rect 2372 21088 2378 21100
rect 3142 21088 3148 21100
rect 3200 21088 3206 21140
rect 4062 21128 4068 21140
rect 4023 21100 4068 21128
rect 4062 21088 4068 21100
rect 4120 21088 4126 21140
rect 4522 21128 4528 21140
rect 4483 21100 4528 21128
rect 4522 21088 4528 21100
rect 4580 21128 4586 21140
rect 4798 21128 4804 21140
rect 4580 21100 4804 21128
rect 4580 21088 4586 21100
rect 4798 21088 4804 21100
rect 4856 21088 4862 21140
rect 7282 21088 7288 21140
rect 7340 21128 7346 21140
rect 7561 21131 7619 21137
rect 7561 21128 7573 21131
rect 7340 21100 7573 21128
rect 7340 21088 7346 21100
rect 7561 21097 7573 21100
rect 7607 21128 7619 21131
rect 8018 21128 8024 21140
rect 7607 21100 8024 21128
rect 7607 21097 7619 21100
rect 7561 21091 7619 21097
rect 8018 21088 8024 21100
rect 8076 21088 8082 21140
rect 9030 21128 9036 21140
rect 8991 21100 9036 21128
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 11057 21131 11115 21137
rect 11057 21128 11069 21131
rect 10980 21100 11069 21128
rect 1765 21063 1823 21069
rect 1765 21029 1777 21063
rect 1811 21060 1823 21063
rect 2406 21060 2412 21072
rect 1811 21032 2412 21060
rect 1811 21029 1823 21032
rect 1765 21023 1823 21029
rect 2406 21020 2412 21032
rect 2464 21020 2470 21072
rect 6089 21063 6147 21069
rect 6089 21029 6101 21063
rect 6135 21060 6147 21063
rect 6362 21060 6368 21072
rect 6135 21032 6368 21060
rect 6135 21029 6147 21032
rect 6089 21023 6147 21029
rect 6362 21020 6368 21032
rect 6420 21020 6426 21072
rect 9674 21020 9680 21072
rect 9732 21060 9738 21072
rect 9922 21063 9980 21069
rect 9922 21060 9934 21063
rect 9732 21032 9934 21060
rect 9732 21020 9738 21032
rect 9922 21029 9934 21032
rect 9968 21029 9980 21063
rect 9922 21023 9980 21029
rect 10980 21060 11008 21100
rect 11057 21097 11069 21100
rect 11103 21097 11115 21131
rect 11057 21091 11115 21097
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12161 21131 12219 21137
rect 12161 21128 12173 21131
rect 12124 21100 12173 21128
rect 12124 21088 12130 21100
rect 12161 21097 12173 21100
rect 12207 21097 12219 21131
rect 12161 21091 12219 21097
rect 13541 21131 13599 21137
rect 13541 21097 13553 21131
rect 13587 21128 13599 21131
rect 13722 21128 13728 21140
rect 13587 21100 13728 21128
rect 13587 21097 13599 21100
rect 13541 21091 13599 21097
rect 13722 21088 13728 21100
rect 13780 21088 13786 21140
rect 14274 21128 14280 21140
rect 14235 21100 14280 21128
rect 14274 21088 14280 21100
rect 14332 21088 14338 21140
rect 14458 21088 14464 21140
rect 14516 21128 14522 21140
rect 14826 21128 14832 21140
rect 14516 21100 14832 21128
rect 14516 21088 14522 21100
rect 14826 21088 14832 21100
rect 14884 21128 14890 21140
rect 15289 21131 15347 21137
rect 15289 21128 15301 21131
rect 14884 21100 15301 21128
rect 14884 21088 14890 21100
rect 15289 21097 15301 21100
rect 15335 21097 15347 21131
rect 16850 21128 16856 21140
rect 16811 21100 16856 21128
rect 15289 21091 15347 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 18049 21131 18107 21137
rect 18049 21128 18061 21131
rect 16991 21100 18061 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 18049 21097 18061 21100
rect 18095 21128 18107 21131
rect 18138 21128 18144 21140
rect 18095 21100 18144 21128
rect 18095 21097 18107 21100
rect 18049 21091 18107 21097
rect 18138 21088 18144 21100
rect 18196 21088 18202 21140
rect 18966 21128 18972 21140
rect 18927 21100 18972 21128
rect 18966 21088 18972 21100
rect 19024 21088 19030 21140
rect 19058 21088 19064 21140
rect 19116 21128 19122 21140
rect 19613 21131 19671 21137
rect 19613 21128 19625 21131
rect 19116 21100 19625 21128
rect 19116 21088 19122 21100
rect 19613 21097 19625 21100
rect 19659 21097 19671 21131
rect 20346 21128 20352 21140
rect 20307 21100 20352 21128
rect 19613 21091 19671 21097
rect 12710 21060 12716 21072
rect 10980 21032 12716 21060
rect 3970 20952 3976 21004
rect 4028 20992 4034 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 4028 20964 4445 20992
rect 4028 20952 4034 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 5997 20995 6055 21001
rect 5997 20961 6009 20995
rect 6043 20992 6055 20995
rect 6270 20992 6276 21004
rect 6043 20964 6276 20992
rect 6043 20961 6055 20964
rect 5997 20955 6055 20961
rect 6270 20952 6276 20964
rect 6328 20952 6334 21004
rect 7101 20995 7159 21001
rect 7101 20961 7113 20995
rect 7147 20992 7159 20995
rect 8294 20992 8300 21004
rect 7147 20964 8300 20992
rect 7147 20961 7159 20964
rect 7101 20955 7159 20961
rect 8294 20952 8300 20964
rect 8352 20992 8358 21004
rect 10980 20992 11008 21032
rect 12710 21020 12716 21032
rect 12768 21020 12774 21072
rect 13630 21020 13636 21072
rect 13688 21060 13694 21072
rect 13817 21063 13875 21069
rect 13817 21060 13829 21063
rect 13688 21032 13829 21060
rect 13688 21020 13694 21032
rect 13817 21029 13829 21032
rect 13863 21029 13875 21063
rect 13817 21023 13875 21029
rect 16574 21020 16580 21072
rect 16632 21060 16638 21072
rect 17313 21063 17371 21069
rect 17313 21060 17325 21063
rect 16632 21032 17325 21060
rect 16632 21020 16638 21032
rect 17313 21029 17325 21032
rect 17359 21060 17371 21063
rect 17862 21060 17868 21072
rect 17359 21032 17868 21060
rect 17359 21029 17371 21032
rect 17313 21023 17371 21029
rect 17862 21020 17868 21032
rect 17920 21020 17926 21072
rect 18417 21063 18475 21069
rect 18417 21029 18429 21063
rect 18463 21060 18475 21063
rect 19242 21060 19248 21072
rect 18463 21032 19248 21060
rect 18463 21029 18475 21032
rect 18417 21023 18475 21029
rect 19242 21020 19248 21032
rect 19300 21060 19306 21072
rect 19518 21060 19524 21072
rect 19300 21032 19524 21060
rect 19300 21020 19306 21032
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 8352 20964 11008 20992
rect 12069 20995 12127 21001
rect 8352 20952 8358 20964
rect 12069 20961 12081 20995
rect 12115 20992 12127 20995
rect 12526 20992 12532 21004
rect 12115 20964 12532 20992
rect 12115 20961 12127 20964
rect 12069 20955 12127 20961
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 12618 20952 12624 21004
rect 12676 20992 12682 21004
rect 14093 20995 14151 21001
rect 12676 20964 12721 20992
rect 12676 20952 12682 20964
rect 14093 20961 14105 20995
rect 14139 20992 14151 20995
rect 14734 20992 14740 21004
rect 14139 20964 14740 20992
rect 14139 20961 14151 20964
rect 14093 20955 14151 20961
rect 14734 20952 14740 20964
rect 14792 20952 14798 21004
rect 15657 20995 15715 21001
rect 15657 20961 15669 20995
rect 15703 20961 15715 20995
rect 15657 20955 15715 20961
rect 16485 20995 16543 21001
rect 16485 20961 16497 20995
rect 16531 20992 16543 20995
rect 16942 20992 16948 21004
rect 16531 20964 16948 20992
rect 16531 20961 16543 20964
rect 16485 20955 16543 20961
rect 2409 20927 2467 20933
rect 2409 20893 2421 20927
rect 2455 20893 2467 20927
rect 2590 20924 2596 20936
rect 2551 20896 2596 20924
rect 2409 20887 2467 20893
rect 2424 20856 2452 20887
rect 2590 20884 2596 20896
rect 2648 20884 2654 20936
rect 3237 20927 3295 20933
rect 3237 20893 3249 20927
rect 3283 20924 3295 20927
rect 4617 20927 4675 20933
rect 4617 20924 4629 20927
rect 3283 20896 4629 20924
rect 3283 20893 3295 20896
rect 3237 20887 3295 20893
rect 4617 20893 4629 20896
rect 4663 20924 4675 20927
rect 5077 20927 5135 20933
rect 5077 20924 5089 20927
rect 4663 20896 5089 20924
rect 4663 20893 4675 20896
rect 4617 20887 4675 20893
rect 5077 20893 5089 20896
rect 5123 20924 5135 20927
rect 5350 20924 5356 20936
rect 5123 20896 5356 20924
rect 5123 20893 5135 20896
rect 5077 20887 5135 20893
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 6181 20927 6239 20933
rect 6181 20893 6193 20927
rect 6227 20924 6239 20927
rect 6454 20924 6460 20936
rect 6227 20896 6460 20924
rect 6227 20893 6239 20896
rect 6181 20887 6239 20893
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 7650 20924 7656 20936
rect 7611 20896 7656 20924
rect 7650 20884 7656 20896
rect 7708 20884 7714 20936
rect 7742 20884 7748 20936
rect 7800 20924 7806 20936
rect 9677 20927 9735 20933
rect 7800 20896 7845 20924
rect 7800 20884 7806 20896
rect 9677 20893 9689 20927
rect 9723 20893 9735 20927
rect 11606 20924 11612 20936
rect 11567 20896 11612 20924
rect 9677 20887 9735 20893
rect 2866 20856 2872 20868
rect 2424 20828 2872 20856
rect 2866 20816 2872 20828
rect 2924 20816 2930 20868
rect 3878 20816 3884 20868
rect 3936 20856 3942 20868
rect 5445 20859 5503 20865
rect 5445 20856 5457 20859
rect 3936 20828 5457 20856
rect 3936 20816 3942 20828
rect 5445 20825 5457 20828
rect 5491 20825 5503 20859
rect 5445 20819 5503 20825
rect 5534 20816 5540 20868
rect 5592 20856 5598 20868
rect 5629 20859 5687 20865
rect 5629 20856 5641 20859
rect 5592 20828 5641 20856
rect 5592 20816 5598 20828
rect 5629 20825 5641 20828
rect 5675 20856 5687 20859
rect 6641 20859 6699 20865
rect 6641 20856 6653 20859
rect 5675 20828 6653 20856
rect 5675 20825 5687 20828
rect 5629 20819 5687 20825
rect 6641 20825 6653 20828
rect 6687 20825 6699 20859
rect 6641 20819 6699 20825
rect 8478 20816 8484 20868
rect 8536 20856 8542 20868
rect 8665 20859 8723 20865
rect 8665 20856 8677 20859
rect 8536 20828 8677 20856
rect 8536 20816 8542 20828
rect 8665 20825 8677 20828
rect 8711 20856 8723 20859
rect 9582 20856 9588 20868
rect 8711 20828 9588 20856
rect 8711 20825 8723 20828
rect 8665 20819 8723 20825
rect 9582 20816 9588 20828
rect 9640 20816 9646 20868
rect 3602 20788 3608 20800
rect 3563 20760 3608 20788
rect 3602 20748 3608 20760
rect 3660 20748 3666 20800
rect 7190 20788 7196 20800
rect 7151 20760 7196 20788
rect 7190 20748 7196 20760
rect 7248 20748 7254 20800
rect 9398 20788 9404 20800
rect 9359 20760 9404 20788
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 9692 20788 9720 20887
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 12710 20884 12716 20936
rect 12768 20924 12774 20936
rect 12768 20896 12813 20924
rect 12768 20884 12774 20896
rect 10042 20788 10048 20800
rect 9692 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 14642 20788 14648 20800
rect 14603 20760 14648 20788
rect 14642 20748 14648 20760
rect 14700 20748 14706 20800
rect 14826 20748 14832 20800
rect 14884 20788 14890 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14884 20760 15025 20788
rect 14884 20748 14890 20760
rect 15013 20757 15025 20760
rect 15059 20788 15071 20791
rect 15672 20788 15700 20955
rect 16942 20952 16948 20964
rect 17000 20952 17006 21004
rect 17405 20995 17463 21001
rect 17405 20961 17417 20995
rect 17451 20992 17463 20995
rect 17586 20992 17592 21004
rect 17451 20964 17592 20992
rect 17451 20961 17463 20964
rect 17405 20955 17463 20961
rect 17586 20952 17592 20964
rect 17644 20952 17650 21004
rect 18138 20952 18144 21004
rect 18196 20992 18202 21004
rect 18506 20992 18512 21004
rect 18196 20964 18512 20992
rect 18196 20952 18202 20964
rect 18506 20952 18512 20964
rect 18564 20952 18570 21004
rect 18874 20992 18880 21004
rect 18835 20964 18880 20992
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 15746 20884 15752 20936
rect 15804 20924 15810 20936
rect 15930 20924 15936 20936
rect 15804 20896 15849 20924
rect 15891 20896 15936 20924
rect 15804 20884 15810 20896
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16206 20884 16212 20936
rect 16264 20884 16270 20936
rect 17494 20924 17500 20936
rect 17455 20896 17500 20924
rect 17494 20884 17500 20896
rect 17552 20884 17558 20936
rect 19058 20924 19064 20936
rect 19019 20896 19064 20924
rect 19058 20884 19064 20896
rect 19116 20884 19122 20936
rect 16224 20856 16252 20884
rect 15948 20828 16252 20856
rect 19628 20856 19656 21091
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 20714 21128 20720 21140
rect 20675 21100 20720 21128
rect 20714 21088 20720 21100
rect 20772 21088 20778 21140
rect 21726 21128 21732 21140
rect 21687 21100 21732 21128
rect 21726 21088 21732 21100
rect 21784 21088 21790 21140
rect 23658 21088 23664 21140
rect 23716 21128 23722 21140
rect 24213 21131 24271 21137
rect 24213 21128 24225 21131
rect 23716 21100 24225 21128
rect 23716 21088 23722 21100
rect 24213 21097 24225 21100
rect 24259 21128 24271 21131
rect 24765 21131 24823 21137
rect 24765 21128 24777 21131
rect 24259 21100 24777 21128
rect 24259 21097 24271 21100
rect 24213 21091 24271 21097
rect 24765 21097 24777 21100
rect 24811 21097 24823 21131
rect 24765 21091 24823 21097
rect 19981 21063 20039 21069
rect 19981 21029 19993 21063
rect 20027 21060 20039 21063
rect 20622 21060 20628 21072
rect 20027 21032 20628 21060
rect 20027 21029 20039 21032
rect 19981 21023 20039 21029
rect 20622 21020 20628 21032
rect 20680 21020 20686 21072
rect 22186 21069 22192 21072
rect 22180 21060 22192 21069
rect 22147 21032 22192 21060
rect 22180 21023 22192 21032
rect 22186 21020 22192 21023
rect 22244 21020 22250 21072
rect 22462 21020 22468 21072
rect 22520 21060 22526 21072
rect 23937 21063 23995 21069
rect 23937 21060 23949 21063
rect 22520 21032 23949 21060
rect 22520 21020 22526 21032
rect 23937 21029 23949 21032
rect 23983 21060 23995 21063
rect 24118 21060 24124 21072
rect 23983 21032 24124 21060
rect 23983 21029 23995 21032
rect 23937 21023 23995 21029
rect 24118 21020 24124 21032
rect 24176 21020 24182 21072
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20893 21971 20927
rect 21913 20887 21971 20893
rect 20806 20856 20812 20868
rect 19628 20828 20812 20856
rect 15948 20800 15976 20828
rect 20806 20816 20812 20828
rect 20864 20856 20870 20868
rect 21928 20856 21956 20887
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 24857 20927 24915 20933
rect 24857 20924 24869 20927
rect 23532 20896 24869 20924
rect 23532 20884 23538 20896
rect 24857 20893 24869 20896
rect 24903 20893 24915 20927
rect 25038 20924 25044 20936
rect 24999 20896 25044 20924
rect 24857 20887 24915 20893
rect 20864 20828 21956 20856
rect 24872 20856 24900 20887
rect 25038 20884 25044 20896
rect 25096 20884 25102 20936
rect 26234 20856 26240 20868
rect 24872 20828 26240 20856
rect 20864 20816 20870 20828
rect 26234 20816 26240 20828
rect 26292 20816 26298 20868
rect 15059 20760 15700 20788
rect 15059 20757 15071 20760
rect 15013 20751 15071 20757
rect 15930 20748 15936 20800
rect 15988 20748 15994 20800
rect 16206 20748 16212 20800
rect 16264 20788 16270 20800
rect 16482 20788 16488 20800
rect 16264 20760 16488 20788
rect 16264 20748 16270 20760
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 18506 20788 18512 20800
rect 18467 20760 18512 20788
rect 18506 20748 18512 20760
rect 18564 20748 18570 20800
rect 19150 20748 19156 20800
rect 19208 20788 19214 20800
rect 19426 20788 19432 20800
rect 19208 20760 19432 20788
rect 19208 20748 19214 20760
rect 19426 20748 19432 20760
rect 19484 20748 19490 20800
rect 21818 20748 21824 20800
rect 21876 20788 21882 20800
rect 23293 20791 23351 20797
rect 23293 20788 23305 20791
rect 21876 20760 23305 20788
rect 21876 20748 21882 20760
rect 23293 20757 23305 20760
rect 23339 20788 23351 20791
rect 23566 20788 23572 20800
rect 23339 20760 23572 20788
rect 23339 20757 23351 20760
rect 23293 20751 23351 20757
rect 23566 20748 23572 20760
rect 23624 20748 23630 20800
rect 24118 20748 24124 20800
rect 24176 20788 24182 20800
rect 24397 20791 24455 20797
rect 24397 20788 24409 20791
rect 24176 20760 24409 20788
rect 24176 20748 24182 20760
rect 24397 20757 24409 20760
rect 24443 20757 24455 20791
rect 24397 20751 24455 20757
rect 1104 20698 26864 20720
rect 1104 20646 5648 20698
rect 5700 20646 5712 20698
rect 5764 20646 5776 20698
rect 5828 20646 5840 20698
rect 5892 20646 14982 20698
rect 15034 20646 15046 20698
rect 15098 20646 15110 20698
rect 15162 20646 15174 20698
rect 15226 20646 24315 20698
rect 24367 20646 24379 20698
rect 24431 20646 24443 20698
rect 24495 20646 24507 20698
rect 24559 20646 26864 20698
rect 1104 20624 26864 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1765 20587 1823 20593
rect 1765 20584 1777 20587
rect 992 20556 1777 20584
rect 992 20544 998 20556
rect 1765 20553 1777 20556
rect 1811 20553 1823 20587
rect 1765 20547 1823 20553
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2130 20584 2136 20596
rect 1995 20556 2136 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 1780 20448 1808 20547
rect 2130 20544 2136 20556
rect 2188 20544 2194 20596
rect 2866 20544 2872 20596
rect 2924 20584 2930 20596
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 2924 20556 3065 20584
rect 2924 20544 2930 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 3694 20584 3700 20596
rect 3099 20556 3700 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 3694 20544 3700 20556
rect 3752 20584 3758 20596
rect 6181 20587 6239 20593
rect 6181 20584 6193 20587
rect 3752 20556 6193 20584
rect 3752 20544 3758 20556
rect 6181 20553 6193 20556
rect 6227 20584 6239 20587
rect 6270 20584 6276 20596
rect 6227 20556 6276 20584
rect 6227 20553 6239 20556
rect 6181 20547 6239 20553
rect 6270 20544 6276 20556
rect 6328 20544 6334 20596
rect 6454 20584 6460 20596
rect 6415 20556 6460 20584
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7377 20587 7435 20593
rect 7377 20584 7389 20587
rect 6972 20556 7389 20584
rect 6972 20544 6978 20556
rect 7377 20553 7389 20556
rect 7423 20584 7435 20587
rect 7742 20584 7748 20596
rect 7423 20556 7748 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 9582 20544 9588 20596
rect 9640 20584 9646 20596
rect 10321 20587 10379 20593
rect 10321 20584 10333 20587
rect 9640 20556 10333 20584
rect 9640 20544 9646 20556
rect 10321 20553 10333 20556
rect 10367 20553 10379 20587
rect 10321 20547 10379 20553
rect 10870 20544 10876 20596
rect 10928 20544 10934 20596
rect 12437 20587 12495 20593
rect 12437 20553 12449 20587
rect 12483 20584 12495 20587
rect 12526 20584 12532 20596
rect 12483 20556 12532 20584
rect 12483 20553 12495 20556
rect 12437 20547 12495 20553
rect 12526 20544 12532 20556
rect 12584 20544 12590 20596
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 13449 20587 13507 20593
rect 13449 20584 13461 20587
rect 12860 20556 13461 20584
rect 12860 20544 12866 20556
rect 13449 20553 13461 20556
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 16209 20587 16267 20593
rect 16209 20584 16221 20587
rect 14424 20556 16221 20584
rect 14424 20544 14430 20556
rect 16209 20553 16221 20556
rect 16255 20553 16267 20587
rect 16209 20547 16267 20553
rect 16393 20587 16451 20593
rect 16393 20553 16405 20587
rect 16439 20584 16451 20587
rect 16482 20584 16488 20596
rect 16439 20556 16488 20584
rect 16439 20553 16451 20556
rect 16393 20547 16451 20553
rect 3142 20476 3148 20528
rect 3200 20516 3206 20528
rect 3329 20519 3387 20525
rect 3329 20516 3341 20519
rect 3200 20488 3341 20516
rect 3200 20476 3206 20488
rect 3329 20485 3341 20488
rect 3375 20516 3387 20519
rect 3510 20516 3516 20528
rect 3375 20488 3516 20516
rect 3375 20485 3387 20488
rect 3329 20479 3387 20485
rect 3510 20476 3516 20488
rect 3568 20476 3574 20528
rect 6472 20516 6500 20544
rect 10229 20519 10287 20525
rect 6472 20488 7880 20516
rect 2406 20448 2412 20460
rect 1780 20420 2412 20448
rect 2406 20408 2412 20420
rect 2464 20408 2470 20460
rect 2590 20448 2596 20460
rect 2551 20420 2596 20448
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 7852 20448 7880 20488
rect 10229 20485 10241 20519
rect 10275 20516 10287 20519
rect 10888 20516 10916 20544
rect 10275 20488 10916 20516
rect 10275 20485 10287 20488
rect 10229 20479 10287 20485
rect 10962 20476 10968 20528
rect 11020 20516 11026 20528
rect 12618 20516 12624 20528
rect 11020 20488 12624 20516
rect 11020 20476 11026 20488
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 13909 20519 13967 20525
rect 13909 20485 13921 20519
rect 13955 20516 13967 20519
rect 13955 20488 14596 20516
rect 13955 20485 13967 20488
rect 13909 20479 13967 20485
rect 14568 20460 14596 20488
rect 14918 20476 14924 20528
rect 14976 20516 14982 20528
rect 15470 20516 15476 20528
rect 14976 20488 15476 20516
rect 14976 20476 14982 20488
rect 15470 20476 15476 20488
rect 15528 20476 15534 20528
rect 7800 20420 7972 20448
rect 7800 20408 7806 20420
rect 3786 20380 3792 20392
rect 3747 20352 3792 20380
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 4056 20383 4114 20389
rect 4056 20349 4068 20383
rect 4102 20380 4114 20383
rect 4614 20380 4620 20392
rect 4102 20352 4620 20380
rect 4102 20349 4114 20352
rect 4056 20343 4114 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20380 5782 20392
rect 6362 20380 6368 20392
rect 5776 20352 6368 20380
rect 5776 20340 5782 20352
rect 6362 20340 6368 20352
rect 6420 20340 6426 20392
rect 7837 20383 7895 20389
rect 7837 20380 7849 20383
rect 7668 20352 7849 20380
rect 7668 20256 7696 20352
rect 7837 20349 7849 20352
rect 7883 20349 7895 20383
rect 7944 20380 7972 20420
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 9732 20420 10885 20448
rect 9732 20408 9738 20420
rect 10873 20417 10885 20420
rect 10919 20448 10931 20451
rect 11333 20451 11391 20457
rect 11333 20448 11345 20451
rect 10919 20420 11345 20448
rect 10919 20417 10931 20420
rect 10873 20411 10931 20417
rect 11333 20417 11345 20420
rect 11379 20448 11391 20451
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11379 20420 11805 20448
rect 11379 20417 11391 20420
rect 11333 20411 11391 20417
rect 11793 20417 11805 20420
rect 11839 20448 11851 20451
rect 11882 20448 11888 20460
rect 11839 20420 11888 20448
rect 11839 20417 11851 20420
rect 11793 20411 11851 20417
rect 11882 20408 11888 20420
rect 11940 20448 11946 20460
rect 12989 20451 13047 20457
rect 12989 20448 13001 20451
rect 11940 20420 13001 20448
rect 11940 20408 11946 20420
rect 12989 20417 13001 20420
rect 13035 20417 13047 20451
rect 14550 20448 14556 20460
rect 14511 20420 14556 20448
rect 12989 20411 13047 20417
rect 14550 20408 14556 20420
rect 14608 20408 14614 20460
rect 8093 20383 8151 20389
rect 8093 20380 8105 20383
rect 7944 20352 8105 20380
rect 7837 20343 7895 20349
rect 8093 20349 8105 20352
rect 8139 20380 8151 20383
rect 8570 20380 8576 20392
rect 8139 20352 8576 20380
rect 8139 20349 8151 20352
rect 8093 20343 8151 20349
rect 8570 20340 8576 20352
rect 8628 20340 8634 20392
rect 10778 20380 10784 20392
rect 10739 20352 10784 20380
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 12618 20380 12624 20392
rect 12176 20352 12624 20380
rect 11514 20312 11520 20324
rect 10704 20284 11520 20312
rect 10704 20256 10732 20284
rect 11514 20272 11520 20284
rect 11572 20272 11578 20324
rect 12176 20256 12204 20352
rect 12618 20340 12624 20352
rect 12676 20340 12682 20392
rect 12894 20380 12900 20392
rect 12855 20352 12900 20380
rect 12894 20340 12900 20352
rect 12952 20340 12958 20392
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 15657 20383 15715 20389
rect 15657 20380 15669 20383
rect 13504 20352 15669 20380
rect 13504 20340 13510 20352
rect 15657 20349 15669 20352
rect 15703 20380 15715 20383
rect 15746 20380 15752 20392
rect 15703 20352 15752 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 15746 20340 15752 20352
rect 15804 20340 15810 20392
rect 14461 20315 14519 20321
rect 14461 20281 14473 20315
rect 14507 20312 14519 20315
rect 14550 20312 14556 20324
rect 14507 20284 14556 20312
rect 14507 20281 14519 20284
rect 14461 20275 14519 20281
rect 14550 20272 14556 20284
rect 14608 20272 14614 20324
rect 16224 20312 16252 20547
rect 16482 20544 16488 20556
rect 16540 20544 16546 20596
rect 17494 20584 17500 20596
rect 17455 20556 17500 20584
rect 17494 20544 17500 20556
rect 17552 20544 17558 20596
rect 18966 20584 18972 20596
rect 18927 20556 18972 20584
rect 18966 20544 18972 20556
rect 19024 20544 19030 20596
rect 21177 20587 21235 20593
rect 21177 20553 21189 20587
rect 21223 20584 21235 20587
rect 21450 20584 21456 20596
rect 21223 20556 21456 20584
rect 21223 20553 21235 20556
rect 21177 20547 21235 20553
rect 21450 20544 21456 20556
rect 21508 20584 21514 20596
rect 22186 20584 22192 20596
rect 21508 20556 22192 20584
rect 21508 20544 21514 20556
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 23474 20584 23480 20596
rect 23435 20556 23480 20584
rect 23474 20544 23480 20556
rect 23532 20584 23538 20596
rect 23532 20556 24164 20584
rect 23532 20544 23538 20556
rect 18233 20519 18291 20525
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 19150 20516 19156 20528
rect 18279 20488 19156 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 19150 20476 19156 20488
rect 19208 20476 19214 20528
rect 20806 20476 20812 20528
rect 20864 20516 20870 20528
rect 22646 20516 22652 20528
rect 20864 20488 22652 20516
rect 20864 20476 20870 20488
rect 22646 20476 22652 20488
rect 22704 20476 22710 20528
rect 22830 20476 22836 20528
rect 22888 20516 22894 20528
rect 23661 20519 23719 20525
rect 23661 20516 23673 20519
rect 22888 20488 23673 20516
rect 22888 20476 22894 20488
rect 23661 20485 23673 20488
rect 23707 20485 23719 20519
rect 23661 20479 23719 20485
rect 16942 20448 16948 20460
rect 16903 20420 16948 20448
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 22278 20448 22284 20460
rect 20588 20420 22284 20448
rect 20588 20408 20594 20420
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 24136 20457 24164 20556
rect 24854 20544 24860 20596
rect 24912 20584 24918 20596
rect 25409 20587 25467 20593
rect 25409 20584 25421 20587
rect 24912 20556 25421 20584
rect 24912 20544 24918 20556
rect 25409 20553 25421 20556
rect 25455 20553 25467 20587
rect 26234 20584 26240 20596
rect 26195 20556 26240 20584
rect 25409 20547 25467 20553
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 24121 20451 24179 20457
rect 24121 20417 24133 20451
rect 24167 20417 24179 20451
rect 24302 20448 24308 20460
rect 24263 20420 24308 20448
rect 24121 20411 24179 20417
rect 16758 20380 16764 20392
rect 16719 20352 16764 20380
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 18046 20380 18052 20392
rect 18007 20352 18052 20380
rect 18046 20340 18052 20352
rect 18104 20380 18110 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18104 20352 18613 20380
rect 18104 20340 18110 20352
rect 18601 20349 18613 20352
rect 18647 20349 18659 20383
rect 18601 20343 18659 20349
rect 19153 20383 19211 20389
rect 19153 20349 19165 20383
rect 19199 20380 19211 20383
rect 19242 20380 19248 20392
rect 19199 20352 19248 20380
rect 19199 20349 19211 20352
rect 19153 20343 19211 20349
rect 19242 20340 19248 20352
rect 19300 20340 19306 20392
rect 21545 20383 21603 20389
rect 21545 20349 21557 20383
rect 21591 20380 21603 20383
rect 21634 20380 21640 20392
rect 21591 20352 21640 20380
rect 21591 20349 21603 20352
rect 21545 20343 21603 20349
rect 21634 20340 21640 20352
rect 21692 20340 21698 20392
rect 21726 20340 21732 20392
rect 21784 20380 21790 20392
rect 22005 20383 22063 20389
rect 22005 20380 22017 20383
rect 21784 20352 22017 20380
rect 21784 20340 21790 20352
rect 22005 20349 22017 20352
rect 22051 20349 22063 20383
rect 22005 20343 22063 20349
rect 22097 20383 22155 20389
rect 22097 20349 22109 20383
rect 22143 20380 22155 20383
rect 22462 20380 22468 20392
rect 22143 20352 22468 20380
rect 22143 20349 22155 20352
rect 22097 20343 22155 20349
rect 22462 20340 22468 20352
rect 22520 20340 22526 20392
rect 24136 20380 24164 20411
rect 24302 20408 24308 20420
rect 24360 20448 24366 20460
rect 24673 20451 24731 20457
rect 24673 20448 24685 20451
rect 24360 20420 24685 20448
rect 24360 20408 24366 20420
rect 24673 20417 24685 20420
rect 24719 20417 24731 20451
rect 24673 20411 24731 20417
rect 25225 20383 25283 20389
rect 25225 20380 25237 20383
rect 24136 20352 25237 20380
rect 25225 20349 25237 20352
rect 25271 20380 25283 20383
rect 25777 20383 25835 20389
rect 25777 20380 25789 20383
rect 25271 20352 25789 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 25777 20349 25789 20352
rect 25823 20349 25835 20383
rect 25777 20343 25835 20349
rect 16850 20312 16856 20324
rect 16224 20284 16856 20312
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 17770 20312 17776 20324
rect 17731 20284 17776 20312
rect 17770 20272 17776 20284
rect 17828 20272 17834 20324
rect 19420 20315 19478 20321
rect 19420 20281 19432 20315
rect 19466 20312 19478 20315
rect 19518 20312 19524 20324
rect 19466 20284 19524 20312
rect 19466 20281 19478 20284
rect 19420 20275 19478 20281
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 23109 20315 23167 20321
rect 23109 20281 23121 20315
rect 23155 20312 23167 20315
rect 24029 20315 24087 20321
rect 24029 20312 24041 20315
rect 23155 20284 24041 20312
rect 23155 20281 23167 20284
rect 23109 20275 23167 20281
rect 24029 20281 24041 20284
rect 24075 20312 24087 20315
rect 24210 20312 24216 20324
rect 24075 20284 24216 20312
rect 24075 20281 24087 20284
rect 24029 20275 24087 20281
rect 24210 20272 24216 20284
rect 24268 20272 24274 20324
rect 2314 20244 2320 20256
rect 2275 20216 2320 20244
rect 2314 20204 2320 20216
rect 2372 20204 2378 20256
rect 4522 20204 4528 20256
rect 4580 20244 4586 20256
rect 5169 20247 5227 20253
rect 5169 20244 5181 20247
rect 4580 20216 5181 20244
rect 4580 20204 4586 20216
rect 5169 20213 5181 20216
rect 5215 20213 5227 20247
rect 7650 20244 7656 20256
rect 7611 20216 7656 20244
rect 5169 20207 5227 20213
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9217 20247 9275 20253
rect 9217 20244 9229 20247
rect 8352 20216 9229 20244
rect 8352 20204 8358 20216
rect 9217 20213 9229 20216
rect 9263 20213 9275 20247
rect 9217 20207 9275 20213
rect 9861 20247 9919 20253
rect 9861 20213 9873 20247
rect 9907 20244 9919 20247
rect 10042 20244 10048 20256
rect 9907 20216 10048 20244
rect 9907 20213 9919 20216
rect 9861 20207 9919 20213
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 10686 20244 10692 20256
rect 10647 20216 10692 20244
rect 10686 20204 10692 20216
rect 10744 20204 10750 20256
rect 12158 20244 12164 20256
rect 12119 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 12805 20247 12863 20253
rect 12805 20244 12817 20247
rect 12676 20216 12817 20244
rect 12676 20204 12682 20216
rect 12805 20213 12817 20216
rect 12851 20244 12863 20247
rect 13170 20244 13176 20256
rect 12851 20216 13176 20244
rect 12851 20213 12863 20216
rect 12805 20207 12863 20213
rect 13170 20204 13176 20216
rect 13228 20204 13234 20256
rect 13998 20244 14004 20256
rect 13959 20216 14004 20244
rect 13998 20204 14004 20216
rect 14056 20204 14062 20256
rect 14366 20244 14372 20256
rect 14327 20216 14372 20244
rect 14366 20204 14372 20216
rect 14424 20204 14430 20256
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15252 20216 15301 20244
rect 15252 20204 15258 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 20530 20244 20536 20256
rect 20491 20216 20536 20244
rect 15289 20207 15347 20213
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 21634 20244 21640 20256
rect 21595 20216 21640 20244
rect 21634 20204 21640 20216
rect 21692 20204 21698 20256
rect 22646 20244 22652 20256
rect 22607 20216 22652 20244
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 25038 20244 25044 20256
rect 24999 20216 25044 20244
rect 25038 20204 25044 20216
rect 25096 20204 25102 20256
rect 1104 20154 26864 20176
rect 1104 20102 10315 20154
rect 10367 20102 10379 20154
rect 10431 20102 10443 20154
rect 10495 20102 10507 20154
rect 10559 20102 19648 20154
rect 19700 20102 19712 20154
rect 19764 20102 19776 20154
rect 19828 20102 19840 20154
rect 19892 20102 26864 20154
rect 1104 20080 26864 20102
rect 1118 20000 1124 20052
rect 1176 20040 1182 20052
rect 1949 20043 2007 20049
rect 1949 20040 1961 20043
rect 1176 20012 1961 20040
rect 1176 20000 1182 20012
rect 1949 20009 1961 20012
rect 1995 20040 2007 20043
rect 2314 20040 2320 20052
rect 1995 20012 2320 20040
rect 1995 20009 2007 20012
rect 1949 20003 2007 20009
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 4614 20000 4620 20052
rect 4672 20040 4678 20052
rect 5077 20043 5135 20049
rect 5077 20040 5089 20043
rect 4672 20012 5089 20040
rect 4672 20000 4678 20012
rect 5077 20009 5089 20012
rect 5123 20040 5135 20043
rect 6914 20040 6920 20052
rect 5123 20012 6920 20040
rect 5123 20009 5135 20012
rect 5077 20003 5135 20009
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7742 20000 7748 20052
rect 7800 20040 7806 20052
rect 7837 20043 7895 20049
rect 7837 20040 7849 20043
rect 7800 20012 7849 20040
rect 7800 20000 7806 20012
rect 7837 20009 7849 20012
rect 7883 20009 7895 20043
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 7837 20003 7895 20009
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 9677 20043 9735 20049
rect 9677 20009 9689 20043
rect 9723 20040 9735 20043
rect 9858 20040 9864 20052
rect 9723 20012 9864 20040
rect 9723 20009 9735 20012
rect 9677 20003 9735 20009
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 11149 20043 11207 20049
rect 11149 20009 11161 20043
rect 11195 20040 11207 20043
rect 11330 20040 11336 20052
rect 11195 20012 11336 20040
rect 11195 20009 11207 20012
rect 11149 20003 11207 20009
rect 11330 20000 11336 20012
rect 11388 20040 11394 20052
rect 11606 20040 11612 20052
rect 11388 20012 11612 20040
rect 11388 20000 11394 20012
rect 11606 20000 11612 20012
rect 11664 20000 11670 20052
rect 12529 20043 12587 20049
rect 12529 20009 12541 20043
rect 12575 20040 12587 20043
rect 12894 20040 12900 20052
rect 12575 20012 12900 20040
rect 12575 20009 12587 20012
rect 12529 20003 12587 20009
rect 12894 20000 12900 20012
rect 12952 20000 12958 20052
rect 13630 20000 13636 20052
rect 13688 20040 13694 20052
rect 14093 20043 14151 20049
rect 14093 20040 14105 20043
rect 13688 20012 14105 20040
rect 13688 20000 13694 20012
rect 14093 20009 14105 20012
rect 14139 20040 14151 20043
rect 14550 20040 14556 20052
rect 14139 20012 14556 20040
rect 14139 20009 14151 20012
rect 14093 20003 14151 20009
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15749 20043 15807 20049
rect 15749 20009 15761 20043
rect 15795 20040 15807 20043
rect 16022 20040 16028 20052
rect 15795 20012 16028 20040
rect 15795 20009 15807 20012
rect 15749 20003 15807 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 16485 20043 16543 20049
rect 16485 20009 16497 20043
rect 16531 20040 16543 20043
rect 16758 20040 16764 20052
rect 16531 20012 16764 20040
rect 16531 20009 16543 20012
rect 16485 20003 16543 20009
rect 16758 20000 16764 20012
rect 16816 20000 16822 20052
rect 18322 20000 18328 20052
rect 18380 20040 18386 20052
rect 18598 20040 18604 20052
rect 18380 20012 18604 20040
rect 18380 20000 18386 20012
rect 18598 20000 18604 20012
rect 18656 20040 18662 20052
rect 19061 20043 19119 20049
rect 19061 20040 19073 20043
rect 18656 20012 19073 20040
rect 18656 20000 18662 20012
rect 19061 20009 19073 20012
rect 19107 20040 19119 20043
rect 19334 20040 19340 20052
rect 19107 20012 19340 20040
rect 19107 20009 19119 20012
rect 19061 20003 19119 20009
rect 19334 20000 19340 20012
rect 19392 20000 19398 20052
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19613 20043 19671 20049
rect 19613 20040 19625 20043
rect 19576 20012 19625 20040
rect 19576 20000 19582 20012
rect 19613 20009 19625 20012
rect 19659 20009 19671 20043
rect 19613 20003 19671 20009
rect 20257 20043 20315 20049
rect 20257 20009 20269 20043
rect 20303 20040 20315 20043
rect 20530 20040 20536 20052
rect 20303 20012 20536 20040
rect 20303 20009 20315 20012
rect 20257 20003 20315 20009
rect 2866 19972 2872 19984
rect 2827 19944 2872 19972
rect 2866 19932 2872 19944
rect 2924 19932 2930 19984
rect 3237 19975 3295 19981
rect 3237 19941 3249 19975
rect 3283 19972 3295 19975
rect 3513 19975 3571 19981
rect 3513 19972 3525 19975
rect 3283 19944 3525 19972
rect 3283 19941 3295 19944
rect 3237 19935 3295 19941
rect 3513 19941 3525 19944
rect 3559 19972 3571 19975
rect 3970 19972 3976 19984
rect 3559 19944 3976 19972
rect 3559 19941 3571 19944
rect 3513 19935 3571 19941
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 4709 19975 4767 19981
rect 4709 19941 4721 19975
rect 4755 19972 4767 19975
rect 4798 19972 4804 19984
rect 4755 19944 4804 19972
rect 4755 19941 4767 19944
rect 4709 19935 4767 19941
rect 4798 19932 4804 19944
rect 4856 19932 4862 19984
rect 5534 19932 5540 19984
rect 5592 19972 5598 19984
rect 5782 19975 5840 19981
rect 5782 19972 5794 19975
rect 5592 19944 5794 19972
rect 5592 19932 5598 19944
rect 5782 19941 5794 19944
rect 5828 19972 5840 19975
rect 6454 19972 6460 19984
rect 5828 19944 6460 19972
rect 5828 19941 5840 19944
rect 5782 19935 5840 19941
rect 6454 19932 6460 19944
rect 6512 19932 6518 19984
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19972 8447 19975
rect 9398 19972 9404 19984
rect 8435 19944 9404 19972
rect 8435 19941 8447 19944
rect 8389 19935 8447 19941
rect 9398 19932 9404 19944
rect 9456 19932 9462 19984
rect 11072 19972 11100 20000
rect 12069 19975 12127 19981
rect 12069 19972 12081 19975
rect 11072 19944 12081 19972
rect 12069 19941 12081 19944
rect 12115 19941 12127 19975
rect 12069 19935 12127 19941
rect 12618 19932 12624 19984
rect 12676 19972 12682 19984
rect 12980 19975 13038 19981
rect 12980 19972 12992 19975
rect 12676 19944 12992 19972
rect 12676 19932 12682 19944
rect 12980 19941 12992 19944
rect 13026 19941 13038 19975
rect 12980 19935 13038 19941
rect 2777 19907 2835 19913
rect 2777 19873 2789 19907
rect 2823 19904 2835 19907
rect 3878 19904 3884 19916
rect 2823 19876 3884 19904
rect 2823 19873 2835 19876
rect 2777 19867 2835 19873
rect 3878 19864 3884 19876
rect 3936 19864 3942 19916
rect 4062 19904 4068 19916
rect 4023 19876 4068 19904
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 6270 19904 6276 19916
rect 5552 19876 6276 19904
rect 1397 19839 1455 19845
rect 1397 19805 1409 19839
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 1412 19768 1440 19799
rect 2590 19796 2596 19848
rect 2648 19836 2654 19848
rect 3053 19839 3111 19845
rect 3053 19836 3065 19839
rect 2648 19808 3065 19836
rect 2648 19796 2654 19808
rect 3053 19805 3065 19808
rect 3099 19836 3111 19839
rect 4522 19836 4528 19848
rect 3099 19808 4528 19836
rect 3099 19805 3111 19808
rect 3053 19799 3111 19805
rect 4522 19796 4528 19808
rect 4580 19796 4586 19848
rect 5552 19845 5580 19876
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 6546 19864 6552 19916
rect 6604 19904 6610 19916
rect 8754 19904 8760 19916
rect 6604 19876 8760 19904
rect 6604 19864 6610 19876
rect 8754 19864 8760 19876
rect 8812 19864 8818 19916
rect 9674 19864 9680 19916
rect 9732 19904 9738 19916
rect 10226 19904 10232 19916
rect 9732 19876 10232 19904
rect 9732 19864 9738 19876
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 11057 19907 11115 19913
rect 11057 19873 11069 19907
rect 11103 19904 11115 19907
rect 12250 19904 12256 19916
rect 11103 19876 12256 19904
rect 11103 19873 11115 19876
rect 11057 19867 11115 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12713 19907 12771 19913
rect 12713 19873 12725 19907
rect 12759 19904 12771 19907
rect 12802 19904 12808 19916
rect 12759 19876 12808 19904
rect 12759 19873 12771 19876
rect 12713 19867 12771 19873
rect 12802 19864 12808 19876
rect 12860 19864 12866 19916
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19904 15715 19907
rect 15930 19904 15936 19916
rect 15703 19876 15936 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 15930 19864 15936 19876
rect 15988 19864 15994 19916
rect 17402 19904 17408 19916
rect 17363 19876 17408 19904
rect 17402 19864 17408 19876
rect 17460 19864 17466 19916
rect 17497 19907 17555 19913
rect 17497 19873 17509 19907
rect 17543 19904 17555 19907
rect 17678 19904 17684 19916
rect 17543 19876 17684 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 17678 19864 17684 19876
rect 17736 19864 17742 19916
rect 18414 19864 18420 19916
rect 18472 19904 18478 19916
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18472 19876 18981 19904
rect 18472 19864 18478 19876
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19805 5595 19839
rect 5537 19799 5595 19805
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 7098 19836 7104 19848
rect 6880 19808 7104 19836
rect 6880 19796 6886 19808
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 8018 19836 8024 19848
rect 7607 19808 8024 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 8018 19796 8024 19808
rect 8076 19836 8082 19848
rect 8481 19839 8539 19845
rect 8481 19836 8493 19839
rect 8076 19808 8493 19836
rect 8076 19796 8082 19808
rect 8481 19805 8493 19808
rect 8527 19805 8539 19839
rect 8481 19799 8539 19805
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19805 8631 19839
rect 11330 19836 11336 19848
rect 11291 19808 11336 19836
rect 8573 19799 8631 19805
rect 3237 19771 3295 19777
rect 3237 19768 3249 19771
rect 1412 19740 3249 19768
rect 3237 19737 3249 19740
rect 3283 19737 3295 19771
rect 3237 19731 3295 19737
rect 3878 19728 3884 19780
rect 3936 19768 3942 19780
rect 3936 19740 5488 19768
rect 3936 19728 3942 19740
rect 5460 19712 5488 19740
rect 8294 19728 8300 19780
rect 8352 19768 8358 19780
rect 8588 19768 8616 19799
rect 11330 19796 11336 19808
rect 11388 19836 11394 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11388 19808 11713 19836
rect 11388 19796 11394 19808
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 15838 19836 15844 19848
rect 15799 19808 15844 19836
rect 11701 19799 11759 19805
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 17589 19839 17647 19845
rect 17589 19805 17601 19839
rect 17635 19805 17647 19839
rect 17589 19799 17647 19805
rect 10689 19771 10747 19777
rect 10689 19768 10701 19771
rect 8352 19740 8616 19768
rect 9692 19740 10701 19768
rect 8352 19728 8358 19740
rect 9692 19712 9720 19740
rect 10689 19737 10701 19740
rect 10735 19737 10747 19771
rect 10689 19731 10747 19737
rect 13814 19728 13820 19780
rect 13872 19768 13878 19780
rect 14366 19768 14372 19780
rect 13872 19740 14372 19768
rect 13872 19728 13878 19740
rect 14366 19728 14372 19740
rect 14424 19768 14430 19780
rect 14645 19771 14703 19777
rect 14645 19768 14657 19771
rect 14424 19740 14657 19768
rect 14424 19728 14430 19740
rect 14645 19737 14657 19740
rect 14691 19737 14703 19771
rect 14645 19731 14703 19737
rect 16850 19728 16856 19780
rect 16908 19768 16914 19780
rect 17604 19768 17632 19799
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19208 19808 19257 19836
rect 19208 19796 19214 19808
rect 19245 19805 19257 19808
rect 19291 19836 19303 19839
rect 20272 19836 20300 20003
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 22278 20000 22284 20052
rect 22336 20040 22342 20052
rect 22833 20043 22891 20049
rect 22833 20040 22845 20043
rect 22336 20012 22845 20040
rect 22336 20000 22342 20012
rect 22833 20009 22845 20012
rect 22879 20009 22891 20043
rect 22833 20003 22891 20009
rect 23566 19932 23572 19984
rect 23624 19981 23630 19984
rect 23624 19975 23688 19981
rect 23624 19941 23642 19975
rect 23676 19972 23688 19975
rect 24302 19972 24308 19984
rect 23676 19944 24308 19972
rect 23676 19941 23688 19944
rect 23624 19935 23688 19941
rect 23624 19932 23630 19935
rect 24302 19932 24308 19944
rect 24360 19932 24366 19984
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 21168 19907 21226 19913
rect 21168 19873 21180 19907
rect 21214 19904 21226 19907
rect 21450 19904 21456 19916
rect 21214 19876 21456 19904
rect 21214 19873 21226 19876
rect 21168 19867 21226 19873
rect 21450 19864 21456 19876
rect 21508 19864 21514 19916
rect 23382 19836 23388 19848
rect 19291 19808 20300 19836
rect 23343 19808 23388 19836
rect 19291 19805 19303 19808
rect 19245 19799 19303 19805
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 16908 19740 17632 19768
rect 18141 19771 18199 19777
rect 16908 19728 16914 19740
rect 18141 19737 18153 19771
rect 18187 19768 18199 19771
rect 18509 19771 18567 19777
rect 18509 19768 18521 19771
rect 18187 19740 18521 19768
rect 18187 19737 18199 19740
rect 18141 19731 18199 19737
rect 18509 19737 18521 19740
rect 18555 19768 18567 19771
rect 18782 19768 18788 19780
rect 18555 19740 18788 19768
rect 18555 19737 18567 19740
rect 18509 19731 18567 19737
rect 18782 19728 18788 19740
rect 18840 19768 18846 19780
rect 19168 19768 19196 19796
rect 18840 19740 19196 19768
rect 18840 19728 18846 19740
rect 22186 19728 22192 19780
rect 22244 19768 22250 19780
rect 22281 19771 22339 19777
rect 22281 19768 22293 19771
rect 22244 19740 22293 19768
rect 22244 19728 22250 19740
rect 22281 19737 22293 19740
rect 22327 19737 22339 19771
rect 22281 19731 22339 19737
rect 22370 19728 22376 19780
rect 22428 19768 22434 19780
rect 22428 19740 23428 19768
rect 22428 19728 22434 19740
rect 2314 19660 2320 19712
rect 2372 19700 2378 19712
rect 2409 19703 2467 19709
rect 2409 19700 2421 19703
rect 2372 19672 2421 19700
rect 2372 19660 2378 19672
rect 2409 19669 2421 19672
rect 2455 19669 2467 19703
rect 3786 19700 3792 19712
rect 3747 19672 3792 19700
rect 2409 19663 2467 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 4246 19700 4252 19712
rect 4207 19672 4252 19700
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 5442 19700 5448 19712
rect 5403 19672 5448 19700
rect 5442 19660 5448 19672
rect 5500 19660 5506 19712
rect 9122 19700 9128 19712
rect 9083 19672 9128 19700
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 9490 19700 9496 19712
rect 9451 19672 9496 19700
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 9674 19660 9680 19712
rect 9732 19660 9738 19712
rect 9766 19660 9772 19712
rect 9824 19700 9830 19712
rect 10321 19703 10379 19709
rect 10321 19700 10333 19703
rect 9824 19672 10333 19700
rect 9824 19660 9830 19672
rect 10321 19669 10333 19672
rect 10367 19700 10379 19703
rect 10594 19700 10600 19712
rect 10367 19672 10600 19700
rect 10367 19669 10379 19672
rect 10321 19663 10379 19669
rect 10594 19660 10600 19672
rect 10652 19660 10658 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 13078 19700 13084 19712
rect 11848 19672 13084 19700
rect 11848 19660 11854 19672
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 15289 19703 15347 19709
rect 15289 19700 15301 19703
rect 14516 19672 15301 19700
rect 14516 19660 14522 19672
rect 15289 19669 15301 19672
rect 15335 19669 15347 19703
rect 16942 19700 16948 19712
rect 16903 19672 16948 19700
rect 15289 19663 15347 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17037 19703 17095 19709
rect 17037 19669 17049 19703
rect 17083 19700 17095 19703
rect 17586 19700 17592 19712
rect 17083 19672 17592 19700
rect 17083 19669 17095 19672
rect 17037 19663 17095 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 19242 19700 19248 19712
rect 18647 19672 19248 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 19242 19660 19248 19672
rect 19300 19660 19306 19712
rect 20717 19703 20775 19709
rect 20717 19669 20729 19703
rect 20763 19700 20775 19703
rect 22002 19700 22008 19712
rect 20763 19672 22008 19700
rect 20763 19669 20775 19672
rect 20717 19663 20775 19669
rect 22002 19660 22008 19672
rect 22060 19660 22066 19712
rect 23290 19700 23296 19712
rect 23251 19672 23296 19700
rect 23290 19660 23296 19672
rect 23348 19660 23354 19712
rect 23400 19700 23428 19740
rect 24765 19703 24823 19709
rect 24765 19700 24777 19703
rect 23400 19672 24777 19700
rect 24765 19669 24777 19672
rect 24811 19669 24823 19703
rect 24765 19663 24823 19669
rect 1104 19610 26864 19632
rect 1104 19558 5648 19610
rect 5700 19558 5712 19610
rect 5764 19558 5776 19610
rect 5828 19558 5840 19610
rect 5892 19558 14982 19610
rect 15034 19558 15046 19610
rect 15098 19558 15110 19610
rect 15162 19558 15174 19610
rect 15226 19558 24315 19610
rect 24367 19558 24379 19610
rect 24431 19558 24443 19610
rect 24495 19558 24507 19610
rect 24559 19558 26864 19610
rect 1104 19536 26864 19558
rect 2866 19496 2872 19508
rect 2779 19468 2872 19496
rect 1578 19388 1584 19440
rect 1636 19428 1642 19440
rect 2038 19428 2044 19440
rect 1636 19400 2044 19428
rect 1636 19388 1642 19400
rect 2038 19388 2044 19400
rect 2096 19388 2102 19440
rect 2682 19320 2688 19372
rect 2740 19360 2746 19372
rect 2792 19360 2820 19468
rect 2866 19456 2872 19468
rect 2924 19496 2930 19508
rect 3513 19499 3571 19505
rect 3513 19496 3525 19499
rect 2924 19468 3525 19496
rect 2924 19456 2930 19468
rect 3513 19465 3525 19468
rect 3559 19465 3571 19499
rect 4062 19496 4068 19508
rect 4023 19468 4068 19496
rect 3513 19459 3571 19465
rect 4062 19456 4068 19468
rect 4120 19456 4126 19508
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 6512 19468 6561 19496
rect 6512 19456 6518 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 6549 19459 6607 19465
rect 9401 19499 9459 19505
rect 9401 19465 9413 19499
rect 9447 19496 9459 19499
rect 9490 19496 9496 19508
rect 9447 19468 9496 19496
rect 9447 19465 9459 19468
rect 9401 19459 9459 19465
rect 9490 19456 9496 19468
rect 9548 19456 9554 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 10962 19496 10968 19508
rect 10744 19468 10968 19496
rect 10744 19456 10750 19468
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11146 19456 11152 19508
rect 11204 19496 11210 19508
rect 11422 19496 11428 19508
rect 11204 19468 11428 19496
rect 11204 19456 11210 19468
rect 11422 19456 11428 19468
rect 11480 19456 11486 19508
rect 11885 19499 11943 19505
rect 11885 19465 11897 19499
rect 11931 19496 11943 19499
rect 12250 19496 12256 19508
rect 11931 19468 12256 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 12250 19456 12256 19468
rect 12308 19456 12314 19508
rect 12618 19496 12624 19508
rect 12360 19468 12624 19496
rect 3786 19428 3792 19440
rect 2740 19332 2820 19360
rect 2884 19400 3792 19428
rect 2740 19320 2746 19332
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1854 19292 1860 19304
rect 1443 19264 1860 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1854 19252 1860 19264
rect 1912 19292 1918 19304
rect 2041 19295 2099 19301
rect 2041 19292 2053 19295
rect 1912 19264 2053 19292
rect 1912 19252 1918 19264
rect 2041 19261 2053 19264
rect 2087 19292 2099 19295
rect 2130 19292 2136 19304
rect 2087 19264 2136 19292
rect 2087 19261 2099 19264
rect 2041 19255 2099 19261
rect 2130 19252 2136 19264
rect 2188 19252 2194 19304
rect 2406 19252 2412 19304
rect 2464 19292 2470 19304
rect 2884 19292 2912 19400
rect 3786 19388 3792 19400
rect 3844 19388 3850 19440
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19397 10839 19431
rect 10781 19391 10839 19397
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 3375 19332 3525 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3513 19329 3525 19332
rect 3559 19360 3571 19363
rect 3878 19360 3884 19372
rect 3559 19332 3884 19360
rect 3559 19329 3571 19332
rect 3513 19323 3571 19329
rect 3878 19320 3884 19332
rect 3936 19320 3942 19372
rect 6270 19360 6276 19372
rect 6183 19332 6276 19360
rect 3050 19292 3056 19304
rect 2464 19264 2912 19292
rect 3011 19264 3056 19292
rect 2464 19252 2470 19264
rect 3050 19252 3056 19264
rect 3108 19252 3114 19304
rect 4522 19301 4528 19304
rect 4249 19295 4307 19301
rect 4249 19261 4261 19295
rect 4295 19261 4307 19295
rect 4516 19292 4528 19301
rect 4483 19264 4528 19292
rect 4249 19255 4307 19261
rect 4516 19255 4528 19264
rect 2593 19227 2651 19233
rect 2593 19193 2605 19227
rect 2639 19224 2651 19227
rect 3068 19224 3096 19252
rect 3786 19224 3792 19236
rect 2639 19196 3096 19224
rect 3699 19196 3792 19224
rect 2639 19193 2651 19196
rect 2593 19187 2651 19193
rect 3786 19184 3792 19196
rect 3844 19224 3850 19236
rect 4264 19224 4292 19255
rect 4522 19252 4528 19255
rect 4580 19252 4586 19304
rect 6196 19224 6224 19332
rect 6270 19320 6276 19332
rect 6328 19360 6334 19372
rect 7650 19360 7656 19372
rect 6328 19332 7656 19360
rect 6328 19320 6334 19332
rect 7650 19320 7656 19332
rect 7708 19360 7714 19372
rect 7837 19363 7895 19369
rect 7837 19360 7849 19363
rect 7708 19332 7849 19360
rect 7708 19320 7714 19332
rect 7837 19329 7849 19332
rect 7883 19360 7895 19363
rect 8021 19363 8079 19369
rect 8021 19360 8033 19363
rect 7883 19332 8033 19360
rect 7883 19329 7895 19332
rect 7837 19323 7895 19329
rect 8021 19329 8033 19332
rect 8067 19329 8079 19363
rect 8021 19323 8079 19329
rect 9398 19320 9404 19372
rect 9456 19360 9462 19372
rect 9456 19332 9628 19360
rect 9456 19320 9462 19332
rect 6825 19295 6883 19301
rect 6825 19261 6837 19295
rect 6871 19292 6883 19295
rect 7006 19292 7012 19304
rect 6871 19264 7012 19292
rect 6871 19261 6883 19264
rect 6825 19255 6883 19261
rect 7006 19252 7012 19264
rect 7064 19292 7070 19304
rect 9600 19292 9628 19332
rect 10796 19292 10824 19391
rect 11606 19388 11612 19440
rect 11664 19428 11670 19440
rect 12161 19431 12219 19437
rect 12161 19428 12173 19431
rect 11664 19400 12173 19428
rect 11664 19388 11670 19400
rect 12161 19397 12173 19400
rect 12207 19397 12219 19431
rect 12161 19391 12219 19397
rect 11330 19360 11336 19372
rect 11291 19332 11336 19360
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 12360 19360 12388 19468
rect 12618 19456 12624 19468
rect 12676 19456 12682 19508
rect 14550 19496 14556 19508
rect 14511 19468 14556 19496
rect 14550 19456 14556 19468
rect 14608 19496 14614 19508
rect 14921 19499 14979 19505
rect 14921 19496 14933 19499
rect 14608 19468 14933 19496
rect 14608 19456 14614 19468
rect 14921 19465 14933 19468
rect 14967 19496 14979 19499
rect 16850 19496 16856 19508
rect 14967 19468 15148 19496
rect 16811 19468 16856 19496
rect 14967 19465 14979 19468
rect 14921 19459 14979 19465
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 12894 19428 12900 19440
rect 12492 19400 12900 19428
rect 12492 19388 12498 19400
rect 12894 19388 12900 19400
rect 12952 19388 12958 19440
rect 13078 19388 13084 19440
rect 13136 19428 13142 19440
rect 13136 19400 14964 19428
rect 13136 19388 13142 19400
rect 14936 19372 14964 19400
rect 12802 19360 12808 19372
rect 12360 19332 12572 19360
rect 12763 19332 12808 19360
rect 12544 19304 12572 19332
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13725 19363 13783 19369
rect 13725 19360 13737 19363
rect 13320 19332 13737 19360
rect 13320 19320 13326 19332
rect 13725 19329 13737 19332
rect 13771 19329 13783 19363
rect 14458 19360 14464 19372
rect 13725 19323 13783 19329
rect 14108 19332 14464 19360
rect 11238 19292 11244 19304
rect 7064 19264 7512 19292
rect 9600 19264 10824 19292
rect 11164 19264 11244 19292
rect 7064 19252 7070 19264
rect 3844 19196 6224 19224
rect 3844 19184 3850 19196
rect 1578 19156 1584 19168
rect 1539 19128 1584 19156
rect 1578 19116 1584 19128
rect 1636 19116 1642 19168
rect 2682 19156 2688 19168
rect 2643 19128 2688 19156
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3326 19156 3332 19168
rect 3191 19128 3332 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3326 19116 3332 19128
rect 3384 19116 3390 19168
rect 5626 19156 5632 19168
rect 5587 19128 5632 19156
rect 5626 19116 5632 19128
rect 5684 19116 5690 19168
rect 6196 19156 6224 19196
rect 7484 19168 7512 19264
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 8266 19227 8324 19233
rect 8266 19224 8278 19227
rect 8168 19196 8278 19224
rect 8168 19184 8174 19196
rect 8266 19193 8278 19196
rect 8312 19193 8324 19227
rect 8266 19187 8324 19193
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11164 19224 11192 19264
rect 11238 19252 11244 19264
rect 11296 19252 11302 19304
rect 12526 19252 12532 19304
rect 12584 19252 12590 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 14108 19292 14136 19332
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 14918 19320 14924 19372
rect 14976 19320 14982 19372
rect 15120 19360 15148 19468
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 20714 19456 20720 19508
rect 20772 19496 20778 19508
rect 21450 19496 21456 19508
rect 20772 19468 21456 19496
rect 20772 19456 20778 19468
rect 21450 19456 21456 19468
rect 21508 19496 21514 19508
rect 21545 19499 21603 19505
rect 21545 19496 21557 19499
rect 21508 19468 21557 19496
rect 21508 19456 21514 19468
rect 21545 19465 21557 19468
rect 21591 19465 21603 19499
rect 21545 19459 21603 19465
rect 24210 19456 24216 19508
rect 24268 19496 24274 19508
rect 24673 19499 24731 19505
rect 24673 19496 24685 19499
rect 24268 19468 24685 19496
rect 24268 19456 24274 19468
rect 24320 19440 24348 19468
rect 24673 19465 24685 19468
rect 24719 19465 24731 19499
rect 24673 19459 24731 19465
rect 20806 19388 20812 19440
rect 20864 19428 20870 19440
rect 21177 19431 21235 19437
rect 21177 19428 21189 19431
rect 20864 19400 21189 19428
rect 20864 19388 20870 19400
rect 21177 19397 21189 19400
rect 21223 19397 21235 19431
rect 21177 19391 21235 19397
rect 24302 19388 24308 19440
rect 24360 19388 24366 19440
rect 15657 19363 15715 19369
rect 15657 19360 15669 19363
rect 15120 19332 15669 19360
rect 15657 19329 15669 19332
rect 15703 19360 15715 19363
rect 15838 19360 15844 19372
rect 15703 19332 15844 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 19245 19363 19303 19369
rect 19245 19329 19257 19363
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 14274 19292 14280 19304
rect 13679 19264 14136 19292
rect 14235 19264 14280 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 14274 19252 14280 19264
rect 14332 19252 14338 19304
rect 15562 19292 15568 19304
rect 15523 19264 15568 19292
rect 15562 19252 15568 19264
rect 15620 19252 15626 19304
rect 16942 19292 16948 19304
rect 16903 19264 16948 19292
rect 16942 19252 16948 19264
rect 17000 19252 17006 19304
rect 13722 19224 13728 19236
rect 10367 19196 11192 19224
rect 13188 19196 13728 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 6270 19156 6276 19168
rect 6196 19128 6276 19156
rect 6270 19116 6276 19128
rect 6328 19116 6334 19168
rect 7006 19156 7012 19168
rect 6967 19128 7012 19156
rect 7006 19116 7012 19128
rect 7064 19116 7070 19168
rect 7466 19156 7472 19168
rect 7427 19128 7472 19156
rect 7466 19116 7472 19128
rect 7524 19116 7530 19168
rect 10689 19159 10747 19165
rect 10689 19125 10701 19159
rect 10735 19156 10747 19159
rect 11149 19159 11207 19165
rect 11149 19156 11161 19159
rect 10735 19128 11161 19156
rect 10735 19125 10747 19128
rect 10689 19119 10747 19125
rect 11149 19125 11161 19128
rect 11195 19156 11207 19159
rect 11514 19156 11520 19168
rect 11195 19128 11520 19156
rect 11195 19125 11207 19128
rect 11149 19119 11207 19125
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 13188 19165 13216 19196
rect 13722 19184 13728 19196
rect 13780 19184 13786 19236
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 14884 19196 15056 19224
rect 14884 19184 14890 19196
rect 13173 19159 13231 19165
rect 13173 19125 13185 19159
rect 13219 19125 13231 19159
rect 13538 19156 13544 19168
rect 13499 19128 13544 19156
rect 13173 19119 13231 19125
rect 13538 19116 13544 19128
rect 13596 19116 13602 19168
rect 15028 19156 15056 19196
rect 15286 19184 15292 19236
rect 15344 19224 15350 19236
rect 15473 19227 15531 19233
rect 15473 19224 15485 19227
rect 15344 19196 15485 19224
rect 15344 19184 15350 19196
rect 15473 19193 15485 19196
rect 15519 19193 15531 19227
rect 15473 19187 15531 19193
rect 17034 19184 17040 19236
rect 17092 19224 17098 19236
rect 17402 19224 17408 19236
rect 17092 19196 17408 19224
rect 17092 19184 17098 19196
rect 17402 19184 17408 19196
rect 17460 19184 17466 19236
rect 19260 19224 19288 19323
rect 20530 19320 20536 19372
rect 20588 19360 20594 19372
rect 20717 19363 20775 19369
rect 20717 19360 20729 19363
rect 20588 19332 20729 19360
rect 20588 19320 20594 19332
rect 20717 19329 20729 19332
rect 20763 19329 20775 19363
rect 20717 19323 20775 19329
rect 22370 19320 22376 19372
rect 22428 19360 22434 19372
rect 22557 19363 22615 19369
rect 22557 19360 22569 19363
rect 22428 19332 22569 19360
rect 22428 19320 22434 19332
rect 22557 19329 22569 19332
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 22646 19320 22652 19372
rect 22704 19360 22710 19372
rect 23382 19360 23388 19372
rect 22704 19332 23388 19360
rect 22704 19320 22710 19332
rect 23382 19320 23388 19332
rect 23440 19320 23446 19372
rect 24210 19360 24216 19372
rect 24171 19332 24216 19360
rect 24210 19320 24216 19332
rect 24268 19320 24274 19372
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19613 19295 19671 19301
rect 19613 19292 19625 19295
rect 19392 19264 19625 19292
rect 19392 19252 19398 19264
rect 19613 19261 19625 19264
rect 19659 19261 19671 19295
rect 19613 19255 19671 19261
rect 19978 19252 19984 19304
rect 20036 19292 20042 19304
rect 22465 19295 22523 19301
rect 20036 19264 20576 19292
rect 20036 19252 20042 19264
rect 20548 19233 20576 19264
rect 22465 19261 22477 19295
rect 22511 19292 22523 19295
rect 23290 19292 23296 19304
rect 22511 19264 23296 19292
rect 22511 19261 22523 19264
rect 22465 19255 22523 19261
rect 23290 19252 23296 19264
rect 23348 19252 23354 19304
rect 23934 19252 23940 19304
rect 23992 19292 23998 19304
rect 24121 19295 24179 19301
rect 24121 19292 24133 19295
rect 23992 19264 24133 19292
rect 23992 19252 23998 19264
rect 24121 19261 24133 19264
rect 24167 19261 24179 19295
rect 24121 19255 24179 19261
rect 25225 19295 25283 19301
rect 25225 19261 25237 19295
rect 25271 19292 25283 19295
rect 25314 19292 25320 19304
rect 25271 19264 25320 19292
rect 25271 19261 25283 19264
rect 25225 19255 25283 19261
rect 25314 19252 25320 19264
rect 25372 19292 25378 19304
rect 25777 19295 25835 19301
rect 25777 19292 25789 19295
rect 25372 19264 25789 19292
rect 25372 19252 25378 19264
rect 25777 19261 25789 19264
rect 25823 19261 25835 19295
rect 25777 19255 25835 19261
rect 20073 19227 20131 19233
rect 19260 19196 19371 19224
rect 19343 19168 19371 19196
rect 20073 19193 20085 19227
rect 20119 19224 20131 19227
rect 20533 19227 20591 19233
rect 20119 19196 20484 19224
rect 20119 19193 20131 19196
rect 20073 19187 20131 19193
rect 15105 19159 15163 19165
rect 15105 19156 15117 19159
rect 15028 19128 15117 19156
rect 15105 19125 15117 19128
rect 15151 19125 15163 19159
rect 15105 19119 15163 19125
rect 15930 19116 15936 19168
rect 15988 19156 15994 19168
rect 16117 19159 16175 19165
rect 16117 19156 16129 19159
rect 15988 19128 16129 19156
rect 15988 19116 15994 19128
rect 16117 19125 16129 19128
rect 16163 19125 16175 19159
rect 16117 19119 16175 19125
rect 17129 19159 17187 19165
rect 17129 19125 17141 19159
rect 17175 19156 17187 19159
rect 17310 19156 17316 19168
rect 17175 19128 17316 19156
rect 17175 19125 17187 19128
rect 17129 19119 17187 19125
rect 17310 19116 17316 19128
rect 17368 19116 17374 19168
rect 17678 19116 17684 19168
rect 17736 19156 17742 19168
rect 17773 19159 17831 19165
rect 17773 19156 17785 19159
rect 17736 19128 17785 19156
rect 17736 19116 17742 19128
rect 17773 19125 17785 19128
rect 17819 19125 17831 19159
rect 18414 19156 18420 19168
rect 18375 19128 18420 19156
rect 17773 19119 17831 19125
rect 18414 19116 18420 19128
rect 18472 19116 18478 19168
rect 18598 19156 18604 19168
rect 18559 19128 18604 19156
rect 18598 19116 18604 19128
rect 18656 19116 18662 19168
rect 18966 19156 18972 19168
rect 18927 19128 18972 19156
rect 18966 19116 18972 19128
rect 19024 19116 19030 19168
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19242 19156 19248 19168
rect 19107 19128 19248 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19242 19116 19248 19128
rect 19300 19116 19306 19168
rect 19334 19116 19340 19168
rect 19392 19116 19398 19168
rect 20165 19159 20223 19165
rect 20165 19125 20177 19159
rect 20211 19156 20223 19159
rect 20254 19156 20260 19168
rect 20211 19128 20260 19156
rect 20211 19125 20223 19128
rect 20165 19119 20223 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20456 19156 20484 19196
rect 20533 19193 20545 19227
rect 20579 19193 20591 19227
rect 24029 19227 24087 19233
rect 24029 19224 24041 19227
rect 20533 19187 20591 19193
rect 22020 19196 24041 19224
rect 20622 19156 20628 19168
rect 20456 19128 20628 19156
rect 20622 19116 20628 19128
rect 20680 19116 20686 19168
rect 22020 19165 22048 19196
rect 24029 19193 24041 19196
rect 24075 19224 24087 19227
rect 25041 19227 25099 19233
rect 25041 19224 25053 19227
rect 24075 19196 25053 19224
rect 24075 19193 24087 19196
rect 24029 19187 24087 19193
rect 25041 19193 25053 19196
rect 25087 19193 25099 19227
rect 25041 19187 25099 19193
rect 22005 19159 22063 19165
rect 22005 19125 22017 19159
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 22152 19128 22385 19156
rect 22152 19116 22158 19128
rect 22373 19125 22385 19128
rect 22419 19156 22431 19159
rect 22830 19156 22836 19168
rect 22419 19128 22836 19156
rect 22419 19125 22431 19128
rect 22373 19119 22431 19125
rect 22830 19116 22836 19128
rect 22888 19116 22894 19168
rect 23014 19156 23020 19168
rect 22975 19128 23020 19156
rect 23014 19116 23020 19128
rect 23072 19116 23078 19168
rect 23658 19156 23664 19168
rect 23619 19128 23664 19156
rect 23658 19116 23664 19128
rect 23716 19116 23722 19168
rect 25409 19159 25467 19165
rect 25409 19125 25421 19159
rect 25455 19156 25467 19159
rect 25498 19156 25504 19168
rect 25455 19128 25504 19156
rect 25455 19125 25467 19128
rect 25409 19119 25467 19125
rect 25498 19116 25504 19128
rect 25556 19116 25562 19168
rect 25590 19116 25596 19168
rect 25648 19156 25654 19168
rect 26326 19156 26332 19168
rect 25648 19128 26332 19156
rect 25648 19116 25654 19128
rect 26326 19116 26332 19128
rect 26384 19116 26390 19168
rect 1104 19066 26864 19088
rect 1104 19014 10315 19066
rect 10367 19014 10379 19066
rect 10431 19014 10443 19066
rect 10495 19014 10507 19066
rect 10559 19014 19648 19066
rect 19700 19014 19712 19066
rect 19764 19014 19776 19066
rect 19828 19014 19840 19066
rect 19892 19014 26864 19066
rect 1104 18992 26864 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18921 1639 18955
rect 1581 18915 1639 18921
rect 1949 18955 2007 18961
rect 1949 18921 1961 18955
rect 1995 18952 2007 18955
rect 2590 18952 2596 18964
rect 1995 18924 2596 18952
rect 1995 18921 2007 18924
rect 1949 18915 2007 18921
rect 1596 18884 1624 18915
rect 2590 18912 2596 18924
rect 2648 18912 2654 18964
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 3142 18952 3148 18964
rect 2915 18924 3148 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 3513 18955 3571 18961
rect 3513 18921 3525 18955
rect 3559 18952 3571 18955
rect 3878 18952 3884 18964
rect 3559 18924 3884 18952
rect 3559 18921 3571 18924
rect 3513 18915 3571 18921
rect 3878 18912 3884 18924
rect 3936 18912 3942 18964
rect 4522 18912 4528 18964
rect 4580 18952 4586 18964
rect 4617 18955 4675 18961
rect 4617 18952 4629 18955
rect 4580 18924 4629 18952
rect 4580 18912 4586 18924
rect 4617 18921 4629 18924
rect 4663 18921 4675 18955
rect 4617 18915 4675 18921
rect 5534 18912 5540 18964
rect 5592 18952 5598 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 5592 18924 6745 18952
rect 5592 18912 5598 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 8018 18952 8024 18964
rect 7979 18924 8024 18952
rect 6733 18915 6791 18921
rect 8018 18912 8024 18924
rect 8076 18912 8082 18964
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 9398 18912 9404 18964
rect 9456 18952 9462 18964
rect 9493 18955 9551 18961
rect 9493 18952 9505 18955
rect 9456 18924 9505 18952
rect 9456 18912 9462 18924
rect 9493 18921 9505 18924
rect 9539 18952 9551 18955
rect 9582 18952 9588 18964
rect 9539 18924 9588 18952
rect 9539 18921 9551 18924
rect 9493 18915 9551 18921
rect 9582 18912 9588 18924
rect 9640 18912 9646 18964
rect 9858 18952 9864 18964
rect 9819 18924 9864 18952
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10505 18955 10563 18961
rect 10505 18921 10517 18955
rect 10551 18952 10563 18955
rect 11330 18952 11336 18964
rect 10551 18924 11336 18952
rect 10551 18921 10563 18924
rect 10505 18915 10563 18921
rect 11330 18912 11336 18924
rect 11388 18952 11394 18964
rect 12161 18955 12219 18961
rect 12161 18952 12173 18955
rect 11388 18924 12173 18952
rect 11388 18912 11394 18924
rect 12161 18921 12173 18924
rect 12207 18921 12219 18955
rect 12161 18915 12219 18921
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12584 18924 12725 18952
rect 12584 18912 12590 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 13262 18952 13268 18964
rect 13223 18924 13268 18952
rect 12713 18915 12771 18921
rect 13262 18912 13268 18924
rect 13320 18912 13326 18964
rect 15105 18955 15163 18961
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15562 18952 15568 18964
rect 15151 18924 15568 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16022 18912 16028 18964
rect 16080 18952 16086 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 16080 18924 16129 18952
rect 16080 18912 16086 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17681 18955 17739 18961
rect 17681 18952 17693 18955
rect 17552 18924 17693 18952
rect 17552 18912 17558 18924
rect 17681 18921 17693 18924
rect 17727 18921 17739 18955
rect 17681 18915 17739 18921
rect 18506 18912 18512 18964
rect 18564 18952 18570 18964
rect 19245 18955 19303 18961
rect 19245 18952 19257 18955
rect 18564 18924 19257 18952
rect 18564 18912 18570 18924
rect 19245 18921 19257 18924
rect 19291 18952 19303 18955
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19291 18924 19809 18952
rect 19291 18921 19303 18924
rect 19245 18915 19303 18921
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 19978 18912 19984 18964
rect 20036 18952 20042 18964
rect 20165 18955 20223 18961
rect 20165 18952 20177 18955
rect 20036 18924 20177 18952
rect 20036 18912 20042 18924
rect 20165 18921 20177 18924
rect 20211 18921 20223 18955
rect 20165 18915 20223 18921
rect 20717 18955 20775 18961
rect 20717 18921 20729 18955
rect 20763 18952 20775 18955
rect 21358 18952 21364 18964
rect 20763 18924 21364 18952
rect 20763 18921 20775 18924
rect 20717 18915 20775 18921
rect 21358 18912 21364 18924
rect 21416 18952 21422 18964
rect 21453 18955 21511 18961
rect 21453 18952 21465 18955
rect 21416 18924 21465 18952
rect 21416 18912 21422 18924
rect 21453 18921 21465 18924
rect 21499 18921 21511 18955
rect 21453 18915 21511 18921
rect 22097 18955 22155 18961
rect 22097 18921 22109 18955
rect 22143 18952 22155 18955
rect 22370 18952 22376 18964
rect 22143 18924 22376 18952
rect 22143 18921 22155 18924
rect 22097 18915 22155 18921
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 23014 18912 23020 18964
rect 23072 18952 23078 18964
rect 23937 18955 23995 18961
rect 23937 18952 23949 18955
rect 23072 18924 23949 18952
rect 23072 18912 23078 18924
rect 23937 18921 23949 18924
rect 23983 18952 23995 18955
rect 24210 18952 24216 18964
rect 23983 18924 24216 18952
rect 23983 18921 23995 18924
rect 23937 18915 23995 18921
rect 24210 18912 24216 18924
rect 24268 18912 24274 18964
rect 24854 18912 24860 18964
rect 24912 18952 24918 18964
rect 25225 18955 25283 18961
rect 25225 18952 25237 18955
rect 24912 18924 25237 18952
rect 24912 18912 24918 18924
rect 25225 18921 25237 18924
rect 25271 18921 25283 18955
rect 25225 18915 25283 18921
rect 5626 18893 5632 18896
rect 5620 18884 5632 18893
rect 1596 18856 4108 18884
rect 5587 18856 5632 18884
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18785 1455 18819
rect 1397 18779 1455 18785
rect 1412 18680 1440 18779
rect 2130 18776 2136 18828
rect 2188 18816 2194 18828
rect 2777 18819 2835 18825
rect 2777 18816 2789 18819
rect 2188 18788 2789 18816
rect 2188 18776 2194 18788
rect 2777 18785 2789 18788
rect 2823 18816 2835 18819
rect 3878 18816 3884 18828
rect 2823 18788 3884 18816
rect 2823 18785 2835 18788
rect 2777 18779 2835 18785
rect 3878 18776 3884 18788
rect 3936 18776 3942 18828
rect 4080 18825 4108 18856
rect 5620 18847 5632 18856
rect 5626 18844 5632 18847
rect 5684 18844 5690 18896
rect 6270 18844 6276 18896
rect 6328 18844 6334 18896
rect 6454 18844 6460 18896
rect 6512 18884 6518 18896
rect 7469 18887 7527 18893
rect 7469 18884 7481 18887
rect 6512 18856 7481 18884
rect 6512 18844 6518 18856
rect 7469 18853 7481 18856
rect 7515 18853 7527 18887
rect 7469 18847 7527 18853
rect 4065 18819 4123 18825
rect 4065 18785 4077 18819
rect 4111 18816 4123 18819
rect 4522 18816 4528 18828
rect 4111 18788 4528 18816
rect 4111 18785 4123 18788
rect 4065 18779 4123 18785
rect 4522 18776 4528 18788
rect 4580 18776 4586 18828
rect 5353 18819 5411 18825
rect 5353 18785 5365 18819
rect 5399 18816 5411 18819
rect 6288 18816 6316 18844
rect 5399 18788 6316 18816
rect 5399 18785 5411 18788
rect 5353 18779 5411 18785
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 2280 18720 2329 18748
rect 2280 18708 2286 18720
rect 2317 18717 2329 18720
rect 2363 18748 2375 18751
rect 2406 18748 2412 18760
rect 2363 18720 2412 18748
rect 2363 18717 2375 18720
rect 2317 18711 2375 18717
rect 2406 18708 2412 18720
rect 2464 18708 2470 18760
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3234 18748 3240 18760
rect 3099 18720 3240 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 3234 18708 3240 18720
rect 3292 18708 3298 18760
rect 4154 18708 4160 18760
rect 4212 18748 4218 18760
rect 5166 18748 5172 18760
rect 4212 18720 5172 18748
rect 4212 18708 4218 18720
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 7484 18748 7512 18847
rect 7926 18844 7932 18896
rect 7984 18884 7990 18896
rect 9033 18887 9091 18893
rect 9033 18884 9045 18887
rect 7984 18856 9045 18884
rect 7984 18844 7990 18856
rect 9033 18853 9045 18856
rect 9079 18853 9091 18887
rect 9033 18847 9091 18853
rect 11048 18887 11106 18893
rect 11048 18853 11060 18887
rect 11094 18884 11106 18887
rect 11146 18884 11152 18896
rect 11094 18856 11152 18884
rect 11094 18853 11106 18856
rect 11048 18847 11106 18853
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 12894 18844 12900 18896
rect 12952 18884 12958 18896
rect 20806 18884 20812 18896
rect 12952 18856 20812 18884
rect 12952 18844 12958 18856
rect 20806 18844 20812 18856
rect 20864 18884 20870 18896
rect 21266 18884 21272 18896
rect 20864 18856 21272 18884
rect 20864 18844 20870 18856
rect 21266 18844 21272 18856
rect 21324 18884 21330 18896
rect 22388 18884 22416 18912
rect 22802 18887 22860 18893
rect 22802 18884 22814 18887
rect 21324 18856 21404 18884
rect 22388 18856 22814 18884
rect 21324 18844 21330 18856
rect 7650 18776 7656 18828
rect 7708 18816 7714 18828
rect 8389 18819 8447 18825
rect 8389 18816 8401 18819
rect 7708 18788 8401 18816
rect 7708 18776 7714 18788
rect 8389 18785 8401 18788
rect 8435 18785 8447 18819
rect 8389 18779 8447 18785
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18816 9735 18819
rect 9858 18816 9864 18828
rect 9723 18788 9864 18816
rect 9723 18785 9735 18788
rect 9677 18779 9735 18785
rect 9858 18776 9864 18788
rect 9916 18776 9922 18828
rect 10042 18776 10048 18828
rect 10100 18816 10106 18828
rect 10781 18819 10839 18825
rect 10781 18816 10793 18819
rect 10100 18788 10793 18816
rect 10100 18776 10106 18788
rect 10781 18785 10793 18788
rect 10827 18816 10839 18819
rect 11514 18816 11520 18828
rect 10827 18788 11520 18816
rect 10827 18785 10839 18788
rect 10781 18779 10839 18785
rect 11514 18776 11520 18788
rect 11572 18816 11578 18828
rect 12802 18816 12808 18828
rect 11572 18788 12808 18816
rect 11572 18776 11578 18788
rect 12802 18776 12808 18788
rect 12860 18776 12866 18828
rect 13078 18776 13084 18828
rect 13136 18816 13142 18828
rect 13725 18819 13783 18825
rect 13725 18816 13737 18819
rect 13136 18788 13737 18816
rect 13136 18776 13142 18788
rect 13725 18785 13737 18788
rect 13771 18785 13783 18819
rect 15286 18816 15292 18828
rect 15247 18788 15292 18816
rect 13725 18779 13783 18785
rect 15286 18776 15292 18788
rect 15344 18776 15350 18828
rect 15470 18776 15476 18828
rect 15528 18816 15534 18828
rect 16301 18819 16359 18825
rect 16301 18816 16313 18819
rect 15528 18788 16313 18816
rect 15528 18776 15534 18788
rect 16301 18785 16313 18788
rect 16347 18785 16359 18819
rect 16301 18779 16359 18785
rect 16568 18819 16626 18825
rect 16568 18785 16580 18819
rect 16614 18816 16626 18819
rect 17402 18816 17408 18828
rect 16614 18788 17408 18816
rect 16614 18785 16626 18788
rect 16568 18779 16626 18785
rect 17402 18776 17408 18788
rect 17460 18776 17466 18828
rect 19153 18819 19211 18825
rect 19153 18785 19165 18819
rect 19199 18816 19211 18819
rect 20254 18816 20260 18828
rect 19199 18788 20260 18816
rect 19199 18785 19211 18788
rect 19153 18779 19211 18785
rect 20254 18776 20260 18788
rect 20312 18776 20318 18828
rect 21376 18825 21404 18856
rect 22802 18853 22814 18856
rect 22848 18853 22860 18887
rect 22802 18847 22860 18853
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18785 21419 18819
rect 21361 18779 21419 18785
rect 22557 18819 22615 18825
rect 22557 18785 22569 18819
rect 22603 18816 22615 18819
rect 22646 18816 22652 18828
rect 22603 18788 22652 18816
rect 22603 18785 22615 18788
rect 22557 18779 22615 18785
rect 22646 18776 22652 18788
rect 22704 18776 22710 18828
rect 23934 18776 23940 18828
rect 23992 18816 23998 18828
rect 24489 18819 24547 18825
rect 24489 18816 24501 18819
rect 23992 18788 24501 18816
rect 23992 18776 23998 18788
rect 24489 18785 24501 18788
rect 24535 18785 24547 18819
rect 24489 18779 24547 18785
rect 24946 18776 24952 18828
rect 25004 18816 25010 18828
rect 25041 18819 25099 18825
rect 25041 18816 25053 18819
rect 25004 18788 25053 18816
rect 25004 18776 25010 18788
rect 25041 18785 25053 18788
rect 25087 18785 25099 18819
rect 25041 18779 25099 18785
rect 8294 18748 8300 18760
rect 7484 18720 8300 18748
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8570 18748 8576 18760
rect 8531 18720 8576 18748
rect 8570 18708 8576 18720
rect 8628 18748 8634 18760
rect 10229 18751 10287 18757
rect 10229 18748 10241 18751
rect 8628 18720 10241 18748
rect 8628 18708 8634 18720
rect 10229 18717 10241 18720
rect 10275 18748 10287 18751
rect 10505 18751 10563 18757
rect 10505 18748 10517 18751
rect 10275 18720 10517 18748
rect 10275 18717 10287 18720
rect 10229 18711 10287 18717
rect 10505 18717 10517 18720
rect 10551 18748 10563 18751
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10551 18720 10609 18748
rect 10551 18717 10563 18720
rect 10505 18711 10563 18717
rect 10597 18717 10609 18720
rect 10643 18717 10655 18751
rect 10597 18711 10655 18717
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 13817 18751 13875 18757
rect 13817 18748 13829 18751
rect 13688 18720 13829 18748
rect 13688 18708 13694 18720
rect 13817 18717 13829 18720
rect 13863 18717 13875 18751
rect 13817 18711 13875 18717
rect 14001 18751 14059 18757
rect 14001 18717 14013 18751
rect 14047 18748 14059 18751
rect 14550 18748 14556 18760
rect 14047 18720 14556 18748
rect 14047 18717 14059 18720
rect 14001 18711 14059 18717
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 17920 18720 18337 18748
rect 17920 18708 17926 18720
rect 18325 18717 18337 18720
rect 18371 18748 18383 18751
rect 19334 18748 19340 18760
rect 18371 18720 19340 18748
rect 18371 18717 18383 18720
rect 18325 18711 18383 18717
rect 19334 18708 19340 18720
rect 19392 18748 19398 18760
rect 19392 18720 19485 18748
rect 19392 18708 19398 18720
rect 21082 18708 21088 18760
rect 21140 18748 21146 18760
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 21140 18720 21557 18748
rect 21140 18708 21146 18720
rect 21545 18717 21557 18720
rect 21591 18748 21603 18751
rect 21818 18748 21824 18760
rect 21591 18720 21824 18748
rect 21591 18717 21603 18720
rect 21545 18711 21603 18717
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 2958 18680 2964 18692
rect 1412 18652 2964 18680
rect 2958 18640 2964 18652
rect 3016 18640 3022 18692
rect 15473 18683 15531 18689
rect 15473 18649 15485 18683
rect 15519 18680 15531 18683
rect 16114 18680 16120 18692
rect 15519 18652 16120 18680
rect 15519 18649 15531 18652
rect 15473 18643 15531 18649
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 18966 18680 18972 18692
rect 18616 18652 18972 18680
rect 2409 18615 2467 18621
rect 2409 18581 2421 18615
rect 2455 18612 2467 18615
rect 3326 18612 3332 18624
rect 2455 18584 3332 18612
rect 2455 18581 2467 18584
rect 2409 18575 2467 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 4062 18572 4068 18624
rect 4120 18612 4126 18624
rect 4249 18615 4307 18621
rect 4249 18612 4261 18615
rect 4120 18584 4261 18612
rect 4120 18572 4126 18584
rect 4249 18581 4261 18584
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8110 18612 8116 18624
rect 7975 18584 8116 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 13357 18615 13415 18621
rect 13357 18581 13369 18615
rect 13403 18612 13415 18615
rect 13538 18612 13544 18624
rect 13403 18584 13544 18612
rect 13403 18581 13415 18584
rect 13357 18575 13415 18581
rect 13538 18572 13544 18584
rect 13596 18612 13602 18624
rect 13722 18612 13728 18624
rect 13596 18584 13728 18612
rect 13596 18572 13602 18584
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14366 18612 14372 18624
rect 14327 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18572 14430 18624
rect 15838 18612 15844 18624
rect 15799 18584 15844 18612
rect 15838 18572 15844 18584
rect 15896 18572 15902 18624
rect 18506 18572 18512 18624
rect 18564 18612 18570 18624
rect 18616 18621 18644 18652
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 20993 18683 21051 18689
rect 20993 18649 21005 18683
rect 21039 18680 21051 18683
rect 21910 18680 21916 18692
rect 21039 18652 21916 18680
rect 21039 18649 21051 18652
rect 20993 18643 21051 18649
rect 21910 18640 21916 18652
rect 21968 18640 21974 18692
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18564 18584 18613 18612
rect 18564 18572 18570 18584
rect 18601 18581 18613 18584
rect 18647 18581 18659 18615
rect 18601 18575 18659 18581
rect 18785 18615 18843 18621
rect 18785 18581 18797 18615
rect 18831 18612 18843 18615
rect 19150 18612 19156 18624
rect 18831 18584 19156 18612
rect 18831 18581 18843 18584
rect 18785 18575 18843 18581
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19518 18572 19524 18624
rect 19576 18612 19582 18624
rect 21726 18612 21732 18624
rect 19576 18584 21732 18612
rect 19576 18572 19582 18584
rect 21726 18572 21732 18584
rect 21784 18572 21790 18624
rect 22186 18572 22192 18624
rect 22244 18612 22250 18624
rect 22373 18615 22431 18621
rect 22373 18612 22385 18615
rect 22244 18584 22385 18612
rect 22244 18572 22250 18584
rect 22373 18581 22385 18584
rect 22419 18581 22431 18615
rect 22373 18575 22431 18581
rect 1104 18522 26864 18544
rect 1104 18470 5648 18522
rect 5700 18470 5712 18522
rect 5764 18470 5776 18522
rect 5828 18470 5840 18522
rect 5892 18470 14982 18522
rect 15034 18470 15046 18522
rect 15098 18470 15110 18522
rect 15162 18470 15174 18522
rect 15226 18470 24315 18522
rect 24367 18470 24379 18522
rect 24431 18470 24443 18522
rect 24495 18470 24507 18522
rect 24559 18470 26864 18522
rect 1104 18448 26864 18470
rect 1765 18411 1823 18417
rect 1765 18377 1777 18411
rect 1811 18408 1823 18411
rect 3142 18408 3148 18420
rect 1811 18380 3148 18408
rect 1811 18377 1823 18380
rect 1765 18371 1823 18377
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3476 18380 3617 18408
rect 3476 18368 3482 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 4522 18408 4528 18420
rect 4483 18380 4528 18408
rect 3605 18371 3663 18377
rect 4522 18368 4528 18380
rect 4580 18368 4586 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5534 18408 5540 18420
rect 5123 18380 5540 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 2130 18340 2136 18352
rect 2091 18312 2136 18340
rect 2130 18300 2136 18312
rect 2188 18300 2194 18352
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 4249 18343 4307 18349
rect 4249 18340 4261 18343
rect 3292 18312 4261 18340
rect 3292 18300 3298 18312
rect 4249 18309 4261 18312
rect 4295 18340 4307 18343
rect 5092 18340 5120 18371
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 6270 18368 6276 18420
rect 6328 18408 6334 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6328 18380 6377 18408
rect 6328 18368 6334 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 8570 18368 8576 18420
rect 8628 18408 8634 18420
rect 8941 18411 8999 18417
rect 8941 18408 8953 18411
rect 8628 18380 8953 18408
rect 8628 18368 8634 18380
rect 8941 18377 8953 18380
rect 8987 18377 8999 18411
rect 9214 18408 9220 18420
rect 9175 18380 9220 18408
rect 8941 18371 8999 18377
rect 9214 18368 9220 18380
rect 9272 18368 9278 18420
rect 9582 18368 9588 18420
rect 9640 18408 9646 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9640 18380 10793 18408
rect 9640 18368 9646 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 11793 18411 11851 18417
rect 11793 18408 11805 18411
rect 11572 18380 11805 18408
rect 11572 18368 11578 18380
rect 11793 18377 11805 18380
rect 11839 18408 11851 18411
rect 11882 18408 11888 18420
rect 11839 18380 11888 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 11882 18368 11888 18380
rect 11940 18368 11946 18420
rect 13078 18408 13084 18420
rect 12544 18380 13084 18408
rect 4295 18312 5120 18340
rect 7101 18343 7159 18349
rect 4295 18309 4307 18312
rect 4249 18303 4307 18309
rect 7101 18309 7113 18343
rect 7147 18340 7159 18343
rect 7147 18312 8248 18340
rect 7147 18309 7159 18312
rect 7101 18303 7159 18309
rect 8220 18284 8248 18312
rect 8386 18300 8392 18352
rect 8444 18340 8450 18352
rect 8444 18312 9812 18340
rect 8444 18300 8450 18312
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 5166 18232 5172 18284
rect 5224 18272 5230 18284
rect 5721 18275 5779 18281
rect 5721 18272 5733 18275
rect 5224 18244 5733 18272
rect 5224 18232 5230 18244
rect 5721 18241 5733 18244
rect 5767 18272 5779 18275
rect 6270 18272 6276 18284
rect 5767 18244 6276 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 6270 18232 6276 18244
rect 6328 18232 6334 18284
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18272 6699 18275
rect 7834 18272 7840 18284
rect 6687 18244 7840 18272
rect 6687 18241 6699 18244
rect 6641 18235 6699 18241
rect 7834 18232 7840 18244
rect 7892 18272 7898 18284
rect 8021 18275 8079 18281
rect 8021 18272 8033 18275
rect 7892 18244 8033 18272
rect 7892 18232 7898 18244
rect 8021 18241 8033 18244
rect 8067 18241 8079 18275
rect 8202 18272 8208 18284
rect 8163 18244 8208 18272
rect 8021 18235 8079 18241
rect 8202 18232 8208 18244
rect 8260 18232 8266 18284
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8536 18244 8585 18272
rect 8536 18232 8542 18244
rect 8573 18241 8585 18244
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 9784 18281 9812 18312
rect 11146 18300 11152 18352
rect 11204 18340 11210 18352
rect 12161 18343 12219 18349
rect 12161 18340 12173 18343
rect 11204 18312 12173 18340
rect 11204 18300 11210 18312
rect 12161 18309 12173 18312
rect 12207 18309 12219 18343
rect 12161 18303 12219 18309
rect 9677 18275 9735 18281
rect 9677 18272 9689 18275
rect 9456 18244 9689 18272
rect 9456 18232 9462 18244
rect 9677 18241 9689 18244
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18241 9827 18275
rect 11330 18272 11336 18284
rect 11291 18244 11336 18272
rect 9769 18235 9827 18241
rect 11330 18232 11336 18244
rect 11388 18232 11394 18284
rect 12544 18281 12572 18380
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 13541 18411 13599 18417
rect 13541 18408 13553 18411
rect 13504 18380 13553 18408
rect 13504 18368 13510 18380
rect 13541 18377 13553 18380
rect 13587 18377 13599 18411
rect 14550 18408 14556 18420
rect 14511 18380 14556 18408
rect 13541 18371 13599 18377
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 17402 18408 17408 18420
rect 17363 18380 17408 18408
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 17862 18408 17868 18420
rect 17823 18380 17868 18408
rect 17862 18368 17868 18380
rect 17920 18368 17926 18420
rect 18601 18411 18659 18417
rect 18601 18377 18613 18411
rect 18647 18408 18659 18411
rect 18782 18408 18788 18420
rect 18647 18380 18788 18408
rect 18647 18377 18659 18380
rect 18601 18371 18659 18377
rect 18782 18368 18788 18380
rect 18840 18368 18846 18420
rect 19334 18368 19340 18420
rect 19392 18408 19398 18420
rect 19702 18408 19708 18420
rect 19392 18380 19708 18408
rect 19392 18368 19398 18380
rect 19702 18368 19708 18380
rect 19760 18408 19766 18420
rect 20441 18411 20499 18417
rect 20441 18408 20453 18411
rect 19760 18380 20453 18408
rect 19760 18368 19766 18380
rect 20441 18377 20453 18380
rect 20487 18377 20499 18411
rect 20441 18371 20499 18377
rect 20806 18368 20812 18420
rect 20864 18408 20870 18420
rect 20993 18411 21051 18417
rect 20993 18408 21005 18411
rect 20864 18380 21005 18408
rect 20864 18368 20870 18380
rect 20993 18377 21005 18380
rect 21039 18377 21051 18411
rect 21358 18408 21364 18420
rect 21319 18380 21364 18408
rect 20993 18371 21051 18377
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 23290 18368 23296 18420
rect 23348 18408 23354 18420
rect 23661 18411 23719 18417
rect 23661 18408 23673 18411
rect 23348 18380 23673 18408
rect 23348 18368 23354 18380
rect 23661 18377 23673 18380
rect 23707 18377 23719 18411
rect 23661 18371 23719 18377
rect 24210 18368 24216 18420
rect 24268 18408 24274 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 24268 18380 24685 18408
rect 24268 18368 24274 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 24673 18371 24731 18377
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 25041 18411 25099 18417
rect 25041 18408 25053 18411
rect 25004 18380 25053 18408
rect 25004 18368 25010 18380
rect 25041 18377 25053 18380
rect 25087 18377 25099 18411
rect 25406 18408 25412 18420
rect 25367 18380 25412 18408
rect 25041 18371 25099 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 13078 18272 13084 18284
rect 12952 18244 13084 18272
rect 12952 18232 12958 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13998 18232 14004 18284
rect 14056 18272 14062 18284
rect 14185 18275 14243 18281
rect 14185 18272 14197 18275
rect 14056 18244 14197 18272
rect 14056 18232 14062 18244
rect 14185 18241 14197 18244
rect 14231 18272 14243 18275
rect 14568 18272 14596 18368
rect 16114 18300 16120 18352
rect 16172 18340 16178 18352
rect 16482 18340 16488 18352
rect 16172 18312 16488 18340
rect 16172 18300 16178 18312
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 14231 18244 14596 18272
rect 17972 18244 18184 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 2492 18207 2550 18213
rect 2492 18173 2504 18207
rect 2538 18204 2550 18207
rect 2866 18204 2872 18216
rect 2538 18176 2872 18204
rect 2538 18173 2550 18176
rect 2492 18167 2550 18173
rect 2866 18164 2872 18176
rect 2924 18164 2930 18216
rect 7469 18207 7527 18213
rect 7469 18173 7481 18207
rect 7515 18204 7527 18207
rect 7650 18204 7656 18216
rect 7515 18176 7656 18204
rect 7515 18173 7527 18176
rect 7469 18167 7527 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7926 18204 7932 18216
rect 7887 18176 7932 18204
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9122 18164 9128 18216
rect 9180 18204 9186 18216
rect 9582 18204 9588 18216
rect 9180 18176 9588 18204
rect 9180 18164 9186 18176
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9858 18164 9864 18216
rect 9916 18204 9922 18216
rect 10321 18207 10379 18213
rect 10321 18204 10333 18207
rect 9916 18176 10333 18204
rect 9916 18164 9922 18176
rect 10321 18173 10333 18176
rect 10367 18204 10379 18207
rect 10962 18204 10968 18216
rect 10367 18176 10968 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 13354 18204 13360 18216
rect 11572 18176 13360 18204
rect 11572 18164 11578 18176
rect 13354 18164 13360 18176
rect 13412 18164 13418 18216
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18204 13967 18207
rect 14274 18204 14280 18216
rect 13955 18176 14280 18204
rect 13955 18173 13967 18176
rect 13909 18167 13967 18173
rect 14274 18164 14280 18176
rect 14332 18164 14338 18216
rect 15102 18204 15108 18216
rect 14936 18176 15108 18204
rect 5534 18136 5540 18148
rect 5495 18108 5540 18136
rect 5534 18096 5540 18108
rect 5592 18096 5598 18148
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 11149 18139 11207 18145
rect 11149 18136 11161 18139
rect 10928 18108 11161 18136
rect 10928 18096 10934 18108
rect 11072 18080 11100 18108
rect 11149 18105 11161 18108
rect 11195 18105 11207 18139
rect 11149 18099 11207 18105
rect 12802 18096 12808 18148
rect 12860 18136 12866 18148
rect 14001 18139 14059 18145
rect 12860 18108 13952 18136
rect 12860 18096 12866 18108
rect 5166 18068 5172 18080
rect 5127 18040 5172 18068
rect 5166 18028 5172 18040
rect 5224 18028 5230 18080
rect 5626 18068 5632 18080
rect 5587 18040 5632 18068
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 6273 18071 6331 18077
rect 6273 18037 6285 18071
rect 6319 18068 6331 18071
rect 6365 18071 6423 18077
rect 6365 18068 6377 18071
rect 6319 18040 6377 18068
rect 6319 18037 6331 18040
rect 6273 18031 6331 18037
rect 6365 18037 6377 18040
rect 6411 18068 6423 18071
rect 6638 18068 6644 18080
rect 6411 18040 6644 18068
rect 6411 18037 6423 18040
rect 6365 18031 6423 18037
rect 6638 18028 6644 18040
rect 6696 18028 6702 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 7561 18071 7619 18077
rect 7561 18068 7573 18071
rect 7524 18040 7573 18068
rect 7524 18028 7530 18040
rect 7561 18037 7573 18040
rect 7607 18037 7619 18071
rect 7561 18031 7619 18037
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 11054 18068 11060 18080
rect 10735 18040 11060 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11054 18028 11060 18040
rect 11112 18028 11118 18080
rect 11238 18068 11244 18080
rect 11199 18040 11244 18068
rect 11238 18028 11244 18040
rect 11296 18028 11302 18080
rect 13354 18068 13360 18080
rect 13315 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18068 13418 18080
rect 13630 18068 13636 18080
rect 13412 18040 13636 18068
rect 13412 18028 13418 18040
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 13924 18068 13952 18108
rect 14001 18105 14013 18139
rect 14047 18136 14059 18139
rect 14090 18136 14096 18148
rect 14047 18108 14096 18136
rect 14047 18105 14059 18108
rect 14001 18099 14059 18105
rect 14090 18096 14096 18108
rect 14148 18096 14154 18148
rect 14936 18077 14964 18176
rect 15102 18164 15108 18176
rect 15160 18164 15166 18216
rect 15372 18207 15430 18213
rect 15372 18173 15384 18207
rect 15418 18204 15430 18207
rect 15838 18204 15844 18216
rect 15418 18176 15844 18204
rect 15418 18173 15430 18176
rect 15372 18167 15430 18173
rect 15838 18164 15844 18176
rect 15896 18164 15902 18216
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 13924 18040 14933 18068
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 14921 18031 14979 18037
rect 15470 18028 15476 18080
rect 15528 18068 15534 18080
rect 17037 18071 17095 18077
rect 17037 18068 17049 18071
rect 15528 18040 17049 18068
rect 15528 18028 15534 18040
rect 17037 18037 17049 18040
rect 17083 18068 17095 18071
rect 17972 18068 18000 18244
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18173 18107 18207
rect 18156 18204 18184 18244
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18414 18272 18420 18284
rect 18288 18244 18420 18272
rect 18288 18232 18294 18244
rect 18414 18232 18420 18244
rect 18472 18232 18478 18284
rect 18800 18272 18828 18368
rect 23477 18343 23535 18349
rect 23477 18309 23489 18343
rect 23523 18340 23535 18343
rect 23566 18340 23572 18352
rect 23523 18312 23572 18340
rect 23523 18309 23535 18312
rect 23477 18303 23535 18309
rect 23566 18300 23572 18312
rect 23624 18300 23630 18352
rect 22186 18272 22192 18284
rect 18800 18244 19196 18272
rect 22147 18244 22192 18272
rect 18877 18207 18935 18213
rect 18877 18204 18889 18207
rect 18156 18176 18889 18204
rect 18049 18167 18107 18173
rect 18877 18173 18889 18176
rect 18923 18204 18935 18207
rect 19061 18207 19119 18213
rect 19061 18204 19073 18207
rect 18923 18176 19073 18204
rect 18923 18173 18935 18176
rect 18877 18167 18935 18173
rect 19061 18173 19073 18176
rect 19107 18173 19119 18207
rect 19168 18204 19196 18244
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 23109 18275 23167 18281
rect 23109 18241 23121 18275
rect 23155 18272 23167 18275
rect 23842 18272 23848 18284
rect 23155 18244 23848 18272
rect 23155 18241 23167 18244
rect 23109 18235 23167 18241
rect 23842 18232 23848 18244
rect 23900 18272 23906 18284
rect 24228 18281 24256 18368
rect 24121 18275 24179 18281
rect 24121 18272 24133 18275
rect 23900 18244 24133 18272
rect 23900 18232 23906 18244
rect 24121 18241 24133 18244
rect 24167 18241 24179 18275
rect 24121 18235 24179 18241
rect 24213 18275 24271 18281
rect 24213 18241 24225 18275
rect 24259 18241 24271 18275
rect 24213 18235 24271 18241
rect 19317 18207 19375 18213
rect 19317 18204 19329 18207
rect 19168 18176 19329 18204
rect 19061 18167 19119 18173
rect 19317 18173 19329 18176
rect 19363 18173 19375 18207
rect 19702 18204 19708 18216
rect 19317 18167 19375 18173
rect 19444 18176 19708 18204
rect 18064 18136 18092 18167
rect 18966 18136 18972 18148
rect 18064 18108 18972 18136
rect 18966 18096 18972 18108
rect 19024 18096 19030 18148
rect 18046 18068 18052 18080
rect 17083 18040 18052 18068
rect 17083 18037 17095 18040
rect 17037 18031 17095 18037
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18230 18068 18236 18080
rect 18191 18040 18236 18068
rect 18230 18028 18236 18040
rect 18288 18028 18294 18080
rect 19334 18028 19340 18080
rect 19392 18068 19398 18080
rect 19444 18068 19472 18176
rect 19702 18164 19708 18176
rect 19760 18164 19766 18216
rect 21358 18164 21364 18216
rect 21416 18204 21422 18216
rect 21913 18207 21971 18213
rect 21913 18204 21925 18207
rect 21416 18176 21925 18204
rect 21416 18164 21422 18176
rect 21913 18173 21925 18176
rect 21959 18173 21971 18207
rect 21913 18167 21971 18173
rect 23566 18164 23572 18216
rect 23624 18204 23630 18216
rect 24029 18207 24087 18213
rect 24029 18204 24041 18207
rect 23624 18176 24041 18204
rect 23624 18164 23630 18176
rect 24029 18173 24041 18176
rect 24075 18173 24087 18207
rect 25222 18204 25228 18216
rect 25183 18176 25228 18204
rect 24029 18167 24087 18173
rect 25222 18164 25228 18176
rect 25280 18204 25286 18216
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25280 18176 25789 18204
rect 25280 18164 25286 18176
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 19610 18096 19616 18148
rect 19668 18136 19674 18148
rect 21266 18136 21272 18148
rect 19668 18108 21272 18136
rect 19668 18096 19674 18108
rect 21266 18096 21272 18108
rect 21324 18096 21330 18148
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 25314 18136 25320 18148
rect 21876 18108 25320 18136
rect 21876 18096 21882 18108
rect 25314 18096 25320 18108
rect 25372 18096 25378 18148
rect 19392 18040 19472 18068
rect 19392 18028 19398 18040
rect 19518 18028 19524 18080
rect 19576 18068 19582 18080
rect 20806 18068 20812 18080
rect 19576 18040 20812 18068
rect 19576 18028 19582 18040
rect 20806 18028 20812 18040
rect 20864 18028 20870 18080
rect 21542 18068 21548 18080
rect 21503 18040 21548 18068
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 21634 18028 21640 18080
rect 21692 18068 21698 18080
rect 22002 18068 22008 18080
rect 21692 18040 22008 18068
rect 21692 18028 21698 18040
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 22649 18071 22707 18077
rect 22649 18037 22661 18071
rect 22695 18068 22707 18071
rect 22738 18068 22744 18080
rect 22695 18040 22744 18068
rect 22695 18037 22707 18040
rect 22649 18031 22707 18037
rect 22738 18028 22744 18040
rect 22796 18028 22802 18080
rect 1104 17978 26864 18000
rect 1104 17926 10315 17978
rect 10367 17926 10379 17978
rect 10431 17926 10443 17978
rect 10495 17926 10507 17978
rect 10559 17926 19648 17978
rect 19700 17926 19712 17978
rect 19764 17926 19776 17978
rect 19828 17926 19840 17978
rect 19892 17926 26864 17978
rect 1104 17904 26864 17926
rect 2958 17824 2964 17876
rect 3016 17864 3022 17876
rect 3878 17864 3884 17876
rect 3016 17836 3884 17864
rect 3016 17824 3022 17836
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4893 17867 4951 17873
rect 4893 17833 4905 17867
rect 4939 17864 4951 17867
rect 5442 17864 5448 17876
rect 4939 17836 5448 17864
rect 4939 17833 4951 17836
rect 4893 17827 4951 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 6270 17864 6276 17876
rect 6231 17836 6276 17864
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 7929 17867 7987 17873
rect 7929 17833 7941 17867
rect 7975 17864 7987 17867
rect 8481 17867 8539 17873
rect 8481 17864 8493 17867
rect 7975 17836 8493 17864
rect 7975 17833 7987 17836
rect 7929 17827 7987 17833
rect 8481 17833 8493 17836
rect 8527 17864 8539 17867
rect 9677 17867 9735 17873
rect 9677 17864 9689 17867
rect 8527 17836 9689 17864
rect 8527 17833 8539 17836
rect 8481 17827 8539 17833
rect 9677 17833 9689 17836
rect 9723 17833 9735 17867
rect 10870 17864 10876 17876
rect 10831 17836 10876 17864
rect 9677 17827 9735 17833
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11480 17836 13768 17864
rect 11480 17824 11486 17836
rect 1756 17799 1814 17805
rect 1756 17765 1768 17799
rect 1802 17796 1814 17799
rect 1802 17768 2820 17796
rect 1802 17765 1814 17768
rect 1756 17759 1814 17765
rect 1489 17731 1547 17737
rect 1489 17697 1501 17731
rect 1535 17728 1547 17731
rect 2222 17728 2228 17740
rect 1535 17700 2228 17728
rect 1535 17697 1547 17700
rect 1489 17691 1547 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 2792 17728 2820 17768
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 2924 17768 3433 17796
rect 2924 17756 2930 17768
rect 3421 17765 3433 17768
rect 3467 17765 3479 17799
rect 3421 17759 3479 17765
rect 5350 17756 5356 17808
rect 5408 17796 5414 17808
rect 6546 17796 6552 17808
rect 5408 17768 6552 17796
rect 5408 17756 5414 17768
rect 6546 17756 6552 17768
rect 6604 17756 6610 17808
rect 8754 17756 8760 17808
rect 8812 17796 8818 17808
rect 9030 17796 9036 17808
rect 8812 17768 9036 17796
rect 8812 17756 8818 17768
rect 9030 17756 9036 17768
rect 9088 17756 9094 17808
rect 11609 17799 11667 17805
rect 11609 17765 11621 17799
rect 11655 17796 11667 17799
rect 12526 17796 12532 17808
rect 11655 17768 12532 17796
rect 11655 17765 11667 17768
rect 11609 17759 11667 17765
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 13740 17796 13768 17836
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 14921 17867 14979 17873
rect 14921 17864 14933 17867
rect 13872 17836 14933 17864
rect 13872 17824 13878 17836
rect 14921 17833 14933 17836
rect 14967 17833 14979 17867
rect 17586 17864 17592 17876
rect 17547 17836 17592 17864
rect 14921 17827 14979 17833
rect 17586 17824 17592 17836
rect 17644 17824 17650 17876
rect 17954 17864 17960 17876
rect 17915 17836 17960 17864
rect 17954 17824 17960 17836
rect 18012 17824 18018 17876
rect 19705 17867 19763 17873
rect 19705 17833 19717 17867
rect 19751 17833 19763 17867
rect 20254 17864 20260 17876
rect 20215 17836 20260 17864
rect 19705 17827 19763 17833
rect 13909 17799 13967 17805
rect 13740 17768 13860 17796
rect 4798 17728 4804 17740
rect 2792 17700 3464 17728
rect 4759 17700 4804 17728
rect 3436 17672 3464 17700
rect 4798 17688 4804 17700
rect 4856 17728 4862 17740
rect 5261 17731 5319 17737
rect 5261 17728 5273 17731
rect 4856 17700 5273 17728
rect 4856 17688 4862 17700
rect 5261 17697 5273 17700
rect 5307 17697 5319 17731
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 5261 17691 5319 17697
rect 6564 17700 6837 17728
rect 6564 17672 6592 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 6825 17691 6883 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8352 17700 8401 17728
rect 8352 17688 8358 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9732 17700 10057 17728
rect 9732 17688 9738 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 11701 17731 11759 17737
rect 11701 17697 11713 17731
rect 11747 17728 11759 17731
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11747 17700 12265 17728
rect 11747 17697 11759 17700
rect 11701 17691 11759 17697
rect 12253 17697 12265 17700
rect 12299 17728 12311 17731
rect 12802 17728 12808 17740
rect 12299 17700 12808 17728
rect 12299 17697 12311 17700
rect 12253 17691 12311 17697
rect 12802 17688 12808 17700
rect 12860 17688 12866 17740
rect 13173 17731 13231 17737
rect 13173 17697 13185 17731
rect 13219 17728 13231 17731
rect 13832 17728 13860 17768
rect 13909 17765 13921 17799
rect 13955 17796 13967 17799
rect 13998 17796 14004 17808
rect 13955 17768 14004 17796
rect 13955 17765 13967 17768
rect 13909 17759 13967 17765
rect 13998 17756 14004 17768
rect 14056 17756 14062 17808
rect 14090 17756 14096 17808
rect 14148 17796 14154 17808
rect 15562 17805 15568 17808
rect 14553 17799 14611 17805
rect 14553 17796 14565 17799
rect 14148 17768 14565 17796
rect 14148 17756 14154 17768
rect 14553 17765 14565 17768
rect 14599 17765 14611 17799
rect 15556 17796 15568 17805
rect 15475 17768 15568 17796
rect 14553 17759 14611 17765
rect 15556 17759 15568 17768
rect 15620 17796 15626 17808
rect 16022 17796 16028 17808
rect 15620 17768 16028 17796
rect 15562 17756 15568 17759
rect 15620 17756 15626 17768
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 18141 17799 18199 17805
rect 18141 17765 18153 17799
rect 18187 17796 18199 17799
rect 19720 17796 19748 17827
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 20717 17867 20775 17873
rect 20717 17833 20729 17867
rect 20763 17864 20775 17867
rect 21082 17864 21088 17876
rect 20763 17836 21088 17864
rect 20763 17833 20775 17836
rect 20717 17827 20775 17833
rect 21082 17824 21088 17836
rect 21140 17824 21146 17876
rect 22370 17824 22376 17876
rect 22428 17864 22434 17876
rect 22557 17867 22615 17873
rect 22557 17864 22569 17867
rect 22428 17836 22569 17864
rect 22428 17824 22434 17836
rect 22557 17833 22569 17836
rect 22603 17833 22615 17867
rect 22557 17827 22615 17833
rect 24854 17824 24860 17876
rect 24912 17864 24918 17876
rect 25409 17867 25467 17873
rect 25409 17864 25421 17867
rect 24912 17836 25421 17864
rect 24912 17824 24918 17836
rect 25409 17833 25421 17836
rect 25455 17833 25467 17867
rect 25409 17827 25467 17833
rect 20622 17796 20628 17808
rect 18187 17768 18736 17796
rect 19720 17768 20628 17796
rect 18187 17765 18199 17768
rect 18141 17759 18199 17765
rect 13219 17700 13768 17728
rect 13832 17700 17816 17728
rect 13219 17697 13231 17700
rect 13173 17691 13231 17697
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 5074 17620 5080 17672
rect 5132 17660 5138 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 5132 17632 5365 17660
rect 5132 17620 5138 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 5445 17663 5503 17669
rect 5445 17629 5457 17663
rect 5491 17629 5503 17663
rect 5445 17623 5503 17629
rect 4433 17595 4491 17601
rect 4433 17561 4445 17595
rect 4479 17592 4491 17595
rect 5460 17592 5488 17623
rect 6546 17620 6552 17672
rect 6604 17620 6610 17672
rect 6914 17660 6920 17672
rect 6875 17632 6920 17660
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17629 7067 17663
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 7009 17623 7067 17629
rect 5534 17592 5540 17604
rect 4479 17564 5540 17592
rect 4479 17561 4491 17564
rect 4433 17555 4491 17561
rect 5534 17552 5540 17564
rect 5592 17592 5598 17604
rect 5905 17595 5963 17601
rect 5905 17592 5917 17595
rect 5592 17564 5917 17592
rect 5592 17552 5598 17564
rect 5905 17561 5917 17564
rect 5951 17592 5963 17595
rect 7024 17592 7052 17623
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 9030 17620 9036 17672
rect 9088 17660 9094 17672
rect 10137 17663 10195 17669
rect 10137 17660 10149 17663
rect 9088 17632 10149 17660
rect 9088 17620 9094 17632
rect 10137 17629 10149 17632
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 10226 17620 10232 17672
rect 10284 17660 10290 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 10284 17632 10329 17660
rect 11716 17632 11805 17660
rect 10284 17620 10290 17632
rect 11716 17604 11744 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 13262 17660 13268 17672
rect 13223 17632 13268 17660
rect 11793 17623 11851 17629
rect 13262 17620 13268 17632
rect 13320 17620 13326 17672
rect 13449 17663 13507 17669
rect 13449 17629 13461 17663
rect 13495 17660 13507 17663
rect 13630 17660 13636 17672
rect 13495 17632 13636 17660
rect 13495 17629 13507 17632
rect 13449 17623 13507 17629
rect 13630 17620 13636 17632
rect 13688 17620 13694 17672
rect 13740 17660 13768 17700
rect 13998 17660 14004 17672
rect 13740 17632 14004 17660
rect 13998 17620 14004 17632
rect 14056 17620 14062 17672
rect 15102 17620 15108 17672
rect 15160 17660 15166 17672
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15160 17632 15301 17660
rect 15160 17620 15166 17632
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 5951 17564 7052 17592
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 8386 17552 8392 17604
rect 8444 17592 8450 17604
rect 9217 17595 9275 17601
rect 9217 17592 9229 17595
rect 8444 17564 9229 17592
rect 8444 17552 8450 17564
rect 9217 17561 9229 17564
rect 9263 17561 9275 17595
rect 9217 17555 9275 17561
rect 11698 17552 11704 17604
rect 11756 17552 11762 17604
rect 12066 17552 12072 17604
rect 12124 17592 12130 17604
rect 14185 17595 14243 17601
rect 14185 17592 14197 17595
rect 12124 17564 14197 17592
rect 12124 17552 12130 17564
rect 14185 17561 14197 17564
rect 14231 17561 14243 17595
rect 14185 17555 14243 17561
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 6454 17524 6460 17536
rect 6415 17496 6460 17524
rect 6454 17484 6460 17496
rect 6512 17484 6518 17536
rect 6638 17484 6644 17536
rect 6696 17524 6702 17536
rect 7469 17527 7527 17533
rect 7469 17524 7481 17527
rect 6696 17496 7481 17524
rect 6696 17484 6702 17496
rect 7469 17493 7481 17496
rect 7515 17493 7527 17527
rect 8018 17524 8024 17536
rect 7979 17496 8024 17524
rect 7469 17487 7527 17493
rect 8018 17484 8024 17496
rect 8076 17484 8082 17536
rect 11238 17524 11244 17536
rect 11199 17496 11244 17524
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 12526 17484 12532 17536
rect 12584 17524 12590 17536
rect 12621 17527 12679 17533
rect 12621 17524 12633 17527
rect 12584 17496 12633 17524
rect 12584 17484 12590 17496
rect 12621 17493 12633 17496
rect 12667 17493 12679 17527
rect 12621 17487 12679 17493
rect 12805 17527 12863 17533
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 14090 17524 14096 17536
rect 12851 17496 14096 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 15304 17524 15332 17623
rect 17788 17592 17816 17700
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 18581 17731 18639 17737
rect 18581 17728 18593 17731
rect 17920 17700 18593 17728
rect 17920 17688 17926 17700
rect 18581 17697 18593 17700
rect 18627 17697 18639 17731
rect 18708 17728 18736 17768
rect 20622 17756 20628 17768
rect 20680 17756 20686 17808
rect 21266 17796 21272 17808
rect 21179 17768 21272 17796
rect 21266 17756 21272 17768
rect 21324 17796 21330 17808
rect 22830 17796 22836 17808
rect 21324 17768 22836 17796
rect 21324 17756 21330 17768
rect 22830 17756 22836 17768
rect 22888 17756 22894 17808
rect 23198 17756 23204 17808
rect 23256 17796 23262 17808
rect 23382 17796 23388 17808
rect 23256 17768 23388 17796
rect 23256 17756 23262 17768
rect 23382 17756 23388 17768
rect 23440 17756 23446 17808
rect 25038 17796 25044 17808
rect 24999 17768 25044 17796
rect 25038 17756 25044 17768
rect 25096 17756 25102 17808
rect 20714 17728 20720 17740
rect 18708 17700 20720 17728
rect 18581 17691 18639 17697
rect 20714 17688 20720 17700
rect 20772 17688 20778 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21082 17728 21088 17740
rect 20956 17700 21088 17728
rect 20956 17688 20962 17700
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 22646 17688 22652 17740
rect 22704 17728 22710 17740
rect 23014 17737 23020 17740
rect 22997 17731 23020 17737
rect 22997 17728 23009 17731
rect 22704 17700 23009 17728
rect 22704 17688 22710 17700
rect 22997 17697 23009 17700
rect 23072 17728 23078 17740
rect 23072 17700 23145 17728
rect 22997 17691 23020 17697
rect 23014 17688 23020 17691
rect 23072 17688 23078 17700
rect 25130 17688 25136 17740
rect 25188 17728 25194 17740
rect 25225 17731 25283 17737
rect 25225 17728 25237 17731
rect 25188 17700 25237 17728
rect 25188 17688 25194 17700
rect 25225 17697 25237 17700
rect 25271 17728 25283 17731
rect 25774 17728 25780 17740
rect 25271 17700 25780 17728
rect 25271 17697 25283 17700
rect 25225 17691 25283 17697
rect 25774 17688 25780 17700
rect 25832 17688 25838 17740
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18104 17632 18337 17660
rect 18104 17620 18110 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20312 17632 21373 17660
rect 20312 17620 20318 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17629 21511 17663
rect 22738 17660 22744 17672
rect 22699 17632 22744 17660
rect 21453 17623 21511 17629
rect 18141 17595 18199 17601
rect 18141 17592 18153 17595
rect 17788 17564 18153 17592
rect 18141 17561 18153 17564
rect 18187 17561 18199 17595
rect 18141 17555 18199 17561
rect 20714 17552 20720 17604
rect 20772 17592 20778 17604
rect 21468 17592 21496 17623
rect 22738 17620 22744 17632
rect 22796 17620 22802 17672
rect 20772 17564 21496 17592
rect 20772 17552 20778 17564
rect 23750 17552 23756 17604
rect 23808 17592 23814 17604
rect 24673 17595 24731 17601
rect 24673 17592 24685 17595
rect 23808 17564 24685 17592
rect 23808 17552 23814 17564
rect 24673 17561 24685 17564
rect 24719 17561 24731 17595
rect 24673 17555 24731 17561
rect 15470 17524 15476 17536
rect 15304 17496 15476 17524
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 17313 17527 17371 17533
rect 17313 17493 17325 17527
rect 17359 17524 17371 17527
rect 17586 17524 17592 17536
rect 17359 17496 17592 17524
rect 17359 17493 17371 17496
rect 17313 17487 17371 17493
rect 17586 17484 17592 17496
rect 17644 17484 17650 17536
rect 20898 17524 20904 17536
rect 20859 17496 20904 17524
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 21542 17484 21548 17536
rect 21600 17524 21606 17536
rect 21913 17527 21971 17533
rect 21913 17524 21925 17527
rect 21600 17496 21925 17524
rect 21600 17484 21606 17496
rect 21913 17493 21925 17496
rect 21959 17524 21971 17527
rect 22002 17524 22008 17536
rect 21959 17496 22008 17524
rect 21959 17493 21971 17496
rect 21913 17487 21971 17493
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 22186 17484 22192 17536
rect 22244 17524 22250 17536
rect 24121 17527 24179 17533
rect 24121 17524 24133 17527
rect 22244 17496 24133 17524
rect 22244 17484 22250 17496
rect 24121 17493 24133 17496
rect 24167 17493 24179 17527
rect 24121 17487 24179 17493
rect 25774 17484 25780 17536
rect 25832 17524 25838 17536
rect 25958 17524 25964 17536
rect 25832 17496 25964 17524
rect 25832 17484 25838 17496
rect 25958 17484 25964 17496
rect 26016 17484 26022 17536
rect 1104 17434 26864 17456
rect 1104 17382 5648 17434
rect 5700 17382 5712 17434
rect 5764 17382 5776 17434
rect 5828 17382 5840 17434
rect 5892 17382 14982 17434
rect 15034 17382 15046 17434
rect 15098 17382 15110 17434
rect 15162 17382 15174 17434
rect 15226 17382 24315 17434
rect 24367 17382 24379 17434
rect 24431 17382 24443 17434
rect 24495 17382 24507 17434
rect 24559 17382 26864 17434
rect 1104 17360 26864 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 2041 17323 2099 17329
rect 2041 17320 2053 17323
rect 1719 17292 2053 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 2041 17289 2053 17292
rect 2087 17320 2099 17323
rect 2130 17320 2136 17332
rect 2087 17292 2136 17320
rect 2087 17289 2099 17292
rect 2041 17283 2099 17289
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 3510 17280 3516 17332
rect 3568 17320 3574 17332
rect 4249 17323 4307 17329
rect 4249 17320 4261 17323
rect 3568 17292 4261 17320
rect 3568 17280 3574 17292
rect 4249 17289 4261 17292
rect 4295 17320 4307 17323
rect 5074 17320 5080 17332
rect 4295 17292 5080 17320
rect 4295 17289 4307 17292
rect 4249 17283 4307 17289
rect 5074 17280 5080 17292
rect 5132 17280 5138 17332
rect 5169 17323 5227 17329
rect 5169 17289 5181 17323
rect 5215 17320 5227 17323
rect 5442 17320 5448 17332
rect 5215 17292 5448 17320
rect 5215 17289 5227 17292
rect 5169 17283 5227 17289
rect 5442 17280 5448 17292
rect 5500 17280 5506 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 8757 17323 8815 17329
rect 8757 17320 8769 17323
rect 8720 17292 8769 17320
rect 8720 17280 8726 17292
rect 8757 17289 8769 17292
rect 8803 17289 8815 17323
rect 8757 17283 8815 17289
rect 9401 17323 9459 17329
rect 9401 17289 9413 17323
rect 9447 17320 9459 17323
rect 10226 17320 10232 17332
rect 9447 17292 10232 17320
rect 9447 17289 9459 17292
rect 9401 17283 9459 17289
rect 10226 17280 10232 17292
rect 10284 17280 10290 17332
rect 11882 17280 11888 17332
rect 11940 17320 11946 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 11940 17292 12173 17320
rect 11940 17280 11946 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 12161 17283 12219 17289
rect 2148 17193 2176 17280
rect 3694 17212 3700 17264
rect 3752 17252 3758 17264
rect 4617 17255 4675 17261
rect 4617 17252 4629 17255
rect 3752 17224 4629 17252
rect 3752 17212 3758 17224
rect 4617 17221 4629 17224
rect 4663 17221 4675 17255
rect 9674 17252 9680 17264
rect 9635 17224 9680 17252
rect 4617 17215 4675 17221
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 2400 17051 2458 17057
rect 2400 17048 2412 17051
rect 2148 17020 2412 17048
rect 2148 16992 2176 17020
rect 2400 17017 2412 17020
rect 2446 17048 2458 17051
rect 2866 17048 2872 17060
rect 2446 17020 2872 17048
rect 2446 17017 2458 17020
rect 2400 17011 2458 17017
rect 2866 17008 2872 17020
rect 2924 17048 2930 17060
rect 3786 17048 3792 17060
rect 2924 17020 3792 17048
rect 2924 17008 2930 17020
rect 3786 17008 3792 17020
rect 3844 17008 3850 17060
rect 4632 17048 4660 17215
rect 9674 17212 9680 17224
rect 9732 17212 9738 17264
rect 5534 17144 5540 17196
rect 5592 17184 5598 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5592 17156 5733 17184
rect 5592 17144 5598 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 12176 17184 12204 17283
rect 16114 17280 16120 17332
rect 16172 17320 16178 17332
rect 16209 17323 16267 17329
rect 16209 17320 16221 17323
rect 16172 17292 16221 17320
rect 16172 17280 16178 17292
rect 16209 17289 16221 17292
rect 16255 17320 16267 17323
rect 17494 17320 17500 17332
rect 16255 17292 16896 17320
rect 17455 17292 17500 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 15289 17255 15347 17261
rect 15289 17221 15301 17255
rect 15335 17252 15347 17255
rect 15562 17252 15568 17264
rect 15335 17224 15568 17252
rect 15335 17221 15347 17224
rect 15289 17215 15347 17221
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12176 17156 12449 17184
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17116 5135 17119
rect 5626 17116 5632 17128
rect 5123 17088 5632 17116
rect 5123 17085 5135 17088
rect 5077 17079 5135 17085
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 6638 17076 6644 17128
rect 6696 17116 6702 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6696 17088 6837 17116
rect 6696 17076 6702 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 9861 17119 9919 17125
rect 9861 17085 9873 17119
rect 9907 17116 9919 17119
rect 9950 17116 9956 17128
rect 9907 17088 9956 17116
rect 9907 17085 9919 17088
rect 9861 17079 9919 17085
rect 9950 17076 9956 17088
rect 10008 17116 10014 17128
rect 12176 17116 12204 17156
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 12437 17147 12495 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 16868 17193 16896 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17862 17320 17868 17332
rect 17823 17292 17868 17320
rect 17862 17280 17868 17292
rect 17920 17320 17926 17332
rect 20441 17323 20499 17329
rect 20441 17320 20453 17323
rect 17920 17292 20453 17320
rect 17920 17280 17926 17292
rect 20441 17289 20453 17292
rect 20487 17320 20499 17323
rect 20622 17320 20628 17332
rect 20487 17292 20628 17320
rect 20487 17289 20499 17292
rect 20441 17283 20499 17289
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 23477 17323 23535 17329
rect 23477 17289 23489 17323
rect 23523 17320 23535 17323
rect 23566 17320 23572 17332
rect 23523 17292 23572 17320
rect 23523 17289 23535 17292
rect 23477 17283 23535 17289
rect 23566 17280 23572 17292
rect 23624 17280 23630 17332
rect 24670 17280 24676 17332
rect 24728 17320 24734 17332
rect 25409 17323 25467 17329
rect 25409 17320 25421 17323
rect 24728 17292 25421 17320
rect 24728 17280 24734 17292
rect 25409 17289 25421 17292
rect 25455 17289 25467 17323
rect 25409 17283 25467 17289
rect 25682 17280 25688 17332
rect 25740 17320 25746 17332
rect 26050 17320 26056 17332
rect 25740 17292 26056 17320
rect 25740 17280 25746 17292
rect 26050 17280 26056 17292
rect 26108 17280 26114 17332
rect 18046 17212 18052 17264
rect 18104 17252 18110 17264
rect 18509 17255 18567 17261
rect 18509 17252 18521 17255
rect 18104 17224 18521 17252
rect 18104 17212 18110 17224
rect 18509 17221 18521 17224
rect 18555 17252 18567 17255
rect 18877 17255 18935 17261
rect 18877 17252 18889 17255
rect 18555 17224 18889 17252
rect 18555 17221 18567 17224
rect 18509 17215 18567 17221
rect 18877 17221 18889 17224
rect 18923 17252 18935 17255
rect 21453 17255 21511 17261
rect 18923 17224 19104 17252
rect 18923 17221 18935 17224
rect 18877 17215 18935 17221
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17153 16911 17187
rect 16853 17147 16911 17153
rect 17037 17187 17095 17193
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17586 17184 17592 17196
rect 17083 17156 17592 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 19076 17193 19104 17224
rect 21453 17221 21465 17255
rect 21499 17252 21511 17255
rect 23014 17252 23020 17264
rect 21499 17224 23020 17252
rect 21499 17221 21511 17224
rect 21453 17215 21511 17221
rect 19061 17187 19119 17193
rect 19061 17153 19073 17187
rect 19107 17153 19119 17187
rect 19061 17147 19119 17153
rect 10008 17088 12204 17116
rect 16761 17119 16819 17125
rect 10008 17076 10014 17088
rect 16761 17085 16773 17119
rect 16807 17116 16819 17119
rect 17494 17116 17500 17128
rect 16807 17088 17500 17116
rect 16807 17085 16819 17088
rect 16761 17079 16819 17085
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 19334 17125 19340 17128
rect 19328 17079 19340 17125
rect 19392 17116 19398 17128
rect 21928 17125 21956 17224
rect 23014 17212 23020 17224
rect 23072 17212 23078 17264
rect 22094 17184 22100 17196
rect 22055 17156 22100 17184
rect 22094 17144 22100 17156
rect 22152 17144 22158 17196
rect 23584 17184 23612 17280
rect 24121 17187 24179 17193
rect 24121 17184 24133 17187
rect 23584 17156 24133 17184
rect 24121 17153 24133 17156
rect 24167 17153 24179 17187
rect 24121 17147 24179 17153
rect 24213 17187 24271 17193
rect 24213 17153 24225 17187
rect 24259 17153 24271 17187
rect 24213 17147 24271 17153
rect 21913 17119 21971 17125
rect 19392 17088 20024 17116
rect 19334 17076 19340 17079
rect 19392 17076 19398 17088
rect 19996 17060 20024 17088
rect 21913 17085 21925 17119
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 22462 17076 22468 17128
rect 22520 17116 22526 17128
rect 23382 17116 23388 17128
rect 22520 17088 23388 17116
rect 22520 17076 22526 17088
rect 23382 17076 23388 17088
rect 23440 17116 23446 17128
rect 24228 17116 24256 17147
rect 24673 17119 24731 17125
rect 24673 17116 24685 17119
rect 23440 17088 24685 17116
rect 23440 17076 23446 17088
rect 24673 17085 24685 17088
rect 24719 17116 24731 17119
rect 24762 17116 24768 17128
rect 24719 17088 24768 17116
rect 24719 17085 24731 17088
rect 24673 17079 24731 17085
rect 24762 17076 24768 17088
rect 24820 17076 24826 17128
rect 25222 17116 25228 17128
rect 25183 17088 25228 17116
rect 25222 17076 25228 17088
rect 25280 17116 25286 17128
rect 25777 17119 25835 17125
rect 25777 17116 25789 17119
rect 25280 17088 25789 17116
rect 25280 17076 25286 17088
rect 25777 17085 25789 17088
rect 25823 17085 25835 17119
rect 25777 17079 25835 17085
rect 5537 17051 5595 17057
rect 5537 17048 5549 17051
rect 4632 17020 5549 17048
rect 5537 17017 5549 17020
rect 5583 17017 5595 17051
rect 5537 17011 5595 17017
rect 6270 17008 6276 17060
rect 6328 17048 6334 17060
rect 7070 17051 7128 17057
rect 7070 17048 7082 17051
rect 6328 17020 7082 17048
rect 6328 17008 6334 17020
rect 7070 17017 7082 17020
rect 7116 17048 7128 17051
rect 7926 17048 7932 17060
rect 7116 17020 7932 17048
rect 7116 17017 7128 17020
rect 7070 17011 7128 17017
rect 7926 17008 7932 17020
rect 7984 17008 7990 17060
rect 9398 17008 9404 17060
rect 9456 17048 9462 17060
rect 10106 17051 10164 17057
rect 10106 17048 10118 17051
rect 9456 17020 10118 17048
rect 9456 17008 9462 17020
rect 10106 17017 10118 17020
rect 10152 17048 10164 17051
rect 11698 17048 11704 17060
rect 10152 17020 11704 17048
rect 10152 17017 10164 17020
rect 10106 17011 10164 17017
rect 11698 17008 11704 17020
rect 11756 17048 11762 17060
rect 11793 17051 11851 17057
rect 11793 17048 11805 17051
rect 11756 17020 11805 17048
rect 11756 17008 11762 17020
rect 11793 17017 11805 17020
rect 11839 17017 11851 17051
rect 11793 17011 11851 17017
rect 12618 17008 12624 17060
rect 12676 17057 12682 17060
rect 12676 17051 12740 17057
rect 12676 17017 12694 17051
rect 12728 17017 12740 17051
rect 12676 17011 12740 17017
rect 12676 17008 12682 17011
rect 13630 17008 13636 17060
rect 13688 17048 13694 17060
rect 14369 17051 14427 17057
rect 14369 17048 14381 17051
rect 13688 17020 14381 17048
rect 13688 17008 13694 17020
rect 14369 17017 14381 17020
rect 14415 17017 14427 17051
rect 14369 17011 14427 17017
rect 19978 17008 19984 17060
rect 20036 17008 20042 17060
rect 22005 17051 22063 17057
rect 22005 17048 22017 17051
rect 21008 17020 22017 17048
rect 2130 16940 2136 16992
rect 2188 16940 2194 16992
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 3513 16983 3571 16989
rect 3513 16980 3525 16983
rect 3476 16952 3525 16980
rect 3476 16940 3482 16952
rect 3513 16949 3525 16952
rect 3559 16949 3571 16983
rect 6546 16980 6552 16992
rect 6507 16952 6552 16980
rect 3513 16943 3571 16949
rect 6546 16940 6552 16952
rect 6604 16940 6610 16992
rect 8202 16980 8208 16992
rect 8163 16952 8208 16980
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11241 16983 11299 16989
rect 11241 16980 11253 16983
rect 11204 16952 11253 16980
rect 11204 16940 11210 16952
rect 11241 16949 11253 16952
rect 11287 16949 11299 16983
rect 13814 16980 13820 16992
rect 13775 16952 13820 16980
rect 11241 16943 11299 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 14921 16983 14979 16989
rect 14921 16949 14933 16983
rect 14967 16980 14979 16983
rect 15102 16980 15108 16992
rect 14967 16952 15108 16980
rect 14967 16949 14979 16952
rect 14921 16943 14979 16949
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 15528 16952 15853 16980
rect 15528 16940 15534 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 16390 16980 16396 16992
rect 16351 16952 16396 16980
rect 15841 16943 15899 16949
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 16942 16940 16948 16992
rect 17000 16980 17006 16992
rect 17678 16980 17684 16992
rect 17000 16952 17684 16980
rect 17000 16940 17006 16952
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 18046 16980 18052 16992
rect 18007 16952 18052 16980
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 20898 16940 20904 16992
rect 20956 16980 20962 16992
rect 21008 16989 21036 17020
rect 22005 17017 22017 17020
rect 22051 17017 22063 17051
rect 22005 17011 22063 17017
rect 22186 17008 22192 17060
rect 22244 17048 22250 17060
rect 23017 17051 23075 17057
rect 23017 17048 23029 17051
rect 22244 17020 23029 17048
rect 22244 17008 22250 17020
rect 23017 17017 23029 17020
rect 23063 17048 23075 17051
rect 24029 17051 24087 17057
rect 24029 17048 24041 17051
rect 23063 17020 24041 17048
rect 23063 17017 23075 17020
rect 23017 17011 23075 17017
rect 24029 17017 24041 17020
rect 24075 17017 24087 17051
rect 24029 17011 24087 17017
rect 20993 16983 21051 16989
rect 20993 16980 21005 16983
rect 20956 16952 21005 16980
rect 20956 16940 20962 16952
rect 20993 16949 21005 16952
rect 21039 16949 21051 16983
rect 20993 16943 21051 16949
rect 21450 16940 21456 16992
rect 21508 16980 21514 16992
rect 21545 16983 21603 16989
rect 21545 16980 21557 16983
rect 21508 16952 21557 16980
rect 21508 16940 21514 16952
rect 21545 16949 21557 16952
rect 21591 16949 21603 16983
rect 22738 16980 22744 16992
rect 22699 16952 22744 16980
rect 21545 16943 21603 16949
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 23658 16980 23664 16992
rect 23619 16952 23664 16980
rect 23658 16940 23664 16952
rect 23716 16940 23722 16992
rect 25130 16980 25136 16992
rect 25091 16952 25136 16980
rect 25130 16940 25136 16952
rect 25188 16940 25194 16992
rect 1104 16890 26864 16912
rect 1104 16838 10315 16890
rect 10367 16838 10379 16890
rect 10431 16838 10443 16890
rect 10495 16838 10507 16890
rect 10559 16838 19648 16890
rect 19700 16838 19712 16890
rect 19764 16838 19776 16890
rect 19828 16838 19840 16890
rect 19892 16838 26864 16890
rect 1104 16816 26864 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 2590 16776 2596 16788
rect 1627 16748 2596 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 2590 16736 2596 16748
rect 2648 16736 2654 16788
rect 2774 16736 2780 16788
rect 2832 16736 2838 16788
rect 3510 16776 3516 16788
rect 3471 16748 3516 16776
rect 3510 16736 3516 16748
rect 3568 16736 3574 16788
rect 3786 16776 3792 16788
rect 3747 16748 3792 16776
rect 3786 16736 3792 16748
rect 3844 16736 3850 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 6365 16779 6423 16785
rect 6365 16776 6377 16779
rect 5592 16748 6377 16776
rect 5592 16736 5598 16748
rect 6365 16745 6377 16748
rect 6411 16745 6423 16779
rect 7926 16776 7932 16788
rect 7887 16748 7932 16776
rect 6365 16739 6423 16745
rect 2133 16711 2191 16717
rect 2133 16677 2145 16711
rect 2179 16708 2191 16711
rect 2498 16708 2504 16720
rect 2179 16680 2504 16708
rect 2179 16677 2191 16680
rect 2133 16671 2191 16677
rect 2498 16668 2504 16680
rect 2556 16708 2562 16720
rect 2792 16708 2820 16736
rect 2556 16680 2820 16708
rect 2869 16711 2927 16717
rect 2556 16668 2562 16680
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 2915 16680 3188 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 2038 16640 2044 16652
rect 1964 16612 2044 16640
rect 1964 16584 1992 16612
rect 2038 16600 2044 16612
rect 2096 16600 2102 16652
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3050 16640 3056 16652
rect 2823 16612 3056 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 1946 16532 1952 16584
rect 2004 16532 2010 16584
rect 2406 16532 2412 16584
rect 2464 16572 2470 16584
rect 2958 16572 2964 16584
rect 2464 16544 2728 16572
rect 2919 16544 2964 16572
rect 2464 16532 2470 16544
rect 2700 16448 2728 16544
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 3160 16572 3188 16680
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 4310 16711 4368 16717
rect 4310 16708 4322 16711
rect 3476 16680 4322 16708
rect 3476 16668 3482 16680
rect 4310 16677 4322 16680
rect 4356 16677 4368 16711
rect 6380 16708 6408 16739
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 8076 16748 8493 16776
rect 8076 16736 8082 16748
rect 8481 16745 8493 16748
rect 8527 16776 8539 16779
rect 8570 16776 8576 16788
rect 8527 16748 8576 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 9398 16776 9404 16788
rect 8720 16748 9404 16776
rect 8720 16736 8726 16748
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 9950 16776 9956 16788
rect 9911 16748 9956 16776
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 11698 16776 11704 16788
rect 11659 16748 11704 16776
rect 11698 16736 11704 16748
rect 11756 16736 11762 16788
rect 12802 16776 12808 16788
rect 12763 16748 12808 16776
rect 12802 16736 12808 16748
rect 12860 16736 12866 16788
rect 14182 16776 14188 16788
rect 14143 16748 14188 16776
rect 14182 16736 14188 16748
rect 14240 16736 14246 16788
rect 14550 16776 14556 16788
rect 14511 16748 14556 16776
rect 14550 16736 14556 16748
rect 14608 16736 14614 16788
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 16022 16776 16028 16788
rect 14884 16748 16028 16776
rect 14884 16736 14890 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16574 16736 16580 16788
rect 16632 16776 16638 16788
rect 17129 16779 17187 16785
rect 17129 16776 17141 16779
rect 16632 16748 17141 16776
rect 16632 16736 16638 16748
rect 17129 16745 17141 16748
rect 17175 16776 17187 16779
rect 17402 16776 17408 16788
rect 17175 16748 17408 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 17862 16736 17868 16788
rect 17920 16776 17926 16788
rect 18322 16776 18328 16788
rect 17920 16748 18328 16776
rect 17920 16736 17926 16748
rect 18322 16736 18328 16748
rect 18380 16776 18386 16788
rect 18693 16779 18751 16785
rect 18693 16776 18705 16779
rect 18380 16748 18705 16776
rect 18380 16736 18386 16748
rect 18693 16745 18705 16748
rect 18739 16745 18751 16779
rect 18693 16739 18751 16745
rect 19242 16736 19248 16788
rect 19300 16776 19306 16788
rect 19705 16779 19763 16785
rect 19705 16776 19717 16779
rect 19300 16748 19717 16776
rect 19300 16736 19306 16748
rect 19705 16745 19717 16748
rect 19751 16745 19763 16779
rect 20254 16776 20260 16788
rect 20215 16748 20260 16776
rect 19705 16739 19763 16745
rect 20254 16736 20260 16748
rect 20312 16736 20318 16788
rect 20622 16776 20628 16788
rect 20583 16748 20628 16776
rect 20622 16736 20628 16748
rect 20680 16736 20686 16788
rect 20898 16776 20904 16788
rect 20859 16748 20904 16776
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 22646 16776 22652 16788
rect 21008 16748 21496 16776
rect 22607 16748 22652 16776
rect 6794 16711 6852 16717
rect 6794 16708 6806 16711
rect 6380 16680 6806 16708
rect 4310 16671 4368 16677
rect 6794 16677 6806 16680
rect 6840 16677 6852 16711
rect 6794 16671 6852 16677
rect 7006 16668 7012 16720
rect 7064 16668 7070 16720
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 4614 16640 4620 16652
rect 4111 16612 4620 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16640 6147 16643
rect 6362 16640 6368 16652
rect 6135 16612 6368 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 6362 16600 6368 16612
rect 6420 16600 6426 16652
rect 6454 16600 6460 16652
rect 6512 16640 6518 16652
rect 7024 16640 7052 16668
rect 6512 16612 7052 16640
rect 6512 16600 6518 16612
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 9030 16640 9036 16652
rect 8536 16612 9036 16640
rect 8536 16600 8542 16612
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9968 16640 9996 16736
rect 10134 16668 10140 16720
rect 10192 16708 10198 16720
rect 10566 16711 10624 16717
rect 10566 16708 10578 16711
rect 10192 16680 10578 16708
rect 10192 16668 10198 16680
rect 10566 16677 10578 16680
rect 10612 16677 10624 16711
rect 10566 16671 10624 16677
rect 13173 16711 13231 16717
rect 13173 16677 13185 16711
rect 13219 16708 13231 16711
rect 13446 16708 13452 16720
rect 13219 16680 13452 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 13446 16668 13452 16680
rect 13504 16668 13510 16720
rect 14918 16708 14924 16720
rect 14879 16680 14924 16708
rect 14918 16668 14924 16680
rect 14976 16668 14982 16720
rect 15657 16711 15715 16717
rect 15657 16677 15669 16711
rect 15703 16708 15715 16711
rect 15703 16680 17448 16708
rect 15703 16677 15715 16680
rect 15657 16671 15715 16677
rect 10318 16640 10324 16652
rect 9968 16612 10324 16640
rect 10318 16600 10324 16612
rect 10376 16600 10382 16652
rect 13814 16640 13820 16652
rect 13775 16612 13820 16640
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 15746 16640 15752 16652
rect 15707 16612 15752 16640
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16500 16612 17233 16640
rect 3602 16572 3608 16584
rect 3160 16544 3608 16572
rect 3602 16532 3608 16544
rect 3660 16532 3666 16584
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6549 16575 6607 16581
rect 6549 16572 6561 16575
rect 6328 16544 6561 16572
rect 6328 16532 6334 16544
rect 6549 16541 6561 16544
rect 6595 16541 6607 16575
rect 13262 16572 13268 16584
rect 13223 16544 13268 16572
rect 6549 16535 6607 16541
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 13449 16575 13507 16581
rect 13449 16541 13461 16575
rect 13495 16572 13507 16575
rect 13722 16572 13728 16584
rect 13495 16544 13728 16572
rect 13495 16541 13507 16544
rect 13449 16535 13507 16541
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 15930 16532 15936 16584
rect 15988 16572 15994 16584
rect 16500 16572 16528 16612
rect 17221 16609 17233 16612
rect 17267 16640 17279 16643
rect 17267 16612 17356 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 15988 16544 16528 16572
rect 15988 16532 15994 16544
rect 5000 16476 6592 16504
rect 5000 16448 5028 16476
rect 2406 16436 2412 16448
rect 2367 16408 2412 16436
rect 2406 16396 2412 16408
rect 2464 16396 2470 16448
rect 2682 16396 2688 16448
rect 2740 16396 2746 16448
rect 4982 16396 4988 16448
rect 5040 16396 5046 16448
rect 5442 16436 5448 16448
rect 5403 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 6564 16436 6592 16476
rect 11422 16464 11428 16516
rect 11480 16504 11486 16516
rect 11698 16504 11704 16516
rect 11480 16476 11704 16504
rect 11480 16464 11486 16476
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 16298 16464 16304 16516
rect 16356 16504 16362 16516
rect 16485 16507 16543 16513
rect 16485 16504 16497 16507
rect 16356 16476 16497 16504
rect 16356 16464 16362 16476
rect 16485 16473 16497 16476
rect 16531 16504 16543 16507
rect 16850 16504 16856 16516
rect 16531 16476 16856 16504
rect 16531 16473 16543 16476
rect 16485 16467 16543 16473
rect 16850 16464 16856 16476
rect 16908 16464 16914 16516
rect 17328 16504 17356 16612
rect 17420 16581 17448 16680
rect 18138 16668 18144 16720
rect 18196 16708 18202 16720
rect 18785 16711 18843 16717
rect 18785 16708 18797 16711
rect 18196 16680 18797 16708
rect 18196 16668 18202 16680
rect 18785 16677 18797 16680
rect 18831 16708 18843 16711
rect 18966 16708 18972 16720
rect 18831 16680 18972 16708
rect 18831 16677 18843 16680
rect 18785 16671 18843 16677
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 19429 16711 19487 16717
rect 19429 16677 19441 16711
rect 19475 16708 19487 16711
rect 19978 16708 19984 16720
rect 19475 16680 19984 16708
rect 19475 16677 19487 16680
rect 19429 16671 19487 16677
rect 19978 16668 19984 16680
rect 20036 16668 20042 16720
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 20272 16640 20300 16736
rect 19392 16612 20300 16640
rect 20640 16640 20668 16736
rect 20806 16668 20812 16720
rect 20864 16708 20870 16720
rect 21008 16708 21036 16748
rect 21358 16708 21364 16720
rect 20864 16680 21036 16708
rect 21319 16680 21364 16708
rect 20864 16668 20870 16680
rect 21358 16668 21364 16680
rect 21416 16668 21422 16720
rect 21266 16640 21272 16652
rect 20640 16612 20760 16640
rect 21227 16612 21272 16640
rect 19392 16600 19398 16612
rect 17405 16575 17463 16581
rect 17405 16541 17417 16575
rect 17451 16572 17463 16575
rect 17678 16572 17684 16584
rect 17451 16544 17684 16572
rect 17451 16541 17463 16544
rect 17405 16535 17463 16541
rect 17678 16532 17684 16544
rect 17736 16572 17742 16584
rect 18969 16575 19027 16581
rect 18969 16572 18981 16575
rect 17736 16544 18981 16572
rect 17736 16532 17742 16544
rect 18969 16541 18981 16544
rect 19015 16572 19027 16575
rect 19150 16572 19156 16584
rect 19015 16544 19156 16572
rect 19015 16541 19027 16544
rect 18969 16535 19027 16541
rect 19150 16532 19156 16544
rect 19208 16532 19214 16584
rect 20732 16572 20760 16612
rect 21266 16600 21272 16612
rect 21324 16600 21330 16652
rect 21468 16640 21496 16748
rect 22646 16736 22652 16748
rect 22704 16736 22710 16788
rect 22830 16736 22836 16788
rect 22888 16776 22894 16788
rect 24673 16779 24731 16785
rect 24673 16776 24685 16779
rect 22888 16748 24685 16776
rect 22888 16736 22894 16748
rect 24673 16745 24685 16748
rect 24719 16745 24731 16779
rect 24673 16739 24731 16745
rect 25409 16779 25467 16785
rect 25409 16745 25421 16779
rect 25455 16776 25467 16779
rect 25590 16776 25596 16788
rect 25455 16748 25596 16776
rect 25455 16745 25467 16748
rect 25409 16739 25467 16745
rect 25590 16736 25596 16748
rect 25648 16736 25654 16788
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 22986 16711 23044 16717
rect 22986 16708 22998 16711
rect 22336 16680 22998 16708
rect 22336 16668 22342 16680
rect 22986 16677 22998 16680
rect 23032 16677 23044 16711
rect 22986 16671 23044 16677
rect 24854 16668 24860 16720
rect 24912 16708 24918 16720
rect 25041 16711 25099 16717
rect 25041 16708 25053 16711
rect 24912 16680 25053 16708
rect 24912 16668 24918 16680
rect 25041 16677 25053 16680
rect 25087 16677 25099 16711
rect 25041 16671 25099 16677
rect 25225 16643 25283 16649
rect 25225 16640 25237 16643
rect 21468 16612 23796 16640
rect 20806 16572 20812 16584
rect 20719 16544 20812 16572
rect 20806 16532 20812 16544
rect 20864 16572 20870 16584
rect 21453 16575 21511 16581
rect 21453 16572 21465 16575
rect 20864 16544 21465 16572
rect 20864 16532 20870 16544
rect 21453 16541 21465 16544
rect 21499 16541 21511 16575
rect 21453 16535 21511 16541
rect 22646 16532 22652 16584
rect 22704 16572 22710 16584
rect 22741 16575 22799 16581
rect 22741 16572 22753 16575
rect 22704 16544 22753 16572
rect 22704 16532 22710 16544
rect 22741 16541 22753 16544
rect 22787 16541 22799 16575
rect 22741 16535 22799 16541
rect 17954 16504 17960 16516
rect 17328 16476 17960 16504
rect 17954 16464 17960 16476
rect 18012 16464 18018 16516
rect 19978 16464 19984 16516
rect 20036 16504 20042 16516
rect 21913 16507 21971 16513
rect 21913 16504 21925 16507
rect 20036 16476 21925 16504
rect 20036 16464 20042 16476
rect 21913 16473 21925 16476
rect 21959 16504 21971 16507
rect 22094 16504 22100 16516
rect 21959 16476 22100 16504
rect 21959 16473 21971 16476
rect 21913 16467 21971 16473
rect 22094 16464 22100 16476
rect 22152 16464 22158 16516
rect 23768 16504 23796 16612
rect 25056 16612 25237 16640
rect 25056 16584 25084 16612
rect 25225 16609 25237 16612
rect 25271 16609 25283 16643
rect 25225 16603 25283 16609
rect 25038 16532 25044 16584
rect 25096 16532 25102 16584
rect 26050 16504 26056 16516
rect 23768 16476 26056 16504
rect 26050 16464 26056 16476
rect 26108 16464 26114 16516
rect 7190 16436 7196 16448
rect 6564 16408 7196 16436
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 12529 16439 12587 16445
rect 12529 16405 12541 16439
rect 12575 16436 12587 16439
rect 12618 16436 12624 16448
rect 12575 16408 12624 16436
rect 12575 16405 12587 16408
rect 12529 16399 12587 16405
rect 12618 16396 12624 16408
rect 12676 16396 12682 16448
rect 16758 16436 16764 16448
rect 16719 16408 16764 16436
rect 16758 16396 16764 16408
rect 16816 16396 16822 16448
rect 18046 16436 18052 16448
rect 18007 16408 18052 16436
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18322 16436 18328 16448
rect 18283 16408 18328 16436
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 23750 16396 23756 16448
rect 23808 16436 23814 16448
rect 23934 16436 23940 16448
rect 23808 16408 23940 16436
rect 23808 16396 23814 16408
rect 23934 16396 23940 16408
rect 23992 16396 23998 16448
rect 24121 16439 24179 16445
rect 24121 16405 24133 16439
rect 24167 16436 24179 16439
rect 24670 16436 24676 16448
rect 24167 16408 24676 16436
rect 24167 16405 24179 16408
rect 24121 16399 24179 16405
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 1104 16346 26864 16368
rect 1104 16294 5648 16346
rect 5700 16294 5712 16346
rect 5764 16294 5776 16346
rect 5828 16294 5840 16346
rect 5892 16294 14982 16346
rect 15034 16294 15046 16346
rect 15098 16294 15110 16346
rect 15162 16294 15174 16346
rect 15226 16294 24315 16346
rect 24367 16294 24379 16346
rect 24431 16294 24443 16346
rect 24495 16294 24507 16346
rect 24559 16294 26864 16346
rect 1104 16272 26864 16294
rect 2958 16192 2964 16244
rect 3016 16232 3022 16244
rect 3053 16235 3111 16241
rect 3053 16232 3065 16235
rect 3016 16204 3065 16232
rect 3016 16192 3022 16204
rect 3053 16201 3065 16204
rect 3099 16201 3111 16235
rect 3053 16195 3111 16201
rect 5077 16235 5135 16241
rect 5077 16201 5089 16235
rect 5123 16232 5135 16235
rect 5534 16232 5540 16244
rect 5123 16204 5540 16232
rect 5123 16201 5135 16204
rect 5077 16195 5135 16201
rect 5534 16192 5540 16204
rect 5592 16232 5598 16244
rect 6181 16235 6239 16241
rect 6181 16232 6193 16235
rect 5592 16204 6193 16232
rect 5592 16192 5598 16204
rect 5169 16167 5227 16173
rect 5169 16164 5181 16167
rect 4080 16136 5181 16164
rect 2498 16056 2504 16108
rect 2556 16096 2562 16108
rect 2685 16099 2743 16105
rect 2685 16096 2697 16099
rect 2556 16068 2697 16096
rect 2556 16056 2562 16068
rect 2685 16065 2697 16068
rect 2731 16096 2743 16099
rect 3050 16096 3056 16108
rect 2731 16068 3056 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 3050 16056 3056 16068
rect 3108 16056 3114 16108
rect 4080 16105 4108 16136
rect 5169 16133 5181 16136
rect 5215 16164 5227 16167
rect 5626 16164 5632 16176
rect 5215 16136 5632 16164
rect 5215 16133 5227 16136
rect 5169 16127 5227 16133
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 5828 16105 5856 16204
rect 6181 16201 6193 16204
rect 6227 16232 6239 16235
rect 6270 16232 6276 16244
rect 6227 16204 6276 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6270 16192 6276 16204
rect 6328 16192 6334 16244
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 8159 16204 8892 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 4065 16099 4123 16105
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 4157 16099 4215 16105
rect 4157 16065 4169 16099
rect 4203 16065 4215 16099
rect 4157 16059 4215 16065
rect 5813 16099 5871 16105
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 8662 16096 8668 16108
rect 8623 16068 8668 16096
rect 5813 16059 5871 16065
rect 1854 15988 1860 16040
rect 1912 15988 1918 16040
rect 1949 16031 2007 16037
rect 1949 15997 1961 16031
rect 1995 16028 2007 16031
rect 1995 16000 2636 16028
rect 1995 15997 2007 16000
rect 1949 15991 2007 15997
rect 1872 15960 1900 15988
rect 2222 15960 2228 15972
rect 1872 15932 2228 15960
rect 2222 15920 2228 15932
rect 2280 15960 2286 15972
rect 2501 15963 2559 15969
rect 2501 15960 2513 15963
rect 2280 15932 2513 15960
rect 2280 15920 2286 15932
rect 2501 15929 2513 15932
rect 2547 15929 2559 15963
rect 2501 15923 2559 15929
rect 2038 15892 2044 15904
rect 1999 15864 2044 15892
rect 2038 15852 2044 15864
rect 2096 15852 2102 15904
rect 2409 15895 2467 15901
rect 2409 15861 2421 15895
rect 2455 15892 2467 15895
rect 2608 15892 2636 16000
rect 3694 15988 3700 16040
rect 3752 16028 3758 16040
rect 3970 16028 3976 16040
rect 3752 16000 3976 16028
rect 3752 15988 3758 16000
rect 3970 15988 3976 16000
rect 4028 16028 4034 16040
rect 4172 16028 4200 16059
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 8864 16105 8892 16204
rect 10318 16192 10324 16244
rect 10376 16232 10382 16244
rect 10778 16232 10784 16244
rect 10376 16204 10784 16232
rect 10376 16192 10382 16204
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 12526 16232 12532 16244
rect 12487 16204 12532 16232
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 13633 16235 13691 16241
rect 13633 16201 13645 16235
rect 13679 16232 13691 16235
rect 13722 16232 13728 16244
rect 13679 16204 13728 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 12161 16167 12219 16173
rect 12161 16164 12173 16167
rect 11164 16136 12173 16164
rect 8849 16099 8907 16105
rect 8849 16065 8861 16099
rect 8895 16096 8907 16099
rect 9214 16096 9220 16108
rect 8895 16068 9220 16096
rect 8895 16065 8907 16068
rect 8849 16059 8907 16065
rect 9214 16056 9220 16068
rect 9272 16056 9278 16108
rect 10134 16056 10140 16108
rect 10192 16096 10198 16108
rect 11164 16105 11192 16136
rect 12161 16133 12173 16136
rect 12207 16164 12219 16167
rect 12207 16136 13216 16164
rect 12207 16133 12219 16136
rect 12161 16127 12219 16133
rect 10321 16099 10379 16105
rect 10321 16096 10333 16099
rect 10192 16068 10333 16096
rect 10192 16056 10198 16068
rect 10321 16065 10333 16068
rect 10367 16096 10379 16099
rect 11149 16099 11207 16105
rect 11149 16096 11161 16099
rect 10367 16068 11161 16096
rect 10367 16065 10379 16068
rect 10321 16059 10379 16065
rect 11149 16065 11161 16068
rect 11195 16065 11207 16099
rect 11149 16059 11207 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16096 11943 16099
rect 12986 16096 12992 16108
rect 11931 16068 12992 16096
rect 11931 16065 11943 16068
rect 11885 16059 11943 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 13188 16105 13216 16136
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16096 13231 16099
rect 13648 16096 13676 16195
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 15930 16232 15936 16244
rect 15891 16204 15936 16232
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 16390 16232 16396 16244
rect 16351 16204 16396 16232
rect 16390 16192 16396 16204
rect 16448 16192 16454 16244
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18966 16192 18972 16244
rect 19024 16232 19030 16244
rect 19061 16235 19119 16241
rect 19061 16232 19073 16235
rect 19024 16204 19073 16232
rect 19024 16192 19030 16204
rect 19061 16201 19073 16204
rect 19107 16201 19119 16235
rect 19061 16195 19119 16201
rect 19518 16192 19524 16244
rect 19576 16232 19582 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 19576 16204 19625 16232
rect 19576 16192 19582 16204
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 20714 16232 20720 16244
rect 20675 16204 20720 16232
rect 19613 16195 19671 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 22278 16192 22284 16244
rect 22336 16232 22342 16244
rect 22373 16235 22431 16241
rect 22373 16232 22385 16235
rect 22336 16204 22385 16232
rect 22336 16192 22342 16204
rect 22373 16201 22385 16204
rect 22419 16201 22431 16235
rect 22373 16195 22431 16201
rect 22646 16192 22652 16244
rect 22704 16232 22710 16244
rect 22741 16235 22799 16241
rect 22741 16232 22753 16235
rect 22704 16204 22753 16232
rect 22704 16192 22710 16204
rect 22741 16201 22753 16204
rect 22787 16201 22799 16235
rect 22741 16195 22799 16201
rect 23293 16235 23351 16241
rect 23293 16201 23305 16235
rect 23339 16232 23351 16235
rect 23382 16232 23388 16244
rect 23339 16204 23388 16232
rect 23339 16201 23351 16204
rect 23293 16195 23351 16201
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23661 16235 23719 16241
rect 23661 16201 23673 16235
rect 23707 16232 23719 16235
rect 23842 16232 23848 16244
rect 23707 16204 23848 16232
rect 23707 16201 23719 16204
rect 23661 16195 23719 16201
rect 23842 16192 23848 16204
rect 23900 16192 23906 16244
rect 24118 16192 24124 16244
rect 24176 16232 24182 16244
rect 24673 16235 24731 16241
rect 24673 16232 24685 16235
rect 24176 16204 24685 16232
rect 24176 16192 24182 16204
rect 24673 16201 24685 16204
rect 24719 16201 24731 16235
rect 25406 16232 25412 16244
rect 25367 16204 25412 16232
rect 24673 16195 24731 16201
rect 25406 16192 25412 16204
rect 25464 16192 25470 16244
rect 17402 16164 17408 16176
rect 13219 16068 13676 16096
rect 13924 16136 17408 16164
rect 13219 16065 13231 16068
rect 13173 16059 13231 16065
rect 4028 16000 4200 16028
rect 6825 16031 6883 16037
rect 4028 15988 4034 16000
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7469 16031 7527 16037
rect 7469 16028 7481 16031
rect 6871 16000 7481 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7469 15997 7481 16000
rect 7515 16028 7527 16031
rect 8386 16028 8392 16040
rect 7515 16000 8392 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 8386 15988 8392 16000
rect 8444 15988 8450 16040
rect 8570 16028 8576 16040
rect 8531 16000 8576 16028
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 9674 16028 9680 16040
rect 9587 16000 9680 16028
rect 9674 15988 9680 16000
rect 9732 16028 9738 16040
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 9732 16000 10241 16028
rect 9732 15988 9738 16000
rect 10229 15997 10241 16000
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 12066 15988 12072 16040
rect 12124 16028 12130 16040
rect 13924 16028 13952 16136
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 21177 16167 21235 16173
rect 21177 16133 21189 16167
rect 21223 16164 21235 16167
rect 21266 16164 21272 16176
rect 21223 16136 21272 16164
rect 21223 16133 21235 16136
rect 21177 16127 21235 16133
rect 21266 16124 21272 16136
rect 21324 16164 21330 16176
rect 26145 16167 26203 16173
rect 26145 16164 26157 16167
rect 21324 16136 26157 16164
rect 21324 16124 21330 16136
rect 26145 16133 26157 16136
rect 26191 16133 26203 16167
rect 26145 16127 26203 16133
rect 13998 16056 14004 16108
rect 14056 16056 14062 16108
rect 14737 16099 14795 16105
rect 14737 16065 14749 16099
rect 14783 16096 14795 16099
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 14783 16068 15485 16096
rect 14783 16065 14795 16068
rect 14737 16059 14795 16065
rect 15473 16065 15485 16068
rect 15519 16096 15531 16099
rect 16298 16096 16304 16108
rect 15519 16068 16304 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 16298 16056 16304 16068
rect 16356 16056 16362 16108
rect 17037 16099 17095 16105
rect 17037 16065 17049 16099
rect 17083 16096 17095 16099
rect 17678 16096 17684 16108
rect 17083 16068 17684 16096
rect 17083 16065 17095 16068
rect 17037 16059 17095 16065
rect 17678 16056 17684 16068
rect 17736 16056 17742 16108
rect 18046 16056 18052 16108
rect 18104 16096 18110 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18104 16068 18521 16096
rect 18104 16056 18110 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18690 16096 18696 16108
rect 18651 16068 18696 16096
rect 18509 16059 18567 16065
rect 18690 16056 18696 16068
rect 18748 16056 18754 16108
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 20073 16099 20131 16105
rect 20073 16096 20085 16099
rect 19484 16068 20085 16096
rect 19484 16056 19490 16068
rect 20073 16065 20085 16068
rect 20119 16065 20131 16099
rect 20073 16059 20131 16065
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16096 20315 16099
rect 20530 16096 20536 16108
rect 20303 16068 20536 16096
rect 20303 16065 20315 16068
rect 20257 16059 20315 16065
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 21910 16096 21916 16108
rect 21867 16068 21916 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 21910 16056 21916 16068
rect 21968 16096 21974 16108
rect 22094 16096 22100 16108
rect 21968 16068 22100 16096
rect 21968 16056 21974 16068
rect 22094 16056 22100 16068
rect 22152 16056 22158 16108
rect 23293 16099 23351 16105
rect 23293 16065 23305 16099
rect 23339 16096 23351 16099
rect 24213 16099 24271 16105
rect 24213 16096 24225 16099
rect 23339 16068 24225 16096
rect 23339 16065 23351 16068
rect 23293 16059 23351 16065
rect 24213 16065 24225 16068
rect 24259 16065 24271 16099
rect 24213 16059 24271 16065
rect 12124 16000 13952 16028
rect 14016 16028 14044 16056
rect 14458 16028 14464 16040
rect 14016 16000 14464 16028
rect 12124 15988 12130 16000
rect 14458 15988 14464 16000
rect 14516 15988 14522 16040
rect 18414 16028 18420 16040
rect 18375 16000 18420 16028
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 19978 16028 19984 16040
rect 19939 16000 19984 16028
rect 19978 15988 19984 16000
rect 20036 15988 20042 16040
rect 20714 15988 20720 16040
rect 20772 16028 20778 16040
rect 21545 16031 21603 16037
rect 21545 16028 21557 16031
rect 20772 16000 21557 16028
rect 20772 15988 20778 16000
rect 21545 15997 21557 16000
rect 21591 15997 21603 16031
rect 24118 16028 24124 16040
rect 24079 16000 24124 16028
rect 21545 15991 21603 15997
rect 24118 15988 24124 16000
rect 24176 15988 24182 16040
rect 25222 16028 25228 16040
rect 25183 16000 25228 16028
rect 25222 15988 25228 16000
rect 25280 16028 25286 16040
rect 25777 16031 25835 16037
rect 25777 16028 25789 16031
rect 25280 16000 25789 16028
rect 25280 15988 25286 16000
rect 25777 15997 25789 16000
rect 25823 15997 25835 16031
rect 25777 15991 25835 15997
rect 5629 15963 5687 15969
rect 5629 15929 5641 15963
rect 5675 15960 5687 15963
rect 8018 15960 8024 15972
rect 5675 15932 8024 15960
rect 5675 15929 5687 15932
rect 5629 15923 5687 15929
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 9309 15963 9367 15969
rect 9309 15929 9321 15963
rect 9355 15960 9367 15963
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 9355 15932 10149 15960
rect 9355 15929 9367 15932
rect 9309 15923 9367 15929
rect 10137 15929 10149 15932
rect 10183 15960 10195 15963
rect 11333 15963 11391 15969
rect 11333 15960 11345 15963
rect 10183 15932 11345 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 11333 15929 11345 15932
rect 11379 15929 11391 15963
rect 11333 15923 11391 15929
rect 12897 15963 12955 15969
rect 12897 15929 12909 15963
rect 12943 15960 12955 15963
rect 13998 15960 14004 15972
rect 12943 15932 14004 15960
rect 12943 15929 12955 15932
rect 12897 15923 12955 15929
rect 13998 15920 14004 15932
rect 14056 15920 14062 15972
rect 15286 15960 15292 15972
rect 15199 15932 15292 15960
rect 15286 15920 15292 15932
rect 15344 15960 15350 15972
rect 15344 15932 18092 15960
rect 15344 15920 15350 15932
rect 2682 15892 2688 15904
rect 2455 15864 2688 15892
rect 2455 15861 2467 15864
rect 2409 15855 2467 15861
rect 2682 15852 2688 15864
rect 2740 15852 2746 15904
rect 3418 15892 3424 15904
rect 3379 15864 3424 15892
rect 3418 15852 3424 15864
rect 3476 15852 3482 15904
rect 3602 15892 3608 15904
rect 3563 15864 3608 15892
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 3973 15895 4031 15901
rect 3973 15892 3985 15895
rect 3936 15864 3985 15892
rect 3936 15852 3942 15864
rect 3973 15861 3985 15864
rect 4019 15861 4031 15895
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 3973 15855 4031 15861
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 5534 15892 5540 15904
rect 5495 15864 5540 15892
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6546 15892 6552 15904
rect 6420 15864 6552 15892
rect 6420 15852 6426 15864
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 7006 15892 7012 15904
rect 6967 15864 7012 15892
rect 7006 15852 7012 15864
rect 7064 15852 7070 15904
rect 8202 15892 8208 15904
rect 8163 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9674 15852 9680 15904
rect 9732 15892 9738 15904
rect 9769 15895 9827 15901
rect 9769 15892 9781 15895
rect 9732 15864 9781 15892
rect 9732 15852 9738 15864
rect 9769 15861 9781 15864
rect 9815 15861 9827 15895
rect 9769 15855 9827 15861
rect 13814 15852 13820 15904
rect 13872 15892 13878 15904
rect 14277 15895 14335 15901
rect 14277 15892 14289 15895
rect 13872 15864 14289 15892
rect 13872 15852 13878 15864
rect 14277 15861 14289 15864
rect 14323 15861 14335 15895
rect 14277 15855 14335 15861
rect 14829 15895 14887 15901
rect 14829 15861 14841 15895
rect 14875 15892 14887 15895
rect 15010 15892 15016 15904
rect 14875 15864 15016 15892
rect 14875 15861 14887 15864
rect 14829 15855 14887 15861
rect 15010 15852 15016 15864
rect 15068 15852 15074 15904
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 16301 15895 16359 15901
rect 16301 15892 16313 15895
rect 16264 15864 16313 15892
rect 16264 15852 16270 15864
rect 16301 15861 16313 15864
rect 16347 15892 16359 15895
rect 16666 15892 16672 15904
rect 16347 15864 16672 15892
rect 16347 15861 16359 15864
rect 16301 15855 16359 15861
rect 16666 15852 16672 15864
rect 16724 15892 16730 15904
rect 16761 15895 16819 15901
rect 16761 15892 16773 15895
rect 16724 15864 16773 15892
rect 16724 15852 16730 15864
rect 16761 15861 16773 15864
rect 16807 15861 16819 15895
rect 16761 15855 16819 15861
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17586 15892 17592 15904
rect 16908 15864 17592 15892
rect 16908 15852 16914 15864
rect 17586 15852 17592 15864
rect 17644 15852 17650 15904
rect 18064 15901 18092 15932
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 21082 15960 21088 15972
rect 20680 15932 21088 15960
rect 20680 15920 20686 15932
rect 21082 15920 21088 15932
rect 21140 15920 21146 15972
rect 23290 15920 23296 15972
rect 23348 15960 23354 15972
rect 25314 15960 25320 15972
rect 23348 15932 25320 15960
rect 23348 15920 23354 15932
rect 25314 15920 25320 15932
rect 25372 15920 25378 15972
rect 18049 15895 18107 15901
rect 18049 15861 18061 15895
rect 18095 15861 18107 15895
rect 18049 15855 18107 15861
rect 19150 15852 19156 15904
rect 19208 15892 19214 15904
rect 19518 15892 19524 15904
rect 19208 15864 19524 15892
rect 19208 15852 19214 15864
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 20898 15852 20904 15904
rect 20956 15892 20962 15904
rect 20993 15895 21051 15901
rect 20993 15892 21005 15895
rect 20956 15864 21005 15892
rect 20956 15852 20962 15864
rect 20993 15861 21005 15864
rect 21039 15892 21051 15895
rect 21637 15895 21695 15901
rect 21637 15892 21649 15895
rect 21039 15864 21649 15892
rect 21039 15861 21051 15864
rect 20993 15855 21051 15861
rect 21637 15861 21649 15864
rect 21683 15861 21695 15895
rect 24026 15892 24032 15904
rect 23987 15864 24032 15892
rect 21637 15855 21695 15861
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 25038 15892 25044 15904
rect 24999 15864 25044 15892
rect 25038 15852 25044 15864
rect 25096 15852 25102 15904
rect 1104 15802 26864 15824
rect 1104 15750 10315 15802
rect 10367 15750 10379 15802
rect 10431 15750 10443 15802
rect 10495 15750 10507 15802
rect 10559 15750 19648 15802
rect 19700 15750 19712 15802
rect 19764 15750 19776 15802
rect 19828 15750 19840 15802
rect 19892 15750 26864 15802
rect 1104 15728 26864 15750
rect 3694 15688 3700 15700
rect 3655 15660 3700 15688
rect 3694 15648 3700 15660
rect 3752 15648 3758 15700
rect 6270 15688 6276 15700
rect 6231 15660 6276 15688
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 7190 15688 7196 15700
rect 7151 15660 7196 15688
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 7929 15691 7987 15697
rect 7929 15657 7941 15691
rect 7975 15688 7987 15691
rect 8110 15688 8116 15700
rect 7975 15660 8116 15688
rect 7975 15657 7987 15660
rect 7929 15651 7987 15657
rect 8110 15648 8116 15660
rect 8168 15648 8174 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8846 15688 8852 15700
rect 8527 15660 8852 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 9398 15688 9404 15700
rect 9359 15660 9404 15688
rect 9398 15648 9404 15660
rect 9456 15648 9462 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9677 15691 9735 15697
rect 9677 15688 9689 15691
rect 9548 15660 9689 15688
rect 9548 15648 9554 15660
rect 9677 15657 9689 15660
rect 9723 15657 9735 15691
rect 10134 15688 10140 15700
rect 10095 15660 10140 15688
rect 9677 15651 9735 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 13538 15688 13544 15700
rect 12492 15660 13544 15688
rect 12492 15648 12498 15660
rect 13538 15648 13544 15660
rect 13596 15688 13602 15700
rect 13817 15691 13875 15697
rect 13817 15688 13829 15691
rect 13596 15660 13829 15688
rect 13596 15648 13602 15660
rect 13817 15657 13829 15660
rect 13863 15657 13875 15691
rect 14366 15688 14372 15700
rect 14327 15660 14372 15688
rect 13817 15651 13875 15657
rect 14366 15648 14372 15660
rect 14424 15648 14430 15700
rect 14734 15688 14740 15700
rect 14695 15660 14740 15688
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15562 15688 15568 15700
rect 15523 15660 15568 15688
rect 15562 15648 15568 15660
rect 15620 15648 15626 15700
rect 17129 15691 17187 15697
rect 17129 15657 17141 15691
rect 17175 15688 17187 15691
rect 17310 15688 17316 15700
rect 17175 15660 17316 15688
rect 17175 15657 17187 15660
rect 17129 15651 17187 15657
rect 17310 15648 17316 15660
rect 17368 15648 17374 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18322 15688 18328 15700
rect 18012 15660 18328 15688
rect 18012 15648 18018 15660
rect 18322 15648 18328 15660
rect 18380 15688 18386 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18380 15660 18705 15688
rect 18380 15648 18386 15660
rect 18693 15657 18705 15660
rect 18739 15657 18751 15691
rect 18693 15651 18751 15657
rect 19981 15691 20039 15697
rect 19981 15657 19993 15691
rect 20027 15688 20039 15691
rect 20162 15688 20168 15700
rect 20027 15660 20168 15688
rect 20027 15657 20039 15660
rect 19981 15651 20039 15657
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 21542 15688 21548 15700
rect 21131 15660 21548 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 21542 15648 21548 15660
rect 21600 15648 21606 15700
rect 22094 15688 22100 15700
rect 21836 15660 22100 15688
rect 2777 15623 2835 15629
rect 2777 15589 2789 15623
rect 2823 15620 2835 15623
rect 3786 15620 3792 15632
rect 2823 15592 3792 15620
rect 2823 15589 2835 15592
rect 2777 15583 2835 15589
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 4801 15623 4859 15629
rect 4801 15589 4813 15623
rect 4847 15620 4859 15623
rect 5160 15623 5218 15629
rect 5160 15620 5172 15623
rect 4847 15592 5172 15620
rect 4847 15589 4859 15592
rect 4801 15583 4859 15589
rect 5160 15589 5172 15592
rect 5206 15620 5218 15623
rect 5442 15620 5448 15632
rect 5206 15592 5448 15620
rect 5206 15589 5218 15592
rect 5160 15583 5218 15589
rect 5442 15580 5448 15592
rect 5500 15580 5506 15632
rect 7561 15623 7619 15629
rect 7561 15589 7573 15623
rect 7607 15620 7619 15623
rect 8662 15620 8668 15632
rect 7607 15592 8668 15620
rect 7607 15589 7619 15592
rect 7561 15583 7619 15589
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 11054 15580 11060 15632
rect 11112 15629 11118 15632
rect 11112 15623 11176 15629
rect 11112 15589 11130 15623
rect 11164 15589 11176 15623
rect 11112 15583 11176 15589
rect 12897 15623 12955 15629
rect 12897 15589 12909 15623
rect 12943 15620 12955 15623
rect 13262 15620 13268 15632
rect 12943 15592 13268 15620
rect 12943 15589 12955 15592
rect 12897 15583 12955 15589
rect 11112 15580 11118 15583
rect 13262 15580 13268 15592
rect 13320 15580 13326 15632
rect 13722 15620 13728 15632
rect 13683 15592 13728 15620
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 18414 15580 18420 15632
rect 18472 15620 18478 15632
rect 19245 15623 19303 15629
rect 19245 15620 19257 15623
rect 18472 15592 19257 15620
rect 18472 15580 18478 15592
rect 19245 15589 19257 15592
rect 19291 15589 19303 15623
rect 19245 15583 19303 15589
rect 19705 15623 19763 15629
rect 19705 15589 19717 15623
rect 19751 15620 19763 15623
rect 20530 15620 20536 15632
rect 19751 15592 20536 15620
rect 19751 15589 19763 15592
rect 19705 15583 19763 15589
rect 20530 15580 20536 15592
rect 20588 15580 20594 15632
rect 20714 15580 20720 15632
rect 20772 15620 20778 15632
rect 21836 15629 21864 15660
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 24486 15688 24492 15700
rect 24447 15660 24492 15688
rect 24486 15648 24492 15660
rect 24544 15648 24550 15700
rect 24854 15648 24860 15700
rect 24912 15688 24918 15700
rect 25501 15691 25559 15697
rect 25501 15688 25513 15691
rect 24912 15660 25513 15688
rect 24912 15648 24918 15660
rect 25501 15657 25513 15660
rect 25547 15657 25559 15691
rect 25501 15651 25559 15657
rect 21821 15623 21879 15629
rect 21821 15620 21833 15623
rect 20772 15592 21833 15620
rect 20772 15580 20778 15592
rect 21821 15589 21833 15592
rect 21867 15589 21879 15623
rect 22646 15620 22652 15632
rect 21821 15583 21879 15589
rect 22020 15592 22652 15620
rect 22020 15564 22048 15592
rect 22646 15580 22652 15592
rect 22704 15580 22710 15632
rect 24026 15580 24032 15632
rect 24084 15620 24090 15632
rect 24305 15623 24363 15629
rect 24305 15620 24317 15623
rect 24084 15592 24317 15620
rect 24084 15580 24090 15592
rect 24305 15589 24317 15592
rect 24351 15589 24363 15623
rect 24946 15620 24952 15632
rect 24305 15583 24363 15589
rect 24872 15592 24952 15620
rect 1397 15555 1455 15561
rect 1397 15521 1409 15555
rect 1443 15552 1455 15555
rect 2406 15552 2412 15564
rect 1443 15524 2412 15552
rect 1443 15521 1455 15524
rect 1397 15515 1455 15521
rect 2406 15512 2412 15524
rect 2464 15512 2470 15564
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15552 2927 15555
rect 2958 15552 2964 15564
rect 2915 15524 2964 15552
rect 2915 15521 2927 15524
rect 2869 15515 2927 15521
rect 2958 15512 2964 15524
rect 3016 15512 3022 15564
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 4893 15555 4951 15561
rect 4893 15552 4905 15555
rect 4672 15524 4905 15552
rect 4672 15512 4678 15524
rect 4893 15521 4905 15524
rect 4939 15552 4951 15555
rect 6546 15552 6552 15564
rect 4939 15524 6552 15552
rect 4939 15521 4951 15524
rect 4893 15515 4951 15521
rect 6546 15512 6552 15524
rect 6604 15512 6610 15564
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15552 8447 15555
rect 8478 15552 8484 15564
rect 8435 15524 8484 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 8478 15512 8484 15524
rect 8536 15512 8542 15564
rect 10778 15512 10784 15564
rect 10836 15552 10842 15564
rect 10873 15555 10931 15561
rect 10873 15552 10885 15555
rect 10836 15524 10885 15552
rect 10836 15512 10842 15524
rect 10873 15521 10885 15524
rect 10919 15521 10931 15555
rect 10873 15515 10931 15521
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 15749 15555 15807 15561
rect 15749 15552 15761 15555
rect 15620 15524 15761 15552
rect 15620 15512 15626 15524
rect 15749 15521 15761 15524
rect 15795 15521 15807 15555
rect 15749 15515 15807 15521
rect 16016 15555 16074 15561
rect 16016 15521 16028 15555
rect 16062 15552 16074 15555
rect 16298 15552 16304 15564
rect 16062 15524 16304 15552
rect 16062 15521 16074 15524
rect 16016 15515 16074 15521
rect 16298 15512 16304 15524
rect 16356 15512 16362 15564
rect 17678 15512 17684 15564
rect 17736 15552 17742 15564
rect 18601 15555 18659 15561
rect 18601 15552 18613 15555
rect 17736 15524 18613 15552
rect 17736 15512 17742 15524
rect 18601 15521 18613 15524
rect 18647 15521 18659 15555
rect 18601 15515 18659 15521
rect 19797 15555 19855 15561
rect 19797 15521 19809 15555
rect 19843 15552 19855 15555
rect 19978 15552 19984 15564
rect 19843 15524 19984 15552
rect 19843 15521 19855 15524
rect 19797 15515 19855 15521
rect 19978 15512 19984 15524
rect 20036 15512 20042 15564
rect 20901 15555 20959 15561
rect 20901 15521 20913 15555
rect 20947 15552 20959 15555
rect 20990 15552 20996 15564
rect 20947 15524 20996 15552
rect 20947 15521 20959 15524
rect 20901 15515 20959 15521
rect 20990 15512 20996 15524
rect 21048 15552 21054 15564
rect 21726 15552 21732 15564
rect 21048 15524 21732 15552
rect 21048 15512 21054 15524
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 22002 15552 22008 15564
rect 21915 15524 22008 15552
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 22272 15555 22330 15561
rect 22272 15521 22284 15555
rect 22318 15552 22330 15555
rect 22830 15552 22836 15564
rect 22318 15524 22836 15552
rect 22318 15521 22330 15524
rect 22272 15515 22330 15521
rect 22830 15512 22836 15524
rect 22888 15512 22894 15564
rect 24872 15561 24900 15592
rect 24946 15580 24952 15592
rect 25004 15580 25010 15632
rect 24857 15555 24915 15561
rect 24857 15521 24869 15555
rect 24903 15521 24915 15555
rect 24857 15515 24915 15521
rect 3050 15484 3056 15496
rect 2963 15456 3056 15484
rect 3050 15444 3056 15456
rect 3108 15484 3114 15496
rect 4062 15484 4068 15496
rect 3108 15456 4068 15484
rect 3108 15444 3114 15456
rect 4062 15444 4068 15456
rect 4120 15444 4126 15496
rect 4341 15487 4399 15493
rect 4341 15453 4353 15487
rect 4387 15484 4399 15487
rect 4706 15484 4712 15496
rect 4387 15456 4712 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 13998 15484 14004 15496
rect 13959 15456 14004 15484
rect 8573 15447 8631 15453
rect 1581 15419 1639 15425
rect 1581 15385 1593 15419
rect 1627 15416 1639 15419
rect 1854 15416 1860 15428
rect 1627 15388 1860 15416
rect 1627 15385 1639 15388
rect 1581 15379 1639 15385
rect 1854 15376 1860 15388
rect 1912 15376 1918 15428
rect 8018 15416 8024 15428
rect 7979 15388 8024 15416
rect 8018 15376 8024 15388
rect 8076 15376 8082 15428
rect 8294 15376 8300 15428
rect 8352 15416 8358 15428
rect 8588 15416 8616 15447
rect 13998 15444 14004 15456
rect 14056 15444 14062 15496
rect 18690 15484 18696 15496
rect 18064 15456 18696 15484
rect 8352 15388 8616 15416
rect 13265 15419 13323 15425
rect 8352 15376 8358 15388
rect 13265 15385 13277 15419
rect 13311 15416 13323 15419
rect 13446 15416 13452 15428
rect 13311 15388 13452 15416
rect 13311 15385 13323 15388
rect 13265 15379 13323 15385
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 18064 15360 18092 15456
rect 18690 15444 18696 15456
rect 18748 15484 18754 15496
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 18748 15456 18797 15484
rect 18748 15444 18754 15456
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 18785 15447 18843 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20806 15484 20812 15496
rect 20763 15456 20812 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20806 15444 20812 15456
rect 20864 15444 20870 15496
rect 24946 15484 24952 15496
rect 24907 15456 24952 15484
rect 24946 15444 24952 15456
rect 25004 15444 25010 15496
rect 25041 15487 25099 15493
rect 25041 15453 25053 15487
rect 25087 15453 25099 15487
rect 25041 15447 25099 15453
rect 18138 15376 18144 15428
rect 18196 15416 18202 15428
rect 18233 15419 18291 15425
rect 18233 15416 18245 15419
rect 18196 15388 18245 15416
rect 18196 15376 18202 15388
rect 18233 15385 18245 15388
rect 18279 15385 18291 15419
rect 18233 15379 18291 15385
rect 19518 15376 19524 15428
rect 19576 15416 19582 15428
rect 21545 15419 21603 15425
rect 19576 15388 20668 15416
rect 19576 15376 19582 15388
rect 20640 15360 20668 15388
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 21910 15416 21916 15428
rect 21591 15388 21916 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 21910 15376 21916 15388
rect 21968 15376 21974 15428
rect 24762 15376 24768 15428
rect 24820 15416 24826 15428
rect 25056 15416 25084 15447
rect 25958 15416 25964 15428
rect 24820 15388 25964 15416
rect 24820 15376 24826 15388
rect 25958 15376 25964 15388
rect 26016 15376 26022 15428
rect 2133 15351 2191 15357
rect 2133 15317 2145 15351
rect 2179 15348 2191 15351
rect 2222 15348 2228 15360
rect 2179 15320 2228 15348
rect 2179 15317 2191 15320
rect 2133 15311 2191 15317
rect 2222 15308 2228 15320
rect 2280 15308 2286 15360
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15348 2467 15351
rect 2590 15348 2596 15360
rect 2455 15320 2596 15348
rect 2455 15317 2467 15320
rect 2409 15311 2467 15317
rect 2590 15308 2596 15320
rect 2648 15308 2654 15360
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8628 15320 9045 15348
rect 8628 15308 8634 15320
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 10502 15348 10508 15360
rect 10463 15320 10508 15348
rect 9033 15311 9091 15317
rect 10502 15308 10508 15320
rect 10560 15308 10566 15360
rect 12250 15348 12256 15360
rect 12211 15320 12256 15348
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 13354 15348 13360 15360
rect 13315 15320 13360 15348
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 20346 15348 20352 15360
rect 20307 15320 20352 15348
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20622 15308 20628 15360
rect 20680 15308 20686 15360
rect 23382 15348 23388 15360
rect 23343 15320 23388 15348
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 24029 15351 24087 15357
rect 24029 15317 24041 15351
rect 24075 15348 24087 15351
rect 24118 15348 24124 15360
rect 24075 15320 24124 15348
rect 24075 15317 24087 15320
rect 24029 15311 24087 15317
rect 24118 15308 24124 15320
rect 24176 15308 24182 15360
rect 1104 15258 26864 15280
rect 1104 15206 5648 15258
rect 5700 15206 5712 15258
rect 5764 15206 5776 15258
rect 5828 15206 5840 15258
rect 5892 15206 14982 15258
rect 15034 15206 15046 15258
rect 15098 15206 15110 15258
rect 15162 15206 15174 15258
rect 15226 15206 24315 15258
rect 24367 15206 24379 15258
rect 24431 15206 24443 15258
rect 24495 15206 24507 15258
rect 24559 15206 26864 15258
rect 1104 15184 26864 15206
rect 2866 15104 2872 15156
rect 2924 15144 2930 15156
rect 6270 15144 6276 15156
rect 2924 15116 6276 15144
rect 2924 15104 2930 15116
rect 1578 15076 1584 15088
rect 1539 15048 1584 15076
rect 1578 15036 1584 15048
rect 1636 15036 1642 15088
rect 3068 15017 3096 15116
rect 6270 15104 6276 15116
rect 6328 15104 6334 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7101 15147 7159 15153
rect 7101 15144 7113 15147
rect 6972 15116 7113 15144
rect 6972 15104 6978 15116
rect 7101 15113 7113 15116
rect 7147 15113 7159 15147
rect 7101 15107 7159 15113
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8478 15144 8484 15156
rect 8251 15116 8484 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 8846 15144 8852 15156
rect 8619 15116 8852 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 8846 15104 8852 15116
rect 8904 15104 8910 15156
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 10873 15147 10931 15153
rect 10873 15144 10885 15147
rect 10836 15116 10885 15144
rect 10836 15104 10842 15116
rect 10873 15113 10885 15116
rect 10919 15113 10931 15147
rect 10873 15107 10931 15113
rect 11146 15104 11152 15156
rect 11204 15144 11210 15156
rect 11422 15144 11428 15156
rect 11204 15116 11428 15144
rect 11204 15104 11210 15116
rect 11422 15104 11428 15116
rect 11480 15104 11486 15156
rect 13538 15144 13544 15156
rect 13499 15116 13544 15144
rect 13538 15104 13544 15116
rect 13596 15104 13602 15156
rect 13906 15104 13912 15156
rect 13964 15144 13970 15156
rect 14277 15147 14335 15153
rect 14277 15144 14289 15147
rect 13964 15116 14289 15144
rect 13964 15104 13970 15116
rect 14277 15113 14289 15116
rect 14323 15113 14335 15147
rect 14277 15107 14335 15113
rect 16758 15104 16764 15156
rect 16816 15144 16822 15156
rect 17405 15147 17463 15153
rect 17405 15144 17417 15147
rect 16816 15116 17417 15144
rect 16816 15104 16822 15116
rect 17405 15113 17417 15116
rect 17451 15144 17463 15147
rect 17678 15144 17684 15156
rect 17451 15116 17684 15144
rect 17451 15113 17463 15116
rect 17405 15107 17463 15113
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 17862 15144 17868 15156
rect 17823 15116 17868 15144
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15144 20867 15147
rect 22462 15144 22468 15156
rect 20855 15116 22468 15144
rect 20855 15113 20867 15116
rect 20809 15107 20867 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 22830 15104 22836 15156
rect 22888 15144 22894 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 22888 15116 22937 15144
rect 22888 15104 22894 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 22925 15107 22983 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24210 15104 24216 15156
rect 24268 15144 24274 15156
rect 25409 15147 25467 15153
rect 25409 15144 25421 15147
rect 24268 15116 25421 15144
rect 24268 15104 24274 15116
rect 25409 15113 25421 15116
rect 25455 15113 25467 15147
rect 25409 15107 25467 15113
rect 25958 15104 25964 15156
rect 26016 15144 26022 15156
rect 26145 15147 26203 15153
rect 26145 15144 26157 15147
rect 26016 15116 26157 15144
rect 26016 15104 26022 15116
rect 26145 15113 26157 15116
rect 26191 15113 26203 15147
rect 26145 15107 26203 15113
rect 3697 15079 3755 15085
rect 3697 15045 3709 15079
rect 3743 15076 3755 15079
rect 3786 15076 3792 15088
rect 3743 15048 3792 15076
rect 3743 15045 3755 15048
rect 3697 15039 3755 15045
rect 3786 15036 3792 15048
rect 3844 15076 3850 15088
rect 4062 15076 4068 15088
rect 3844 15048 4068 15076
rect 3844 15036 3850 15048
rect 4062 15036 4068 15048
rect 4120 15036 4126 15088
rect 13998 15036 14004 15088
rect 14056 15076 14062 15088
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 14056 15048 14565 15076
rect 14056 15036 14062 15048
rect 14553 15045 14565 15048
rect 14599 15045 14611 15079
rect 14553 15039 14611 15045
rect 21821 15079 21879 15085
rect 21821 15045 21833 15079
rect 21867 15076 21879 15079
rect 22002 15076 22008 15088
rect 21867 15048 22008 15076
rect 21867 15045 21879 15048
rect 21821 15039 21879 15045
rect 22002 15036 22008 15048
rect 22060 15036 22066 15088
rect 22278 15036 22284 15088
rect 22336 15076 22342 15088
rect 22646 15076 22652 15088
rect 22336 15048 22652 15076
rect 22336 15036 22342 15048
rect 22646 15036 22652 15048
rect 22704 15036 22710 15088
rect 3053 15011 3111 15017
rect 3053 14977 3065 15011
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 3237 15011 3295 15017
rect 3237 14977 3249 15011
rect 3283 15008 3295 15011
rect 3510 15008 3516 15020
rect 3283 14980 3516 15008
rect 3283 14977 3295 14980
rect 3237 14971 3295 14977
rect 3510 14968 3516 14980
rect 3568 14968 3574 15020
rect 7466 14968 7472 15020
rect 7524 15008 7530 15020
rect 7653 15011 7711 15017
rect 7653 15008 7665 15011
rect 7524 14980 7665 15008
rect 7524 14968 7530 14980
rect 7653 14977 7665 14980
rect 7699 15008 7711 15011
rect 8294 15008 8300 15020
rect 7699 14980 8300 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 8294 14968 8300 14980
rect 8352 14968 8358 15020
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11701 15011 11759 15017
rect 11701 15008 11713 15011
rect 11112 14980 11713 15008
rect 11112 14968 11118 14980
rect 11701 14977 11713 14980
rect 11747 15008 11759 15011
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 11747 14980 12265 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 12253 14977 12265 14980
rect 12299 15008 12311 15011
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12299 14980 13093 15008
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 13081 14977 13093 14980
rect 13127 15008 13139 15011
rect 13446 15008 13452 15020
rect 13127 14980 13452 15008
rect 13127 14977 13139 14980
rect 13081 14971 13139 14977
rect 13446 14968 13452 14980
rect 13504 14968 13510 15020
rect 13814 14968 13820 15020
rect 13872 15008 13878 15020
rect 13909 15011 13967 15017
rect 13909 15008 13921 15011
rect 13872 14980 13921 15008
rect 13872 14968 13878 14980
rect 13909 14977 13921 14980
rect 13955 14977 13967 15011
rect 13909 14971 13967 14977
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21361 15011 21419 15017
rect 21361 15008 21373 15011
rect 20772 14980 21373 15008
rect 20772 14968 20778 14980
rect 21361 14977 21373 14980
rect 21407 15008 21419 15011
rect 21637 15011 21695 15017
rect 21637 15008 21649 15011
rect 21407 14980 21649 15008
rect 21407 14977 21419 14980
rect 21361 14971 21419 14977
rect 21637 14977 21649 14980
rect 21683 14977 21695 15011
rect 21637 14971 21695 14977
rect 22557 15011 22615 15017
rect 22557 14977 22569 15011
rect 22603 14977 22615 15011
rect 23492 15008 23520 15104
rect 24854 15036 24860 15088
rect 24912 15076 24918 15088
rect 25041 15079 25099 15085
rect 25041 15076 25053 15079
rect 24912 15048 25053 15076
rect 24912 15036 24918 15048
rect 25041 15045 25053 15048
rect 25087 15045 25099 15079
rect 25041 15039 25099 15045
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23492 14980 24225 15008
rect 22557 14971 22615 14977
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 24213 14971 24271 14977
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 2958 14940 2964 14952
rect 1443 14912 2084 14940
rect 2919 14912 2964 14940
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 2056 14816 2084 14912
rect 2958 14900 2964 14912
rect 3016 14900 3022 14952
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4424 14943 4482 14949
rect 4424 14909 4436 14943
rect 4470 14940 4482 14943
rect 4706 14940 4712 14952
rect 4470 14912 4712 14940
rect 4470 14909 4482 14912
rect 4424 14903 4482 14909
rect 2501 14875 2559 14881
rect 2501 14841 2513 14875
rect 2547 14872 2559 14875
rect 3050 14872 3056 14884
rect 2547 14844 3056 14872
rect 2547 14841 2559 14844
rect 2501 14835 2559 14841
rect 3050 14832 3056 14844
rect 3108 14832 3114 14884
rect 4065 14875 4123 14881
rect 4065 14841 4077 14875
rect 4111 14872 4123 14875
rect 4172 14872 4200 14903
rect 4706 14900 4712 14912
rect 4764 14900 4770 14952
rect 7190 14900 7196 14952
rect 7248 14940 7254 14952
rect 7561 14943 7619 14949
rect 7561 14940 7573 14943
rect 7248 14912 7573 14940
rect 7248 14900 7254 14912
rect 7561 14909 7573 14912
rect 7607 14940 7619 14943
rect 8018 14940 8024 14952
rect 7607 14912 8024 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8665 14943 8723 14949
rect 8665 14909 8677 14943
rect 8711 14940 8723 14943
rect 14093 14943 14151 14949
rect 8711 14912 9076 14940
rect 8711 14909 8723 14912
rect 8665 14903 8723 14909
rect 9048 14884 9076 14912
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14182 14940 14188 14952
rect 14139 14912 14188 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14182 14900 14188 14912
rect 14240 14940 14246 14952
rect 14458 14940 14464 14952
rect 14240 14912 14464 14940
rect 14240 14900 14246 14912
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 15381 14943 15439 14949
rect 15381 14909 15393 14943
rect 15427 14940 15439 14943
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 15427 14912 15485 14940
rect 15427 14909 15439 14912
rect 15381 14903 15439 14909
rect 15473 14909 15485 14912
rect 15519 14940 15531 14943
rect 15562 14940 15568 14952
rect 15519 14912 15568 14940
rect 15519 14909 15531 14912
rect 15473 14903 15531 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 18230 14900 18236 14952
rect 18288 14940 18294 14952
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18288 14912 18337 14940
rect 18288 14900 18294 14912
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 19334 14940 19340 14952
rect 19247 14912 19340 14940
rect 18325 14903 18383 14909
rect 19334 14900 19340 14912
rect 19392 14940 19398 14952
rect 19429 14943 19487 14949
rect 19429 14940 19441 14943
rect 19392 14912 19441 14940
rect 19392 14900 19398 14912
rect 19429 14909 19441 14912
rect 19475 14940 19487 14943
rect 19518 14940 19524 14952
rect 19475 14912 19524 14940
rect 19475 14909 19487 14912
rect 19429 14903 19487 14909
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 22094 14900 22100 14952
rect 22152 14940 22158 14952
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 22152 14912 22385 14940
rect 22152 14900 22158 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 4522 14872 4528 14884
rect 4111 14844 4528 14872
rect 4111 14841 4123 14844
rect 4065 14835 4123 14841
rect 4522 14832 4528 14844
rect 4580 14832 4586 14884
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7374 14872 7380 14884
rect 6687 14844 7380 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7374 14832 7380 14844
rect 7432 14872 7438 14884
rect 7469 14875 7527 14881
rect 7469 14872 7481 14875
rect 7432 14844 7481 14872
rect 7432 14832 7438 14844
rect 7469 14841 7481 14844
rect 7515 14872 7527 14875
rect 7742 14872 7748 14884
rect 7515 14844 7748 14872
rect 7515 14841 7527 14844
rect 7469 14835 7527 14841
rect 7742 14832 7748 14844
rect 7800 14832 7806 14884
rect 8570 14832 8576 14884
rect 8628 14872 8634 14884
rect 8910 14875 8968 14881
rect 8910 14872 8922 14875
rect 8628 14844 8922 14872
rect 8628 14832 8634 14844
rect 8910 14841 8922 14844
rect 8956 14841 8968 14875
rect 8910 14835 8968 14841
rect 9030 14832 9036 14884
rect 9088 14872 9094 14884
rect 10778 14872 10784 14884
rect 9088 14844 10784 14872
rect 9088 14832 9094 14844
rect 10778 14832 10784 14844
rect 10836 14832 10842 14884
rect 12897 14875 12955 14881
rect 12897 14841 12909 14875
rect 12943 14872 12955 14875
rect 13354 14872 13360 14884
rect 12943 14844 13360 14872
rect 12943 14841 12955 14844
rect 12897 14835 12955 14841
rect 13354 14832 13360 14844
rect 13412 14872 13418 14884
rect 13722 14872 13728 14884
rect 13412 14844 13728 14872
rect 13412 14832 13418 14844
rect 13722 14832 13728 14844
rect 13780 14832 13786 14884
rect 15013 14875 15071 14881
rect 15013 14841 15025 14875
rect 15059 14872 15071 14875
rect 15740 14875 15798 14881
rect 15740 14872 15752 14875
rect 15059 14844 15752 14872
rect 15059 14841 15071 14844
rect 15013 14835 15071 14841
rect 15740 14841 15752 14844
rect 15786 14872 15798 14875
rect 16482 14872 16488 14884
rect 15786 14844 16488 14872
rect 15786 14841 15798 14844
rect 15740 14835 15798 14841
rect 16482 14832 16488 14844
rect 16540 14832 16546 14884
rect 18046 14832 18052 14884
rect 18104 14872 18110 14884
rect 18874 14872 18880 14884
rect 18104 14844 18880 14872
rect 18104 14832 18110 14844
rect 18874 14832 18880 14844
rect 18932 14832 18938 14884
rect 19696 14875 19754 14881
rect 19696 14841 19708 14875
rect 19742 14872 19754 14875
rect 20346 14872 20352 14884
rect 19742 14844 20352 14872
rect 19742 14841 19754 14844
rect 19696 14835 19754 14841
rect 20346 14832 20352 14844
rect 20404 14832 20410 14884
rect 21637 14875 21695 14881
rect 21637 14841 21649 14875
rect 21683 14872 21695 14875
rect 22572 14872 22600 14971
rect 23934 14900 23940 14952
rect 23992 14940 23998 14952
rect 24673 14943 24731 14949
rect 24673 14940 24685 14943
rect 23992 14912 24685 14940
rect 23992 14900 23998 14912
rect 24673 14909 24685 14912
rect 24719 14940 24731 14943
rect 24946 14940 24952 14952
rect 24719 14912 24952 14940
rect 24719 14909 24731 14912
rect 24673 14903 24731 14909
rect 24946 14900 24952 14912
rect 25004 14940 25010 14952
rect 25225 14943 25283 14949
rect 25225 14940 25237 14943
rect 25004 14912 25237 14940
rect 25004 14900 25010 14912
rect 25225 14909 25237 14912
rect 25271 14940 25283 14943
rect 25777 14943 25835 14949
rect 25777 14940 25789 14943
rect 25271 14912 25789 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 25777 14909 25789 14912
rect 25823 14909 25835 14943
rect 25777 14903 25835 14909
rect 24026 14872 24032 14884
rect 21683 14844 22600 14872
rect 23987 14844 24032 14872
rect 21683 14841 21695 14844
rect 21637 14835 21695 14841
rect 24026 14832 24032 14844
rect 24084 14832 24090 14884
rect 2038 14804 2044 14816
rect 1999 14776 2044 14804
rect 2038 14764 2044 14776
rect 2096 14764 2102 14816
rect 2593 14807 2651 14813
rect 2593 14773 2605 14807
rect 2639 14804 2651 14807
rect 2866 14804 2872 14816
rect 2639 14776 2872 14804
rect 2639 14773 2651 14776
rect 2593 14767 2651 14773
rect 2866 14764 2872 14776
rect 2924 14764 2930 14816
rect 5534 14804 5540 14816
rect 5495 14776 5540 14804
rect 5534 14764 5540 14776
rect 5592 14764 5598 14816
rect 6181 14807 6239 14813
rect 6181 14773 6193 14807
rect 6227 14804 6239 14807
rect 6546 14804 6552 14816
rect 6227 14776 6552 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 9490 14764 9496 14816
rect 9548 14804 9554 14816
rect 10045 14807 10103 14813
rect 10045 14804 10057 14807
rect 9548 14776 10057 14804
rect 9548 14764 9554 14776
rect 10045 14773 10057 14776
rect 10091 14773 10103 14807
rect 11146 14804 11152 14816
rect 11107 14776 11152 14804
rect 10045 14767 10103 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 12526 14804 12532 14816
rect 12487 14776 12532 14804
rect 12526 14764 12532 14776
rect 12584 14764 12590 14816
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13078 14804 13084 14816
rect 13035 14776 13084 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13078 14764 13084 14776
rect 13136 14764 13142 14816
rect 16850 14804 16856 14816
rect 16811 14776 16856 14804
rect 16850 14764 16856 14776
rect 16908 14764 16914 14816
rect 18506 14804 18512 14816
rect 18467 14776 18512 14804
rect 18506 14764 18512 14776
rect 18564 14764 18570 14816
rect 21910 14804 21916 14816
rect 21871 14776 21916 14804
rect 21910 14764 21916 14776
rect 21968 14764 21974 14816
rect 22278 14804 22284 14816
rect 22239 14776 22284 14804
rect 22278 14764 22284 14776
rect 22336 14764 22342 14816
rect 23658 14804 23664 14816
rect 23619 14776 23664 14804
rect 23658 14764 23664 14776
rect 23716 14764 23722 14816
rect 24118 14804 24124 14816
rect 24079 14776 24124 14804
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 1104 14714 26864 14736
rect 1104 14662 10315 14714
rect 10367 14662 10379 14714
rect 10431 14662 10443 14714
rect 10495 14662 10507 14714
rect 10559 14662 19648 14714
rect 19700 14662 19712 14714
rect 19764 14662 19776 14714
rect 19828 14662 19840 14714
rect 19892 14662 26864 14714
rect 1104 14640 26864 14662
rect 1949 14603 2007 14609
rect 1949 14569 1961 14603
rect 1995 14600 2007 14603
rect 2314 14600 2320 14612
rect 1995 14572 2320 14600
rect 1995 14569 2007 14572
rect 1949 14563 2007 14569
rect 1397 14467 1455 14473
rect 1397 14433 1409 14467
rect 1443 14464 1455 14467
rect 1964 14464 1992 14563
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 2406 14560 2412 14612
rect 2464 14600 2470 14612
rect 2464 14572 2509 14600
rect 2464 14560 2470 14572
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3384 14572 3801 14600
rect 3384 14560 3390 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 3789 14563 3847 14569
rect 4522 14560 4528 14612
rect 4580 14560 4586 14612
rect 6270 14600 6276 14612
rect 6231 14572 6276 14600
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 7466 14600 7472 14612
rect 7427 14572 7472 14600
rect 7466 14560 7472 14572
rect 7524 14600 7530 14612
rect 7837 14603 7895 14609
rect 7837 14600 7849 14603
rect 7524 14572 7849 14600
rect 7524 14560 7530 14572
rect 7837 14569 7849 14572
rect 7883 14569 7895 14603
rect 11054 14600 11060 14612
rect 11015 14572 11060 14600
rect 7837 14563 7895 14569
rect 2866 14532 2872 14544
rect 2827 14504 2872 14532
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 3510 14532 3516 14544
rect 3471 14504 3516 14532
rect 3510 14492 3516 14504
rect 3568 14492 3574 14544
rect 1443 14436 1992 14464
rect 1443 14433 1455 14436
rect 1397 14427 1455 14433
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 4341 14467 4399 14473
rect 2832 14436 2877 14464
rect 2832 14424 2838 14436
rect 4341 14433 4353 14467
rect 4387 14464 4399 14467
rect 4540 14464 4568 14560
rect 4608 14535 4666 14541
rect 4608 14501 4620 14535
rect 4654 14532 4666 14535
rect 4706 14532 4712 14544
rect 4654 14504 4712 14532
rect 4654 14501 4666 14504
rect 4608 14495 4666 14501
rect 4706 14492 4712 14504
rect 4764 14532 4770 14544
rect 5534 14532 5540 14544
rect 4764 14504 5540 14532
rect 4764 14492 4770 14504
rect 5534 14492 5540 14504
rect 5592 14492 5598 14544
rect 7852 14532 7880 14563
rect 11054 14560 11060 14572
rect 11112 14560 11118 14612
rect 11330 14600 11336 14612
rect 11291 14572 11336 14600
rect 11330 14560 11336 14572
rect 11388 14560 11394 14612
rect 12986 14560 12992 14612
rect 13044 14600 13050 14612
rect 13354 14600 13360 14612
rect 13044 14572 13360 14600
rect 13044 14560 13050 14572
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 13538 14600 13544 14612
rect 13499 14572 13544 14600
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 14090 14600 14096 14612
rect 14051 14572 14096 14600
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14826 14600 14832 14612
rect 14787 14572 14832 14600
rect 14826 14560 14832 14572
rect 14884 14560 14890 14612
rect 16298 14600 16304 14612
rect 16211 14572 16304 14600
rect 16298 14560 16304 14572
rect 16356 14600 16362 14612
rect 16850 14600 16856 14612
rect 16356 14572 16856 14600
rect 16356 14560 16362 14572
rect 16850 14560 16856 14572
rect 16908 14560 16914 14612
rect 18782 14600 18788 14612
rect 18743 14572 18788 14600
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 21082 14600 21088 14612
rect 21043 14572 21088 14600
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 21818 14560 21824 14612
rect 21876 14600 21882 14612
rect 21913 14603 21971 14609
rect 21913 14600 21925 14603
rect 21876 14572 21925 14600
rect 21876 14560 21882 14572
rect 21913 14569 21925 14572
rect 21959 14600 21971 14603
rect 22278 14600 22284 14612
rect 21959 14572 22284 14600
rect 21959 14569 21971 14572
rect 21913 14563 21971 14569
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 22830 14560 22836 14612
rect 22888 14600 22894 14612
rect 23106 14600 23112 14612
rect 22888 14572 23112 14600
rect 22888 14560 22894 14572
rect 23106 14560 23112 14572
rect 23164 14600 23170 14612
rect 23385 14603 23443 14609
rect 23385 14600 23397 14603
rect 23164 14572 23397 14600
rect 23164 14560 23170 14572
rect 23385 14569 23397 14572
rect 23431 14569 23443 14603
rect 24946 14600 24952 14612
rect 24907 14572 24952 14600
rect 23385 14563 23443 14569
rect 24946 14560 24952 14572
rect 25004 14560 25010 14612
rect 7852 14504 8524 14532
rect 4387 14436 4568 14464
rect 4387 14433 4399 14436
rect 4341 14427 4399 14433
rect 5626 14424 5632 14476
rect 5684 14464 5690 14476
rect 6822 14464 6828 14476
rect 5684 14436 6828 14464
rect 5684 14424 5690 14436
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 8386 14464 8392 14476
rect 8347 14436 8392 14464
rect 8386 14424 8392 14436
rect 8444 14424 8450 14476
rect 8496 14464 8524 14504
rect 12250 14492 12256 14544
rect 12308 14532 12314 14544
rect 12434 14541 12440 14544
rect 12428 14532 12440 14541
rect 12308 14504 12440 14532
rect 12308 14492 12314 14504
rect 12428 14495 12440 14504
rect 12492 14532 12498 14544
rect 14550 14532 14556 14544
rect 12492 14504 12576 14532
rect 14463 14504 14556 14532
rect 12434 14492 12440 14495
rect 12492 14492 12498 14504
rect 14550 14492 14556 14504
rect 14608 14532 14614 14544
rect 15102 14532 15108 14544
rect 14608 14504 15108 14532
rect 14608 14492 14614 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 16752 14535 16810 14541
rect 16752 14501 16764 14535
rect 16798 14532 16810 14535
rect 17770 14532 17776 14544
rect 16798 14504 17776 14532
rect 16798 14501 16810 14504
rect 16752 14495 16810 14501
rect 17770 14492 17776 14504
rect 17828 14492 17834 14544
rect 10321 14467 10379 14473
rect 8496 14436 8616 14464
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 8588 14405 8616 14436
rect 10321 14433 10333 14467
rect 10367 14464 10379 14467
rect 10778 14464 10784 14476
rect 10367 14436 10784 14464
rect 10367 14433 10379 14436
rect 10321 14427 10379 14433
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 11698 14464 11704 14476
rect 11659 14436 11704 14464
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 16390 14464 16396 14476
rect 15620 14436 16396 14464
rect 15620 14424 15626 14436
rect 16390 14424 16396 14436
rect 16448 14464 16454 14476
rect 16485 14467 16543 14473
rect 16485 14464 16497 14467
rect 16448 14436 16497 14464
rect 16448 14424 16454 14436
rect 16485 14433 16497 14436
rect 16531 14433 16543 14467
rect 18800 14464 18828 14560
rect 18874 14492 18880 14544
rect 18932 14532 18938 14544
rect 20717 14535 20775 14541
rect 18932 14504 19564 14532
rect 18932 14492 18938 14504
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 18800 14436 19349 14464
rect 16485 14427 16543 14433
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2188 14368 2973 14396
rect 2188 14356 2194 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 8573 14399 8631 14405
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 8754 14396 8760 14408
rect 8619 14368 8760 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 7006 14328 7012 14340
rect 6967 14300 7012 14328
rect 7006 14288 7012 14300
rect 7064 14288 7070 14340
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8021 14331 8079 14337
rect 8021 14328 8033 14331
rect 7892 14300 8033 14328
rect 7892 14288 7898 14300
rect 8021 14297 8033 14300
rect 8067 14297 8079 14331
rect 8496 14328 8524 14359
rect 8754 14356 8760 14368
rect 8812 14356 8818 14408
rect 10042 14356 10048 14408
rect 10100 14396 10106 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10100 14368 10425 14396
rect 10100 14356 10106 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10597 14399 10655 14405
rect 10597 14365 10609 14399
rect 10643 14396 10655 14399
rect 11054 14396 11060 14408
rect 10643 14368 11060 14396
rect 10643 14365 10655 14368
rect 10597 14359 10655 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 12158 14396 12164 14408
rect 12119 14368 12164 14396
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 17586 14356 17592 14408
rect 17644 14396 17650 14408
rect 18782 14396 18788 14408
rect 17644 14368 18788 14396
rect 17644 14356 17650 14368
rect 18782 14356 18788 14368
rect 18840 14356 18846 14408
rect 19242 14356 19248 14408
rect 19300 14396 19306 14408
rect 19536 14405 19564 14504
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 20990 14532 20996 14544
rect 20763 14504 20996 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 20990 14492 20996 14504
rect 21048 14492 21054 14544
rect 22462 14492 22468 14544
rect 22520 14492 22526 14544
rect 19610 14424 19616 14476
rect 19668 14464 19674 14476
rect 20073 14467 20131 14473
rect 20073 14464 20085 14467
rect 19668 14436 20085 14464
rect 19668 14424 19674 14436
rect 20073 14433 20085 14436
rect 20119 14464 20131 14467
rect 20901 14467 20959 14473
rect 20119 14436 20852 14464
rect 20119 14433 20131 14436
rect 20073 14427 20131 14433
rect 19429 14399 19487 14405
rect 19429 14396 19441 14399
rect 19300 14368 19441 14396
rect 19300 14356 19306 14368
rect 19429 14365 19441 14368
rect 19475 14365 19487 14399
rect 19429 14359 19487 14365
rect 19521 14399 19579 14405
rect 19521 14365 19533 14399
rect 19567 14365 19579 14399
rect 19521 14359 19579 14365
rect 20254 14356 20260 14408
rect 20312 14396 20318 14408
rect 20438 14396 20444 14408
rect 20312 14368 20444 14396
rect 20312 14356 20318 14368
rect 20438 14356 20444 14368
rect 20496 14356 20502 14408
rect 20824 14396 20852 14436
rect 20901 14433 20913 14467
rect 20947 14464 20959 14467
rect 21082 14464 21088 14476
rect 20947 14436 21088 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21082 14424 21088 14436
rect 21140 14424 21146 14476
rect 22002 14464 22008 14476
rect 21963 14436 22008 14464
rect 22002 14424 22008 14436
rect 22060 14424 22066 14476
rect 22272 14467 22330 14473
rect 22272 14433 22284 14467
rect 22318 14464 22330 14467
rect 22480 14464 22508 14492
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 22318 14436 23949 14464
rect 22318 14433 22330 14436
rect 22272 14427 22330 14433
rect 23937 14433 23949 14436
rect 23983 14464 23995 14467
rect 24210 14464 24216 14476
rect 23983 14436 24216 14464
rect 23983 14433 23995 14436
rect 23937 14427 23995 14433
rect 24210 14424 24216 14436
rect 24268 14424 24274 14476
rect 24854 14464 24860 14476
rect 24815 14436 24860 14464
rect 24854 14424 24860 14436
rect 24912 14464 24918 14476
rect 25222 14464 25228 14476
rect 24912 14436 25228 14464
rect 24912 14424 24918 14436
rect 25222 14424 25228 14436
rect 25280 14424 25286 14476
rect 22020 14396 22048 14424
rect 20824 14368 22048 14396
rect 24228 14396 24256 14424
rect 24670 14396 24676 14408
rect 24228 14368 24676 14396
rect 24670 14356 24676 14368
rect 24728 14396 24734 14408
rect 25041 14399 25099 14405
rect 25041 14396 25053 14399
rect 24728 14368 25053 14396
rect 24728 14356 24734 14368
rect 25041 14365 25053 14368
rect 25087 14365 25099 14399
rect 25041 14359 25099 14365
rect 9214 14328 9220 14340
rect 8496 14300 9220 14328
rect 8021 14291 8079 14297
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 15838 14328 15844 14340
rect 14332 14300 15844 14328
rect 14332 14288 14338 14300
rect 15838 14288 15844 14300
rect 15896 14288 15902 14340
rect 18969 14331 19027 14337
rect 18969 14297 18981 14331
rect 19015 14328 19027 14331
rect 21453 14331 21511 14337
rect 21453 14328 21465 14331
rect 19015 14300 21465 14328
rect 19015 14297 19027 14300
rect 18969 14291 19027 14297
rect 21453 14297 21465 14300
rect 21499 14328 21511 14331
rect 22002 14328 22008 14340
rect 21499 14300 22008 14328
rect 21499 14297 21511 14300
rect 21453 14291 21511 14297
rect 22002 14288 22008 14300
rect 22060 14288 22066 14340
rect 23474 14288 23480 14340
rect 23532 14328 23538 14340
rect 24026 14328 24032 14340
rect 23532 14300 24032 14328
rect 23532 14288 23538 14300
rect 24026 14288 24032 14300
rect 24084 14328 24090 14340
rect 24305 14331 24363 14337
rect 24305 14328 24317 14331
rect 24084 14300 24317 14328
rect 24084 14288 24090 14300
rect 24305 14297 24317 14300
rect 24351 14297 24363 14331
rect 24946 14328 24952 14340
rect 24305 14291 24363 14297
rect 24412 14300 24952 14328
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 1854 14260 1860 14272
rect 1627 14232 1860 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 1854 14220 1860 14232
rect 1912 14220 1918 14272
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14260 2375 14263
rect 4154 14260 4160 14272
rect 2363 14232 4160 14260
rect 2363 14229 2375 14232
rect 2317 14223 2375 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5592 14232 5733 14260
rect 5592 14220 5598 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 5721 14223 5779 14229
rect 6270 14220 6276 14272
rect 6328 14260 6334 14272
rect 6641 14263 6699 14269
rect 6641 14260 6653 14263
rect 6328 14232 6653 14260
rect 6328 14220 6334 14232
rect 6641 14229 6653 14232
rect 6687 14229 6699 14263
rect 9030 14260 9036 14272
rect 8991 14232 9036 14260
rect 6641 14223 6699 14229
rect 9030 14220 9036 14232
rect 9088 14220 9094 14272
rect 9490 14260 9496 14272
rect 9451 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9950 14260 9956 14272
rect 9911 14232 9956 14260
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 17862 14260 17868 14272
rect 17823 14232 17868 14260
rect 17862 14220 17868 14232
rect 17920 14220 17926 14272
rect 18509 14263 18567 14269
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 19518 14260 19524 14272
rect 18555 14232 19524 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20438 14260 20444 14272
rect 20128 14232 20444 14260
rect 20128 14220 20134 14232
rect 20438 14220 20444 14232
rect 20496 14220 20502 14272
rect 20530 14220 20536 14272
rect 20588 14260 20594 14272
rect 24412 14260 24440 14300
rect 24946 14288 24952 14300
rect 25004 14288 25010 14340
rect 20588 14232 24440 14260
rect 24489 14263 24547 14269
rect 20588 14220 20594 14232
rect 24489 14229 24501 14263
rect 24535 14260 24547 14263
rect 24670 14260 24676 14272
rect 24535 14232 24676 14260
rect 24535 14229 24547 14232
rect 24489 14223 24547 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 25222 14220 25228 14272
rect 25280 14260 25286 14272
rect 25501 14263 25559 14269
rect 25501 14260 25513 14263
rect 25280 14232 25513 14260
rect 25280 14220 25286 14232
rect 25501 14229 25513 14232
rect 25547 14229 25559 14263
rect 25501 14223 25559 14229
rect 1104 14170 26864 14192
rect 1104 14118 5648 14170
rect 5700 14118 5712 14170
rect 5764 14118 5776 14170
rect 5828 14118 5840 14170
rect 5892 14118 14982 14170
rect 15034 14118 15046 14170
rect 15098 14118 15110 14170
rect 15162 14118 15174 14170
rect 15226 14118 24315 14170
rect 24367 14118 24379 14170
rect 24431 14118 24443 14170
rect 24495 14118 24507 14170
rect 24559 14118 26864 14170
rect 1104 14096 26864 14118
rect 2774 14016 2780 14068
rect 2832 14056 2838 14068
rect 3234 14056 3240 14068
rect 2832 14028 3240 14056
rect 2832 14016 2838 14028
rect 3234 14016 3240 14028
rect 3292 14056 3298 14068
rect 3421 14059 3479 14065
rect 3421 14056 3433 14059
rect 3292 14028 3433 14056
rect 3292 14016 3298 14028
rect 3421 14025 3433 14028
rect 3467 14025 3479 14059
rect 3421 14019 3479 14025
rect 3694 14016 3700 14068
rect 3752 14056 3758 14068
rect 5166 14056 5172 14068
rect 3752 14028 5172 14056
rect 3752 14016 3758 14028
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 9214 14056 9220 14068
rect 9175 14028 9220 14056
rect 9214 14016 9220 14028
rect 9272 14016 9278 14068
rect 9769 14059 9827 14065
rect 9769 14025 9781 14059
rect 9815 14056 9827 14059
rect 9815 14028 10824 14056
rect 9815 14025 9827 14028
rect 9769 14019 9827 14025
rect 1581 13991 1639 13997
rect 1581 13957 1593 13991
rect 1627 13988 1639 13991
rect 2222 13988 2228 14000
rect 1627 13960 2228 13988
rect 1627 13957 1639 13960
rect 1581 13951 1639 13957
rect 2222 13948 2228 13960
rect 2280 13948 2286 14000
rect 3329 13991 3387 13997
rect 3329 13957 3341 13991
rect 3375 13988 3387 13991
rect 3510 13988 3516 14000
rect 3375 13960 3516 13988
rect 3375 13957 3387 13960
rect 3329 13951 3387 13957
rect 3510 13948 3516 13960
rect 3568 13948 3574 14000
rect 4982 13988 4988 14000
rect 3896 13960 4988 13988
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13920 2194 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2188 13892 2605 13920
rect 2188 13880 2194 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 1946 13812 1952 13864
rect 2004 13852 2010 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 2004 13824 2053 13852
rect 2004 13812 2010 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 3528 13852 3556 13948
rect 3896 13929 3924 13960
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 8570 13988 8576 14000
rect 8531 13960 8576 13988
rect 8570 13948 8576 13960
rect 8628 13948 8634 14000
rect 10796 13988 10824 14028
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11112 14028 11253 14056
rect 11112 14016 11118 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 11241 14019 11299 14025
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 12437 14059 12495 14065
rect 12437 14025 12449 14059
rect 12483 14056 12495 14059
rect 12894 14056 12900 14068
rect 12483 14028 12900 14056
rect 12483 14025 12495 14028
rect 12437 14019 12495 14025
rect 12894 14016 12900 14028
rect 12952 14016 12958 14068
rect 13446 14056 13452 14068
rect 13407 14028 13452 14056
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 16206 14056 16212 14068
rect 15795 14028 16212 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16206 14016 16212 14028
rect 16264 14016 16270 14068
rect 16390 14016 16396 14068
rect 16448 14056 16454 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16448 14028 16865 14056
rect 16448 14016 16454 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 17313 14059 17371 14065
rect 17313 14025 17325 14059
rect 17359 14056 17371 14059
rect 17770 14056 17776 14068
rect 17359 14028 17776 14056
rect 17359 14025 17371 14028
rect 17313 14019 17371 14025
rect 12176 13988 12204 14016
rect 10796 13960 12204 13988
rect 3881 13923 3939 13929
rect 3881 13889 3893 13923
rect 3927 13889 3939 13923
rect 3881 13883 3939 13889
rect 3973 13923 4031 13929
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 3988 13852 4016 13883
rect 4154 13880 4160 13932
rect 4212 13920 4218 13932
rect 5629 13923 5687 13929
rect 5629 13920 5641 13923
rect 4212 13892 5641 13920
rect 4212 13880 4218 13892
rect 5629 13889 5641 13892
rect 5675 13920 5687 13923
rect 5997 13923 6055 13929
rect 5997 13920 6009 13923
rect 5675 13892 6009 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5997 13889 6009 13892
rect 6043 13889 6055 13923
rect 5997 13883 6055 13889
rect 6917 13923 6975 13929
rect 6917 13889 6929 13923
rect 6963 13920 6975 13923
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6963 13892 7205 13920
rect 6963 13889 6975 13892
rect 6917 13883 6975 13889
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 9030 13880 9036 13932
rect 9088 13880 9094 13932
rect 3528 13824 4016 13852
rect 4893 13855 4951 13861
rect 2041 13815 2099 13821
rect 4893 13821 4905 13855
rect 4939 13852 4951 13855
rect 5442 13852 5448 13864
rect 4939 13824 5448 13852
rect 4939 13821 4951 13824
rect 4893 13815 4951 13821
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 6270 13812 6276 13864
rect 6328 13852 6334 13864
rect 7449 13855 7507 13861
rect 7449 13852 7461 13855
rect 6328 13824 7461 13852
rect 6328 13812 6334 13824
rect 7449 13821 7461 13824
rect 7495 13852 7507 13855
rect 7834 13852 7840 13864
rect 7495 13824 7840 13852
rect 7495 13821 7507 13824
rect 7449 13815 7507 13821
rect 7834 13812 7840 13824
rect 7892 13812 7898 13864
rect 9048 13852 9076 13880
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 7944 13824 9873 13852
rect 4525 13787 4583 13793
rect 4525 13753 4537 13787
rect 4571 13784 4583 13787
rect 4614 13784 4620 13796
rect 4571 13756 4620 13784
rect 4571 13753 4583 13756
rect 4525 13747 4583 13753
rect 4614 13744 4620 13756
rect 4672 13784 4678 13796
rect 5350 13784 5356 13796
rect 4672 13756 5356 13784
rect 4672 13744 4678 13756
rect 5350 13744 5356 13756
rect 5408 13744 5414 13796
rect 6454 13744 6460 13796
rect 6512 13784 6518 13796
rect 6917 13787 6975 13793
rect 6917 13784 6929 13787
rect 6512 13756 6929 13784
rect 6512 13744 6518 13756
rect 6917 13753 6929 13756
rect 6963 13784 6975 13787
rect 7009 13787 7067 13793
rect 7009 13784 7021 13787
rect 6963 13756 7021 13784
rect 6963 13753 6975 13756
rect 6917 13747 6975 13753
rect 7009 13753 7021 13756
rect 7055 13784 7067 13787
rect 7944 13784 7972 13824
rect 9861 13821 9873 13824
rect 9907 13852 9919 13855
rect 10888 13852 10916 13960
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12434 13920 12440 13932
rect 11931 13892 12440 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12434 13880 12440 13892
rect 12492 13920 12498 13932
rect 12986 13920 12992 13932
rect 12492 13892 12992 13920
rect 12492 13880 12498 13892
rect 12986 13880 12992 13892
rect 13044 13920 13050 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 13044 13892 13093 13920
rect 13044 13880 13050 13892
rect 13081 13889 13093 13892
rect 13127 13889 13139 13923
rect 13081 13883 13139 13889
rect 13446 13880 13452 13932
rect 13504 13920 13510 13932
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 13504 13892 14565 13920
rect 13504 13880 13510 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 15427 13892 16405 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 16393 13889 16405 13892
rect 16439 13920 16451 13923
rect 17328 13920 17356 14019
rect 17770 14016 17776 14028
rect 17828 14016 17834 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 19242 14056 19248 14068
rect 19107 14028 19248 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 19242 14016 19248 14028
rect 19300 14016 19306 14068
rect 20530 14056 20536 14068
rect 19352 14028 20536 14056
rect 19352 13988 19380 14028
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 20622 14016 20628 14068
rect 20680 14056 20686 14068
rect 20717 14059 20775 14065
rect 20717 14056 20729 14059
rect 20680 14028 20729 14056
rect 20680 14016 20686 14028
rect 20717 14025 20729 14028
rect 20763 14025 20775 14059
rect 20717 14019 20775 14025
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21269 14059 21327 14065
rect 21269 14056 21281 14059
rect 21140 14028 21281 14056
rect 21140 14016 21146 14028
rect 21269 14025 21281 14028
rect 21315 14025 21327 14059
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 21269 14019 21327 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 22094 14016 22100 14068
rect 22152 14056 22158 14068
rect 22833 14059 22891 14065
rect 22833 14056 22845 14059
rect 22152 14028 22845 14056
rect 22152 14016 22158 14028
rect 22833 14025 22845 14028
rect 22879 14025 22891 14059
rect 22833 14019 22891 14025
rect 23290 14016 23296 14068
rect 23348 14056 23354 14068
rect 23385 14059 23443 14065
rect 23385 14056 23397 14059
rect 23348 14028 23397 14056
rect 23348 14016 23354 14028
rect 23385 14025 23397 14028
rect 23431 14025 23443 14059
rect 23385 14019 23443 14025
rect 16439 13892 17356 13920
rect 17972 13960 19380 13988
rect 16439 13889 16451 13892
rect 16393 13883 16451 13889
rect 12894 13852 12900 13864
rect 9907 13824 10916 13852
rect 12855 13824 12900 13852
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 12894 13812 12900 13824
rect 12952 13812 12958 13864
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 14461 13855 14519 13861
rect 14461 13852 14473 13855
rect 13872 13824 14473 13852
rect 13872 13812 13878 13824
rect 14461 13821 14473 13824
rect 14507 13852 14519 13855
rect 14918 13852 14924 13864
rect 14507 13824 14924 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15838 13812 15844 13864
rect 15896 13852 15902 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15896 13824 16221 13852
rect 15896 13812 15902 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16298 13812 16304 13864
rect 16356 13852 16362 13864
rect 16356 13824 16401 13852
rect 16356 13812 16362 13824
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 16540 13824 17785 13852
rect 16540 13812 16546 13824
rect 17773 13821 17785 13824
rect 17819 13852 17831 13855
rect 17862 13852 17868 13864
rect 17819 13824 17868 13852
rect 17819 13821 17831 13824
rect 17773 13815 17831 13821
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 17972 13796 18000 13960
rect 19334 13920 19340 13932
rect 19295 13892 19340 13920
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21729 13923 21787 13929
rect 21729 13920 21741 13923
rect 20772 13892 21741 13920
rect 20772 13880 20778 13892
rect 21729 13889 21741 13892
rect 21775 13920 21787 13923
rect 22373 13923 22431 13929
rect 22373 13920 22385 13923
rect 21775 13892 22385 13920
rect 21775 13889 21787 13892
rect 21729 13883 21787 13889
rect 22373 13889 22385 13892
rect 22419 13889 22431 13923
rect 22373 13883 22431 13889
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22189 13855 22247 13861
rect 22189 13852 22201 13855
rect 22152 13824 22201 13852
rect 22152 13812 22158 13824
rect 22189 13821 22201 13824
rect 22235 13821 22247 13855
rect 22189 13815 22247 13821
rect 22830 13812 22836 13864
rect 22888 13852 22894 13864
rect 23400 13852 23428 14019
rect 24026 14016 24032 14068
rect 24084 14056 24090 14068
rect 24673 14059 24731 14065
rect 24673 14056 24685 14059
rect 24084 14028 24685 14056
rect 24084 14016 24090 14028
rect 24673 14025 24685 14028
rect 24719 14056 24731 14059
rect 24854 14056 24860 14068
rect 24719 14028 24860 14056
rect 24719 14025 24731 14028
rect 24673 14019 24731 14025
rect 24854 14016 24860 14028
rect 24912 14016 24918 14068
rect 24946 14016 24952 14068
rect 25004 14056 25010 14068
rect 25041 14059 25099 14065
rect 25041 14056 25053 14059
rect 25004 14028 25053 14056
rect 25004 14016 25010 14028
rect 25041 14025 25053 14028
rect 25087 14025 25099 14059
rect 25041 14019 25099 14025
rect 25409 14059 25467 14065
rect 25409 14025 25421 14059
rect 25455 14056 25467 14059
rect 25498 14056 25504 14068
rect 25455 14028 25504 14056
rect 25455 14025 25467 14028
rect 25409 14019 25467 14025
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 23474 13948 23480 14000
rect 23532 13988 23538 14000
rect 23661 13991 23719 13997
rect 23661 13988 23673 13991
rect 23532 13960 23673 13988
rect 23532 13948 23538 13960
rect 23661 13957 23673 13960
rect 23707 13957 23719 13991
rect 23661 13951 23719 13957
rect 24210 13920 24216 13932
rect 24171 13892 24216 13920
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 24121 13855 24179 13861
rect 24121 13852 24133 13855
rect 22888 13824 24133 13852
rect 22888 13812 22894 13824
rect 24121 13821 24133 13824
rect 24167 13821 24179 13855
rect 24121 13815 24179 13821
rect 24854 13812 24860 13864
rect 24912 13852 24918 13864
rect 25225 13855 25283 13861
rect 25225 13852 25237 13855
rect 24912 13824 25237 13852
rect 24912 13812 24918 13824
rect 25225 13821 25237 13824
rect 25271 13852 25283 13855
rect 25777 13855 25835 13861
rect 25777 13852 25789 13855
rect 25271 13824 25789 13852
rect 25271 13821 25283 13824
rect 25225 13815 25283 13821
rect 25777 13821 25789 13824
rect 25823 13821 25835 13855
rect 26234 13852 26240 13864
rect 26195 13824 26240 13852
rect 25777 13815 25835 13821
rect 26234 13812 26240 13824
rect 26292 13812 26298 13864
rect 7055 13756 7972 13784
rect 7055 13753 7067 13756
rect 7009 13747 7067 13753
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 10106 13787 10164 13793
rect 10106 13784 10118 13787
rect 9548 13756 10118 13784
rect 9548 13744 9554 13756
rect 10106 13753 10118 13756
rect 10152 13753 10164 13787
rect 10106 13747 10164 13753
rect 10594 13744 10600 13796
rect 10652 13784 10658 13796
rect 11054 13784 11060 13796
rect 10652 13756 11060 13784
rect 10652 13744 10658 13756
rect 11054 13744 11060 13756
rect 11112 13744 11118 13796
rect 12526 13744 12532 13796
rect 12584 13784 12590 13796
rect 12805 13787 12863 13793
rect 12805 13784 12817 13787
rect 12584 13756 12817 13784
rect 12584 13744 12590 13756
rect 12805 13753 12817 13756
rect 12851 13784 12863 13787
rect 13722 13784 13728 13796
rect 12851 13756 13728 13784
rect 12851 13753 12863 13756
rect 12805 13747 12863 13753
rect 13722 13744 13728 13756
rect 13780 13744 13786 13796
rect 14369 13787 14427 13793
rect 14369 13784 14381 13787
rect 13924 13756 14381 13784
rect 13924 13728 13952 13756
rect 14369 13753 14381 13756
rect 14415 13753 14427 13787
rect 14369 13747 14427 13753
rect 16022 13744 16028 13796
rect 16080 13784 16086 13796
rect 17954 13784 17960 13796
rect 16080 13756 17960 13784
rect 16080 13744 16086 13756
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 19518 13744 19524 13796
rect 19576 13793 19582 13796
rect 19576 13787 19640 13793
rect 19576 13753 19594 13787
rect 19628 13753 19640 13787
rect 19576 13747 19640 13753
rect 22281 13787 22339 13793
rect 22281 13753 22293 13787
rect 22327 13784 22339 13787
rect 22370 13784 22376 13796
rect 22327 13756 22376 13784
rect 22327 13753 22339 13756
rect 22281 13747 22339 13753
rect 19576 13744 19582 13747
rect 22370 13744 22376 13756
rect 22428 13744 22434 13796
rect 23014 13744 23020 13796
rect 23072 13784 23078 13796
rect 23072 13756 25268 13784
rect 23072 13744 23078 13756
rect 25240 13728 25268 13756
rect 1762 13676 1768 13728
rect 1820 13716 1826 13728
rect 1949 13719 2007 13725
rect 1949 13716 1961 13719
rect 1820 13688 1961 13716
rect 1820 13676 1826 13688
rect 1949 13685 1961 13688
rect 1995 13716 2007 13719
rect 2314 13716 2320 13728
rect 1995 13688 2320 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 2590 13676 2596 13728
rect 2648 13716 2654 13728
rect 3786 13716 3792 13728
rect 2648 13688 3792 13716
rect 2648 13676 2654 13688
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 6546 13716 6552 13728
rect 6507 13688 6552 13716
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 13262 13676 13268 13728
rect 13320 13716 13326 13728
rect 13906 13716 13912 13728
rect 13320 13688 13912 13716
rect 13320 13676 13326 13688
rect 13906 13676 13912 13688
rect 13964 13676 13970 13728
rect 14001 13719 14059 13725
rect 14001 13685 14013 13719
rect 14047 13716 14059 13719
rect 14182 13716 14188 13728
rect 14047 13688 14188 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 14182 13676 14188 13688
rect 14240 13676 14246 13728
rect 15838 13716 15844 13728
rect 15799 13688 15844 13716
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 18322 13716 18328 13728
rect 18283 13688 18328 13716
rect 18322 13676 18328 13688
rect 18380 13676 18386 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 21910 13716 21916 13728
rect 19208 13688 21916 13716
rect 19208 13676 19214 13688
rect 21910 13676 21916 13688
rect 21968 13676 21974 13728
rect 22094 13676 22100 13728
rect 22152 13716 22158 13728
rect 22462 13716 22468 13728
rect 22152 13688 22468 13716
rect 22152 13676 22158 13688
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 23566 13676 23572 13728
rect 23624 13716 23630 13728
rect 24029 13719 24087 13725
rect 24029 13716 24041 13719
rect 23624 13688 24041 13716
rect 23624 13676 23630 13688
rect 24029 13685 24041 13688
rect 24075 13685 24087 13719
rect 24029 13679 24087 13685
rect 25222 13676 25228 13728
rect 25280 13676 25286 13728
rect 1104 13626 26864 13648
rect 1104 13574 10315 13626
rect 10367 13574 10379 13626
rect 10431 13574 10443 13626
rect 10495 13574 10507 13626
rect 10559 13574 19648 13626
rect 19700 13574 19712 13626
rect 19764 13574 19776 13626
rect 19828 13574 19840 13626
rect 19892 13574 26864 13626
rect 1104 13552 26864 13574
rect 1673 13515 1731 13521
rect 1673 13481 1685 13515
rect 1719 13512 1731 13515
rect 2130 13512 2136 13524
rect 1719 13484 2136 13512
rect 1719 13481 1731 13484
rect 1673 13475 1731 13481
rect 2130 13472 2136 13484
rect 2188 13472 2194 13524
rect 2317 13515 2375 13521
rect 2317 13481 2329 13515
rect 2363 13512 2375 13515
rect 2406 13512 2412 13524
rect 2363 13484 2412 13512
rect 2363 13481 2375 13484
rect 2317 13475 2375 13481
rect 2406 13472 2412 13484
rect 2464 13472 2470 13524
rect 3234 13512 3240 13524
rect 3195 13484 3240 13512
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 4706 13512 4712 13524
rect 4667 13484 4712 13512
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 4890 13512 4896 13524
rect 4851 13484 4896 13512
rect 4890 13472 4896 13484
rect 4948 13472 4954 13524
rect 7834 13512 7840 13524
rect 7795 13484 7840 13512
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8754 13512 8760 13524
rect 8715 13484 8760 13512
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 9490 13512 9496 13524
rect 9451 13484 9496 13512
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 11330 13512 11336 13524
rect 10008 13484 11336 13512
rect 10008 13472 10014 13484
rect 11330 13472 11336 13484
rect 11388 13512 11394 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11388 13484 11621 13512
rect 11388 13472 11394 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 13630 13512 13636 13524
rect 11609 13475 11667 13481
rect 11808 13484 13636 13512
rect 2682 13404 2688 13456
rect 2740 13444 2746 13456
rect 2961 13447 3019 13453
rect 2961 13444 2973 13447
rect 2740 13416 2973 13444
rect 2740 13404 2746 13416
rect 2961 13413 2973 13416
rect 3007 13444 3019 13447
rect 4724 13444 4752 13472
rect 3007 13416 4752 13444
rect 3007 13413 3019 13416
rect 2961 13407 3019 13413
rect 4982 13404 4988 13456
rect 5040 13444 5046 13456
rect 5353 13447 5411 13453
rect 5353 13444 5365 13447
rect 5040 13416 5365 13444
rect 5040 13404 5046 13416
rect 5353 13413 5365 13416
rect 5399 13413 5411 13447
rect 5353 13407 5411 13413
rect 6546 13404 6552 13456
rect 6604 13444 6610 13456
rect 6702 13447 6760 13453
rect 6702 13444 6714 13447
rect 6604 13416 6714 13444
rect 6604 13404 6610 13416
rect 6702 13413 6714 13416
rect 6748 13413 6760 13447
rect 9508 13444 9536 13472
rect 9508 13416 10180 13444
rect 6702 13407 6760 13413
rect 2222 13376 2228 13388
rect 2183 13348 2228 13376
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 3602 13336 3608 13388
rect 3660 13376 3666 13388
rect 5258 13376 5264 13388
rect 3660 13348 5264 13376
rect 3660 13336 3666 13348
rect 5258 13336 5264 13348
rect 5316 13336 5322 13388
rect 5994 13376 6000 13388
rect 5368 13348 6000 13376
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 3050 13308 3056 13320
rect 2547 13280 3056 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 3050 13268 3056 13280
rect 3108 13308 3114 13320
rect 3418 13308 3424 13320
rect 3108 13280 3424 13308
rect 3108 13268 3114 13280
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4522 13308 4528 13320
rect 4212 13280 4528 13308
rect 4212 13268 4218 13280
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4706 13268 4712 13320
rect 4764 13308 4770 13320
rect 5368 13308 5396 13348
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 10045 13379 10103 13385
rect 10045 13376 10057 13379
rect 9824 13348 10057 13376
rect 9824 13336 9830 13348
rect 10045 13345 10057 13348
rect 10091 13345 10103 13379
rect 10152 13376 10180 13416
rect 10594 13376 10600 13388
rect 10152 13348 10600 13376
rect 10045 13339 10103 13345
rect 4764 13280 5396 13308
rect 4764 13268 4770 13280
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 6454 13308 6460 13320
rect 5500 13280 5545 13308
rect 6415 13280 6460 13308
rect 5500 13268 5506 13280
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 9582 13268 9588 13320
rect 9640 13308 9646 13320
rect 10244 13317 10272 13348
rect 10594 13336 10600 13348
rect 10652 13376 10658 13388
rect 10689 13379 10747 13385
rect 10689 13376 10701 13379
rect 10652 13348 10701 13376
rect 10652 13336 10658 13348
rect 10689 13345 10701 13348
rect 10735 13376 10747 13379
rect 11057 13379 11115 13385
rect 11057 13376 11069 13379
rect 10735 13348 11069 13376
rect 10735 13345 10747 13348
rect 10689 13339 10747 13345
rect 11057 13345 11069 13348
rect 11103 13376 11115 13379
rect 11103 13348 11560 13376
rect 11103 13345 11115 13348
rect 11057 13339 11115 13345
rect 10137 13311 10195 13317
rect 10137 13308 10149 13311
rect 9640 13280 10149 13308
rect 9640 13268 9646 13280
rect 10137 13277 10149 13280
rect 10183 13277 10195 13311
rect 10137 13271 10195 13277
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 1394 13200 1400 13252
rect 1452 13240 1458 13252
rect 1857 13243 1915 13249
rect 1857 13240 1869 13243
rect 1452 13212 1869 13240
rect 1452 13200 1458 13212
rect 1857 13209 1869 13212
rect 1903 13209 1915 13243
rect 1857 13203 1915 13209
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 3605 13243 3663 13249
rect 3605 13240 3617 13243
rect 2004 13212 3617 13240
rect 2004 13200 2010 13212
rect 3605 13209 3617 13212
rect 3651 13209 3663 13243
rect 3605 13203 3663 13209
rect 4433 13243 4491 13249
rect 4433 13209 4445 13243
rect 4479 13240 4491 13243
rect 6472 13240 6500 13268
rect 4479 13212 6500 13240
rect 4479 13209 4491 13212
rect 4433 13203 4491 13209
rect 8386 13200 8392 13252
rect 8444 13240 8450 13252
rect 8481 13243 8539 13249
rect 8481 13240 8493 13243
rect 8444 13212 8493 13240
rect 8444 13200 8450 13212
rect 8481 13209 8493 13212
rect 8527 13240 8539 13243
rect 9030 13240 9036 13252
rect 8527 13212 9036 13240
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 9030 13200 9036 13212
rect 9088 13200 9094 13252
rect 11238 13240 11244 13252
rect 11199 13212 11244 13240
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 11532 13240 11560 13348
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11808 13317 11836 13484
rect 13630 13472 13636 13484
rect 13688 13512 13694 13524
rect 13909 13515 13967 13521
rect 13909 13512 13921 13515
rect 13688 13484 13921 13512
rect 13688 13472 13694 13484
rect 13909 13481 13921 13484
rect 13955 13512 13967 13515
rect 14090 13512 14096 13524
rect 13955 13484 14096 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14090 13472 14096 13484
rect 14148 13472 14154 13524
rect 14550 13512 14556 13524
rect 14511 13484 14556 13512
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 15838 13512 15844 13524
rect 15799 13484 15844 13512
rect 15838 13472 15844 13484
rect 15896 13512 15902 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 15896 13484 16405 13512
rect 15896 13472 15902 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 17310 13512 17316 13524
rect 17271 13484 17316 13512
rect 16393 13475 16451 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 17862 13512 17868 13524
rect 17823 13484 17868 13512
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 18230 13512 18236 13524
rect 18191 13484 18236 13512
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 20898 13512 20904 13524
rect 20859 13484 20904 13512
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 21542 13512 21548 13524
rect 21407 13484 21548 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 12529 13447 12587 13453
rect 12529 13413 12541 13447
rect 12575 13444 12587 13447
rect 12986 13444 12992 13456
rect 12575 13416 12992 13444
rect 12575 13413 12587 13416
rect 12529 13407 12587 13413
rect 12986 13404 12992 13416
rect 13044 13444 13050 13456
rect 20349 13447 20407 13453
rect 13044 13416 14596 13444
rect 13044 13404 13050 13416
rect 14568 13388 14596 13416
rect 20349 13413 20361 13447
rect 20395 13444 20407 13447
rect 21376 13444 21404 13475
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 22557 13515 22615 13521
rect 22557 13481 22569 13515
rect 22603 13512 22615 13515
rect 23382 13512 23388 13524
rect 22603 13484 23388 13512
rect 22603 13481 22615 13484
rect 22557 13475 22615 13481
rect 23382 13472 23388 13484
rect 23440 13472 23446 13524
rect 23750 13472 23756 13524
rect 23808 13512 23814 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 23808 13484 24593 13512
rect 23808 13472 23814 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 23014 13444 23020 13456
rect 20395 13416 21404 13444
rect 22975 13416 23020 13444
rect 20395 13413 20407 13416
rect 20349 13407 20407 13413
rect 23014 13404 23020 13416
rect 23072 13404 23078 13456
rect 23566 13404 23572 13456
rect 23624 13444 23630 13456
rect 23661 13447 23719 13453
rect 23661 13444 23673 13447
rect 23624 13416 23673 13444
rect 23624 13404 23630 13416
rect 23661 13413 23673 13416
rect 23707 13413 23719 13447
rect 23661 13407 23719 13413
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 12802 13376 12808 13388
rect 12492 13348 12808 13376
rect 12492 13336 12498 13348
rect 12802 13336 12808 13348
rect 12860 13336 12866 13388
rect 13173 13379 13231 13385
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 14090 13376 14096 13388
rect 13219 13348 14096 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14550 13336 14556 13388
rect 14608 13336 14614 13388
rect 16298 13376 16304 13388
rect 16259 13348 16304 13376
rect 16298 13336 16304 13348
rect 16356 13336 16362 13388
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 18581 13379 18639 13385
rect 18581 13376 18593 13379
rect 18472 13348 18593 13376
rect 18472 13336 18478 13348
rect 18581 13345 18593 13348
rect 18627 13345 18639 13379
rect 18581 13339 18639 13345
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21266 13376 21272 13388
rect 20680 13348 21272 13376
rect 20680 13336 20686 13348
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 21542 13336 21548 13388
rect 21600 13376 21606 13388
rect 22186 13376 22192 13388
rect 21600 13348 22192 13376
rect 21600 13336 21606 13348
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 22370 13376 22376 13388
rect 22331 13348 22376 13376
rect 22370 13336 22376 13348
rect 22428 13336 22434 13388
rect 22830 13336 22836 13388
rect 22888 13376 22894 13388
rect 22925 13379 22983 13385
rect 22925 13376 22937 13379
rect 22888 13348 22937 13376
rect 22888 13336 22894 13348
rect 22925 13345 22937 13348
rect 22971 13376 22983 13379
rect 23474 13376 23480 13388
rect 22971 13348 23480 13376
rect 22971 13345 22983 13348
rect 22925 13339 22983 13345
rect 23474 13336 23480 13348
rect 23532 13336 23538 13388
rect 24489 13379 24547 13385
rect 24489 13345 24501 13379
rect 24535 13376 24547 13379
rect 24762 13376 24768 13388
rect 24535 13348 24768 13376
rect 24535 13345 24547 13348
rect 24489 13339 24547 13345
rect 24762 13336 24768 13348
rect 24820 13336 24826 13388
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13277 11851 13311
rect 11793 13271 11851 13277
rect 11808 13240 11836 13271
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12986 13308 12992 13320
rect 12676 13280 12992 13308
rect 12676 13268 12682 13280
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13262 13308 13268 13320
rect 13223 13280 13268 13308
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 13446 13308 13452 13320
rect 13407 13280 13452 13308
rect 13446 13268 13452 13280
rect 13504 13268 13510 13320
rect 16482 13308 16488 13320
rect 16443 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 18046 13268 18052 13320
rect 18104 13308 18110 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 18104 13280 18337 13308
rect 18104 13268 18110 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 20806 13268 20812 13320
rect 20864 13308 20870 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 20864 13280 21465 13308
rect 20864 13268 20870 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 22646 13268 22652 13320
rect 22704 13268 22710 13320
rect 23106 13308 23112 13320
rect 23067 13280 23112 13308
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 24210 13268 24216 13320
rect 24268 13308 24274 13320
rect 24673 13311 24731 13317
rect 24673 13308 24685 13311
rect 24268 13280 24685 13308
rect 24268 13268 24274 13280
rect 24673 13277 24685 13280
rect 24719 13308 24731 13311
rect 25133 13311 25191 13317
rect 25133 13308 25145 13311
rect 24719 13280 25145 13308
rect 24719 13277 24731 13280
rect 24673 13271 24731 13277
rect 25133 13277 25145 13280
rect 25179 13277 25191 13311
rect 25590 13308 25596 13320
rect 25133 13271 25191 13277
rect 25332 13280 25596 13308
rect 11532 13212 11836 13240
rect 12342 13200 12348 13252
rect 12400 13240 12406 13252
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 12400 13212 14197 13240
rect 12400 13200 12406 13212
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 14826 13240 14832 13252
rect 14185 13203 14243 13209
rect 14568 13212 14832 13240
rect 5994 13172 6000 13184
rect 5907 13144 6000 13172
rect 5994 13132 6000 13144
rect 6052 13172 6058 13184
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 6052 13144 6285 13172
rect 6052 13132 6058 13144
rect 6273 13141 6285 13144
rect 6319 13141 6331 13175
rect 6273 13135 6331 13141
rect 9677 13175 9735 13181
rect 9677 13141 9689 13175
rect 9723 13172 9735 13175
rect 10778 13172 10784 13184
rect 9723 13144 10784 13172
rect 9723 13141 9735 13144
rect 9677 13135 9735 13141
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 12805 13175 12863 13181
rect 12805 13141 12817 13175
rect 12851 13172 12863 13175
rect 14568 13172 14596 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 15930 13240 15936 13252
rect 15891 13212 15936 13240
rect 15930 13200 15936 13212
rect 15988 13200 15994 13252
rect 22664 13240 22692 13268
rect 23014 13240 23020 13252
rect 22664 13212 23020 13240
rect 23014 13200 23020 13212
rect 23072 13200 23078 13252
rect 12851 13144 14596 13172
rect 12851 13141 12863 13144
rect 12805 13135 12863 13141
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14700 13144 14933 13172
rect 14700 13132 14706 13144
rect 14921 13141 14933 13144
rect 14967 13141 14979 13175
rect 17034 13172 17040 13184
rect 16995 13144 17040 13172
rect 14921 13135 14979 13141
rect 17034 13132 17040 13144
rect 17092 13132 17098 13184
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 19702 13172 19708 13184
rect 19576 13144 19708 13172
rect 19576 13132 19582 13144
rect 19702 13132 19708 13144
rect 19760 13132 19766 13184
rect 20714 13172 20720 13184
rect 20675 13144 20720 13172
rect 20714 13132 20720 13144
rect 20772 13132 20778 13184
rect 22094 13172 22100 13184
rect 22055 13144 22100 13172
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 22646 13132 22652 13184
rect 22704 13172 22710 13184
rect 24121 13175 24179 13181
rect 24121 13172 24133 13175
rect 22704 13144 24133 13172
rect 22704 13132 22710 13144
rect 24121 13141 24133 13144
rect 24167 13141 24179 13175
rect 24121 13135 24179 13141
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 25332 13172 25360 13280
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 25498 13172 25504 13184
rect 25096 13144 25360 13172
rect 25459 13144 25504 13172
rect 25096 13132 25102 13144
rect 25498 13132 25504 13144
rect 25556 13132 25562 13184
rect 25590 13132 25596 13184
rect 25648 13172 25654 13184
rect 25869 13175 25927 13181
rect 25869 13172 25881 13175
rect 25648 13144 25881 13172
rect 25648 13132 25654 13144
rect 25869 13141 25881 13144
rect 25915 13141 25927 13175
rect 26234 13172 26240 13184
rect 26195 13144 26240 13172
rect 25869 13135 25927 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 1104 13082 26864 13104
rect 1104 13030 5648 13082
rect 5700 13030 5712 13082
rect 5764 13030 5776 13082
rect 5828 13030 5840 13082
rect 5892 13030 14982 13082
rect 15034 13030 15046 13082
rect 15098 13030 15110 13082
rect 15162 13030 15174 13082
rect 15226 13030 24315 13082
rect 24367 13030 24379 13082
rect 24431 13030 24443 13082
rect 24495 13030 24507 13082
rect 24559 13030 26864 13082
rect 1104 13008 26864 13030
rect 290 12928 296 12980
rect 348 12968 354 12980
rect 1857 12971 1915 12977
rect 1857 12968 1869 12971
rect 348 12940 1869 12968
rect 348 12928 354 12940
rect 1857 12937 1869 12940
rect 1903 12937 1915 12971
rect 2038 12968 2044 12980
rect 1999 12940 2044 12968
rect 1857 12931 1915 12937
rect 1872 12832 1900 12931
rect 2038 12928 2044 12940
rect 2096 12968 2102 12980
rect 2774 12968 2780 12980
rect 2096 12940 2780 12968
rect 2096 12928 2102 12940
rect 2774 12928 2780 12940
rect 2832 12928 2838 12980
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 3602 12968 3608 12980
rect 3563 12940 3608 12968
rect 3602 12928 3608 12940
rect 3660 12928 3666 12980
rect 4893 12971 4951 12977
rect 4893 12968 4905 12971
rect 3712 12940 4905 12968
rect 3712 12900 3740 12940
rect 4893 12937 4905 12940
rect 4939 12968 4951 12971
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4939 12940 4997 12968
rect 4939 12937 4951 12940
rect 4893 12931 4951 12937
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 8386 12968 8392 12980
rect 8347 12940 8392 12968
rect 4985 12931 5043 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8478 12928 8484 12980
rect 8536 12968 8542 12980
rect 8846 12968 8852 12980
rect 8536 12940 8852 12968
rect 8536 12928 8542 12940
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 9950 12968 9956 12980
rect 9911 12940 9956 12968
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 11333 12971 11391 12977
rect 11333 12937 11345 12971
rect 11379 12968 11391 12971
rect 11422 12968 11428 12980
rect 11379 12940 11428 12968
rect 11379 12937 11391 12940
rect 11333 12931 11391 12937
rect 11422 12928 11428 12940
rect 11480 12968 11486 12980
rect 11698 12968 11704 12980
rect 11480 12940 11704 12968
rect 11480 12928 11486 12940
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12894 12968 12900 12980
rect 12807 12940 12900 12968
rect 12894 12928 12900 12940
rect 12952 12968 12958 12980
rect 13262 12968 13268 12980
rect 12952 12940 13268 12968
rect 12952 12928 12958 12940
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 13814 12968 13820 12980
rect 13372 12940 13820 12968
rect 2516 12872 3740 12900
rect 4709 12903 4767 12909
rect 2516 12841 2544 12872
rect 4709 12869 4721 12903
rect 4755 12900 4767 12903
rect 5442 12900 5448 12912
rect 4755 12872 5448 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 5442 12860 5448 12872
rect 5500 12860 5506 12912
rect 5552 12872 5764 12900
rect 2501 12835 2559 12841
rect 2501 12832 2513 12835
rect 1872 12804 2513 12832
rect 2501 12801 2513 12804
rect 2547 12801 2559 12835
rect 2682 12832 2688 12844
rect 2643 12804 2688 12832
rect 2501 12795 2559 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 3970 12792 3976 12844
rect 4028 12832 4034 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 4028 12804 4077 12832
rect 4028 12792 4034 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12764 3571 12767
rect 3878 12764 3884 12776
rect 3559 12736 3884 12764
rect 3559 12733 3571 12736
rect 3513 12727 3571 12733
rect 3878 12724 3884 12736
rect 3936 12764 3942 12776
rect 4172 12764 4200 12795
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4982 12832 4988 12844
rect 4304 12804 4988 12832
rect 4304 12792 4310 12804
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5552 12832 5580 12872
rect 5224 12804 5580 12832
rect 5224 12792 5230 12804
rect 3936 12736 4200 12764
rect 4893 12767 4951 12773
rect 3936 12724 3942 12736
rect 4893 12733 4905 12767
rect 4939 12764 4951 12767
rect 5736 12764 5764 12872
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 6454 12900 6460 12912
rect 6236 12872 6460 12900
rect 6236 12860 6242 12872
rect 6454 12860 6460 12872
rect 6512 12860 6518 12912
rect 7190 12860 7196 12912
rect 7248 12860 7254 12912
rect 8113 12903 8171 12909
rect 8113 12869 8125 12903
rect 8159 12900 8171 12903
rect 9401 12903 9459 12909
rect 9401 12900 9413 12903
rect 8159 12872 9413 12900
rect 8159 12869 8171 12872
rect 8113 12863 8171 12869
rect 9401 12869 9413 12872
rect 9447 12900 9459 12903
rect 9582 12900 9588 12912
rect 9447 12872 9588 12900
rect 9447 12869 9459 12872
rect 9401 12863 9459 12869
rect 9582 12860 9588 12872
rect 9640 12860 9646 12912
rect 12989 12903 13047 12909
rect 12989 12869 13001 12903
rect 13035 12900 13047 12903
rect 13372 12900 13400 12940
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 14090 12968 14096 12980
rect 14003 12940 14096 12968
rect 14090 12928 14096 12940
rect 14148 12968 14154 12980
rect 15286 12968 15292 12980
rect 14148 12940 15292 12968
rect 14148 12928 14154 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 15562 12968 15568 12980
rect 15523 12940 15568 12968
rect 15562 12928 15568 12940
rect 15620 12928 15626 12980
rect 16022 12968 16028 12980
rect 15935 12940 16028 12968
rect 16022 12928 16028 12940
rect 16080 12968 16086 12980
rect 16298 12968 16304 12980
rect 16080 12940 16304 12968
rect 16080 12928 16086 12940
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 19978 12968 19984 12980
rect 18656 12940 19984 12968
rect 18656 12928 18662 12940
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 20901 12971 20959 12977
rect 20901 12968 20913 12971
rect 20864 12940 20913 12968
rect 20864 12928 20870 12940
rect 20901 12937 20913 12940
rect 20947 12937 20959 12971
rect 21726 12968 21732 12980
rect 21687 12940 21732 12968
rect 20901 12931 20959 12937
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 22833 12971 22891 12977
rect 22833 12937 22845 12971
rect 22879 12968 22891 12971
rect 23106 12968 23112 12980
rect 22879 12940 23112 12968
rect 22879 12937 22891 12940
rect 22833 12931 22891 12937
rect 13035 12872 13400 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 13446 12860 13452 12912
rect 13504 12900 13510 12912
rect 14369 12903 14427 12909
rect 14369 12900 14381 12903
rect 13504 12872 14381 12900
rect 13504 12860 13510 12872
rect 14369 12869 14381 12872
rect 14415 12869 14427 12903
rect 14369 12863 14427 12869
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5994 12832 6000 12844
rect 5859 12804 6000 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 5994 12792 6000 12804
rect 6052 12832 6058 12844
rect 7208 12832 7236 12860
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6052 12804 7389 12832
rect 6052 12792 6058 12804
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 8938 12832 8944 12844
rect 8899 12804 8944 12832
rect 7377 12795 7435 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 10594 12832 10600 12844
rect 9876 12804 10364 12832
rect 10555 12804 10600 12832
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 4939 12736 5571 12764
rect 5736 12736 7205 12764
rect 4939 12733 4951 12736
rect 4893 12727 4951 12733
rect 2130 12656 2136 12708
rect 2188 12696 2194 12708
rect 5442 12696 5448 12708
rect 2188 12668 4200 12696
rect 2188 12656 2194 12668
rect 2406 12628 2412 12640
rect 2367 12600 2412 12628
rect 2406 12588 2412 12600
rect 2464 12588 2470 12640
rect 3970 12628 3976 12640
rect 3931 12600 3976 12628
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4172 12628 4200 12668
rect 5184 12668 5448 12696
rect 4890 12628 4896 12640
rect 4172 12600 4896 12628
rect 4890 12588 4896 12600
rect 4948 12588 4954 12640
rect 5184 12637 5212 12668
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 5543 12696 5571 12736
rect 7193 12733 7205 12736
rect 7239 12764 7251 12767
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7239 12736 7849 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7837 12733 7849 12736
rect 7883 12764 7895 12767
rect 9876 12764 9904 12804
rect 7883 12736 9904 12764
rect 7883 12733 7895 12736
rect 7837 12727 7895 12733
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10226 12764 10232 12776
rect 10008 12736 10232 12764
rect 10008 12724 10014 12736
rect 10226 12724 10232 12736
rect 10284 12724 10290 12776
rect 10336 12764 10364 12804
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 11330 12792 11336 12844
rect 11388 12832 11394 12844
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 11388 12804 11621 12832
rect 11388 12792 11394 12804
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 13630 12832 13636 12844
rect 13591 12804 13636 12832
rect 11609 12795 11667 12801
rect 13630 12792 13636 12804
rect 13688 12792 13694 12844
rect 14642 12792 14648 12844
rect 14700 12832 14706 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 14700 12804 15117 12832
rect 14700 12792 14706 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15580 12832 15608 12928
rect 17218 12860 17224 12912
rect 17276 12900 17282 12912
rect 17586 12900 17592 12912
rect 17276 12872 17592 12900
rect 17276 12860 17282 12872
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 15580 12804 16865 12832
rect 15105 12795 15163 12801
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 17034 12832 17040 12844
rect 16947 12804 17040 12832
rect 16853 12795 16911 12801
rect 17034 12792 17040 12804
rect 17092 12832 17098 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17092 12804 17877 12832
rect 17092 12792 17098 12804
rect 17865 12801 17877 12804
rect 17911 12832 17923 12835
rect 17911 12804 18828 12832
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 10502 12764 10508 12776
rect 10336 12736 10508 12764
rect 10502 12724 10508 12736
rect 10560 12724 10566 12776
rect 10870 12724 10876 12776
rect 10928 12764 10934 12776
rect 12250 12764 12256 12776
rect 10928 12736 12256 12764
rect 10928 12724 10934 12736
rect 12250 12724 12256 12736
rect 12308 12724 12314 12776
rect 14826 12724 14832 12776
rect 14884 12764 14890 12776
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14884 12736 14933 12764
rect 14884 12724 14890 12736
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 16758 12764 16764 12776
rect 16719 12736 16764 12764
rect 14921 12727 14979 12733
rect 16758 12724 16764 12736
rect 16816 12764 16822 12776
rect 17405 12767 17463 12773
rect 17405 12764 17417 12767
rect 16816 12736 17417 12764
rect 16816 12724 16822 12736
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 18046 12724 18052 12776
rect 18104 12764 18110 12776
rect 18693 12767 18751 12773
rect 18693 12764 18705 12767
rect 18104 12736 18705 12764
rect 18104 12724 18110 12736
rect 18693 12733 18705 12736
rect 18739 12733 18751 12767
rect 18693 12727 18751 12733
rect 5629 12699 5687 12705
rect 5629 12696 5641 12699
rect 5543 12668 5641 12696
rect 5629 12665 5641 12668
rect 5675 12665 5687 12699
rect 5629 12659 5687 12665
rect 5169 12631 5227 12637
rect 5169 12597 5181 12631
rect 5215 12597 5227 12631
rect 5169 12591 5227 12597
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 5537 12631 5595 12637
rect 5537 12628 5549 12631
rect 5408 12600 5549 12628
rect 5408 12588 5414 12600
rect 5537 12597 5549 12600
rect 5583 12597 5595 12631
rect 5644 12628 5672 12659
rect 5810 12656 5816 12708
rect 5868 12696 5874 12708
rect 8113 12699 8171 12705
rect 8113 12696 8125 12699
rect 5868 12668 8125 12696
rect 5868 12656 5874 12668
rect 8113 12665 8125 12668
rect 8159 12665 8171 12699
rect 8113 12659 8171 12665
rect 8297 12699 8355 12705
rect 8297 12665 8309 12699
rect 8343 12696 8355 12699
rect 8757 12699 8815 12705
rect 8757 12696 8769 12699
rect 8343 12668 8769 12696
rect 8343 12665 8355 12668
rect 8297 12659 8355 12665
rect 8757 12665 8769 12668
rect 8803 12696 8815 12699
rect 9490 12696 9496 12708
rect 8803 12668 9496 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 9490 12656 9496 12668
rect 9548 12656 9554 12708
rect 10413 12699 10471 12705
rect 10413 12696 10425 12699
rect 9784 12668 10425 12696
rect 5994 12628 6000 12640
rect 5644 12600 6000 12628
rect 5537 12591 5595 12597
rect 5994 12588 6000 12600
rect 6052 12588 6058 12640
rect 6546 12628 6552 12640
rect 6507 12600 6552 12628
rect 6546 12588 6552 12600
rect 6604 12588 6610 12640
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 7282 12628 7288 12640
rect 7243 12600 7288 12628
rect 7282 12588 7288 12600
rect 7340 12588 7346 12640
rect 8846 12588 8852 12640
rect 8904 12628 8910 12640
rect 8904 12600 8949 12628
rect 8904 12588 8910 12600
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9784 12637 9812 12668
rect 10413 12665 10425 12668
rect 10459 12696 10471 12699
rect 10686 12696 10692 12708
rect 10459 12668 10692 12696
rect 10459 12665 10471 12668
rect 10413 12659 10471 12665
rect 10686 12656 10692 12668
rect 10744 12656 10750 12708
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 11698 12696 11704 12708
rect 11020 12668 11704 12696
rect 11020 12656 11026 12668
rect 11698 12656 11704 12668
rect 11756 12656 11762 12708
rect 12161 12699 12219 12705
rect 12161 12665 12173 12699
rect 12207 12696 12219 12699
rect 12207 12668 13492 12696
rect 12207 12665 12219 12668
rect 12161 12659 12219 12665
rect 9769 12631 9827 12637
rect 9769 12628 9781 12631
rect 9272 12600 9781 12628
rect 9272 12588 9278 12600
rect 9769 12597 9781 12600
rect 9815 12597 9827 12631
rect 9769 12591 9827 12597
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9916 12600 10333 12628
rect 9916 12588 9922 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 10870 12588 10876 12640
rect 10928 12628 10934 12640
rect 11146 12628 11152 12640
rect 10928 12600 11152 12628
rect 10928 12588 10934 12600
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 11330 12588 11336 12640
rect 11388 12628 11394 12640
rect 11514 12628 11520 12640
rect 11388 12600 11520 12628
rect 11388 12588 11394 12600
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 12176 12628 12204 12659
rect 13464 12640 13492 12668
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 14240 12668 15056 12696
rect 14240 12656 14246 12668
rect 15028 12640 15056 12668
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 18598 12696 18604 12708
rect 16724 12668 18604 12696
rect 16724 12656 16730 12668
rect 18598 12656 18604 12668
rect 18656 12656 18662 12708
rect 18800 12696 18828 12804
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 20990 12832 20996 12844
rect 20128 12804 20996 12832
rect 20128 12792 20134 12804
rect 20990 12792 20996 12804
rect 21048 12792 21054 12844
rect 21637 12835 21695 12841
rect 21637 12801 21649 12835
rect 21683 12832 21695 12835
rect 22373 12835 22431 12841
rect 22373 12832 22385 12835
rect 21683 12804 22385 12832
rect 21683 12801 21695 12804
rect 21637 12795 21695 12801
rect 22373 12801 22385 12804
rect 22419 12832 22431 12835
rect 22848 12832 22876 12931
rect 23106 12928 23112 12940
rect 23164 12928 23170 12980
rect 23474 12968 23480 12980
rect 23435 12940 23480 12968
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 23661 12971 23719 12977
rect 23661 12937 23673 12971
rect 23707 12968 23719 12971
rect 23934 12968 23940 12980
rect 23707 12940 23940 12968
rect 23707 12937 23719 12940
rect 23661 12931 23719 12937
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 24210 12928 24216 12980
rect 24268 12968 24274 12980
rect 24673 12971 24731 12977
rect 24673 12968 24685 12971
rect 24268 12940 24685 12968
rect 24268 12928 24274 12940
rect 24673 12937 24685 12940
rect 24719 12937 24731 12971
rect 25406 12968 25412 12980
rect 25367 12940 25412 12968
rect 24673 12931 24731 12937
rect 25406 12928 25412 12940
rect 25464 12928 25470 12980
rect 26237 12971 26295 12977
rect 26237 12937 26249 12971
rect 26283 12968 26295 12971
rect 26326 12968 26332 12980
rect 26283 12940 26332 12968
rect 26283 12937 26295 12940
rect 26237 12931 26295 12937
rect 26326 12928 26332 12940
rect 26384 12928 26390 12980
rect 22419 12804 22876 12832
rect 23492 12832 23520 12928
rect 23750 12860 23756 12912
rect 23808 12900 23814 12912
rect 24302 12900 24308 12912
rect 23808 12872 24308 12900
rect 23808 12860 23814 12872
rect 24302 12860 24308 12872
rect 24360 12860 24366 12912
rect 24213 12835 24271 12841
rect 24213 12832 24225 12835
rect 23492 12804 24225 12832
rect 22419 12801 22431 12804
rect 22373 12795 22431 12801
rect 24213 12801 24225 12804
rect 24259 12801 24271 12835
rect 24213 12795 24271 12801
rect 19426 12724 19432 12776
rect 19484 12764 19490 12776
rect 20806 12764 20812 12776
rect 19484 12736 20812 12764
rect 19484 12724 19490 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 22738 12724 22744 12776
rect 22796 12764 22802 12776
rect 23106 12764 23112 12776
rect 22796 12736 23112 12764
rect 22796 12724 22802 12736
rect 23106 12724 23112 12736
rect 23164 12724 23170 12776
rect 23474 12724 23480 12776
rect 23532 12764 23538 12776
rect 24762 12764 24768 12776
rect 23532 12736 24768 12764
rect 23532 12724 23538 12736
rect 24762 12724 24768 12736
rect 24820 12764 24826 12776
rect 25041 12767 25099 12773
rect 25041 12764 25053 12767
rect 24820 12736 25053 12764
rect 24820 12724 24826 12736
rect 25041 12733 25053 12736
rect 25087 12733 25099 12767
rect 25222 12764 25228 12776
rect 25135 12736 25228 12764
rect 25041 12727 25099 12733
rect 25222 12724 25228 12736
rect 25280 12764 25286 12776
rect 25406 12764 25412 12776
rect 25280 12736 25412 12764
rect 25280 12724 25286 12736
rect 25406 12724 25412 12736
rect 25464 12764 25470 12776
rect 25777 12767 25835 12773
rect 25777 12764 25789 12767
rect 25464 12736 25789 12764
rect 25464 12724 25470 12736
rect 25777 12733 25789 12736
rect 25823 12733 25835 12767
rect 25777 12727 25835 12733
rect 18960 12699 19018 12705
rect 18960 12696 18972 12699
rect 18800 12668 18972 12696
rect 18960 12665 18972 12668
rect 19006 12696 19018 12699
rect 19334 12696 19340 12708
rect 19006 12668 19340 12696
rect 19006 12665 19018 12668
rect 18960 12659 19018 12665
rect 19334 12656 19340 12668
rect 19392 12656 19398 12708
rect 22189 12699 22247 12705
rect 22189 12665 22201 12699
rect 22235 12696 22247 12699
rect 22646 12696 22652 12708
rect 22235 12668 22652 12696
rect 22235 12665 22247 12668
rect 22189 12659 22247 12665
rect 22646 12656 22652 12668
rect 22704 12656 22710 12708
rect 24029 12699 24087 12705
rect 24029 12665 24041 12699
rect 24075 12696 24087 12699
rect 24302 12696 24308 12708
rect 24075 12668 24308 12696
rect 24075 12665 24087 12668
rect 24029 12659 24087 12665
rect 24302 12656 24308 12668
rect 24360 12656 24366 12708
rect 25590 12696 25596 12708
rect 24688 12668 25596 12696
rect 11664 12600 12204 12628
rect 11664 12588 11670 12600
rect 13170 12588 13176 12640
rect 13228 12628 13234 12640
rect 13357 12631 13415 12637
rect 13357 12628 13369 12631
rect 13228 12600 13369 12628
rect 13228 12588 13234 12600
rect 13357 12597 13369 12600
rect 13403 12597 13415 12631
rect 13357 12591 13415 12597
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 13504 12600 13549 12628
rect 13504 12588 13510 12600
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14553 12631 14611 12637
rect 14553 12628 14565 12631
rect 14424 12600 14565 12628
rect 14424 12588 14430 12600
rect 14553 12597 14565 12600
rect 14599 12597 14611 12631
rect 15010 12628 15016 12640
rect 14971 12600 15016 12628
rect 14553 12591 14611 12597
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 16390 12628 16396 12640
rect 16351 12600 16396 12628
rect 16390 12588 16396 12600
rect 16448 12588 16454 12640
rect 18046 12588 18052 12640
rect 18104 12628 18110 12640
rect 18325 12631 18383 12637
rect 18325 12628 18337 12631
rect 18104 12600 18337 12628
rect 18104 12588 18110 12600
rect 18325 12597 18337 12600
rect 18371 12597 18383 12631
rect 18325 12591 18383 12597
rect 18414 12588 18420 12640
rect 18472 12628 18478 12640
rect 20073 12631 20131 12637
rect 20073 12628 20085 12631
rect 18472 12600 20085 12628
rect 18472 12588 18478 12600
rect 20073 12597 20085 12600
rect 20119 12628 20131 12631
rect 20806 12628 20812 12640
rect 20119 12600 20812 12628
rect 20119 12597 20131 12600
rect 20073 12591 20131 12597
rect 20806 12588 20812 12600
rect 20864 12588 20870 12640
rect 22002 12588 22008 12640
rect 22060 12628 22066 12640
rect 22097 12631 22155 12637
rect 22097 12628 22109 12631
rect 22060 12600 22109 12628
rect 22060 12588 22066 12600
rect 22097 12597 22109 12600
rect 22143 12597 22155 12631
rect 22097 12591 22155 12597
rect 23934 12588 23940 12640
rect 23992 12628 23998 12640
rect 24121 12631 24179 12637
rect 24121 12628 24133 12631
rect 23992 12600 24133 12628
rect 23992 12588 23998 12600
rect 24121 12597 24133 12600
rect 24167 12628 24179 12631
rect 24688 12628 24716 12668
rect 25590 12656 25596 12668
rect 25648 12656 25654 12708
rect 24167 12600 24716 12628
rect 24167 12597 24179 12600
rect 24121 12591 24179 12597
rect 1104 12538 26864 12560
rect 1104 12486 10315 12538
rect 10367 12486 10379 12538
rect 10431 12486 10443 12538
rect 10495 12486 10507 12538
rect 10559 12486 19648 12538
rect 19700 12486 19712 12538
rect 19764 12486 19776 12538
rect 19828 12486 19840 12538
rect 19892 12486 26864 12538
rect 1104 12464 26864 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1670 12424 1676 12436
rect 1627 12396 1676 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1670 12384 1676 12396
rect 1728 12384 1734 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 2869 12427 2927 12433
rect 2869 12424 2881 12427
rect 2832 12396 2881 12424
rect 2832 12384 2838 12396
rect 2869 12393 2881 12396
rect 2915 12393 2927 12427
rect 2869 12387 2927 12393
rect 4154 12384 4160 12436
rect 4212 12424 4218 12436
rect 4249 12427 4307 12433
rect 4249 12424 4261 12427
rect 4212 12396 4261 12424
rect 4212 12384 4218 12396
rect 4249 12393 4261 12396
rect 4295 12393 4307 12427
rect 4249 12387 4307 12393
rect 4890 12384 4896 12436
rect 4948 12424 4954 12436
rect 6825 12427 6883 12433
rect 6825 12424 6837 12427
rect 4948 12396 6837 12424
rect 4948 12384 4954 12396
rect 6825 12393 6837 12396
rect 6871 12424 6883 12427
rect 7006 12424 7012 12436
rect 6871 12396 7012 12424
rect 6871 12393 6883 12396
rect 6825 12387 6883 12393
rect 7006 12384 7012 12396
rect 7064 12424 7070 12436
rect 7282 12424 7288 12436
rect 7064 12396 7288 12424
rect 7064 12384 7070 12396
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 8110 12384 8116 12436
rect 8168 12384 8174 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8757 12427 8815 12433
rect 8757 12424 8769 12427
rect 8628 12396 8769 12424
rect 8628 12384 8634 12396
rect 8757 12393 8769 12396
rect 8803 12393 8815 12427
rect 8757 12387 8815 12393
rect 9493 12427 9551 12433
rect 9493 12393 9505 12427
rect 9539 12424 9551 12427
rect 9766 12424 9772 12436
rect 9539 12396 9772 12424
rect 9539 12393 9551 12396
rect 9493 12387 9551 12393
rect 14 12316 20 12368
rect 72 12356 78 12368
rect 2041 12359 2099 12365
rect 2041 12356 2053 12359
rect 72 12328 2053 12356
rect 72 12316 78 12328
rect 2041 12325 2053 12328
rect 2087 12356 2099 12359
rect 2406 12356 2412 12368
rect 2087 12328 2412 12356
rect 2087 12325 2099 12328
rect 2041 12319 2099 12325
rect 2406 12316 2412 12328
rect 2464 12316 2470 12368
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2556 12328 4108 12356
rect 2556 12316 2562 12328
rect 1394 12288 1400 12300
rect 1355 12260 1400 12288
rect 1394 12248 1400 12260
rect 1452 12248 1458 12300
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 3142 12288 3148 12300
rect 2823 12260 3148 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 3142 12248 3148 12260
rect 3200 12248 3206 12300
rect 4080 12297 4108 12328
rect 4706 12316 4712 12368
rect 4764 12356 4770 12368
rect 5353 12359 5411 12365
rect 5353 12356 5365 12359
rect 4764 12328 5365 12356
rect 4764 12316 4770 12328
rect 5353 12325 5365 12328
rect 5399 12325 5411 12359
rect 5353 12319 5411 12325
rect 5442 12316 5448 12368
rect 5500 12356 5506 12368
rect 5500 12328 5764 12356
rect 5500 12316 5506 12328
rect 4065 12291 4123 12297
rect 4065 12257 4077 12291
rect 4111 12288 4123 12291
rect 4617 12291 4675 12297
rect 4617 12288 4629 12291
rect 4111 12260 4629 12288
rect 4111 12257 4123 12260
rect 4065 12251 4123 12257
rect 4617 12257 4629 12260
rect 4663 12257 4675 12291
rect 5626 12288 5632 12300
rect 4617 12251 4675 12257
rect 5184 12260 5632 12288
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2464 12192 3065 12220
rect 2464 12180 2470 12192
rect 3053 12189 3065 12192
rect 3099 12220 3111 12223
rect 3510 12220 3516 12232
rect 3099 12192 3516 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3510 12180 3516 12192
rect 3568 12220 3574 12232
rect 5184 12220 5212 12260
rect 5626 12248 5632 12260
rect 5684 12248 5690 12300
rect 3568 12192 5212 12220
rect 5353 12223 5411 12229
rect 3568 12180 3574 12192
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 5534 12220 5540 12232
rect 5399 12192 5540 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 5534 12180 5540 12192
rect 5592 12180 5598 12232
rect 5736 12220 5764 12328
rect 6638 12316 6644 12368
rect 6696 12356 6702 12368
rect 7650 12356 7656 12368
rect 6696 12328 7227 12356
rect 6696 12316 6702 12328
rect 5905 12291 5963 12297
rect 5905 12257 5917 12291
rect 5951 12288 5963 12291
rect 6822 12288 6828 12300
rect 5951 12260 6828 12288
rect 5951 12257 5963 12260
rect 5905 12251 5963 12257
rect 6822 12248 6828 12260
rect 6880 12248 6886 12300
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5736 12192 6009 12220
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6270 12220 6276 12232
rect 6227 12192 6276 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 2372 12124 3801 12152
rect 2372 12112 2378 12124
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 5810 12152 5816 12164
rect 4212 12124 5816 12152
rect 4212 12112 4218 12124
rect 5810 12112 5816 12124
rect 5868 12112 5874 12164
rect 6012 12152 6040 12183
rect 6270 12180 6276 12192
rect 6328 12220 6334 12232
rect 6638 12220 6644 12232
rect 6328 12192 6644 12220
rect 6328 12180 6334 12192
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7098 12180 7104 12232
rect 7156 12180 7162 12232
rect 7199 12220 7227 12328
rect 7300 12328 7656 12356
rect 7300 12300 7328 12328
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 8128 12356 8156 12384
rect 8294 12356 8300 12368
rect 8128 12328 8300 12356
rect 8294 12316 8300 12328
rect 8352 12316 8358 12368
rect 7282 12248 7288 12300
rect 7340 12248 7346 12300
rect 7466 12288 7472 12300
rect 7427 12260 7472 12288
rect 7466 12248 7472 12260
rect 7524 12248 7530 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 7742 12288 7748 12300
rect 7607 12260 7748 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 7650 12220 7656 12232
rect 7199 12192 7656 12220
rect 7650 12180 7656 12192
rect 7708 12220 7714 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7708 12192 8401 12220
rect 7708 12180 7714 12192
rect 8389 12189 8401 12192
rect 8435 12220 8447 12223
rect 8938 12220 8944 12232
rect 8435 12192 8944 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 6730 12152 6736 12164
rect 6012 12124 6736 12152
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 7116 12152 7144 12180
rect 9508 12152 9536 12387
rect 9766 12384 9772 12396
rect 9824 12384 9830 12436
rect 9858 12384 9864 12436
rect 9916 12424 9922 12436
rect 9953 12427 10011 12433
rect 9953 12424 9965 12427
rect 9916 12396 9965 12424
rect 9916 12384 9922 12396
rect 9953 12393 9965 12396
rect 9999 12393 10011 12427
rect 14642 12424 14648 12436
rect 14603 12396 14648 12424
rect 9953 12387 10011 12393
rect 14642 12384 14648 12396
rect 14700 12384 14706 12436
rect 14826 12384 14832 12436
rect 14884 12424 14890 12436
rect 15746 12424 15752 12436
rect 14884 12396 15752 12424
rect 14884 12384 14890 12396
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 16025 12427 16083 12433
rect 16025 12393 16037 12427
rect 16071 12424 16083 12427
rect 16482 12424 16488 12436
rect 16071 12396 16488 12424
rect 16071 12393 16083 12396
rect 16025 12387 16083 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16666 12424 16672 12436
rect 16579 12396 16672 12424
rect 16666 12384 16672 12396
rect 16724 12424 16730 12436
rect 17678 12424 17684 12436
rect 16724 12396 17684 12424
rect 16724 12384 16730 12396
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 18414 12424 18420 12436
rect 18375 12396 18420 12424
rect 18414 12384 18420 12396
rect 18472 12384 18478 12436
rect 20346 12424 20352 12436
rect 20307 12396 20352 12424
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 20772 12396 21557 12424
rect 20772 12384 20778 12396
rect 21545 12393 21557 12396
rect 21591 12424 21603 12427
rect 22002 12424 22008 12436
rect 21591 12396 22008 12424
rect 21591 12393 21603 12396
rect 21545 12387 21603 12393
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 22646 12424 22652 12436
rect 22607 12396 22652 12424
rect 22646 12384 22652 12396
rect 22704 12384 22710 12436
rect 23014 12424 23020 12436
rect 22975 12396 23020 12424
rect 23014 12384 23020 12396
rect 23072 12384 23078 12436
rect 23109 12427 23167 12433
rect 23109 12393 23121 12427
rect 23155 12424 23167 12427
rect 23382 12424 23388 12436
rect 23155 12396 23388 12424
rect 23155 12393 23167 12396
rect 23109 12387 23167 12393
rect 23382 12384 23388 12396
rect 23440 12384 23446 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24489 12427 24547 12433
rect 24489 12424 24501 12427
rect 24268 12396 24501 12424
rect 24268 12384 24274 12396
rect 24489 12393 24501 12396
rect 24535 12393 24547 12427
rect 24489 12387 24547 12393
rect 24673 12427 24731 12433
rect 24673 12393 24685 12427
rect 24719 12393 24731 12427
rect 24673 12387 24731 12393
rect 11882 12356 11888 12368
rect 9876 12328 11888 12356
rect 9876 12300 9904 12328
rect 11882 12316 11888 12328
rect 11940 12316 11946 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 14185 12359 14243 12365
rect 14185 12356 14197 12359
rect 13780 12328 14197 12356
rect 13780 12316 13786 12328
rect 14185 12325 14197 12328
rect 14231 12325 14243 12359
rect 14185 12319 14243 12325
rect 16390 12316 16396 12368
rect 16448 12356 16454 12368
rect 17589 12359 17647 12365
rect 17589 12356 17601 12359
rect 16448 12328 17601 12356
rect 16448 12316 16454 12328
rect 17589 12325 17601 12328
rect 17635 12325 17647 12359
rect 17589 12319 17647 12325
rect 19981 12359 20039 12365
rect 19981 12325 19993 12359
rect 20027 12356 20039 12359
rect 20622 12356 20628 12368
rect 20027 12328 20628 12356
rect 20027 12325 20039 12328
rect 19981 12319 20039 12325
rect 20622 12316 20628 12328
rect 20680 12316 20686 12368
rect 21453 12359 21511 12365
rect 21453 12325 21465 12359
rect 21499 12356 21511 12359
rect 22094 12356 22100 12368
rect 21499 12328 22100 12356
rect 21499 12325 21511 12328
rect 21453 12319 21511 12325
rect 22094 12316 22100 12328
rect 22152 12356 22158 12368
rect 22152 12328 22232 12356
rect 22152 12316 22158 12328
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 9766 12288 9772 12300
rect 9640 12260 9772 12288
rect 9640 12248 9646 12260
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 9858 12248 9864 12300
rect 9916 12248 9922 12300
rect 10680 12291 10738 12297
rect 10680 12257 10692 12291
rect 10726 12288 10738 12291
rect 11054 12288 11060 12300
rect 10726 12260 11060 12288
rect 10726 12257 10738 12260
rect 10680 12251 10738 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 13538 12288 13544 12300
rect 13499 12260 13544 12288
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 16577 12291 16635 12297
rect 16577 12257 16589 12291
rect 16623 12257 16635 12291
rect 17218 12288 17224 12300
rect 17179 12260 17224 12288
rect 16577 12251 16635 12257
rect 10410 12220 10416 12232
rect 10371 12192 10416 12220
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12216 12192 13093 12220
rect 12216 12180 12222 12192
rect 13081 12189 13093 12192
rect 13127 12220 13139 12223
rect 13170 12220 13176 12232
rect 13127 12192 13176 12220
rect 13127 12189 13139 12192
rect 13081 12183 13139 12189
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13630 12220 13636 12232
rect 13591 12192 13636 12220
rect 13630 12180 13636 12192
rect 13688 12180 13694 12232
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12189 13783 12223
rect 13725 12183 13783 12189
rect 7116 12124 9536 12152
rect 12713 12155 12771 12161
rect 12713 12121 12725 12155
rect 12759 12152 12771 12155
rect 13740 12152 13768 12183
rect 14090 12152 14096 12164
rect 12759 12124 14096 12152
rect 12759 12121 12771 12124
rect 12713 12115 12771 12121
rect 14090 12112 14096 12124
rect 14148 12112 14154 12164
rect 16592 12152 16620 12251
rect 17218 12248 17224 12260
rect 17276 12248 17282 12300
rect 18966 12248 18972 12300
rect 19024 12288 19030 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19024 12260 19257 12288
rect 19024 12248 19030 12260
rect 19245 12257 19257 12260
rect 19291 12288 19303 12291
rect 20070 12288 20076 12300
rect 19291 12260 20076 12288
rect 19291 12257 19303 12260
rect 19245 12251 19303 12257
rect 20070 12248 20076 12260
rect 20128 12248 20134 12300
rect 21726 12248 21732 12300
rect 21784 12288 21790 12300
rect 21913 12291 21971 12297
rect 21913 12288 21925 12291
rect 21784 12260 21925 12288
rect 21784 12248 21790 12260
rect 21913 12257 21925 12260
rect 21959 12257 21971 12291
rect 21913 12251 21971 12257
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 17402 12220 17408 12232
rect 16899 12192 17408 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17862 12220 17868 12232
rect 17823 12192 17868 12220
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 19337 12223 19395 12229
rect 19337 12220 19349 12223
rect 18984 12192 19349 12220
rect 18984 12164 19012 12192
rect 19337 12189 19349 12192
rect 19383 12189 19395 12223
rect 19337 12183 19395 12189
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 20717 12223 20775 12229
rect 19484 12192 19529 12220
rect 19484 12180 19490 12192
rect 20717 12189 20729 12223
rect 20763 12220 20775 12223
rect 21634 12220 21640 12232
rect 20763 12192 21640 12220
rect 20763 12189 20775 12192
rect 20717 12183 20775 12189
rect 21634 12180 21640 12192
rect 21692 12220 21698 12232
rect 22204 12229 22232 12328
rect 22462 12316 22468 12368
rect 22520 12356 22526 12368
rect 23032 12356 23060 12384
rect 22520 12328 23612 12356
rect 22520 12316 22526 12328
rect 23106 12248 23112 12300
rect 23164 12288 23170 12300
rect 23474 12288 23480 12300
rect 23164 12260 23480 12288
rect 23164 12248 23170 12260
rect 23474 12248 23480 12260
rect 23532 12248 23538 12300
rect 23584 12288 23612 12328
rect 23842 12316 23848 12368
rect 23900 12356 23906 12368
rect 24688 12356 24716 12387
rect 26053 12359 26111 12365
rect 26053 12356 26065 12359
rect 23900 12328 24716 12356
rect 24872 12328 26065 12356
rect 23900 12316 23906 12328
rect 23584 12260 23704 12288
rect 23676 12229 23704 12260
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 24872 12288 24900 12328
rect 26053 12325 26065 12328
rect 26099 12325 26111 12359
rect 26053 12319 26111 12325
rect 24360 12260 24900 12288
rect 24360 12248 24366 12260
rect 24946 12248 24952 12300
rect 25004 12288 25010 12300
rect 25041 12291 25099 12297
rect 25041 12288 25053 12291
rect 25004 12260 25053 12288
rect 25004 12248 25010 12260
rect 25041 12257 25053 12260
rect 25087 12257 25099 12291
rect 25041 12251 25099 12257
rect 25133 12291 25191 12297
rect 25133 12257 25145 12291
rect 25179 12288 25191 12291
rect 25590 12288 25596 12300
rect 25179 12260 25596 12288
rect 25179 12257 25191 12260
rect 25133 12251 25191 12257
rect 25590 12248 25596 12260
rect 25648 12248 25654 12300
rect 22005 12223 22063 12229
rect 22005 12220 22017 12223
rect 21692 12192 22017 12220
rect 21692 12180 21698 12192
rect 22005 12189 22017 12192
rect 22051 12189 22063 12223
rect 22005 12183 22063 12189
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12189 22247 12223
rect 23569 12223 23627 12229
rect 23569 12220 23581 12223
rect 22189 12183 22247 12189
rect 23032 12192 23581 12220
rect 23032 12164 23060 12192
rect 23569 12189 23581 12192
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 23661 12223 23719 12229
rect 23661 12189 23673 12223
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 24213 12223 24271 12229
rect 24213 12189 24225 12223
rect 24259 12220 24271 12223
rect 24259 12192 24900 12220
rect 24259 12189 24271 12192
rect 24213 12183 24271 12189
rect 17494 12152 17500 12164
rect 16592 12124 17500 12152
rect 17494 12112 17500 12124
rect 17552 12112 17558 12164
rect 18966 12112 18972 12164
rect 19024 12112 19030 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 23014 12152 23020 12164
rect 19760 12124 23020 12152
rect 19760 12112 19766 12124
rect 23014 12112 23020 12124
rect 23072 12112 23078 12164
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 23842 12152 23848 12164
rect 23348 12124 23848 12152
rect 23348 12112 23354 12124
rect 23842 12112 23848 12124
rect 23900 12112 23906 12164
rect 24578 12112 24584 12164
rect 24636 12152 24642 12164
rect 24762 12152 24768 12164
rect 24636 12124 24768 12152
rect 24636 12112 24642 12124
rect 24762 12112 24768 12124
rect 24820 12112 24826 12164
rect 24872 12152 24900 12192
rect 25222 12180 25228 12232
rect 25280 12220 25286 12232
rect 25280 12192 25325 12220
rect 25280 12180 25286 12192
rect 25240 12152 25268 12180
rect 24872 12124 25268 12152
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2682 12084 2688 12096
rect 2455 12056 2688 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2682 12044 2688 12056
rect 2740 12044 2746 12096
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 5261 12087 5319 12093
rect 5261 12084 5273 12087
rect 3200 12056 5273 12084
rect 3200 12044 3206 12056
rect 5261 12053 5273 12056
rect 5307 12084 5319 12087
rect 5350 12084 5356 12096
rect 5307 12056 5356 12084
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 6638 12084 6644 12096
rect 5583 12056 6644 12084
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 6638 12044 6644 12056
rect 6696 12044 6702 12096
rect 7098 12084 7104 12096
rect 7059 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 11793 12087 11851 12093
rect 11793 12053 11805 12087
rect 11839 12084 11851 12087
rect 12434 12084 12440 12096
rect 11839 12056 12440 12084
rect 11839 12053 11851 12056
rect 11793 12047 11851 12053
rect 12434 12044 12440 12056
rect 12492 12044 12498 12096
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 14274 12044 14280 12096
rect 14332 12084 14338 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14332 12056 14933 12084
rect 14332 12044 14338 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15565 12087 15623 12093
rect 15565 12053 15577 12087
rect 15611 12084 15623 12087
rect 15654 12084 15660 12096
rect 15611 12056 15660 12084
rect 15611 12053 15623 12056
rect 15565 12047 15623 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16206 12084 16212 12096
rect 16167 12056 16212 12084
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 17218 12084 17224 12096
rect 16632 12056 17224 12084
rect 16632 12044 16638 12056
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18693 12087 18751 12093
rect 18693 12084 18705 12087
rect 18104 12056 18705 12084
rect 18104 12044 18110 12056
rect 18693 12053 18705 12056
rect 18739 12053 18751 12087
rect 18874 12084 18880 12096
rect 18835 12056 18880 12084
rect 18693 12047 18751 12053
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 22738 12084 22744 12096
rect 20128 12056 22744 12084
rect 20128 12044 20134 12056
rect 22738 12044 22744 12056
rect 22796 12044 22802 12096
rect 24854 12044 24860 12096
rect 24912 12084 24918 12096
rect 25685 12087 25743 12093
rect 25685 12084 25697 12087
rect 24912 12056 25697 12084
rect 24912 12044 24918 12056
rect 25685 12053 25697 12056
rect 25731 12053 25743 12087
rect 25685 12047 25743 12053
rect 1104 11994 26864 12016
rect 1104 11942 5648 11994
rect 5700 11942 5712 11994
rect 5764 11942 5776 11994
rect 5828 11942 5840 11994
rect 5892 11942 14982 11994
rect 15034 11942 15046 11994
rect 15098 11942 15110 11994
rect 15162 11942 15174 11994
rect 15226 11942 24315 11994
rect 24367 11942 24379 11994
rect 24431 11942 24443 11994
rect 24495 11942 24507 11994
rect 24559 11942 26864 11994
rect 1104 11920 26864 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 1452 11852 1593 11880
rect 1452 11840 1458 11852
rect 1581 11849 1593 11852
rect 1627 11880 1639 11883
rect 2869 11883 2927 11889
rect 1627 11852 2268 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2240 11753 2268 11852
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 3142 11880 3148 11892
rect 2915 11852 3148 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 3142 11840 3148 11852
rect 3200 11840 3206 11892
rect 5629 11883 5687 11889
rect 5629 11849 5641 11883
rect 5675 11880 5687 11883
rect 6270 11880 6276 11892
rect 5675 11852 6276 11880
rect 5675 11849 5687 11852
rect 5629 11843 5687 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 8754 11880 8760 11892
rect 8715 11852 8760 11880
rect 8754 11840 8760 11852
rect 8812 11840 8818 11892
rect 9401 11883 9459 11889
rect 9401 11849 9413 11883
rect 9447 11880 9459 11883
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 9447 11852 9689 11880
rect 9447 11849 9459 11852
rect 9401 11843 9459 11849
rect 9677 11849 9689 11852
rect 9723 11880 9735 11883
rect 10410 11880 10416 11892
rect 9723 11852 10416 11880
rect 9723 11849 9735 11852
rect 9677 11843 9735 11849
rect 4614 11772 4620 11824
rect 4672 11812 4678 11824
rect 4890 11812 4896 11824
rect 4672 11784 4896 11812
rect 4672 11772 4678 11784
rect 4890 11772 4896 11784
rect 4948 11772 4954 11824
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11713 2283 11747
rect 2406 11744 2412 11756
rect 2367 11716 2412 11744
rect 2225 11707 2283 11713
rect 2406 11704 2412 11716
rect 2464 11704 2470 11756
rect 9784 11753 9812 11852
rect 10410 11840 10416 11852
rect 10468 11880 10474 11892
rect 10468 11852 12112 11880
rect 10468 11840 10474 11852
rect 12084 11824 12112 11852
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 13596 11852 14749 11880
rect 13596 11840 13602 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 16850 11880 16856 11892
rect 14737 11843 14795 11849
rect 15488 11852 16856 11880
rect 12066 11772 12072 11824
rect 12124 11812 12130 11824
rect 12124 11784 12480 11812
rect 12124 11772 12130 11784
rect 12452 11753 12480 11784
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 15488 11812 15516 11852
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 20070 11880 20076 11892
rect 20031 11852 20076 11880
rect 20070 11840 20076 11852
rect 20128 11840 20134 11892
rect 20809 11883 20867 11889
rect 20809 11849 20821 11883
rect 20855 11880 20867 11883
rect 21358 11880 21364 11892
rect 20855 11852 21364 11880
rect 20855 11849 20867 11852
rect 20809 11843 20867 11849
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 21634 11880 21640 11892
rect 21595 11852 21640 11880
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 22741 11883 22799 11889
rect 22741 11849 22753 11883
rect 22787 11880 22799 11883
rect 23474 11880 23480 11892
rect 22787 11852 23480 11880
rect 22787 11849 22799 11852
rect 22741 11843 22799 11849
rect 23474 11840 23480 11852
rect 23532 11840 23538 11892
rect 25314 11840 25320 11892
rect 25372 11880 25378 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 25372 11852 25421 11880
rect 25372 11840 25378 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 26234 11880 26240 11892
rect 26195 11852 26240 11880
rect 25409 11843 25467 11849
rect 26234 11840 26240 11852
rect 26292 11840 26298 11892
rect 19426 11812 19432 11824
rect 14240 11784 15516 11812
rect 19339 11784 19432 11812
rect 14240 11772 14246 11784
rect 19426 11772 19432 11784
rect 19484 11772 19490 11824
rect 19978 11772 19984 11824
rect 20036 11812 20042 11824
rect 23661 11815 23719 11821
rect 23661 11812 23673 11815
rect 20036 11784 23673 11812
rect 20036 11772 20042 11784
rect 23661 11781 23673 11784
rect 23707 11781 23719 11815
rect 23661 11775 23719 11781
rect 24578 11772 24584 11824
rect 24636 11812 24642 11824
rect 25777 11815 25835 11821
rect 25777 11812 25789 11815
rect 24636 11784 25789 11812
rect 24636 11772 24642 11784
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 17126 11704 17132 11756
rect 17184 11744 17190 11756
rect 17678 11744 17684 11756
rect 17184 11716 17684 11744
rect 17184 11704 17190 11716
rect 17678 11704 17684 11716
rect 17736 11744 17742 11756
rect 19444 11744 19472 11772
rect 22281 11747 22339 11753
rect 17736 11716 18184 11744
rect 19444 11716 20392 11744
rect 17736 11704 17742 11716
rect 2130 11676 2136 11688
rect 2091 11648 2136 11676
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11676 3295 11679
rect 3326 11676 3332 11688
rect 3283 11648 3332 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3326 11636 3332 11648
rect 3384 11676 3390 11688
rect 5626 11676 5632 11688
rect 3384 11648 5632 11676
rect 3384 11636 3390 11648
rect 5626 11636 5632 11648
rect 5684 11676 5690 11688
rect 6546 11676 6552 11688
rect 5684 11648 6552 11676
rect 5684 11636 5690 11648
rect 6546 11636 6552 11648
rect 6604 11676 6610 11688
rect 6641 11679 6699 11685
rect 6641 11676 6653 11679
rect 6604 11648 6653 11676
rect 6604 11636 6610 11648
rect 6641 11645 6653 11648
rect 6687 11676 6699 11679
rect 6825 11679 6883 11685
rect 6825 11676 6837 11679
rect 6687 11648 6837 11676
rect 6687 11645 6699 11648
rect 6641 11639 6699 11645
rect 6825 11645 6837 11648
rect 6871 11676 6883 11679
rect 15381 11679 15439 11685
rect 6871 11648 8616 11676
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 3596 11611 3654 11617
rect 3596 11577 3608 11611
rect 3642 11608 3654 11611
rect 3970 11608 3976 11620
rect 3642 11580 3976 11608
rect 3642 11577 3654 11580
rect 3596 11571 3654 11577
rect 3970 11568 3976 11580
rect 4028 11568 4034 11620
rect 7092 11611 7150 11617
rect 7092 11577 7104 11611
rect 7138 11608 7150 11611
rect 7190 11608 7196 11620
rect 7138 11580 7196 11608
rect 7138 11577 7150 11580
rect 7092 11571 7150 11577
rect 7190 11568 7196 11580
rect 7248 11568 7254 11620
rect 8588 11552 8616 11648
rect 15381 11645 15393 11679
rect 15427 11676 15439 11679
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 15427 11648 15485 11676
rect 15427 11645 15439 11648
rect 15381 11639 15439 11645
rect 15473 11645 15485 11648
rect 15519 11676 15531 11679
rect 15562 11676 15568 11688
rect 15519 11648 15568 11676
rect 15519 11645 15531 11648
rect 15473 11639 15531 11645
rect 15562 11636 15568 11648
rect 15620 11636 15626 11688
rect 16758 11636 16764 11688
rect 16816 11676 16822 11688
rect 17773 11679 17831 11685
rect 17773 11676 17785 11679
rect 16816 11648 17785 11676
rect 16816 11636 16822 11648
rect 17773 11645 17785 11648
rect 17819 11676 17831 11679
rect 18046 11676 18052 11688
rect 17819 11648 18052 11676
rect 17819 11645 17831 11648
rect 17773 11639 17831 11645
rect 18046 11636 18052 11648
rect 18104 11636 18110 11688
rect 18156 11676 18184 11716
rect 19702 11676 19708 11688
rect 18156 11648 19708 11676
rect 19702 11636 19708 11648
rect 19760 11636 19766 11688
rect 9582 11568 9588 11620
rect 9640 11608 9646 11620
rect 10014 11611 10072 11617
rect 10014 11608 10026 11611
rect 9640 11580 10026 11608
rect 9640 11568 9646 11580
rect 10014 11577 10026 11580
rect 10060 11577 10072 11611
rect 10014 11571 10072 11577
rect 12526 11568 12532 11620
rect 12584 11608 12590 11620
rect 12682 11611 12740 11617
rect 12682 11608 12694 11611
rect 12584 11580 12694 11608
rect 12584 11568 12590 11580
rect 12682 11577 12694 11580
rect 12728 11577 12740 11611
rect 12682 11571 12740 11577
rect 13630 11568 13636 11620
rect 13688 11608 13694 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 13688 11580 14381 11608
rect 13688 11568 13694 11580
rect 14369 11577 14381 11580
rect 14415 11577 14427 11611
rect 14369 11571 14427 11577
rect 15654 11568 15660 11620
rect 15712 11617 15718 11620
rect 20364 11617 20392 11716
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22462 11744 22468 11756
rect 22327 11716 22468 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22462 11704 22468 11716
rect 22520 11704 22526 11756
rect 23014 11744 23020 11756
rect 22975 11716 23020 11744
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23106 11704 23112 11756
rect 23164 11744 23170 11756
rect 24305 11747 24363 11753
rect 24305 11744 24317 11747
rect 23164 11716 24317 11744
rect 23164 11704 23170 11716
rect 24305 11713 24317 11716
rect 24351 11744 24363 11747
rect 25130 11744 25136 11756
rect 24351 11716 25136 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 20622 11676 20628 11688
rect 20583 11648 20628 11676
rect 20622 11636 20628 11648
rect 20680 11636 20686 11688
rect 20714 11636 20720 11688
rect 20772 11676 20778 11688
rect 21542 11676 21548 11688
rect 20772 11648 21548 11676
rect 20772 11636 20778 11648
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 24946 11636 24952 11688
rect 25004 11676 25010 11688
rect 25240 11685 25268 11784
rect 25777 11781 25789 11784
rect 25823 11781 25835 11815
rect 25777 11775 25835 11781
rect 25041 11679 25099 11685
rect 25041 11676 25053 11679
rect 25004 11648 25053 11676
rect 25004 11636 25010 11648
rect 25041 11645 25053 11648
rect 25087 11645 25099 11679
rect 25041 11639 25099 11645
rect 25225 11679 25283 11685
rect 25225 11645 25237 11679
rect 25271 11645 25283 11679
rect 25225 11639 25283 11645
rect 15712 11611 15776 11617
rect 15712 11577 15730 11611
rect 15764 11577 15776 11611
rect 18294 11611 18352 11617
rect 18294 11608 18306 11611
rect 15712 11571 15776 11577
rect 17420 11580 18306 11608
rect 15712 11568 15718 11571
rect 17420 11552 17448 11580
rect 18294 11577 18306 11580
rect 18340 11577 18352 11611
rect 18294 11571 18352 11577
rect 20349 11611 20407 11617
rect 20349 11577 20361 11611
rect 20395 11608 20407 11611
rect 20806 11608 20812 11620
rect 20395 11580 20812 11608
rect 20395 11577 20407 11580
rect 20349 11571 20407 11577
rect 20806 11568 20812 11580
rect 20864 11568 20870 11620
rect 21450 11608 21456 11620
rect 21411 11580 21456 11608
rect 21450 11568 21456 11580
rect 21508 11608 21514 11620
rect 22005 11611 22063 11617
rect 22005 11608 22017 11611
rect 21508 11580 22017 11608
rect 21508 11568 21514 11580
rect 22005 11577 22017 11580
rect 22051 11577 22063 11611
rect 22005 11571 22063 11577
rect 1762 11540 1768 11552
rect 1723 11512 1768 11540
rect 1762 11500 1768 11512
rect 1820 11500 1826 11552
rect 4614 11500 4620 11552
rect 4672 11540 4678 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4672 11512 4721 11540
rect 4672 11500 4678 11512
rect 4709 11509 4721 11512
rect 4755 11509 4767 11543
rect 4709 11503 4767 11509
rect 7650 11500 7656 11552
rect 7708 11540 7714 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 7708 11512 8217 11540
rect 7708 11500 7714 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 8205 11503 8263 11509
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8628 11512 9229 11540
rect 8628 11500 8634 11512
rect 9217 11509 9229 11512
rect 9263 11540 9275 11543
rect 9401 11543 9459 11549
rect 9401 11540 9413 11543
rect 9263 11512 9413 11540
rect 9263 11509 9275 11512
rect 9217 11503 9275 11509
rect 9401 11509 9413 11512
rect 9447 11509 9459 11543
rect 9401 11503 9459 11509
rect 10870 11500 10876 11552
rect 10928 11540 10934 11552
rect 11054 11540 11060 11552
rect 10928 11512 11060 11540
rect 10928 11500 10934 11512
rect 11054 11500 11060 11512
rect 11112 11540 11118 11552
rect 11149 11543 11207 11549
rect 11149 11540 11161 11543
rect 11112 11512 11161 11540
rect 11112 11500 11118 11512
rect 11149 11509 11161 11512
rect 11195 11540 11207 11543
rect 11701 11543 11759 11549
rect 11701 11540 11713 11543
rect 11195 11512 11713 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11701 11509 11713 11512
rect 11747 11509 11759 11543
rect 11701 11503 11759 11509
rect 12066 11500 12072 11552
rect 12124 11540 12130 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 12124 11512 12265 11540
rect 12124 11500 12130 11512
rect 12253 11509 12265 11512
rect 12299 11509 12311 11543
rect 13814 11540 13820 11552
rect 13775 11512 13820 11540
rect 12253 11503 12311 11509
rect 13814 11500 13820 11512
rect 13872 11500 13878 11552
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 19334 11500 19340 11552
rect 19392 11540 19398 11552
rect 20438 11540 20444 11552
rect 19392 11512 20444 11540
rect 19392 11500 19398 11512
rect 20438 11500 20444 11512
rect 20496 11540 20502 11552
rect 21085 11543 21143 11549
rect 21085 11540 21097 11543
rect 20496 11512 21097 11540
rect 20496 11500 20502 11512
rect 21085 11509 21097 11512
rect 21131 11540 21143 11543
rect 21726 11540 21732 11552
rect 21131 11512 21732 11540
rect 21131 11509 21143 11512
rect 21085 11503 21143 11509
rect 21726 11500 21732 11512
rect 21784 11500 21790 11552
rect 21910 11500 21916 11552
rect 21968 11540 21974 11552
rect 22097 11543 22155 11549
rect 22097 11540 22109 11543
rect 21968 11512 22109 11540
rect 21968 11500 21974 11512
rect 22097 11509 22109 11512
rect 22143 11509 22155 11543
rect 23474 11540 23480 11552
rect 23435 11512 23480 11540
rect 22097 11503 22155 11509
rect 23474 11500 23480 11512
rect 23532 11540 23538 11552
rect 24029 11543 24087 11549
rect 24029 11540 24041 11543
rect 23532 11512 24041 11540
rect 23532 11500 23538 11512
rect 24029 11509 24041 11512
rect 24075 11509 24087 11543
rect 24029 11503 24087 11509
rect 24121 11543 24179 11549
rect 24121 11509 24133 11543
rect 24167 11540 24179 11543
rect 24210 11540 24216 11552
rect 24167 11512 24216 11540
rect 24167 11509 24179 11512
rect 24121 11503 24179 11509
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 24765 11543 24823 11549
rect 24765 11509 24777 11543
rect 24811 11540 24823 11543
rect 25590 11540 25596 11552
rect 24811 11512 25596 11540
rect 24811 11509 24823 11512
rect 24765 11503 24823 11509
rect 25590 11500 25596 11512
rect 25648 11500 25654 11552
rect 1104 11450 26864 11472
rect 1104 11398 10315 11450
rect 10367 11398 10379 11450
rect 10431 11398 10443 11450
rect 10495 11398 10507 11450
rect 10559 11398 19648 11450
rect 19700 11398 19712 11450
rect 19764 11398 19776 11450
rect 19828 11398 19840 11450
rect 19892 11398 26864 11450
rect 1104 11376 26864 11398
rect 1949 11339 2007 11345
rect 1949 11305 1961 11339
rect 1995 11336 2007 11339
rect 2130 11336 2136 11348
rect 1995 11308 2136 11336
rect 1995 11305 2007 11308
rect 1949 11299 2007 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2317 11339 2375 11345
rect 2317 11305 2329 11339
rect 2363 11336 2375 11339
rect 2774 11336 2780 11348
rect 2363 11308 2780 11336
rect 2363 11305 2375 11308
rect 2317 11299 2375 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 3510 11336 3516 11348
rect 2924 11308 2969 11336
rect 3471 11308 3516 11336
rect 2924 11296 2930 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4341 11339 4399 11345
rect 4341 11305 4353 11339
rect 4387 11336 4399 11339
rect 4430 11336 4436 11348
rect 4387 11308 4436 11336
rect 4387 11305 4399 11308
rect 4341 11299 4399 11305
rect 4430 11296 4436 11308
rect 4488 11296 4494 11348
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 6604 11308 6929 11336
rect 6604 11296 6610 11308
rect 6917 11305 6929 11308
rect 6963 11336 6975 11339
rect 7282 11336 7288 11348
rect 6963 11308 7288 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7282 11296 7288 11308
rect 7340 11296 7346 11348
rect 7745 11339 7803 11345
rect 7745 11305 7757 11339
rect 7791 11336 7803 11339
rect 8202 11336 8208 11348
rect 7791 11308 8208 11336
rect 7791 11305 7803 11308
rect 7745 11299 7803 11305
rect 8202 11296 8208 11308
rect 8260 11336 8266 11348
rect 8297 11339 8355 11345
rect 8297 11336 8309 11339
rect 8260 11308 8309 11336
rect 8260 11296 8266 11308
rect 8297 11305 8309 11308
rect 8343 11305 8355 11339
rect 8297 11299 8355 11305
rect 9674 11296 9680 11348
rect 9732 11336 9738 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 9732 11308 10241 11336
rect 9732 11296 9738 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 11514 11336 11520 11348
rect 11475 11308 11520 11336
rect 10229 11299 10287 11305
rect 11514 11296 11520 11308
rect 11572 11296 11578 11348
rect 11882 11336 11888 11348
rect 11843 11308 11888 11336
rect 11882 11296 11888 11308
rect 11940 11296 11946 11348
rect 14090 11336 14096 11348
rect 14051 11308 14096 11336
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 14734 11296 14740 11348
rect 14792 11336 14798 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 14792 11308 15485 11336
rect 14792 11296 14798 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15746 11336 15752 11348
rect 15707 11308 15752 11336
rect 15473 11299 15531 11305
rect 15746 11296 15752 11308
rect 15804 11296 15810 11348
rect 16301 11339 16359 11345
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 17402 11336 17408 11348
rect 16347 11308 17408 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 17402 11296 17408 11308
rect 17460 11336 17466 11348
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 17460 11308 17969 11336
rect 17460 11296 17466 11308
rect 17957 11305 17969 11308
rect 18003 11305 18015 11339
rect 18506 11336 18512 11348
rect 18467 11308 18512 11336
rect 17957 11299 18015 11305
rect 18506 11296 18512 11308
rect 18564 11296 18570 11348
rect 19426 11296 19432 11348
rect 19484 11336 19490 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 19484 11308 19533 11336
rect 19484 11296 19490 11308
rect 19521 11305 19533 11308
rect 19567 11336 19579 11339
rect 20070 11336 20076 11348
rect 19567 11308 20076 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 20070 11296 20076 11308
rect 20128 11296 20134 11348
rect 20901 11339 20959 11345
rect 20901 11305 20913 11339
rect 20947 11336 20959 11339
rect 21082 11336 21088 11348
rect 20947 11308 21088 11336
rect 20947 11305 20959 11308
rect 20901 11299 20959 11305
rect 21082 11296 21088 11308
rect 21140 11296 21146 11348
rect 21269 11339 21327 11345
rect 21269 11305 21281 11339
rect 21315 11336 21327 11339
rect 21542 11336 21548 11348
rect 21315 11308 21548 11336
rect 21315 11305 21327 11308
rect 21269 11299 21327 11305
rect 21542 11296 21548 11308
rect 21600 11296 21606 11348
rect 21910 11336 21916 11348
rect 21871 11308 21916 11336
rect 21910 11296 21916 11308
rect 21968 11296 21974 11348
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 22465 11339 22523 11345
rect 22465 11336 22477 11339
rect 22428 11308 22477 11336
rect 22428 11296 22434 11308
rect 22465 11305 22477 11308
rect 22511 11305 22523 11339
rect 22922 11336 22928 11348
rect 22883 11308 22928 11336
rect 22465 11299 22523 11305
rect 22922 11296 22928 11308
rect 22980 11296 22986 11348
rect 23014 11296 23020 11348
rect 23072 11336 23078 11348
rect 23290 11336 23296 11348
rect 23072 11308 23296 11336
rect 23072 11296 23078 11308
rect 23290 11296 23296 11308
rect 23348 11296 23354 11348
rect 23934 11296 23940 11348
rect 23992 11336 23998 11348
rect 24029 11339 24087 11345
rect 24029 11336 24041 11339
rect 23992 11308 24041 11336
rect 23992 11296 23998 11308
rect 24029 11305 24041 11308
rect 24075 11305 24087 11339
rect 24029 11299 24087 11305
rect 24118 11296 24124 11348
rect 24176 11336 24182 11348
rect 24397 11339 24455 11345
rect 24397 11336 24409 11339
rect 24176 11308 24409 11336
rect 24176 11296 24182 11308
rect 24397 11305 24409 11308
rect 24443 11305 24455 11339
rect 24397 11299 24455 11305
rect 24489 11339 24547 11345
rect 24489 11305 24501 11339
rect 24535 11336 24547 11339
rect 24762 11336 24768 11348
rect 24535 11308 24768 11336
rect 24535 11305 24547 11308
rect 24489 11299 24547 11305
rect 2498 11228 2504 11280
rect 2556 11268 2562 11280
rect 2884 11268 2912 11296
rect 5626 11268 5632 11280
rect 2556 11240 2912 11268
rect 4540 11240 5632 11268
rect 2556 11228 2562 11240
rect 1394 11200 1400 11212
rect 1355 11172 1400 11200
rect 1394 11160 1400 11172
rect 1452 11160 1458 11212
rect 4430 11160 4436 11212
rect 4488 11200 4494 11212
rect 4540 11209 4568 11240
rect 5626 11228 5632 11240
rect 5684 11228 5690 11280
rect 7190 11228 7196 11280
rect 7248 11268 7254 11280
rect 7926 11268 7932 11280
rect 7248 11240 7932 11268
rect 7248 11228 7254 11240
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 10778 11268 10784 11280
rect 9692 11240 10784 11268
rect 9692 11212 9720 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 12066 11228 12072 11280
rect 12124 11268 12130 11280
rect 12980 11271 13038 11277
rect 12124 11240 12756 11268
rect 12124 11228 12130 11240
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4488 11172 4537 11200
rect 4488 11160 4494 11172
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 4614 11160 4620 11212
rect 4672 11200 4678 11212
rect 4781 11203 4839 11209
rect 4781 11200 4793 11203
rect 4672 11172 4793 11200
rect 4672 11160 4678 11172
rect 4781 11169 4793 11172
rect 4827 11200 4839 11203
rect 5350 11200 5356 11212
rect 4827 11172 5356 11200
rect 4827 11169 4839 11172
rect 4781 11163 4839 11169
rect 5350 11160 5356 11172
rect 5408 11160 5414 11212
rect 7558 11160 7564 11212
rect 7616 11200 7622 11212
rect 8110 11200 8116 11212
rect 7616 11172 8116 11200
rect 7616 11160 7622 11172
rect 8110 11160 8116 11172
rect 8168 11200 8174 11212
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 8168 11172 8217 11200
rect 8168 11160 8174 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 9582 11160 9588 11212
rect 9640 11160 9646 11212
rect 9674 11160 9680 11212
rect 9732 11160 9738 11212
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11200 10931 11203
rect 12526 11200 12532 11212
rect 10919 11172 12532 11200
rect 10919 11169 10931 11172
rect 10873 11163 10931 11169
rect 12526 11160 12532 11172
rect 12584 11160 12590 11212
rect 12728 11209 12756 11240
rect 12980 11237 12992 11271
rect 13026 11268 13038 11271
rect 13078 11268 13084 11280
rect 13026 11240 13084 11268
rect 13026 11237 13038 11240
rect 12980 11231 13038 11237
rect 13078 11228 13084 11240
rect 13136 11268 13142 11280
rect 13814 11268 13820 11280
rect 13136 11240 13820 11268
rect 13136 11228 13142 11240
rect 13814 11228 13820 11240
rect 13872 11228 13878 11280
rect 14642 11268 14648 11280
rect 14603 11240 14648 11268
rect 14642 11228 14648 11240
rect 14700 11228 14706 11280
rect 15562 11228 15568 11280
rect 15620 11268 15626 11280
rect 16758 11268 16764 11280
rect 15620 11240 16764 11268
rect 15620 11228 15626 11240
rect 12713 11203 12771 11209
rect 12713 11169 12725 11203
rect 12759 11200 12771 11203
rect 13538 11200 13544 11212
rect 12759 11172 13544 11200
rect 12759 11169 12771 11172
rect 12713 11163 12771 11169
rect 13538 11160 13544 11172
rect 13596 11160 13602 11212
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 15286 11200 15292 11212
rect 14792 11172 15292 11200
rect 14792 11160 14798 11172
rect 15286 11160 15292 11172
rect 15344 11160 15350 11212
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 3510 11132 3516 11144
rect 3099 11104 3516 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 3510 11092 3516 11104
rect 3568 11132 3574 11144
rect 4062 11132 4068 11144
rect 3568 11104 4068 11132
rect 3568 11092 3574 11104
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 7282 11092 7288 11144
rect 7340 11132 7346 11144
rect 8386 11132 8392 11144
rect 7340 11104 8392 11132
rect 7340 11092 7346 11104
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9600 11132 9628 11160
rect 9600 11104 9996 11132
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 1854 11064 1860 11076
rect 1627 11036 1860 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 1854 11024 1860 11036
rect 1912 11024 1918 11076
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2409 11067 2467 11073
rect 2409 11064 2421 11067
rect 2188 11036 2421 11064
rect 2188 11024 2194 11036
rect 2409 11033 2421 11036
rect 2455 11033 2467 11067
rect 2409 11027 2467 11033
rect 5905 11067 5963 11073
rect 5905 11033 5917 11067
rect 5951 11064 5963 11067
rect 6362 11064 6368 11076
rect 5951 11036 6368 11064
rect 5951 11033 5963 11036
rect 5905 11027 5963 11033
rect 6362 11024 6368 11036
rect 6420 11024 6426 11076
rect 7834 11064 7840 11076
rect 7795 11036 7840 11064
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 3881 10999 3939 11005
rect 3881 10965 3893 10999
rect 3927 10996 3939 10999
rect 3970 10996 3976 11008
rect 3927 10968 3976 10996
rect 3927 10965 3939 10968
rect 3881 10959 3939 10965
rect 3970 10956 3976 10968
rect 4028 10956 4034 11008
rect 5442 10956 5448 11008
rect 5500 10996 5506 11008
rect 6270 10996 6276 11008
rect 5500 10968 6276 10996
rect 5500 10956 5506 10968
rect 6270 10956 6276 10968
rect 6328 10956 6334 11008
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 8202 10996 8208 11008
rect 7616 10968 8208 10996
rect 7616 10956 7622 10968
rect 8202 10956 8208 10968
rect 8260 10956 8266 11008
rect 9217 10999 9275 11005
rect 9217 10965 9229 10999
rect 9263 10996 9275 10999
rect 9674 10996 9680 11008
rect 9263 10968 9680 10996
rect 9263 10965 9275 10968
rect 9217 10959 9275 10965
rect 9674 10956 9680 10968
rect 9732 10956 9738 11008
rect 9968 11005 9996 11104
rect 10778 11092 10784 11144
rect 10836 11132 10842 11144
rect 10965 11135 11023 11141
rect 10965 11132 10977 11135
rect 10836 11104 10977 11132
rect 10836 11092 10842 11104
rect 10965 11101 10977 11104
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11238 11132 11244 11144
rect 11195 11104 11244 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11238 11092 11244 11104
rect 11296 11132 11302 11144
rect 12434 11132 12440 11144
rect 11296 11104 12440 11132
rect 11296 11092 11302 11104
rect 12434 11092 12440 11104
rect 12492 11132 12498 11144
rect 16577 11135 16635 11141
rect 12492 11104 12585 11132
rect 12492 11092 12498 11104
rect 16577 11101 16589 11135
rect 16623 11132 16635 11135
rect 16684 11132 16712 11240
rect 16758 11228 16764 11240
rect 16816 11228 16822 11280
rect 18156 11240 19564 11268
rect 16850 11209 16856 11212
rect 16844 11200 16856 11209
rect 16811 11172 16856 11200
rect 16844 11163 16856 11172
rect 16850 11160 16856 11163
rect 16908 11160 16914 11212
rect 16623 11104 16712 11132
rect 16623 11101 16635 11104
rect 16577 11095 16635 11101
rect 10502 11064 10508 11076
rect 10463 11036 10508 11064
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 13780 11036 15025 11064
rect 13780 11024 13786 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15013 11027 15071 11033
rect 9953 10999 10011 11005
rect 9953 10965 9965 10999
rect 9999 10996 10011 10999
rect 11514 10996 11520 11008
rect 9999 10968 11520 10996
rect 9999 10965 10011 10968
rect 9953 10959 10011 10965
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14366 10996 14372 11008
rect 13872 10968 14372 10996
rect 13872 10956 13878 10968
rect 14366 10956 14372 10968
rect 14424 10996 14430 11008
rect 18156 10996 18184 11240
rect 19426 11200 19432 11212
rect 19387 11172 19432 11200
rect 19426 11160 19432 11172
rect 19484 11160 19490 11212
rect 19536 11200 19564 11240
rect 20990 11228 20996 11280
rect 21048 11268 21054 11280
rect 21361 11271 21419 11277
rect 21361 11268 21373 11271
rect 21048 11240 21373 11268
rect 21048 11228 21054 11240
rect 21361 11237 21373 11240
rect 21407 11237 21419 11271
rect 21560 11268 21588 11296
rect 22094 11268 22100 11280
rect 21560 11240 22100 11268
rect 21361 11231 21419 11237
rect 22094 11228 22100 11240
rect 22152 11228 22158 11280
rect 24412 11268 24440 11299
rect 24762 11296 24768 11308
rect 24820 11296 24826 11348
rect 25130 11336 25136 11348
rect 25091 11308 25136 11336
rect 25130 11296 25136 11308
rect 25188 11296 25194 11348
rect 25774 11336 25780 11348
rect 25735 11308 25780 11336
rect 25774 11296 25780 11308
rect 25832 11296 25838 11348
rect 25222 11268 25228 11280
rect 22204 11240 23520 11268
rect 24412 11240 25228 11268
rect 22204 11200 22232 11240
rect 19536 11172 22232 11200
rect 22373 11203 22431 11209
rect 22373 11169 22385 11203
rect 22419 11200 22431 11203
rect 22462 11200 22468 11212
rect 22419 11172 22468 11200
rect 22419 11169 22431 11172
rect 22373 11163 22431 11169
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22830 11200 22836 11212
rect 22791 11172 22836 11200
rect 22830 11160 22836 11172
rect 22888 11160 22894 11212
rect 23492 11200 23520 11240
rect 25222 11228 25228 11240
rect 25280 11228 25286 11280
rect 25406 11268 25412 11280
rect 25367 11240 25412 11268
rect 25406 11228 25412 11240
rect 25464 11228 25470 11280
rect 25590 11200 25596 11212
rect 23492 11172 25596 11200
rect 25590 11160 25596 11172
rect 25648 11200 25654 11212
rect 25774 11200 25780 11212
rect 25648 11172 25780 11200
rect 25648 11160 25654 11172
rect 25774 11160 25780 11172
rect 25832 11160 25838 11212
rect 18690 11092 18696 11144
rect 18748 11132 18754 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 18748 11104 19625 11132
rect 18748 11092 18754 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 20714 11092 20720 11144
rect 20772 11132 20778 11144
rect 21453 11135 21511 11141
rect 21453 11132 21465 11135
rect 20772 11104 21465 11132
rect 20772 11092 20778 11104
rect 21453 11101 21465 11104
rect 21499 11132 21511 11135
rect 23106 11132 23112 11144
rect 21499 11104 23112 11132
rect 21499 11101 21511 11104
rect 21453 11095 21511 11101
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24581 11135 24639 11141
rect 24581 11132 24593 11135
rect 24176 11104 24593 11132
rect 24176 11092 24182 11104
rect 24581 11101 24593 11104
rect 24627 11101 24639 11135
rect 24581 11095 24639 11101
rect 25314 11092 25320 11144
rect 25372 11092 25378 11144
rect 18874 11064 18880 11076
rect 18835 11036 18880 11064
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 19061 11067 19119 11073
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 19150 11064 19156 11076
rect 19107 11036 19156 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 19150 11024 19156 11036
rect 19208 11024 19214 11076
rect 19978 11024 19984 11076
rect 20036 11064 20042 11076
rect 25332 11064 25360 11092
rect 20036 11036 25360 11064
rect 20036 11024 20042 11036
rect 14424 10968 18184 10996
rect 14424 10956 14430 10968
rect 18414 10956 18420 11008
rect 18472 10996 18478 11008
rect 20073 10999 20131 11005
rect 20073 10996 20085 10999
rect 18472 10968 20085 10996
rect 18472 10956 18478 10968
rect 20073 10965 20085 10968
rect 20119 10996 20131 10999
rect 20254 10996 20260 11008
rect 20119 10968 20260 10996
rect 20119 10965 20131 10968
rect 20073 10959 20131 10965
rect 20254 10956 20260 10968
rect 20312 10956 20318 11008
rect 20717 10999 20775 11005
rect 20717 10965 20729 10999
rect 20763 10996 20775 10999
rect 20806 10996 20812 11008
rect 20763 10968 20812 10996
rect 20763 10965 20775 10968
rect 20717 10959 20775 10965
rect 20806 10956 20812 10968
rect 20864 10996 20870 11008
rect 21634 10996 21640 11008
rect 20864 10968 21640 10996
rect 20864 10956 20870 10968
rect 21634 10956 21640 10968
rect 21692 10956 21698 11008
rect 23753 10999 23811 11005
rect 23753 10965 23765 10999
rect 23799 10996 23811 10999
rect 24210 10996 24216 11008
rect 23799 10968 24216 10996
rect 23799 10965 23811 10968
rect 23753 10959 23811 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 25314 10956 25320 11008
rect 25372 10996 25378 11008
rect 26145 10999 26203 11005
rect 26145 10996 26157 10999
rect 25372 10968 26157 10996
rect 25372 10956 25378 10968
rect 26145 10965 26157 10968
rect 26191 10965 26203 10999
rect 26145 10959 26203 10965
rect 1104 10906 26864 10928
rect 1104 10854 5648 10906
rect 5700 10854 5712 10906
rect 5764 10854 5776 10906
rect 5828 10854 5840 10906
rect 5892 10854 14982 10906
rect 15034 10854 15046 10906
rect 15098 10854 15110 10906
rect 15162 10854 15174 10906
rect 15226 10854 24315 10906
rect 24367 10854 24379 10906
rect 24431 10854 24443 10906
rect 24495 10854 24507 10906
rect 24559 10854 26864 10906
rect 1104 10832 26864 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 4985 10795 5043 10801
rect 4985 10792 4997 10795
rect 4580 10764 4997 10792
rect 4580 10752 4586 10764
rect 4985 10761 4997 10764
rect 5031 10761 5043 10795
rect 4985 10755 5043 10761
rect 5169 10795 5227 10801
rect 5169 10761 5181 10795
rect 5215 10792 5227 10795
rect 5258 10792 5264 10804
rect 5215 10764 5264 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 4430 10684 4436 10736
rect 4488 10724 4494 10736
rect 4617 10727 4675 10733
rect 4617 10724 4629 10727
rect 4488 10696 4629 10724
rect 4488 10684 4494 10696
rect 4617 10693 4629 10696
rect 4663 10693 4675 10727
rect 4617 10687 4675 10693
rect 5000 10656 5028 10755
rect 5258 10752 5264 10764
rect 5316 10752 5322 10804
rect 5350 10752 5356 10804
rect 5408 10792 5414 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 5408 10764 6193 10792
rect 5408 10752 5414 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6546 10792 6552 10804
rect 6507 10764 6552 10792
rect 6181 10755 6239 10761
rect 6546 10752 6552 10764
rect 6604 10752 6610 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 11146 10792 11152 10804
rect 9171 10764 11152 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 12437 10795 12495 10801
rect 12437 10761 12449 10795
rect 12483 10792 12495 10795
rect 12618 10792 12624 10804
rect 12483 10764 12624 10792
rect 12483 10761 12495 10764
rect 12437 10755 12495 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 16758 10792 16764 10804
rect 16715 10764 16764 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 16758 10752 16764 10764
rect 16816 10752 16822 10804
rect 18322 10752 18328 10804
rect 18380 10792 18386 10804
rect 20717 10795 20775 10801
rect 18380 10764 20300 10792
rect 18380 10752 18386 10764
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5000 10628 5641 10656
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 5776 10628 5825 10656
rect 5776 10616 5782 10628
rect 5813 10625 5825 10628
rect 5859 10656 5871 10659
rect 6270 10656 6276 10668
rect 5859 10628 6276 10656
rect 5859 10625 5871 10628
rect 5813 10619 5871 10625
rect 6270 10616 6276 10628
rect 6328 10616 6334 10668
rect 6564 10656 6592 10752
rect 7285 10727 7343 10733
rect 7285 10693 7297 10727
rect 7331 10724 7343 10727
rect 7466 10724 7472 10736
rect 7331 10696 7472 10724
rect 7331 10693 7343 10696
rect 7285 10687 7343 10693
rect 7466 10684 7472 10696
rect 7524 10724 7530 10736
rect 8202 10724 8208 10736
rect 7524 10696 8208 10724
rect 7524 10684 7530 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 11698 10684 11704 10736
rect 11756 10724 11762 10736
rect 13814 10724 13820 10736
rect 11756 10696 13820 10724
rect 11756 10684 11762 10696
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 15654 10724 15660 10736
rect 15567 10696 15660 10724
rect 15654 10684 15660 10696
rect 15712 10724 15718 10736
rect 15712 10696 17080 10724
rect 15712 10684 15718 10696
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 6564 10628 7849 10656
rect 1397 10591 1455 10597
rect 1397 10557 1409 10591
rect 1443 10588 1455 10591
rect 2593 10591 2651 10597
rect 1443 10560 2084 10588
rect 1443 10557 1455 10560
rect 1397 10551 1455 10557
rect 2056 10464 2084 10560
rect 2593 10557 2605 10591
rect 2639 10588 2651 10591
rect 2685 10591 2743 10597
rect 2685 10588 2697 10591
rect 2639 10560 2697 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 2685 10557 2697 10560
rect 2731 10588 2743 10591
rect 3326 10588 3332 10600
rect 2731 10560 3332 10588
rect 2731 10557 2743 10560
rect 2685 10551 2743 10557
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 4798 10548 4804 10600
rect 4856 10588 4862 10600
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 4856 10560 5549 10588
rect 4856 10548 4862 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 2958 10529 2964 10532
rect 2952 10520 2964 10529
rect 2919 10492 2964 10520
rect 2952 10483 2964 10492
rect 2958 10480 2964 10483
rect 3016 10480 3022 10532
rect 6270 10480 6276 10532
rect 6328 10520 6334 10532
rect 6564 10520 6592 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 9674 10656 9680 10668
rect 9635 10628 9680 10656
rect 7837 10619 7895 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10229 10659 10287 10665
rect 10229 10625 10241 10659
rect 10275 10656 10287 10659
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 10275 10628 10609 10656
rect 10275 10625 10287 10628
rect 10229 10619 10287 10625
rect 10597 10625 10609 10628
rect 10643 10656 10655 10659
rect 11238 10656 11244 10668
rect 10643 10628 11244 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 13078 10656 13084 10668
rect 12115 10628 13084 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 13538 10656 13544 10668
rect 13451 10628 13544 10656
rect 13538 10616 13544 10628
rect 13596 10656 13602 10668
rect 13596 10628 13860 10656
rect 13596 10616 13602 10628
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10588 7251 10591
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7239 10560 7757 10588
rect 7239 10557 7251 10560
rect 7193 10551 7251 10557
rect 7745 10557 7757 10560
rect 7791 10588 7803 10591
rect 7926 10588 7932 10600
rect 7791 10560 7932 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 7926 10548 7932 10560
rect 7984 10548 7990 10600
rect 8938 10588 8944 10600
rect 8851 10560 8944 10588
rect 8938 10548 8944 10560
rect 8996 10588 9002 10600
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 8996 10560 9597 10588
rect 8996 10548 9002 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 11146 10588 11152 10600
rect 11107 10560 11152 10588
rect 9585 10551 9643 10557
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10588 12955 10591
rect 13722 10588 13728 10600
rect 12943 10560 13728 10588
rect 12943 10557 12955 10560
rect 12897 10551 12955 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 13832 10588 13860 10628
rect 14090 10616 14096 10668
rect 14148 10656 14154 10668
rect 14148 10628 14412 10656
rect 14148 10616 14154 10628
rect 14185 10591 14243 10597
rect 14185 10588 14197 10591
rect 13832 10560 14197 10588
rect 14185 10557 14197 10560
rect 14231 10588 14243 10591
rect 14277 10591 14335 10597
rect 14277 10588 14289 10591
rect 14231 10560 14289 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14277 10557 14289 10560
rect 14323 10557 14335 10591
rect 14384 10588 14412 10628
rect 17052 10600 17080 10696
rect 19426 10684 19432 10736
rect 19484 10724 19490 10736
rect 19613 10727 19671 10733
rect 19613 10724 19625 10727
rect 19484 10696 19625 10724
rect 19484 10684 19490 10696
rect 19613 10693 19625 10696
rect 19659 10724 19671 10727
rect 20070 10724 20076 10736
rect 19659 10696 20076 10724
rect 19659 10693 19671 10696
rect 19613 10687 19671 10693
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 20272 10724 20300 10764
rect 20717 10761 20729 10795
rect 20763 10792 20775 10795
rect 20990 10792 20996 10804
rect 20763 10764 20996 10792
rect 20763 10761 20775 10764
rect 20717 10755 20775 10761
rect 20990 10752 20996 10764
rect 21048 10752 21054 10804
rect 22094 10752 22100 10804
rect 22152 10792 22158 10804
rect 22189 10795 22247 10801
rect 22189 10792 22201 10795
rect 22152 10764 22201 10792
rect 22152 10752 22158 10764
rect 22189 10761 22201 10764
rect 22235 10761 22247 10795
rect 22189 10755 22247 10761
rect 22649 10795 22707 10801
rect 22649 10761 22661 10795
rect 22695 10792 22707 10795
rect 22922 10792 22928 10804
rect 22695 10764 22928 10792
rect 22695 10761 22707 10764
rect 22649 10755 22707 10761
rect 22922 10752 22928 10764
rect 22980 10752 22986 10804
rect 23106 10752 23112 10804
rect 23164 10792 23170 10804
rect 23293 10795 23351 10801
rect 23293 10792 23305 10795
rect 23164 10764 23305 10792
rect 23164 10752 23170 10764
rect 23293 10761 23305 10764
rect 23339 10761 23351 10795
rect 23293 10755 23351 10761
rect 23474 10752 23480 10804
rect 23532 10792 23538 10804
rect 24397 10795 24455 10801
rect 24397 10792 24409 10795
rect 23532 10764 24409 10792
rect 23532 10752 23538 10764
rect 24397 10761 24409 10764
rect 24443 10761 24455 10795
rect 24397 10755 24455 10761
rect 25222 10752 25228 10804
rect 25280 10792 25286 10804
rect 25501 10795 25559 10801
rect 25501 10792 25513 10795
rect 25280 10764 25513 10792
rect 25280 10752 25286 10764
rect 25501 10761 25513 10764
rect 25547 10761 25559 10795
rect 25501 10755 25559 10761
rect 21910 10724 21916 10736
rect 20272 10696 21916 10724
rect 21910 10684 21916 10696
rect 21968 10684 21974 10736
rect 24026 10684 24032 10736
rect 24084 10724 24090 10736
rect 24765 10727 24823 10733
rect 24765 10724 24777 10727
rect 24084 10696 24777 10724
rect 24084 10684 24090 10696
rect 24765 10693 24777 10696
rect 24811 10693 24823 10727
rect 24765 10687 24823 10693
rect 18506 10656 18512 10668
rect 18467 10628 18512 10656
rect 18506 10616 18512 10628
rect 18564 10616 18570 10668
rect 18690 10656 18696 10668
rect 18651 10628 18696 10656
rect 18690 10616 18696 10628
rect 18748 10616 18754 10668
rect 19518 10656 19524 10668
rect 19479 10628 19524 10656
rect 19518 10616 19524 10628
rect 19576 10656 19582 10668
rect 20254 10656 20260 10668
rect 19576 10628 20024 10656
rect 20215 10628 20260 10656
rect 19576 10616 19582 10628
rect 14550 10597 14556 10600
rect 14533 10591 14556 10597
rect 14533 10588 14545 10591
rect 14384 10560 14545 10588
rect 14277 10551 14335 10557
rect 14533 10557 14545 10560
rect 14608 10588 14614 10600
rect 14608 10560 14681 10588
rect 14533 10551 14556 10557
rect 6328 10492 6592 10520
rect 7653 10523 7711 10529
rect 6328 10480 6334 10492
rect 7653 10489 7665 10523
rect 7699 10520 7711 10523
rect 7834 10520 7840 10532
rect 7699 10492 7840 10520
rect 7699 10489 7711 10492
rect 7653 10483 7711 10489
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 8110 10480 8116 10532
rect 8168 10520 8174 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 8168 10492 8401 10520
rect 8168 10480 8174 10492
rect 8389 10489 8401 10492
rect 8435 10520 8447 10523
rect 9030 10520 9036 10532
rect 8435 10492 9036 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 9306 10480 9312 10532
rect 9364 10480 9370 10532
rect 12805 10523 12863 10529
rect 12805 10520 12817 10523
rect 10704 10492 12817 10520
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 3970 10412 3976 10464
rect 4028 10452 4034 10464
rect 4065 10455 4123 10461
rect 4065 10452 4077 10455
rect 4028 10424 4077 10452
rect 4028 10412 4034 10424
rect 4065 10421 4077 10424
rect 4111 10421 4123 10455
rect 4065 10415 4123 10421
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 7558 10452 7564 10464
rect 4304 10424 7564 10452
rect 4304 10412 4310 10424
rect 7558 10412 7564 10424
rect 7616 10412 7622 10464
rect 8846 10412 8852 10464
rect 8904 10452 8910 10464
rect 9324 10452 9352 10480
rect 10704 10461 10732 10492
rect 12805 10489 12817 10492
rect 12851 10520 12863 10523
rect 14292 10520 14320 10551
rect 14550 10548 14556 10551
rect 14608 10548 14614 10560
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16632 10560 16773 10588
rect 16632 10548 16638 10560
rect 16761 10557 16773 10560
rect 16807 10557 16819 10591
rect 16761 10551 16819 10557
rect 17034 10548 17040 10600
rect 17092 10588 17098 10600
rect 17497 10591 17555 10597
rect 17497 10588 17509 10591
rect 17092 10560 17509 10588
rect 17092 10548 17098 10560
rect 17497 10557 17509 10560
rect 17543 10588 17555 10591
rect 18708 10588 18736 10616
rect 19996 10597 20024 10628
rect 20254 10616 20260 10628
rect 20312 10616 20318 10668
rect 21634 10616 21640 10668
rect 21692 10656 21698 10668
rect 21729 10659 21787 10665
rect 21729 10656 21741 10659
rect 21692 10628 21741 10656
rect 21692 10616 21698 10628
rect 21729 10625 21741 10628
rect 21775 10625 21787 10659
rect 21729 10619 21787 10625
rect 23106 10616 23112 10668
rect 23164 10656 23170 10668
rect 23290 10656 23296 10668
rect 23164 10628 23296 10656
rect 23164 10616 23170 10628
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 25869 10659 25927 10665
rect 25869 10656 25881 10659
rect 23400 10628 25881 10656
rect 17543 10560 18736 10588
rect 19981 10591 20039 10597
rect 17543 10557 17555 10560
rect 17497 10551 17555 10557
rect 19981 10557 19993 10591
rect 20027 10557 20039 10591
rect 21542 10588 21548 10600
rect 21503 10560 21548 10588
rect 19981 10551 20039 10557
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 23400 10588 23428 10628
rect 25869 10625 25881 10628
rect 25915 10625 25927 10659
rect 25869 10619 25927 10625
rect 21744 10560 23428 10588
rect 21744 10532 21772 10560
rect 23934 10548 23940 10600
rect 23992 10588 23998 10600
rect 24581 10591 24639 10597
rect 24581 10588 24593 10591
rect 23992 10560 24593 10588
rect 23992 10548 23998 10560
rect 24581 10557 24593 10560
rect 24627 10588 24639 10591
rect 25133 10591 25191 10597
rect 25133 10588 25145 10591
rect 24627 10560 25145 10588
rect 24627 10557 24639 10560
rect 24581 10551 24639 10557
rect 25133 10557 25145 10560
rect 25179 10557 25191 10591
rect 25133 10551 25191 10557
rect 15562 10520 15568 10532
rect 12851 10492 13768 10520
rect 14292 10492 15568 10520
rect 12851 10489 12863 10492
rect 12805 10483 12863 10489
rect 13740 10464 13768 10492
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 16022 10480 16028 10532
rect 16080 10520 16086 10532
rect 17773 10523 17831 10529
rect 17773 10520 17785 10523
rect 16080 10492 17785 10520
rect 16080 10480 16086 10492
rect 17773 10489 17785 10492
rect 17819 10520 17831 10523
rect 17954 10520 17960 10532
rect 17819 10492 17960 10520
rect 17819 10489 17831 10492
rect 17773 10483 17831 10489
rect 17954 10480 17960 10492
rect 18012 10520 18018 10532
rect 18417 10523 18475 10529
rect 18417 10520 18429 10523
rect 18012 10492 18429 10520
rect 18012 10480 18018 10492
rect 18417 10489 18429 10492
rect 18463 10489 18475 10523
rect 18417 10483 18475 10489
rect 20898 10480 20904 10532
rect 20956 10520 20962 10532
rect 21082 10520 21088 10532
rect 20956 10492 21088 10520
rect 20956 10480 20962 10492
rect 21082 10480 21088 10492
rect 21140 10520 21146 10532
rect 21637 10523 21695 10529
rect 21637 10520 21649 10523
rect 21140 10492 21649 10520
rect 21140 10480 21146 10492
rect 21637 10489 21649 10492
rect 21683 10489 21695 10523
rect 21637 10483 21695 10489
rect 21726 10480 21732 10532
rect 21784 10480 21790 10532
rect 22002 10480 22008 10532
rect 22060 10520 22066 10532
rect 24029 10523 24087 10529
rect 24029 10520 24041 10523
rect 22060 10492 24041 10520
rect 22060 10480 22066 10492
rect 24029 10489 24041 10492
rect 24075 10520 24087 10523
rect 24118 10520 24124 10532
rect 24075 10492 24124 10520
rect 24075 10489 24087 10492
rect 24029 10483 24087 10489
rect 24118 10480 24124 10492
rect 24176 10480 24182 10532
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 8904 10424 9505 10452
rect 8904 10412 8910 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10421 10747 10455
rect 11054 10452 11060 10464
rect 11015 10424 11060 10452
rect 10689 10415 10747 10421
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11885 10455 11943 10461
rect 11885 10421 11897 10455
rect 11931 10452 11943 10455
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11931 10424 12081 10452
rect 11931 10421 11943 10424
rect 11885 10415 11943 10421
rect 12069 10421 12081 10424
rect 12115 10452 12127 10455
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 12115 10424 12173 10452
rect 12115 10421 12127 10424
rect 12069 10415 12127 10421
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 13722 10412 13728 10464
rect 13780 10412 13786 10464
rect 16206 10452 16212 10464
rect 16167 10424 16212 10452
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 18046 10452 18052 10464
rect 18007 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 18230 10412 18236 10464
rect 18288 10452 18294 10464
rect 19058 10452 19064 10464
rect 18288 10424 19064 10452
rect 18288 10412 18294 10424
rect 19058 10412 19064 10424
rect 19116 10452 19122 10464
rect 20073 10455 20131 10461
rect 20073 10452 20085 10455
rect 19116 10424 20085 10452
rect 19116 10412 19122 10424
rect 20073 10421 20085 10424
rect 20119 10421 20131 10455
rect 21174 10452 21180 10464
rect 21135 10424 21180 10452
rect 20073 10415 20131 10421
rect 21174 10412 21180 10424
rect 21232 10412 21238 10464
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 22925 10455 22983 10461
rect 22925 10452 22937 10455
rect 22888 10424 22937 10452
rect 22888 10412 22894 10424
rect 22925 10421 22937 10424
rect 22971 10421 22983 10455
rect 22925 10415 22983 10421
rect 23934 10412 23940 10464
rect 23992 10452 23998 10464
rect 25406 10452 25412 10464
rect 23992 10424 25412 10452
rect 23992 10412 23998 10424
rect 25406 10412 25412 10424
rect 25464 10412 25470 10464
rect 26326 10452 26332 10464
rect 26287 10424 26332 10452
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 1104 10362 26864 10384
rect 1104 10310 10315 10362
rect 10367 10310 10379 10362
rect 10431 10310 10443 10362
rect 10495 10310 10507 10362
rect 10559 10310 19648 10362
rect 19700 10310 19712 10362
rect 19764 10310 19776 10362
rect 19828 10310 19840 10362
rect 19892 10310 26864 10362
rect 1104 10288 26864 10310
rect 2317 10251 2375 10257
rect 2317 10217 2329 10251
rect 2363 10248 2375 10251
rect 2498 10248 2504 10260
rect 2363 10220 2504 10248
rect 2363 10217 2375 10220
rect 2317 10211 2375 10217
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 2590 10208 2596 10260
rect 2648 10248 2654 10260
rect 2866 10248 2872 10260
rect 2648 10220 2872 10248
rect 2648 10208 2654 10220
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3142 10208 3148 10260
rect 3200 10248 3206 10260
rect 3694 10248 3700 10260
rect 3200 10220 3700 10248
rect 3200 10208 3206 10220
rect 3694 10208 3700 10220
rect 3752 10248 3758 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3752 10220 4077 10248
rect 3752 10208 3758 10220
rect 4065 10217 4077 10220
rect 4111 10217 4123 10251
rect 4065 10211 4123 10217
rect 4338 10208 4344 10260
rect 4396 10248 4402 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 4396 10220 4445 10248
rect 4396 10208 4402 10220
rect 4433 10217 4445 10220
rect 4479 10217 4491 10251
rect 4433 10211 4491 10217
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10248 4583 10251
rect 4706 10248 4712 10260
rect 4571 10220 4712 10248
rect 4571 10217 4583 10220
rect 4525 10211 4583 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 5169 10251 5227 10257
rect 5169 10248 5181 10251
rect 4856 10220 5181 10248
rect 4856 10208 4862 10220
rect 5169 10217 5181 10220
rect 5215 10217 5227 10251
rect 5169 10211 5227 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10248 5687 10251
rect 5718 10248 5724 10260
rect 5675 10220 5724 10248
rect 5675 10217 5687 10220
rect 5629 10211 5687 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 5902 10248 5908 10260
rect 5863 10220 5908 10248
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 7742 10248 7748 10260
rect 7703 10220 7748 10248
rect 7742 10208 7748 10220
rect 7800 10208 7806 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8110 10248 8116 10260
rect 7984 10220 8116 10248
rect 7984 10208 7990 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8754 10248 8760 10260
rect 8715 10220 8760 10248
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 9861 10251 9919 10257
rect 9861 10217 9873 10251
rect 9907 10248 9919 10251
rect 9950 10248 9956 10260
rect 9907 10220 9956 10248
rect 9907 10217 9919 10220
rect 9861 10211 9919 10217
rect 9950 10208 9956 10220
rect 10008 10208 10014 10260
rect 10134 10248 10140 10260
rect 10095 10220 10140 10248
rect 10134 10208 10140 10220
rect 10192 10208 10198 10260
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 12437 10251 12495 10257
rect 12437 10217 12449 10251
rect 12483 10248 12495 10251
rect 12526 10248 12532 10260
rect 12483 10220 12532 10248
rect 12483 10217 12495 10220
rect 12437 10211 12495 10217
rect 12526 10208 12532 10220
rect 12584 10248 12590 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 12584 10220 13829 10248
rect 12584 10208 12590 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 14550 10208 14556 10260
rect 14608 10248 14614 10260
rect 14645 10251 14703 10257
rect 14645 10248 14657 10251
rect 14608 10220 14657 10248
rect 14608 10208 14614 10220
rect 14645 10217 14657 10220
rect 14691 10217 14703 10251
rect 14645 10211 14703 10217
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15473 10251 15531 10257
rect 15473 10248 15485 10251
rect 15252 10220 15485 10248
rect 15252 10208 15258 10220
rect 15473 10217 15485 10220
rect 15519 10217 15531 10251
rect 16942 10248 16948 10260
rect 16903 10220 16948 10248
rect 15473 10211 15531 10217
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 17770 10208 17776 10260
rect 17828 10248 17834 10260
rect 17957 10251 18015 10257
rect 17957 10248 17969 10251
rect 17828 10220 17969 10248
rect 17828 10208 17834 10220
rect 17957 10217 17969 10220
rect 18003 10217 18015 10251
rect 17957 10211 18015 10217
rect 18414 10208 18420 10260
rect 18472 10248 18478 10260
rect 18509 10251 18567 10257
rect 18509 10248 18521 10251
rect 18472 10220 18521 10248
rect 18472 10208 18478 10220
rect 18509 10217 18521 10220
rect 18555 10217 18567 10251
rect 18509 10211 18567 10217
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18748 10220 18889 10248
rect 18748 10208 18754 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 19426 10248 19432 10260
rect 19339 10220 19432 10248
rect 18877 10211 18935 10217
rect 19426 10208 19432 10220
rect 19484 10248 19490 10260
rect 21358 10248 21364 10260
rect 19484 10220 21364 10248
rect 19484 10208 19490 10220
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 21913 10251 21971 10257
rect 21913 10248 21925 10251
rect 21600 10220 21925 10248
rect 21600 10208 21606 10220
rect 21913 10217 21925 10220
rect 21959 10217 21971 10251
rect 22278 10248 22284 10260
rect 22239 10220 22284 10248
rect 21913 10211 21971 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 23014 10248 23020 10260
rect 22975 10220 23020 10248
rect 23014 10208 23020 10220
rect 23072 10208 23078 10260
rect 23474 10248 23480 10260
rect 23435 10220 23480 10248
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 23566 10208 23572 10260
rect 23624 10248 23630 10260
rect 23753 10251 23811 10257
rect 23753 10248 23765 10251
rect 23624 10220 23765 10248
rect 23624 10208 23630 10220
rect 23753 10217 23765 10220
rect 23799 10217 23811 10251
rect 23753 10211 23811 10217
rect 24489 10251 24547 10257
rect 24489 10217 24501 10251
rect 24535 10248 24547 10251
rect 24762 10248 24768 10260
rect 24535 10220 24768 10248
rect 24535 10217 24547 10220
rect 24489 10211 24547 10217
rect 24762 10208 24768 10220
rect 24820 10208 24826 10260
rect 25130 10208 25136 10260
rect 25188 10248 25194 10260
rect 25501 10251 25559 10257
rect 25501 10248 25513 10251
rect 25188 10220 25513 10248
rect 25188 10208 25194 10220
rect 25501 10217 25513 10220
rect 25547 10217 25559 10251
rect 25501 10211 25559 10217
rect 25682 10208 25688 10260
rect 25740 10248 25746 10260
rect 25869 10251 25927 10257
rect 25869 10248 25881 10251
rect 25740 10220 25881 10248
rect 25740 10208 25746 10220
rect 25869 10217 25881 10220
rect 25915 10217 25927 10251
rect 26326 10248 26332 10260
rect 26287 10220 26332 10248
rect 25869 10211 25927 10217
rect 26326 10208 26332 10220
rect 26384 10208 26390 10260
rect 2777 10183 2835 10189
rect 2777 10149 2789 10183
rect 2823 10180 2835 10183
rect 3878 10180 3884 10192
rect 2823 10152 3884 10180
rect 2823 10149 2835 10152
rect 2777 10143 2835 10149
rect 3878 10140 3884 10152
rect 3936 10140 3942 10192
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 6236 10152 6684 10180
rect 6236 10140 6242 10152
rect 2869 10115 2927 10121
rect 2869 10081 2881 10115
rect 2915 10112 2927 10115
rect 3050 10112 3056 10124
rect 2915 10084 3056 10112
rect 2915 10081 2927 10084
rect 2869 10075 2927 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 6546 10112 6552 10124
rect 6507 10084 6552 10112
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6656 10112 6684 10152
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 7340 10152 7389 10180
rect 7340 10140 7346 10152
rect 7377 10149 7389 10152
rect 7423 10180 7435 10183
rect 7834 10180 7840 10192
rect 7423 10152 7840 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 7834 10140 7840 10152
rect 7892 10140 7898 10192
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 10689 10183 10747 10189
rect 10689 10180 10701 10183
rect 9640 10152 10701 10180
rect 9640 10140 9646 10152
rect 10689 10149 10701 10152
rect 10735 10180 10747 10183
rect 10870 10180 10876 10192
rect 10735 10152 10876 10180
rect 10735 10149 10747 10152
rect 10689 10143 10747 10149
rect 10870 10140 10876 10152
rect 10928 10180 10934 10192
rect 10928 10152 13124 10180
rect 10928 10140 10934 10152
rect 9674 10112 9680 10124
rect 6656 10084 6776 10112
rect 9635 10084 9680 10112
rect 2958 10044 2964 10056
rect 2871 10016 2964 10044
rect 2958 10004 2964 10016
rect 3016 10044 3022 10056
rect 3016 10016 3096 10044
rect 3016 10004 3022 10016
rect 2406 9976 2412 9988
rect 2367 9948 2412 9976
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 3068 9920 3096 10016
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4617 10047 4675 10053
rect 4617 10044 4629 10047
rect 4212 10016 4629 10044
rect 4212 10004 4218 10016
rect 4617 10013 4629 10016
rect 4663 10013 4675 10047
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 4617 10007 4675 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 6748 10053 6776 10084
rect 9674 10072 9680 10084
rect 9732 10072 9738 10124
rect 11238 10112 11244 10124
rect 11199 10084 11244 10112
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11348 10112 11376 10152
rect 11882 10112 11888 10124
rect 11348 10084 11468 10112
rect 11843 10084 11888 10112
rect 6733 10047 6791 10053
rect 6733 10013 6745 10047
rect 6779 10013 6791 10047
rect 8202 10044 8208 10056
rect 8163 10016 8208 10044
rect 6733 10007 6791 10013
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 8386 10044 8392 10056
rect 8347 10016 8392 10044
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9306 10004 9312 10056
rect 9364 10044 9370 10056
rect 11146 10044 11152 10056
rect 9364 10016 11152 10044
rect 9364 10004 9370 10016
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11440 10053 11468 10084
rect 11882 10072 11888 10084
rect 11940 10072 11946 10124
rect 12526 10072 12532 10124
rect 12584 10112 12590 10124
rect 12802 10112 12808 10124
rect 12584 10084 12808 10112
rect 12584 10072 12590 10084
rect 12802 10072 12808 10084
rect 12860 10072 12866 10124
rect 13096 10056 13124 10152
rect 16206 10140 16212 10192
rect 16264 10180 16270 10192
rect 16850 10180 16856 10192
rect 16264 10152 16856 10180
rect 16264 10140 16270 10152
rect 16850 10140 16856 10152
rect 16908 10180 16914 10192
rect 17313 10183 17371 10189
rect 17313 10180 17325 10183
rect 16908 10152 17325 10180
rect 16908 10140 16914 10152
rect 17313 10149 17325 10152
rect 17359 10180 17371 10183
rect 24026 10180 24032 10192
rect 17359 10152 18092 10180
rect 23987 10152 24032 10180
rect 17359 10149 17371 10152
rect 17313 10143 17371 10149
rect 14185 10115 14243 10121
rect 14185 10081 14197 10115
rect 14231 10112 14243 10115
rect 16298 10112 16304 10124
rect 14231 10084 16304 10112
rect 14231 10081 14243 10084
rect 14185 10075 14243 10081
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 17862 10112 17868 10124
rect 17823 10084 17868 10112
rect 17862 10072 17868 10084
rect 17920 10072 17926 10124
rect 11425 10047 11483 10053
rect 11425 10013 11437 10047
rect 11471 10013 11483 10047
rect 11425 10007 11483 10013
rect 12345 10047 12403 10053
rect 12345 10013 12357 10047
rect 12391 10044 12403 10047
rect 12434 10044 12440 10056
rect 12391 10016 12440 10044
rect 12391 10013 12403 10016
rect 12345 10007 12403 10013
rect 12434 10004 12440 10016
rect 12492 10044 12498 10056
rect 12897 10047 12955 10053
rect 12897 10044 12909 10047
rect 12492 10016 12909 10044
rect 12492 10004 12498 10016
rect 12897 10013 12909 10016
rect 12943 10013 12955 10047
rect 13078 10044 13084 10056
rect 13039 10016 13084 10044
rect 12897 10007 12955 10013
rect 13078 10004 13084 10016
rect 13136 10004 13142 10056
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 15746 10044 15752 10056
rect 14516 10016 15752 10044
rect 14516 10004 14522 10016
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16390 10044 16396 10056
rect 16351 10016 16396 10044
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 17034 10044 17040 10056
rect 16623 10016 17040 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6181 9979 6239 9985
rect 6181 9976 6193 9979
rect 5868 9948 6193 9976
rect 5868 9936 5874 9948
rect 6181 9945 6193 9948
rect 6227 9945 6239 9979
rect 6181 9939 6239 9945
rect 8110 9936 8116 9988
rect 8168 9976 8174 9988
rect 8404 9976 8432 10004
rect 8168 9948 8432 9976
rect 10873 9979 10931 9985
rect 8168 9936 8174 9948
rect 10873 9945 10885 9979
rect 10919 9976 10931 9979
rect 11054 9976 11060 9988
rect 10919 9948 11060 9976
rect 10919 9945 10931 9948
rect 10873 9939 10931 9945
rect 11054 9936 11060 9948
rect 11112 9976 11118 9988
rect 15013 9979 15071 9985
rect 15013 9976 15025 9979
rect 11112 9948 15025 9976
rect 11112 9936 11118 9948
rect 15013 9945 15025 9948
rect 15059 9945 15071 9979
rect 15013 9939 15071 9945
rect 15933 9979 15991 9985
rect 15933 9945 15945 9979
rect 15979 9976 15991 9979
rect 17880 9976 17908 10072
rect 18064 10053 18092 10152
rect 24026 10140 24032 10152
rect 24084 10140 24090 10192
rect 20898 10072 20904 10124
rect 20956 10112 20962 10124
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 20956 10084 21281 10112
rect 20956 10072 20962 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 22002 10112 22008 10124
rect 21407 10084 22008 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 22002 10072 22008 10084
rect 22060 10072 22066 10124
rect 22186 10072 22192 10124
rect 22244 10112 22250 10124
rect 22557 10115 22615 10121
rect 22557 10112 22569 10115
rect 22244 10084 22569 10112
rect 22244 10072 22250 10084
rect 22557 10081 22569 10084
rect 22603 10112 22615 10115
rect 22922 10112 22928 10124
rect 22603 10084 22928 10112
rect 22603 10081 22615 10084
rect 22557 10075 22615 10081
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 23569 10115 23627 10121
rect 23569 10081 23581 10115
rect 23615 10112 23627 10115
rect 23658 10112 23664 10124
rect 23615 10084 23664 10112
rect 23615 10081 23627 10084
rect 23569 10075 23627 10081
rect 23658 10072 23664 10084
rect 23716 10072 23722 10124
rect 23750 10072 23756 10124
rect 23808 10112 23814 10124
rect 24118 10112 24124 10124
rect 23808 10084 24124 10112
rect 23808 10072 23814 10084
rect 24118 10072 24124 10084
rect 24176 10112 24182 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 24176 10084 24593 10112
rect 24176 10072 24182 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 24946 10072 24952 10124
rect 25004 10112 25010 10124
rect 25133 10115 25191 10121
rect 25133 10112 25145 10115
rect 25004 10084 25145 10112
rect 25004 10072 25010 10084
rect 25133 10081 25145 10084
rect 25179 10081 25191 10115
rect 25133 10075 25191 10081
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10044 19579 10047
rect 19610 10044 19616 10056
rect 19567 10016 19616 10044
rect 19567 10013 19579 10016
rect 19521 10007 19579 10013
rect 19610 10004 19616 10016
rect 19668 10004 19674 10056
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10044 19763 10047
rect 20254 10044 20260 10056
rect 19751 10016 20260 10044
rect 19751 10013 19763 10016
rect 19705 10007 19763 10013
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21634 10044 21640 10056
rect 21591 10016 21640 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21634 10004 21640 10016
rect 21692 10044 21698 10056
rect 22646 10044 22652 10056
rect 21692 10016 22652 10044
rect 21692 10004 21698 10016
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 15979 9948 17908 9976
rect 15979 9945 15991 9948
rect 15933 9939 15991 9945
rect 20438 9936 20444 9988
rect 20496 9976 20502 9988
rect 21726 9976 21732 9988
rect 20496 9948 21732 9976
rect 20496 9936 20502 9948
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 22741 9979 22799 9985
rect 22741 9945 22753 9979
rect 22787 9976 22799 9979
rect 23382 9976 23388 9988
rect 22787 9948 23388 9976
rect 22787 9945 22799 9948
rect 22741 9939 22799 9945
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 24765 9979 24823 9985
rect 24765 9945 24777 9979
rect 24811 9976 24823 9979
rect 25958 9976 25964 9988
rect 24811 9948 25964 9976
rect 24811 9945 24823 9948
rect 24765 9939 24823 9945
rect 25958 9936 25964 9948
rect 26016 9936 26022 9988
rect 1946 9908 1952 9920
rect 1907 9880 1952 9908
rect 1946 9868 1952 9880
rect 2004 9868 2010 9920
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3513 9911 3571 9917
rect 3513 9908 3525 9911
rect 3108 9880 3525 9908
rect 3108 9868 3114 9880
rect 3513 9877 3525 9880
rect 3559 9877 3571 9911
rect 3513 9871 3571 9877
rect 3602 9868 3608 9920
rect 3660 9908 3666 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3660 9880 3801 9908
rect 3660 9868 3666 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 8846 9908 8852 9920
rect 8444 9880 8852 9908
rect 8444 9868 8450 9880
rect 8846 9868 8852 9880
rect 8904 9908 8910 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 8904 9880 9137 9908
rect 8904 9868 8910 9880
rect 9125 9877 9137 9880
rect 9171 9877 9183 9911
rect 13446 9908 13452 9920
rect 13407 9880 13452 9908
rect 9125 9871 9183 9877
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13630 9868 13636 9920
rect 13688 9908 13694 9920
rect 18782 9908 18788 9920
rect 13688 9880 18788 9908
rect 13688 9868 13694 9880
rect 18782 9868 18788 9880
rect 18840 9868 18846 9920
rect 19058 9908 19064 9920
rect 19019 9880 19064 9908
rect 19058 9868 19064 9880
rect 19116 9868 19122 9920
rect 20070 9908 20076 9920
rect 20031 9880 20076 9908
rect 20070 9868 20076 9880
rect 20128 9868 20134 9920
rect 20714 9908 20720 9920
rect 20675 9880 20720 9908
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 20901 9911 20959 9917
rect 20901 9877 20913 9911
rect 20947 9908 20959 9911
rect 21634 9908 21640 9920
rect 20947 9880 21640 9908
rect 20947 9877 20959 9880
rect 20901 9871 20959 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 22278 9868 22284 9920
rect 22336 9908 22342 9920
rect 22830 9908 22836 9920
rect 22336 9880 22836 9908
rect 22336 9868 22342 9880
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 1104 9818 26864 9840
rect 1104 9766 5648 9818
rect 5700 9766 5712 9818
rect 5764 9766 5776 9818
rect 5828 9766 5840 9818
rect 5892 9766 14982 9818
rect 15034 9766 15046 9818
rect 15098 9766 15110 9818
rect 15162 9766 15174 9818
rect 15226 9766 24315 9818
rect 24367 9766 24379 9818
rect 24431 9766 24443 9818
rect 24495 9766 24507 9818
rect 24559 9766 26864 9818
rect 1104 9744 26864 9766
rect 5905 9707 5963 9713
rect 5905 9673 5917 9707
rect 5951 9704 5963 9707
rect 6178 9704 6184 9716
rect 5951 9676 6184 9704
rect 5951 9673 5963 9676
rect 5905 9667 5963 9673
rect 6178 9664 6184 9676
rect 6236 9664 6242 9716
rect 6454 9664 6460 9716
rect 6512 9704 6518 9716
rect 6914 9704 6920 9716
rect 6512 9676 6920 9704
rect 6512 9664 6518 9676
rect 6914 9664 6920 9676
rect 6972 9664 6978 9716
rect 8202 9704 8208 9716
rect 8163 9676 8208 9704
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 11057 9707 11115 9713
rect 11057 9673 11069 9707
rect 11103 9704 11115 9707
rect 11146 9704 11152 9716
rect 11103 9676 11152 9704
rect 11103 9673 11115 9676
rect 11057 9667 11115 9673
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 11333 9707 11391 9713
rect 11333 9704 11345 9707
rect 11296 9676 11345 9704
rect 11296 9664 11302 9676
rect 11333 9673 11345 9676
rect 11379 9673 11391 9707
rect 12342 9704 12348 9716
rect 11333 9667 11391 9673
rect 12268 9676 12348 9704
rect 7101 9639 7159 9645
rect 7101 9605 7113 9639
rect 7147 9636 7159 9639
rect 8018 9636 8024 9648
rect 7147 9608 8024 9636
rect 7147 9605 7159 9608
rect 7101 9599 7159 9605
rect 8018 9596 8024 9608
rect 8076 9596 8082 9648
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2222 9568 2228 9580
rect 1719 9540 2228 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2222 9528 2228 9540
rect 2280 9568 2286 9580
rect 2409 9571 2467 9577
rect 2409 9568 2421 9571
rect 2280 9540 2421 9568
rect 2280 9528 2286 9540
rect 2409 9537 2421 9540
rect 2455 9568 2467 9571
rect 3050 9568 3056 9580
rect 2455 9540 3056 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 3050 9528 3056 9540
rect 3108 9528 3114 9580
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3326 9568 3332 9580
rect 3283 9540 3332 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 7190 9528 7196 9580
rect 7248 9568 7254 9580
rect 7650 9568 7656 9580
rect 7248 9540 7656 9568
rect 7248 9528 7254 9540
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 7984 9540 8493 9568
rect 7984 9528 7990 9540
rect 8481 9537 8493 9540
rect 8527 9568 8539 9571
rect 8846 9568 8852 9580
rect 8527 9540 8852 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 8956 9540 9168 9568
rect 2130 9460 2136 9512
rect 2188 9460 2194 9512
rect 3142 9500 3148 9512
rect 2424 9472 3148 9500
rect 2148 9432 2176 9460
rect 2225 9435 2283 9441
rect 2225 9432 2237 9435
rect 2148 9404 2237 9432
rect 2225 9401 2237 9404
rect 2271 9401 2283 9435
rect 2225 9395 2283 9401
rect 1762 9364 1768 9376
rect 1723 9336 1768 9364
rect 1762 9324 1768 9336
rect 1820 9324 1826 9376
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2424 9364 2452 9472
rect 3142 9460 3148 9472
rect 3200 9460 3206 9512
rect 6273 9503 6331 9509
rect 6273 9469 6285 9503
rect 6319 9500 6331 9503
rect 7469 9503 7527 9509
rect 7469 9500 7481 9503
rect 6319 9472 7481 9500
rect 6319 9469 6331 9472
rect 6273 9463 6331 9469
rect 7469 9469 7481 9472
rect 7515 9500 7527 9503
rect 8662 9500 8668 9512
rect 7515 9472 8668 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 8662 9460 8668 9472
rect 8720 9460 8726 9512
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2777 9435 2835 9441
rect 2777 9432 2789 9435
rect 2556 9404 2789 9432
rect 2556 9392 2562 9404
rect 2777 9401 2789 9404
rect 2823 9432 2835 9435
rect 2958 9432 2964 9444
rect 2823 9404 2964 9432
rect 2823 9401 2835 9404
rect 2777 9395 2835 9401
rect 2958 9392 2964 9404
rect 3016 9432 3022 9444
rect 3596 9435 3654 9441
rect 3596 9432 3608 9435
rect 3016 9404 3608 9432
rect 3016 9392 3022 9404
rect 3596 9401 3608 9404
rect 3642 9432 3654 9435
rect 4154 9432 4160 9444
rect 3642 9404 4160 9432
rect 3642 9401 3654 9404
rect 3596 9395 3654 9401
rect 4154 9392 4160 9404
rect 4212 9432 4218 9444
rect 5261 9435 5319 9441
rect 5261 9432 5273 9435
rect 4212 9404 5273 9432
rect 4212 9392 4218 9404
rect 5261 9401 5273 9404
rect 5307 9401 5319 9435
rect 8956 9432 8984 9540
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9140 9500 9168 9540
rect 9582 9500 9588 9512
rect 9140 9472 9588 9500
rect 9033 9463 9091 9469
rect 5261 9395 5319 9401
rect 7576 9404 8984 9432
rect 2179 9336 2452 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 3050 9324 3056 9376
rect 3108 9364 3114 9376
rect 4706 9364 4712 9376
rect 3108 9336 4712 9364
rect 3108 9324 3114 9336
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 7576 9373 7604 9404
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 5960 9336 6561 9364
rect 5960 9324 5966 9336
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 6595 9336 7573 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7561 9327 7619 9333
rect 7650 9324 7656 9376
rect 7708 9364 7714 9376
rect 8570 9364 8576 9376
rect 7708 9336 8576 9364
rect 7708 9324 7714 9336
rect 8570 9324 8576 9336
rect 8628 9364 8634 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8628 9336 8861 9364
rect 8628 9324 8634 9336
rect 8849 9333 8861 9336
rect 8895 9364 8907 9367
rect 9048 9364 9076 9463
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 11348 9500 11376 9667
rect 12069 9639 12127 9645
rect 12069 9605 12081 9639
rect 12115 9636 12127 9639
rect 12268 9636 12296 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12434 9664 12440 9716
rect 12492 9704 12498 9716
rect 12492 9676 12537 9704
rect 12492 9664 12498 9676
rect 13078 9664 13084 9716
rect 13136 9704 13142 9716
rect 15197 9707 15255 9713
rect 13136 9676 13768 9704
rect 13136 9664 13142 9676
rect 12115 9608 12296 9636
rect 13740 9636 13768 9676
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15286 9704 15292 9716
rect 15243 9676 15292 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15286 9664 15292 9676
rect 15344 9704 15350 9716
rect 15654 9704 15660 9716
rect 15344 9676 15660 9704
rect 15344 9664 15350 9676
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 18049 9707 18107 9713
rect 16356 9676 16528 9704
rect 16356 9664 16362 9676
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13740 9608 13829 9636
rect 12115 9605 12127 9608
rect 12069 9599 12127 9605
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 15930 9596 15936 9648
rect 15988 9636 15994 9648
rect 16500 9636 16528 9676
rect 18049 9673 18061 9707
rect 18095 9704 18107 9707
rect 18506 9704 18512 9716
rect 18095 9676 18512 9704
rect 18095 9673 18107 9676
rect 18049 9667 18107 9673
rect 18506 9664 18512 9676
rect 18564 9664 18570 9716
rect 19610 9704 19616 9716
rect 19260 9676 19616 9704
rect 16669 9639 16727 9645
rect 16669 9636 16681 9639
rect 15988 9608 16344 9636
rect 16500 9608 16681 9636
rect 15988 9596 15994 9608
rect 16316 9580 16344 9608
rect 16669 9605 16681 9608
rect 16715 9605 16727 9639
rect 16669 9599 16727 9605
rect 18966 9596 18972 9648
rect 19024 9636 19030 9648
rect 19260 9645 19288 9676
rect 19610 9664 19616 9676
rect 19668 9704 19674 9716
rect 20622 9704 20628 9716
rect 19668 9676 20628 9704
rect 19668 9664 19674 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 20898 9704 20904 9716
rect 20859 9676 20904 9704
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 22646 9704 22652 9716
rect 22607 9676 22652 9704
rect 22646 9664 22652 9676
rect 22704 9664 22710 9716
rect 22922 9704 22928 9716
rect 22883 9676 22928 9704
rect 22922 9664 22928 9676
rect 22980 9664 22986 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23716 9676 23857 9704
rect 23716 9664 23722 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 24176 9676 24409 9704
rect 24176 9664 24182 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 24397 9667 24455 9673
rect 19061 9639 19119 9645
rect 19061 9636 19073 9639
rect 19024 9608 19073 9636
rect 19024 9596 19030 9608
rect 19061 9605 19073 9608
rect 19107 9605 19119 9639
rect 19061 9599 19119 9605
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9605 19303 9639
rect 19426 9636 19432 9648
rect 19387 9608 19432 9636
rect 19245 9599 19303 9605
rect 19426 9596 19432 9608
rect 19484 9596 19490 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 21177 9639 21235 9645
rect 19576 9608 20576 9636
rect 19576 9596 19582 9608
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12526 9568 12532 9580
rect 11931 9540 12532 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12676 9540 13001 9568
rect 12676 9528 12682 9540
rect 12989 9537 13001 9540
rect 13035 9568 13047 9571
rect 13449 9571 13507 9577
rect 13449 9568 13461 9571
rect 13035 9540 13461 9568
rect 13035 9537 13047 9540
rect 12989 9531 13047 9537
rect 13449 9537 13461 9540
rect 13495 9568 13507 9571
rect 13722 9568 13728 9580
rect 13495 9540 13728 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14829 9571 14887 9577
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 15841 9571 15899 9577
rect 15841 9568 15853 9571
rect 14875 9540 15853 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 15841 9537 15853 9540
rect 15887 9568 15899 9571
rect 16206 9568 16212 9580
rect 15887 9540 16212 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 16206 9528 16212 9540
rect 16264 9528 16270 9580
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 16390 9528 16396 9580
rect 16448 9568 16454 9580
rect 16448 9540 16493 9568
rect 16448 9528 16454 9540
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 18601 9571 18659 9577
rect 18601 9568 18613 9571
rect 18472 9540 18613 9568
rect 18472 9528 18478 9540
rect 18601 9537 18613 9540
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 19886 9568 19892 9580
rect 19668 9540 19892 9568
rect 19668 9528 19674 9540
rect 19886 9528 19892 9540
rect 19944 9528 19950 9580
rect 20254 9568 20260 9580
rect 20215 9540 20260 9568
rect 20254 9528 20260 9540
rect 20312 9528 20318 9580
rect 20548 9568 20576 9608
rect 21177 9605 21189 9639
rect 21223 9636 21235 9639
rect 21266 9636 21272 9648
rect 21223 9608 21272 9636
rect 21223 9605 21235 9608
rect 21177 9599 21235 9605
rect 21266 9596 21272 9608
rect 21324 9596 21330 9648
rect 24670 9596 24676 9648
rect 24728 9636 24734 9648
rect 24765 9639 24823 9645
rect 24765 9636 24777 9639
rect 24728 9608 24777 9636
rect 24728 9596 24734 9608
rect 24765 9605 24777 9608
rect 24811 9605 24823 9639
rect 24765 9599 24823 9605
rect 25590 9596 25596 9648
rect 25648 9636 25654 9648
rect 25869 9639 25927 9645
rect 25869 9636 25881 9639
rect 25648 9608 25881 9636
rect 25648 9596 25654 9608
rect 25869 9605 25881 9608
rect 25915 9605 25927 9639
rect 26326 9636 26332 9648
rect 26287 9608 26332 9636
rect 25869 9599 25927 9605
rect 26326 9596 26332 9608
rect 26384 9596 26390 9648
rect 20622 9568 20628 9580
rect 20548 9540 20628 9568
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 21634 9568 21640 9580
rect 21595 9540 21640 9568
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9537 21879 9571
rect 22186 9568 22192 9580
rect 22147 9540 22192 9568
rect 21821 9531 21879 9537
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 11348 9472 14013 9500
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 15378 9500 15384 9512
rect 14001 9463 14059 9469
rect 14844 9472 15384 9500
rect 9300 9435 9358 9441
rect 9300 9401 9312 9435
rect 9346 9432 9358 9435
rect 9398 9432 9404 9444
rect 9346 9404 9404 9432
rect 9346 9401 9358 9404
rect 9300 9395 9358 9401
rect 9398 9392 9404 9404
rect 9456 9392 9462 9444
rect 12897 9435 12955 9441
rect 12897 9432 12909 9435
rect 12176 9404 12909 9432
rect 8895 9336 9076 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 10413 9367 10471 9373
rect 10413 9364 10425 9367
rect 9640 9336 10425 9364
rect 9640 9324 9646 9336
rect 10413 9333 10425 9336
rect 10459 9364 10471 9367
rect 11514 9364 11520 9376
rect 10459 9336 11520 9364
rect 10459 9333 10471 9336
rect 10413 9327 10471 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11606 9324 11612 9376
rect 11664 9364 11670 9376
rect 12176 9373 12204 9404
rect 12897 9401 12909 9404
rect 12943 9432 12955 9435
rect 14844 9432 14872 9472
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9500 16911 9503
rect 19981 9503 20039 9509
rect 19981 9500 19993 9503
rect 16899 9472 19993 9500
rect 16899 9469 16911 9472
rect 16853 9463 16911 9469
rect 19981 9469 19993 9472
rect 20027 9500 20039 9503
rect 20070 9500 20076 9512
rect 20027 9472 20076 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 21545 9503 21603 9509
rect 21545 9500 21557 9503
rect 21232 9472 21557 9500
rect 21232 9460 21238 9472
rect 21545 9469 21557 9472
rect 21591 9469 21603 9503
rect 21836 9500 21864 9531
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 25133 9571 25191 9577
rect 25133 9568 25145 9571
rect 24596 9540 25145 9568
rect 21910 9500 21916 9512
rect 21836 9472 21916 9500
rect 21545 9463 21603 9469
rect 21910 9460 21916 9472
rect 21968 9460 21974 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 24596 9509 24624 9540
rect 25133 9537 25145 9540
rect 25179 9537 25191 9571
rect 25133 9531 25191 9537
rect 24581 9503 24639 9509
rect 24581 9500 24593 9503
rect 23440 9472 24593 9500
rect 23440 9460 23446 9472
rect 24581 9469 24593 9472
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 24854 9460 24860 9512
rect 24912 9500 24918 9512
rect 25501 9503 25559 9509
rect 25501 9500 25513 9503
rect 24912 9472 25513 9500
rect 24912 9460 24918 9472
rect 25501 9469 25513 9472
rect 25547 9469 25559 9503
rect 25501 9463 25559 9469
rect 16482 9432 16488 9444
rect 12943 9404 14872 9432
rect 15304 9404 16488 9432
rect 12943 9401 12955 9404
rect 12897 9395 12955 9401
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11664 9336 12081 9364
rect 11664 9324 11670 9336
rect 12069 9333 12081 9336
rect 12115 9364 12127 9367
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 12115 9336 12173 9364
rect 12115 9333 12127 9336
rect 12069 9327 12127 9333
rect 12161 9333 12173 9336
rect 12207 9333 12219 9367
rect 12802 9364 12808 9376
rect 12763 9336 12808 9364
rect 12161 9327 12219 9333
rect 12802 9324 12808 9336
rect 12860 9364 12866 9376
rect 13262 9364 13268 9376
rect 12860 9336 13268 9364
rect 12860 9324 12866 9336
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 15304 9373 15332 9404
rect 16482 9392 16488 9404
rect 16540 9392 16546 9444
rect 17865 9435 17923 9441
rect 17865 9401 17877 9435
rect 17911 9432 17923 9435
rect 17911 9404 18552 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 18524 9376 18552 9404
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 19484 9404 20116 9432
rect 19484 9392 19490 9404
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9333 15347 9367
rect 15654 9364 15660 9376
rect 15615 9336 15660 9364
rect 15289 9327 15347 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 15838 9364 15844 9376
rect 15795 9336 15844 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 17402 9364 17408 9376
rect 17363 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 18414 9364 18420 9376
rect 17460 9336 18420 9364
rect 17460 9324 17466 9336
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 18564 9336 18609 9364
rect 18564 9324 18570 9336
rect 19058 9324 19064 9376
rect 19116 9364 19122 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 19116 9336 19257 9364
rect 19116 9324 19122 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19245 9327 19303 9333
rect 19613 9367 19671 9373
rect 19613 9333 19625 9367
rect 19659 9364 19671 9367
rect 19978 9364 19984 9376
rect 19659 9336 19984 9364
rect 19659 9333 19671 9336
rect 19613 9327 19671 9333
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20088 9373 20116 9404
rect 20073 9367 20131 9373
rect 20073 9333 20085 9367
rect 20119 9333 20131 9367
rect 23290 9364 23296 9376
rect 23251 9336 23296 9364
rect 20073 9327 20131 9333
rect 23290 9324 23296 9336
rect 23348 9324 23354 9376
rect 1104 9274 26864 9296
rect 1104 9222 10315 9274
rect 10367 9222 10379 9274
rect 10431 9222 10443 9274
rect 10495 9222 10507 9274
rect 10559 9222 19648 9274
rect 19700 9222 19712 9274
rect 19764 9222 19776 9274
rect 19828 9222 19840 9274
rect 19892 9222 26864 9274
rect 1104 9200 26864 9222
rect 2222 9160 2228 9172
rect 2183 9132 2228 9160
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2682 9160 2688 9172
rect 2455 9132 2688 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2682 9120 2688 9132
rect 2740 9120 2746 9172
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 4614 9160 4620 9172
rect 4575 9132 4620 9160
rect 4614 9120 4620 9132
rect 4672 9120 4678 9172
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5353 9163 5411 9169
rect 5353 9160 5365 9163
rect 5132 9132 5365 9160
rect 5132 9120 5138 9132
rect 5353 9129 5365 9132
rect 5399 9129 5411 9163
rect 5353 9123 5411 9129
rect 8110 9120 8116 9172
rect 8168 9160 8174 9172
rect 8389 9163 8447 9169
rect 8389 9160 8401 9163
rect 8168 9132 8401 9160
rect 8168 9120 8174 9132
rect 8389 9129 8401 9132
rect 8435 9129 8447 9163
rect 8389 9123 8447 9129
rect 9125 9163 9183 9169
rect 9125 9129 9137 9163
rect 9171 9160 9183 9163
rect 9306 9160 9312 9172
rect 9171 9132 9312 9160
rect 9171 9129 9183 9132
rect 9125 9123 9183 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 10778 9160 10784 9172
rect 10244 9132 10784 9160
rect 10244 9104 10272 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 13170 9120 13176 9172
rect 13228 9160 13234 9172
rect 13633 9163 13691 9169
rect 13633 9160 13645 9163
rect 13228 9132 13645 9160
rect 13228 9120 13234 9132
rect 13633 9129 13645 9132
rect 13679 9129 13691 9163
rect 13633 9123 13691 9129
rect 13998 9120 14004 9172
rect 14056 9160 14062 9172
rect 14553 9163 14611 9169
rect 14553 9160 14565 9163
rect 14056 9132 14565 9160
rect 14056 9120 14062 9132
rect 14553 9129 14565 9132
rect 14599 9129 14611 9163
rect 14553 9123 14611 9129
rect 15105 9163 15163 9169
rect 15105 9129 15117 9163
rect 15151 9160 15163 9163
rect 15286 9160 15292 9172
rect 15151 9132 15292 9160
rect 15151 9129 15163 9132
rect 15105 9123 15163 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 20714 9160 20720 9172
rect 20675 9132 20720 9160
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 21174 9160 21180 9172
rect 20947 9132 21180 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21174 9120 21180 9132
rect 21232 9120 21238 9172
rect 21358 9160 21364 9172
rect 21319 9132 21364 9160
rect 21358 9120 21364 9132
rect 21416 9120 21422 9172
rect 21910 9160 21916 9172
rect 21871 9132 21916 9160
rect 21910 9120 21916 9132
rect 21968 9120 21974 9172
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 22704 9132 23305 9160
rect 22704 9120 22710 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 24394 9160 24400 9172
rect 24355 9132 24400 9160
rect 23293 9123 23351 9129
rect 24394 9120 24400 9132
rect 24452 9120 24458 9172
rect 24762 9160 24768 9172
rect 24723 9132 24768 9160
rect 24762 9120 24768 9132
rect 24820 9120 24826 9172
rect 25866 9160 25872 9172
rect 25827 9132 25872 9160
rect 25866 9120 25872 9132
rect 25924 9120 25930 9172
rect 2590 9052 2596 9104
rect 2648 9092 2654 9104
rect 2777 9095 2835 9101
rect 2777 9092 2789 9095
rect 2648 9064 2789 9092
rect 2648 9052 2654 9064
rect 2777 9061 2789 9064
rect 2823 9092 2835 9095
rect 4798 9092 4804 9104
rect 2823 9064 4804 9092
rect 2823 9061 2835 9064
rect 2777 9055 2835 9061
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 5258 9092 5264 9104
rect 5219 9064 5264 9092
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 8294 9052 8300 9104
rect 8352 9092 8358 9104
rect 9401 9095 9459 9101
rect 9401 9092 9413 9095
rect 8352 9064 9413 9092
rect 8352 9052 8358 9064
rect 9401 9061 9413 9064
rect 9447 9061 9459 9095
rect 9401 9055 9459 9061
rect 10226 9052 10232 9104
rect 10284 9052 10290 9104
rect 10934 9095 10992 9101
rect 10934 9092 10946 9095
rect 10612 9064 10946 9092
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2556 8996 2881 9024
rect 2556 8984 2562 8996
rect 2869 8993 2881 8996
rect 2915 9024 2927 9027
rect 4246 9024 4252 9036
rect 2915 8996 4252 9024
rect 2915 8993 2927 8996
rect 2869 8987 2927 8993
rect 4246 8984 4252 8996
rect 4304 8984 4310 9036
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6546 9024 6552 9036
rect 6503 8996 6552 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6730 9033 6736 9036
rect 6724 9024 6736 9033
rect 6691 8996 6736 9024
rect 6724 8987 6736 8996
rect 6730 8984 6736 8987
rect 6788 8984 6794 9036
rect 10134 8984 10140 9036
rect 10192 9024 10198 9036
rect 10612 9024 10640 9064
rect 10934 9061 10946 9064
rect 10980 9061 10992 9095
rect 13538 9092 13544 9104
rect 13499 9064 13544 9092
rect 10934 9055 10992 9061
rect 13538 9052 13544 9064
rect 13596 9052 13602 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 14185 9095 14243 9101
rect 14185 9092 14197 9095
rect 13872 9064 14197 9092
rect 13872 9052 13878 9064
rect 14185 9061 14197 9064
rect 14231 9061 14243 9095
rect 14185 9055 14243 9061
rect 15470 9052 15476 9104
rect 15528 9101 15534 9104
rect 15528 9095 15592 9101
rect 15528 9061 15546 9095
rect 15580 9061 15592 9095
rect 17954 9092 17960 9104
rect 17867 9064 17960 9092
rect 15528 9055 15592 9061
rect 15528 9052 15534 9055
rect 10192 8996 10640 9024
rect 10689 9027 10747 9033
rect 10192 8984 10198 8996
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 11238 9024 11244 9036
rect 10735 8996 11244 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 11238 8984 11244 8996
rect 11296 8984 11302 9036
rect 14642 8984 14648 9036
rect 14700 9024 14706 9036
rect 17880 9024 17908 9064
rect 17954 9052 17960 9064
rect 18012 9092 18018 9104
rect 18012 9064 20668 9092
rect 18012 9052 18018 9064
rect 18138 9024 18144 9036
rect 14700 8996 17908 9024
rect 18099 8996 18144 9024
rect 14700 8984 14706 8996
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 20070 9024 20076 9036
rect 19751 8996 20076 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20070 8984 20076 8996
rect 20128 8984 20134 9036
rect 20640 9024 20668 9064
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 21269 9095 21327 9101
rect 21269 9092 21281 9095
rect 20864 9064 21281 9092
rect 20864 9052 20870 9064
rect 21269 9061 21281 9064
rect 21315 9092 21327 9095
rect 21542 9092 21548 9104
rect 21315 9064 21548 9092
rect 21315 9061 21327 9064
rect 21269 9055 21327 9061
rect 21542 9052 21548 9064
rect 21600 9052 21606 9104
rect 23842 9092 23848 9104
rect 23584 9064 23848 9092
rect 22002 9024 22008 9036
rect 20640 8996 22008 9024
rect 22002 8984 22008 8996
rect 22060 8984 22066 9036
rect 22465 9027 22523 9033
rect 22465 8993 22477 9027
rect 22511 9024 22523 9027
rect 23014 9024 23020 9036
rect 22511 8996 23020 9024
rect 22511 8993 22523 8996
rect 22465 8987 22523 8993
rect 23014 8984 23020 8996
rect 23072 8984 23078 9036
rect 23584 9033 23612 9064
rect 23842 9052 23848 9064
rect 23900 9092 23906 9104
rect 24029 9095 24087 9101
rect 24029 9092 24041 9095
rect 23900 9064 24041 9092
rect 23900 9052 23906 9064
rect 24029 9061 24041 9064
rect 24075 9061 24087 9095
rect 24029 9055 24087 9061
rect 23569 9027 23627 9033
rect 23569 8993 23581 9027
rect 23615 8993 23627 9027
rect 24118 9024 24124 9036
rect 23569 8987 23627 8993
rect 23768 8996 24124 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 2038 8956 2044 8968
rect 1443 8928 2044 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2958 8956 2964 8968
rect 2919 8928 2964 8956
rect 2958 8916 2964 8928
rect 3016 8956 3022 8968
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 3016 8928 3433 8956
rect 3016 8916 3022 8928
rect 3421 8925 3433 8928
rect 3467 8956 3479 8959
rect 3510 8956 3516 8968
rect 3467 8928 3516 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3510 8916 3516 8928
rect 3568 8916 3574 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 9674 8956 9680 8968
rect 5583 8928 6040 8956
rect 9635 8928 9680 8956
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 1670 8848 1676 8900
rect 1728 8888 1734 8900
rect 5902 8888 5908 8900
rect 1728 8860 5908 8888
rect 1728 8848 1734 8860
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6012 8897 6040 8928
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 12621 8959 12679 8965
rect 12621 8956 12633 8959
rect 12492 8928 12633 8956
rect 12492 8916 12498 8928
rect 12621 8925 12633 8928
rect 12667 8956 12679 8959
rect 12802 8956 12808 8968
rect 12667 8928 12808 8956
rect 12667 8925 12679 8928
rect 12621 8919 12679 8925
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 13722 8956 13728 8968
rect 13683 8928 13728 8956
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 15289 8959 15347 8965
rect 15289 8925 15301 8959
rect 15335 8925 15347 8959
rect 15289 8919 15347 8925
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8956 17371 8959
rect 17770 8956 17776 8968
rect 17359 8928 17776 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 5997 8891 6055 8897
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 6043 8860 6500 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1820 8792 1869 8820
rect 1820 8780 1826 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 3878 8820 3884 8832
rect 3839 8792 3884 8820
rect 1857 8783 1915 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4893 8823 4951 8829
rect 4893 8789 4905 8823
rect 4939 8820 4951 8823
rect 5258 8820 5264 8832
rect 4939 8792 5264 8820
rect 4939 8789 4951 8792
rect 4893 8783 4951 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 6270 8820 6276 8832
rect 6231 8792 6276 8820
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6472 8820 6500 8860
rect 12342 8848 12348 8900
rect 12400 8888 12406 8900
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12400 8860 13185 8888
rect 12400 8848 12406 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 7742 8820 7748 8832
rect 6472 8792 7748 8820
rect 7742 8780 7748 8792
rect 7800 8820 7806 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7800 8792 7849 8820
rect 7800 8780 7806 8792
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 10321 8823 10379 8829
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 10870 8820 10876 8832
rect 10367 8792 10876 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 12066 8820 12072 8832
rect 12027 8792 12072 8820
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 13081 8823 13139 8829
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13722 8820 13728 8832
rect 13127 8792 13728 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13722 8780 13728 8792
rect 13780 8780 13786 8832
rect 15304 8820 15332 8919
rect 17770 8916 17776 8928
rect 17828 8956 17834 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 17828 8928 18245 8956
rect 17828 8916 17834 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18380 8928 19441 8956
rect 18380 8916 18386 8928
rect 19429 8925 19441 8928
rect 19475 8956 19487 8959
rect 20254 8956 20260 8968
rect 19475 8928 20260 8956
rect 19475 8925 19487 8928
rect 19429 8919 19487 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 21453 8959 21511 8965
rect 21453 8925 21465 8959
rect 21499 8925 21511 8959
rect 22922 8956 22928 8968
rect 22883 8928 22928 8956
rect 21453 8919 21511 8925
rect 17681 8891 17739 8897
rect 17681 8857 17693 8891
rect 17727 8888 17739 8891
rect 18340 8888 18368 8916
rect 17727 8860 18368 8888
rect 17727 8857 17739 8860
rect 17681 8851 17739 8857
rect 19242 8848 19248 8900
rect 19300 8888 19306 8900
rect 21468 8888 21496 8919
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 21542 8888 21548 8900
rect 19300 8860 21548 8888
rect 19300 8848 19306 8860
rect 21542 8848 21548 8860
rect 21600 8848 21606 8900
rect 22649 8891 22707 8897
rect 22649 8857 22661 8891
rect 22695 8888 22707 8891
rect 23382 8888 23388 8900
rect 22695 8860 23388 8888
rect 22695 8857 22707 8860
rect 22649 8851 22707 8857
rect 23382 8848 23388 8860
rect 23440 8848 23446 8900
rect 23768 8897 23796 8996
rect 24118 8984 24124 8996
rect 24176 9024 24182 9036
rect 24581 9027 24639 9033
rect 24581 9024 24593 9027
rect 24176 8996 24593 9024
rect 24176 8984 24182 8996
rect 24581 8993 24593 8996
rect 24627 8993 24639 9027
rect 24581 8987 24639 8993
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 25133 9027 25191 9033
rect 25133 9024 25145 9027
rect 24912 8996 25145 9024
rect 24912 8984 24918 8996
rect 25133 8993 25145 8996
rect 25179 8993 25191 9027
rect 25133 8987 25191 8993
rect 25958 8916 25964 8968
rect 26016 8956 26022 8968
rect 26142 8956 26148 8968
rect 26016 8928 26148 8956
rect 26016 8916 26022 8928
rect 26142 8916 26148 8928
rect 26200 8916 26206 8968
rect 23753 8891 23811 8897
rect 23753 8857 23765 8891
rect 23799 8857 23811 8891
rect 23753 8851 23811 8857
rect 15562 8820 15568 8832
rect 15304 8792 15568 8820
rect 15562 8780 15568 8792
rect 15620 8780 15626 8832
rect 16669 8823 16727 8829
rect 16669 8789 16681 8823
rect 16715 8820 16727 8823
rect 16758 8820 16764 8832
rect 16715 8792 16764 8820
rect 16715 8789 16727 8792
rect 16669 8783 16727 8789
rect 16758 8780 16764 8792
rect 16816 8780 16822 8832
rect 17773 8823 17831 8829
rect 17773 8789 17785 8823
rect 17819 8820 17831 8823
rect 17862 8820 17868 8832
rect 17819 8792 17868 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 17862 8780 17868 8792
rect 17920 8780 17926 8832
rect 19058 8820 19064 8832
rect 19019 8792 19064 8820
rect 19058 8780 19064 8792
rect 19116 8780 19122 8832
rect 19886 8820 19892 8832
rect 19847 8792 19892 8820
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 22186 8780 22192 8832
rect 22244 8820 22250 8832
rect 22281 8823 22339 8829
rect 22281 8820 22293 8823
rect 22244 8792 22293 8820
rect 22244 8780 22250 8792
rect 22281 8789 22293 8792
rect 22327 8789 22339 8823
rect 25590 8820 25596 8832
rect 25551 8792 25596 8820
rect 22281 8783 22339 8789
rect 25590 8780 25596 8792
rect 25648 8780 25654 8832
rect 26142 8780 26148 8832
rect 26200 8820 26206 8832
rect 26237 8823 26295 8829
rect 26237 8820 26249 8823
rect 26200 8792 26249 8820
rect 26200 8780 26206 8792
rect 26237 8789 26249 8792
rect 26283 8789 26295 8823
rect 26237 8783 26295 8789
rect 1104 8730 26864 8752
rect 1104 8678 5648 8730
rect 5700 8678 5712 8730
rect 5764 8678 5776 8730
rect 5828 8678 5840 8730
rect 5892 8678 14982 8730
rect 15034 8678 15046 8730
rect 15098 8678 15110 8730
rect 15162 8678 15174 8730
rect 15226 8678 24315 8730
rect 24367 8678 24379 8730
rect 24431 8678 24443 8730
rect 24495 8678 24507 8730
rect 24559 8678 26864 8730
rect 1104 8656 26864 8678
rect 1486 8576 1492 8628
rect 1544 8616 1550 8628
rect 1581 8619 1639 8625
rect 1581 8616 1593 8619
rect 1544 8588 1593 8616
rect 1544 8576 1550 8588
rect 1581 8585 1593 8588
rect 1627 8585 1639 8619
rect 1581 8579 1639 8585
rect 2869 8619 2927 8625
rect 2869 8585 2881 8619
rect 2915 8616 2927 8619
rect 3234 8616 3240 8628
rect 2915 8588 3240 8616
rect 2915 8585 2927 8588
rect 2869 8579 2927 8585
rect 3234 8576 3240 8588
rect 3292 8616 3298 8628
rect 3418 8616 3424 8628
rect 3292 8588 3424 8616
rect 3292 8576 3298 8588
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4249 8619 4307 8625
rect 4249 8616 4261 8619
rect 4212 8588 4261 8616
rect 4212 8576 4218 8588
rect 4249 8585 4261 8588
rect 4295 8616 4307 8619
rect 7190 8616 7196 8628
rect 4295 8588 4651 8616
rect 7151 8588 7196 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 566 8508 572 8560
rect 624 8548 630 8560
rect 2501 8551 2559 8557
rect 2501 8548 2513 8551
rect 624 8520 2513 8548
rect 624 8508 630 8520
rect 2501 8517 2513 8520
rect 2547 8548 2559 8551
rect 2590 8548 2596 8560
rect 2547 8520 2596 8548
rect 2547 8517 2559 8520
rect 2501 8511 2559 8517
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 4522 8548 4528 8560
rect 4479 8520 4528 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 4522 8508 4528 8520
rect 4580 8508 4586 8560
rect 3326 8480 3332 8492
rect 3287 8452 3332 8480
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3510 8480 3516 8492
rect 3471 8452 3516 8480
rect 3510 8440 3516 8452
rect 3568 8440 3574 8492
rect 1394 8412 1400 8424
rect 1355 8384 1400 8412
rect 1394 8372 1400 8384
rect 1452 8372 1458 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 4623 8412 4651 8588
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9306 8616 9312 8628
rect 9079 8588 9312 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9677 8619 9735 8625
rect 9677 8585 9689 8619
rect 9723 8616 9735 8619
rect 9950 8616 9956 8628
rect 9723 8588 9956 8616
rect 9723 8585 9735 8588
rect 9677 8579 9735 8585
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10226 8616 10232 8628
rect 10187 8588 10232 8616
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 11238 8616 11244 8628
rect 11199 8588 11244 8616
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11572 8588 12173 8616
rect 11572 8576 11578 8588
rect 12161 8585 12173 8588
rect 12207 8616 12219 8619
rect 12618 8616 12624 8628
rect 12207 8588 12624 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12805 8619 12863 8625
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 13170 8616 13176 8628
rect 12851 8588 13176 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13538 8616 13544 8628
rect 13280 8588 13544 8616
rect 13081 8551 13139 8557
rect 13081 8517 13093 8551
rect 13127 8548 13139 8551
rect 13280 8548 13308 8588
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14516 8588 14657 8616
rect 14516 8576 14522 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 15746 8616 15752 8628
rect 15707 8588 15752 8616
rect 15746 8576 15752 8588
rect 15804 8576 15810 8628
rect 15838 8576 15844 8628
rect 15896 8616 15902 8628
rect 16390 8616 16396 8628
rect 15896 8588 16396 8616
rect 15896 8576 15902 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 20070 8616 20076 8628
rect 20031 8588 20076 8616
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 20312 8588 20545 8616
rect 20312 8576 20318 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 21542 8616 21548 8628
rect 21503 8588 21548 8616
rect 20533 8579 20591 8585
rect 21542 8576 21548 8588
rect 21600 8576 21606 8628
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24489 8619 24547 8625
rect 24489 8616 24501 8619
rect 24176 8588 24501 8616
rect 24176 8576 24182 8588
rect 24489 8585 24501 8588
rect 24535 8585 24547 8619
rect 25498 8616 25504 8628
rect 25459 8588 25504 8616
rect 24489 8579 24547 8585
rect 25498 8576 25504 8588
rect 25556 8576 25562 8628
rect 25961 8619 26019 8625
rect 25961 8585 25973 8619
rect 26007 8616 26019 8619
rect 26050 8616 26056 8628
rect 26007 8588 26056 8616
rect 26007 8585 26019 8588
rect 25961 8579 26019 8585
rect 26050 8576 26056 8588
rect 26108 8576 26114 8628
rect 26326 8616 26332 8628
rect 26287 8588 26332 8616
rect 26326 8576 26332 8588
rect 26384 8576 26390 8628
rect 13127 8520 13308 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4985 8483 5043 8489
rect 4985 8480 4997 8483
rect 4764 8452 4997 8480
rect 4764 8440 4770 8452
rect 4985 8449 4997 8452
rect 5031 8480 5043 8483
rect 5445 8483 5503 8489
rect 5445 8480 5457 8483
rect 5031 8452 5457 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 5445 8449 5457 8452
rect 5491 8449 5503 8483
rect 6546 8480 6552 8492
rect 5445 8443 5503 8449
rect 6472 8452 6552 8480
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 2096 8384 3280 8412
rect 4623 8384 4813 8412
rect 2096 8372 2102 8384
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 3142 8344 3148 8356
rect 2179 8316 3148 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 3252 8288 3280 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 4948 8384 4993 8412
rect 4948 8372 4954 8384
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 6472 8421 6500 8452
rect 6546 8440 6552 8452
rect 6604 8480 6610 8492
rect 7469 8483 7527 8489
rect 7469 8480 7481 8483
rect 6604 8452 7481 8480
rect 6604 8440 6610 8452
rect 7469 8449 7481 8452
rect 7515 8480 7527 8483
rect 7650 8480 7656 8492
rect 7515 8452 7656 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7650 8440 7656 8452
rect 7708 8440 7714 8492
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 9950 8480 9956 8492
rect 9824 8452 9956 8480
rect 9824 8440 9830 8452
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10778 8480 10784 8492
rect 10739 8452 10784 8480
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 15304 8480 15332 8576
rect 15562 8508 15568 8560
rect 15620 8548 15626 8560
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 15620 8520 16773 8548
rect 15620 8508 15626 8520
rect 16761 8517 16773 8520
rect 16807 8548 16819 8551
rect 17773 8551 17831 8557
rect 17773 8548 17785 8551
rect 16807 8520 17785 8548
rect 16807 8517 16819 8520
rect 16761 8511 16819 8517
rect 17773 8517 17785 8520
rect 17819 8517 17831 8551
rect 17773 8511 17831 8517
rect 16301 8483 16359 8489
rect 16301 8480 16313 8483
rect 15304 8452 16313 8480
rect 16301 8449 16313 8452
rect 16347 8449 16359 8483
rect 17788 8480 17816 8511
rect 19334 8508 19340 8560
rect 19392 8548 19398 8560
rect 19429 8551 19487 8557
rect 19429 8548 19441 8551
rect 19392 8520 19441 8548
rect 19392 8508 19398 8520
rect 19429 8517 19441 8520
rect 19475 8548 19487 8551
rect 20349 8551 20407 8557
rect 20349 8548 20361 8551
rect 19475 8520 20361 8548
rect 19475 8517 19487 8520
rect 19429 8511 19487 8517
rect 20349 8517 20361 8520
rect 20395 8548 20407 8551
rect 22281 8551 22339 8557
rect 20395 8520 21128 8548
rect 20395 8517 20407 8520
rect 20349 8511 20407 8517
rect 18049 8483 18107 8489
rect 18049 8480 18061 8483
rect 17788 8452 18061 8480
rect 16301 8443 16359 8449
rect 18049 8449 18061 8452
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 21100 8489 21128 8520
rect 22281 8517 22293 8551
rect 22327 8548 22339 8551
rect 22646 8548 22652 8560
rect 22327 8520 22652 8548
rect 22327 8517 22339 8520
rect 22281 8511 22339 8517
rect 22646 8508 22652 8520
rect 22704 8508 22710 8560
rect 24854 8548 24860 8560
rect 24815 8520 24860 8548
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 20993 8483 21051 8489
rect 20993 8480 21005 8483
rect 20772 8452 21005 8480
rect 20772 8440 20778 8452
rect 20993 8449 21005 8452
rect 21039 8449 21051 8483
rect 20993 8443 21051 8449
rect 21085 8483 21143 8489
rect 21085 8449 21097 8483
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 23566 8480 23572 8492
rect 23523 8452 23572 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 5408 8384 6469 8412
rect 5408 8372 5414 8384
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10962 8412 10968 8424
rect 10643 8384 10968 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8412 13323 8415
rect 16114 8412 16120 8424
rect 13311 8384 13492 8412
rect 13311 8381 13323 8384
rect 13265 8375 13323 8381
rect 3973 8347 4031 8353
rect 3973 8313 3985 8347
rect 4019 8344 4031 8347
rect 4246 8344 4252 8356
rect 4019 8316 4252 8344
rect 4019 8313 4031 8316
rect 3973 8307 4031 8313
rect 4246 8304 4252 8316
rect 4304 8344 4310 8356
rect 5442 8344 5448 8356
rect 4304 8316 5448 8344
rect 4304 8304 4310 8316
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 6730 8344 6736 8356
rect 6288 8316 6736 8344
rect 6288 8288 6316 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 7898 8347 7956 8353
rect 7898 8344 7910 8347
rect 7800 8316 7910 8344
rect 7800 8304 7806 8316
rect 7898 8313 7910 8316
rect 7944 8313 7956 8347
rect 7898 8307 7956 8313
rect 9766 8304 9772 8356
rect 9824 8344 9830 8356
rect 10689 8347 10747 8353
rect 10689 8344 10701 8347
rect 9824 8316 10701 8344
rect 9824 8304 9830 8316
rect 10689 8313 10701 8316
rect 10735 8344 10747 8347
rect 11609 8347 11667 8353
rect 11609 8344 11621 8347
rect 10735 8316 11621 8344
rect 10735 8313 10747 8316
rect 10689 8307 10747 8313
rect 11609 8313 11621 8316
rect 11655 8313 11667 8347
rect 11609 8307 11667 8313
rect 13464 8288 13492 8384
rect 15212 8384 16120 8412
rect 13532 8347 13590 8353
rect 13532 8313 13544 8347
rect 13578 8344 13590 8347
rect 13722 8344 13728 8356
rect 13578 8316 13728 8344
rect 13578 8313 13590 8316
rect 13532 8307 13590 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 15212 8353 15240 8384
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20901 8415 20959 8421
rect 20901 8412 20913 8415
rect 20036 8384 20913 8412
rect 20036 8372 20042 8384
rect 20901 8381 20913 8384
rect 20947 8412 20959 8415
rect 21913 8415 21971 8421
rect 21913 8412 21925 8415
rect 20947 8384 21925 8412
rect 20947 8381 20959 8384
rect 20901 8375 20959 8381
rect 21913 8381 21925 8384
rect 21959 8381 21971 8415
rect 21913 8375 21971 8381
rect 22097 8415 22155 8421
rect 22097 8381 22109 8415
rect 22143 8412 22155 8415
rect 22649 8415 22707 8421
rect 22649 8412 22661 8415
rect 22143 8384 22661 8412
rect 22143 8381 22155 8384
rect 22097 8375 22155 8381
rect 22649 8381 22661 8384
rect 22695 8381 22707 8415
rect 23014 8412 23020 8424
rect 22975 8384 23020 8412
rect 22649 8375 22707 8381
rect 15197 8347 15255 8353
rect 15197 8344 15209 8347
rect 15028 8316 15209 8344
rect 3234 8276 3240 8288
rect 3195 8248 3240 8276
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 6181 8279 6239 8285
rect 6181 8245 6193 8279
rect 6227 8276 6239 8279
rect 6270 8276 6276 8288
rect 6227 8248 6276 8276
rect 6227 8245 6239 8248
rect 6181 8239 6239 8245
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 10134 8276 10140 8288
rect 10095 8248 10140 8276
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 10778 8236 10784 8288
rect 10836 8276 10842 8288
rect 11146 8276 11152 8288
rect 10836 8248 11152 8276
rect 10836 8236 10842 8248
rect 11146 8236 11152 8248
rect 11204 8236 11210 8288
rect 13446 8236 13452 8288
rect 13504 8236 13510 8288
rect 13630 8236 13636 8288
rect 13688 8276 13694 8288
rect 15028 8276 15056 8316
rect 15197 8313 15209 8316
rect 15243 8313 15255 8347
rect 15562 8344 15568 8356
rect 15523 8316 15568 8344
rect 15197 8307 15255 8313
rect 15562 8304 15568 8316
rect 15620 8344 15626 8356
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 15620 8316 16221 8344
rect 15620 8304 15626 8316
rect 16209 8313 16221 8316
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 16666 8304 16672 8356
rect 16724 8344 16730 8356
rect 18322 8353 18328 8356
rect 17497 8347 17555 8353
rect 17497 8344 17509 8347
rect 16724 8316 17509 8344
rect 16724 8304 16730 8316
rect 17497 8313 17509 8316
rect 17543 8344 17555 8347
rect 18316 8344 18328 8353
rect 17543 8316 18328 8344
rect 17543 8313 17555 8316
rect 17497 8307 17555 8313
rect 18316 8307 18328 8316
rect 18322 8304 18328 8307
rect 18380 8304 18386 8356
rect 21726 8344 21732 8356
rect 20732 8316 21732 8344
rect 20732 8288 20760 8316
rect 21726 8304 21732 8316
rect 21784 8344 21790 8356
rect 22112 8344 22140 8375
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 23658 8412 23664 8424
rect 23619 8384 23664 8412
rect 23658 8372 23664 8384
rect 23716 8412 23722 8424
rect 24121 8415 24179 8421
rect 24121 8412 24133 8415
rect 23716 8384 24133 8412
rect 23716 8372 23722 8384
rect 24121 8381 24133 8384
rect 24167 8381 24179 8415
rect 24121 8375 24179 8381
rect 24673 8415 24731 8421
rect 24673 8381 24685 8415
rect 24719 8381 24731 8415
rect 24673 8375 24731 8381
rect 23198 8344 23204 8356
rect 21784 8316 22140 8344
rect 22204 8316 23204 8344
rect 21784 8304 21790 8316
rect 13688 8248 15056 8276
rect 13688 8236 13694 8248
rect 18598 8236 18604 8288
rect 18656 8276 18662 8288
rect 19150 8276 19156 8288
rect 18656 8248 19156 8276
rect 18656 8236 18662 8248
rect 19150 8236 19156 8248
rect 19208 8236 19214 8288
rect 20714 8236 20720 8288
rect 20772 8236 20778 8288
rect 21818 8236 21824 8288
rect 21876 8276 21882 8288
rect 22204 8276 22232 8316
rect 23198 8304 23204 8316
rect 23256 8304 23262 8356
rect 23474 8304 23480 8356
rect 23532 8344 23538 8356
rect 24688 8344 24716 8375
rect 25133 8347 25191 8353
rect 25133 8344 25145 8347
rect 23532 8316 25145 8344
rect 23532 8304 23538 8316
rect 25133 8313 25145 8316
rect 25179 8313 25191 8347
rect 25133 8307 25191 8313
rect 23842 8276 23848 8288
rect 21876 8248 22232 8276
rect 23803 8248 23848 8276
rect 21876 8236 21882 8248
rect 23842 8236 23848 8248
rect 23900 8236 23906 8288
rect 1104 8186 26864 8208
rect 1104 8134 10315 8186
rect 10367 8134 10379 8186
rect 10431 8134 10443 8186
rect 10495 8134 10507 8186
rect 10559 8134 19648 8186
rect 19700 8134 19712 8186
rect 19764 8134 19776 8186
rect 19828 8134 19840 8186
rect 19892 8134 26864 8186
rect 1104 8112 26864 8134
rect 1946 8032 1952 8084
rect 2004 8072 2010 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 2004 8044 2237 8072
rect 2004 8032 2010 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2406 8072 2412 8084
rect 2367 8044 2412 8072
rect 2225 8035 2283 8041
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 2832 8044 2877 8072
rect 2832 8032 2838 8044
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3292 8044 3433 8072
rect 3292 8032 3298 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 4249 8075 4307 8081
rect 4249 8072 4261 8075
rect 3844 8044 4261 8072
rect 3844 8032 3850 8044
rect 4249 8041 4261 8044
rect 4295 8041 4307 8075
rect 4249 8035 4307 8041
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 4890 8072 4896 8084
rect 4755 8044 4896 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7558 8072 7564 8084
rect 7248 8044 7564 8072
rect 7248 8032 7254 8044
rect 7558 8032 7564 8044
rect 7616 8032 7622 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9582 8072 9588 8084
rect 9539 8044 9588 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9766 8072 9772 8084
rect 9727 8044 9772 8072
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10008 8044 10149 8072
rect 10008 8032 10014 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10229 8075 10287 8081
rect 10229 8041 10241 8075
rect 10275 8072 10287 8075
rect 10686 8072 10692 8084
rect 10275 8044 10692 8072
rect 10275 8041 10287 8044
rect 10229 8035 10287 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11112 8044 11621 8072
rect 11112 8032 11118 8044
rect 11609 8041 11621 8044
rect 11655 8072 11667 8075
rect 12342 8072 12348 8084
rect 11655 8044 12348 8072
rect 11655 8041 11667 8044
rect 11609 8035 11667 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13817 8075 13875 8081
rect 13817 8072 13829 8075
rect 13504 8044 13829 8072
rect 13504 8032 13510 8044
rect 13817 8041 13829 8044
rect 13863 8041 13875 8075
rect 13817 8035 13875 8041
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13964 8044 14197 8072
rect 13964 8032 13970 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 15102 8072 15108 8084
rect 15063 8044 15108 8072
rect 14185 8035 14243 8041
rect 15102 8032 15108 8044
rect 15160 8032 15166 8084
rect 15562 8032 15568 8084
rect 15620 8072 15626 8084
rect 16206 8072 16212 8084
rect 15620 8044 16212 8072
rect 15620 8032 15626 8044
rect 16206 8032 16212 8044
rect 16264 8032 16270 8084
rect 16666 8072 16672 8084
rect 16627 8044 16672 8072
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 17770 8072 17776 8084
rect 17731 8044 17776 8072
rect 17770 8032 17776 8044
rect 17828 8032 17834 8084
rect 18138 8032 18144 8084
rect 18196 8072 18202 8084
rect 19153 8075 19211 8081
rect 19153 8072 19165 8075
rect 18196 8044 19165 8072
rect 18196 8032 18202 8044
rect 19153 8041 19165 8044
rect 19199 8041 19211 8075
rect 19153 8035 19211 8041
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 20257 8075 20315 8081
rect 20257 8072 20269 8075
rect 19484 8044 20269 8072
rect 19484 8032 19490 8044
rect 20257 8041 20269 8044
rect 20303 8041 20315 8075
rect 20257 8035 20315 8041
rect 22554 8032 22560 8084
rect 22612 8072 22618 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22612 8044 22937 8072
rect 22612 8032 22618 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 2869 8007 2927 8013
rect 2869 7973 2881 8007
rect 2915 8004 2927 8007
rect 2958 8004 2964 8016
rect 2915 7976 2964 8004
rect 2915 7973 2927 7976
rect 2869 7967 2927 7973
rect 2958 7964 2964 7976
rect 3016 7964 3022 8016
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 4985 8007 5043 8013
rect 4985 8004 4997 8007
rect 3568 7976 4997 8004
rect 3568 7964 3574 7976
rect 4724 7948 4752 7976
rect 4985 7973 4997 7976
rect 5031 7973 5043 8007
rect 4985 7967 5043 7973
rect 5528 8007 5586 8013
rect 5528 7973 5540 8007
rect 5574 8004 5586 8007
rect 6362 8004 6368 8016
rect 5574 7976 6368 8004
rect 5574 7973 5586 7976
rect 5528 7967 5586 7973
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 7742 8004 7748 8016
rect 7703 7976 7748 8004
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 4062 7936 4068 7948
rect 4023 7908 4068 7936
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 4706 7896 4712 7948
rect 4764 7896 4770 7948
rect 5261 7939 5319 7945
rect 5261 7905 5273 7939
rect 5307 7936 5319 7939
rect 5350 7936 5356 7948
rect 5307 7908 5356 7936
rect 5307 7905 5319 7908
rect 5261 7899 5319 7905
rect 5350 7896 5356 7908
rect 5408 7896 5414 7948
rect 8389 7939 8447 7945
rect 8389 7905 8401 7939
rect 8435 7936 8447 7939
rect 8662 7936 8668 7948
rect 8435 7908 8668 7936
rect 8435 7905 8447 7908
rect 8389 7899 8447 7905
rect 8662 7896 8668 7908
rect 8720 7896 8726 7948
rect 1394 7868 1400 7880
rect 1355 7840 1400 7868
rect 1394 7828 1400 7840
rect 1452 7828 1458 7880
rect 2961 7871 3019 7877
rect 2961 7837 2973 7871
rect 3007 7868 3019 7871
rect 3970 7868 3976 7880
rect 3007 7840 3976 7868
rect 3007 7837 3019 7840
rect 2961 7831 3019 7837
rect 2590 7760 2596 7812
rect 2648 7800 2654 7812
rect 2976 7800 3004 7831
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 7466 7828 7472 7880
rect 7524 7868 7530 7880
rect 8481 7871 8539 7877
rect 8481 7868 8493 7871
rect 7524 7840 8493 7868
rect 7524 7828 7530 7840
rect 8404 7812 8432 7840
rect 8481 7837 8493 7840
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9600 7868 9628 8032
rect 9674 7964 9680 8016
rect 9732 8004 9738 8016
rect 10781 8007 10839 8013
rect 10781 8004 10793 8007
rect 9732 7976 10793 8004
rect 9732 7964 9738 7976
rect 10781 7973 10793 7976
rect 10827 8004 10839 8007
rect 11146 8004 11152 8016
rect 10827 7976 11152 8004
rect 10827 7973 10839 7976
rect 10781 7967 10839 7973
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 12066 7964 12072 8016
rect 12124 8013 12130 8016
rect 12124 8007 12188 8013
rect 12124 7973 12142 8007
rect 12176 7973 12188 8007
rect 15654 8004 15660 8016
rect 12124 7967 12188 7973
rect 15304 7976 15660 8004
rect 12124 7964 12130 7967
rect 11238 7896 11244 7948
rect 11296 7936 11302 7948
rect 11882 7936 11888 7948
rect 11296 7908 11888 7936
rect 11296 7896 11302 7908
rect 11882 7896 11888 7908
rect 11940 7896 11946 7948
rect 15304 7945 15332 7976
rect 15654 7964 15660 7976
rect 15712 7964 15718 8016
rect 18690 7964 18696 8016
rect 18748 8004 18754 8016
rect 18966 8004 18972 8016
rect 18748 7976 18972 8004
rect 18748 7964 18754 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 20346 8004 20352 8016
rect 19352 7976 20352 8004
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 15556 7939 15614 7945
rect 15556 7905 15568 7939
rect 15602 7936 15614 7939
rect 16114 7936 16120 7948
rect 15602 7908 16120 7936
rect 15602 7905 15614 7908
rect 15556 7899 15614 7905
rect 16114 7896 16120 7908
rect 16172 7936 16178 7948
rect 17589 7939 17647 7945
rect 17589 7936 17601 7939
rect 16172 7908 17601 7936
rect 16172 7896 16178 7908
rect 17589 7905 17601 7908
rect 17635 7905 17647 7939
rect 17589 7899 17647 7905
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 8628 7840 8673 7868
rect 9600 7840 10333 7868
rect 8628 7828 8634 7840
rect 10321 7837 10333 7840
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 2648 7772 3004 7800
rect 7377 7803 7435 7809
rect 2648 7760 2654 7772
rect 7377 7769 7389 7803
rect 7423 7800 7435 7803
rect 8110 7800 8116 7812
rect 7423 7772 8116 7800
rect 7423 7769 7435 7772
rect 7377 7763 7435 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8386 7760 8392 7812
rect 8444 7760 8450 7812
rect 9125 7803 9183 7809
rect 9125 7769 9137 7803
rect 9171 7800 9183 7803
rect 9582 7800 9588 7812
rect 9171 7772 9588 7800
rect 9171 7769 9183 7772
rect 9125 7763 9183 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 14182 7760 14188 7812
rect 14240 7800 14246 7812
rect 14366 7800 14372 7812
rect 14240 7772 14372 7800
rect 14240 7760 14246 7772
rect 14366 7760 14372 7772
rect 14424 7760 14430 7812
rect 17604 7800 17632 7899
rect 17678 7896 17684 7948
rect 17736 7936 17742 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17736 7908 18153 7936
rect 17736 7896 17742 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 18233 7939 18291 7945
rect 18233 7905 18245 7939
rect 18279 7936 18291 7939
rect 18598 7936 18604 7948
rect 18279 7908 18604 7936
rect 18279 7905 18291 7908
rect 18233 7899 18291 7905
rect 18598 7896 18604 7908
rect 18656 7936 18662 7948
rect 19352 7945 19380 7976
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 22462 8004 22468 8016
rect 20824 7976 22468 8004
rect 19337 7939 19395 7945
rect 18656 7908 19288 7936
rect 18656 7896 18662 7908
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 19260 7868 19288 7908
rect 19337 7905 19349 7939
rect 19383 7936 19395 7939
rect 19518 7936 19524 7948
rect 19383 7908 19524 7936
rect 19383 7905 19395 7908
rect 19337 7899 19395 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 19886 7936 19892 7948
rect 19847 7908 19892 7936
rect 19886 7896 19892 7908
rect 19944 7896 19950 7948
rect 19978 7896 19984 7948
rect 20036 7936 20042 7948
rect 20438 7936 20444 7948
rect 20036 7908 20444 7936
rect 20036 7896 20042 7908
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 20714 7868 20720 7880
rect 19260 7840 20720 7868
rect 18325 7831 18383 7837
rect 18340 7800 18368 7831
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 18690 7800 18696 7812
rect 17604 7772 18696 7800
rect 18690 7760 18696 7772
rect 18748 7800 18754 7812
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 18748 7772 18797 7800
rect 18748 7760 18754 7772
rect 18785 7769 18797 7772
rect 18831 7769 18843 7803
rect 18785 7763 18843 7769
rect 20070 7760 20076 7812
rect 20128 7800 20134 7812
rect 20824 7800 20852 7976
rect 22462 7964 22468 7976
rect 22520 7964 22526 8016
rect 21174 7896 21180 7948
rect 21232 7936 21238 7948
rect 21269 7939 21327 7945
rect 21269 7936 21281 7939
rect 21232 7908 21281 7936
rect 21232 7896 21238 7908
rect 21269 7905 21281 7908
rect 21315 7905 21327 7939
rect 21269 7899 21327 7905
rect 22189 7939 22247 7945
rect 22189 7905 22201 7939
rect 22235 7936 22247 7939
rect 22370 7936 22376 7948
rect 22235 7908 22376 7936
rect 22235 7905 22247 7908
rect 22189 7899 22247 7905
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 22738 7896 22744 7948
rect 22796 7936 22802 7948
rect 22833 7939 22891 7945
rect 22833 7936 22845 7939
rect 22796 7908 22845 7936
rect 22796 7896 22802 7908
rect 22833 7905 22845 7908
rect 22879 7905 22891 7939
rect 22833 7899 22891 7905
rect 23290 7896 23296 7948
rect 23348 7936 23354 7948
rect 24029 7939 24087 7945
rect 24029 7936 24041 7939
rect 23348 7908 24041 7936
rect 23348 7896 23354 7908
rect 24029 7905 24041 7908
rect 24075 7936 24087 7939
rect 24762 7936 24768 7948
rect 24075 7908 24768 7936
rect 24075 7905 24087 7908
rect 24029 7899 24087 7905
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 25038 7896 25044 7948
rect 25096 7936 25102 7948
rect 25133 7939 25191 7945
rect 25133 7936 25145 7939
rect 25096 7908 25145 7936
rect 25096 7896 25102 7908
rect 25133 7905 25145 7908
rect 25179 7905 25191 7939
rect 25133 7899 25191 7905
rect 21082 7828 21088 7880
rect 21140 7868 21146 7880
rect 21358 7868 21364 7880
rect 21140 7840 21364 7868
rect 21140 7828 21146 7840
rect 21358 7828 21364 7840
rect 21416 7828 21422 7880
rect 21542 7868 21548 7880
rect 21503 7840 21548 7868
rect 21542 7828 21548 7840
rect 21600 7868 21606 7880
rect 23014 7868 23020 7880
rect 21600 7840 23020 7868
rect 21600 7828 21606 7840
rect 23014 7828 23020 7840
rect 23072 7828 23078 7880
rect 20128 7772 20852 7800
rect 20901 7803 20959 7809
rect 20128 7760 20134 7772
rect 20901 7769 20913 7803
rect 20947 7800 20959 7803
rect 22189 7803 22247 7809
rect 22189 7800 22201 7803
rect 20947 7772 22201 7800
rect 20947 7769 20959 7772
rect 20901 7763 20959 7769
rect 22189 7769 22201 7772
rect 22235 7769 22247 7803
rect 22189 7763 22247 7769
rect 22830 7760 22836 7812
rect 22888 7800 22894 7812
rect 23308 7800 23336 7896
rect 23474 7828 23480 7880
rect 23532 7868 23538 7880
rect 24581 7871 24639 7877
rect 24581 7868 24593 7871
rect 23532 7840 24593 7868
rect 23532 7828 23538 7840
rect 24581 7837 24593 7840
rect 24627 7837 24639 7871
rect 24581 7831 24639 7837
rect 22888 7772 23336 7800
rect 24213 7803 24271 7809
rect 22888 7760 22894 7772
rect 24213 7769 24225 7803
rect 24259 7800 24271 7803
rect 25498 7800 25504 7812
rect 24259 7772 25504 7800
rect 24259 7769 24271 7772
rect 24213 7763 24271 7769
rect 25498 7760 25504 7772
rect 25556 7760 25562 7812
rect 1486 7692 1492 7744
rect 1544 7732 1550 7744
rect 1857 7735 1915 7741
rect 1857 7732 1869 7735
rect 1544 7704 1869 7732
rect 1544 7692 1550 7704
rect 1857 7701 1869 7704
rect 1903 7701 1915 7735
rect 1857 7695 1915 7701
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3568 7704 3801 7732
rect 3568 7692 3574 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 6270 7692 6276 7744
rect 6328 7732 6334 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 6328 7704 6653 7732
rect 6328 7692 6334 7704
rect 6641 7701 6653 7704
rect 6687 7701 6699 7735
rect 6641 7695 6699 7701
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8202 7732 8208 7744
rect 8067 7704 8208 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 11241 7735 11299 7741
rect 11241 7701 11253 7735
rect 11287 7732 11299 7735
rect 11698 7732 11704 7744
rect 11287 7704 11704 7732
rect 11287 7701 11299 7704
rect 11241 7695 11299 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 13265 7735 13323 7741
rect 13265 7701 13277 7735
rect 13311 7732 13323 7735
rect 13446 7732 13452 7744
rect 13311 7704 13452 7732
rect 13311 7701 13323 7704
rect 13265 7695 13323 7701
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14645 7735 14703 7741
rect 14645 7732 14657 7735
rect 13872 7704 14657 7732
rect 13872 7692 13878 7704
rect 14645 7701 14657 7704
rect 14691 7701 14703 7735
rect 14645 7695 14703 7701
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 16264 7704 17233 7732
rect 16264 7692 16270 7704
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 17221 7695 17279 7701
rect 19521 7735 19579 7741
rect 19521 7701 19533 7735
rect 19567 7732 19579 7735
rect 20438 7732 20444 7744
rect 19567 7704 20444 7732
rect 19567 7701 19579 7704
rect 19521 7695 19579 7701
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 20714 7732 20720 7744
rect 20675 7704 20720 7732
rect 20714 7692 20720 7704
rect 20772 7732 20778 7744
rect 21542 7732 21548 7744
rect 20772 7704 21548 7732
rect 20772 7692 20778 7704
rect 21542 7692 21548 7704
rect 21600 7692 21606 7744
rect 21726 7692 21732 7744
rect 21784 7732 21790 7744
rect 21913 7735 21971 7741
rect 21913 7732 21925 7735
rect 21784 7704 21925 7732
rect 21784 7692 21790 7704
rect 21913 7701 21925 7704
rect 21959 7701 21971 7735
rect 21913 7695 21971 7701
rect 22465 7735 22523 7741
rect 22465 7701 22477 7735
rect 22511 7732 22523 7735
rect 23198 7732 23204 7744
rect 22511 7704 23204 7732
rect 22511 7701 22523 7704
rect 22465 7695 22523 7701
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 23290 7692 23296 7744
rect 23348 7732 23354 7744
rect 23477 7735 23535 7741
rect 23477 7732 23489 7735
rect 23348 7704 23489 7732
rect 23348 7692 23354 7704
rect 23477 7701 23489 7704
rect 23523 7701 23535 7735
rect 23477 7695 23535 7701
rect 23937 7735 23995 7741
rect 23937 7701 23949 7735
rect 23983 7732 23995 7735
rect 24026 7732 24032 7744
rect 23983 7704 24032 7732
rect 23983 7701 23995 7704
rect 23937 7695 23995 7701
rect 24026 7692 24032 7704
rect 24084 7692 24090 7744
rect 24946 7732 24952 7744
rect 24907 7704 24952 7732
rect 24946 7692 24952 7704
rect 25004 7692 25010 7744
rect 25314 7732 25320 7744
rect 25275 7704 25320 7732
rect 25314 7692 25320 7704
rect 25372 7692 25378 7744
rect 25682 7732 25688 7744
rect 25643 7704 25688 7732
rect 25682 7692 25688 7704
rect 25740 7692 25746 7744
rect 26050 7732 26056 7744
rect 26011 7704 26056 7732
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 1104 7642 26864 7664
rect 1104 7590 5648 7642
rect 5700 7590 5712 7642
rect 5764 7590 5776 7642
rect 5828 7590 5840 7642
rect 5892 7590 14982 7642
rect 15034 7590 15046 7642
rect 15098 7590 15110 7642
rect 15162 7590 15174 7642
rect 15226 7590 24315 7642
rect 24367 7590 24379 7642
rect 24431 7590 24443 7642
rect 24495 7590 24507 7642
rect 24559 7590 26864 7642
rect 1104 7568 26864 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 5166 7528 5172 7540
rect 4663 7500 5172 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6362 7528 6368 7540
rect 6227 7500 6368 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 7650 7528 7656 7540
rect 7611 7500 7656 7528
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 8662 7528 8668 7540
rect 8623 7500 8668 7528
rect 8662 7488 8668 7500
rect 8720 7488 8726 7540
rect 10321 7531 10379 7537
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 10686 7528 10692 7540
rect 10367 7500 10692 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 10686 7488 10692 7500
rect 10744 7488 10750 7540
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 11882 7488 11888 7500
rect 11940 7528 11946 7540
rect 13081 7531 13139 7537
rect 13081 7528 13093 7531
rect 11940 7500 13093 7528
rect 11940 7488 11946 7500
rect 13081 7497 13093 7500
rect 13127 7528 13139 7531
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 13127 7500 13277 7528
rect 13127 7497 13139 7500
rect 13081 7491 13139 7497
rect 13265 7497 13277 7500
rect 13311 7528 13323 7531
rect 13538 7528 13544 7540
rect 13311 7500 13544 7528
rect 13311 7497 13323 7500
rect 13265 7491 13323 7497
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7528 15439 7531
rect 15654 7528 15660 7540
rect 15427 7500 15660 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 15654 7488 15660 7500
rect 15712 7488 15718 7540
rect 15838 7528 15844 7540
rect 15799 7500 15844 7528
rect 15838 7488 15844 7500
rect 15896 7488 15902 7540
rect 17129 7531 17187 7537
rect 17129 7497 17141 7531
rect 17175 7528 17187 7531
rect 17678 7528 17684 7540
rect 17175 7500 17684 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18138 7528 18144 7540
rect 18099 7500 18144 7528
rect 18138 7488 18144 7500
rect 18196 7488 18202 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19518 7528 19524 7540
rect 19475 7500 19524 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 19705 7531 19763 7537
rect 19705 7497 19717 7531
rect 19751 7528 19763 7531
rect 20622 7528 20628 7540
rect 19751 7500 20628 7528
rect 19751 7497 19763 7500
rect 19705 7491 19763 7497
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 22554 7488 22560 7540
rect 22612 7528 22618 7540
rect 22833 7531 22891 7537
rect 22833 7528 22845 7531
rect 22612 7500 22845 7528
rect 22612 7488 22618 7500
rect 22833 7497 22845 7500
rect 22879 7497 22891 7531
rect 22833 7491 22891 7497
rect 23014 7488 23020 7540
rect 23072 7528 23078 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 23072 7500 23213 7528
rect 23072 7488 23078 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23201 7491 23259 7497
rect 24673 7531 24731 7537
rect 24673 7497 24685 7531
rect 24719 7528 24731 7531
rect 24762 7528 24768 7540
rect 24719 7500 24768 7528
rect 24719 7497 24731 7500
rect 24673 7491 24731 7497
rect 24762 7488 24768 7500
rect 24820 7488 24826 7540
rect 25038 7488 25044 7540
rect 25096 7528 25102 7540
rect 25317 7531 25375 7537
rect 25317 7528 25329 7531
rect 25096 7500 25329 7528
rect 25096 7488 25102 7500
rect 25317 7497 25329 7500
rect 25363 7497 25375 7531
rect 25774 7528 25780 7540
rect 25735 7500 25780 7528
rect 25317 7491 25375 7497
rect 25774 7488 25780 7500
rect 25832 7488 25838 7540
rect 25866 7488 25872 7540
rect 25924 7528 25930 7540
rect 26053 7531 26111 7537
rect 26053 7528 26065 7531
rect 25924 7500 26065 7528
rect 25924 7488 25930 7500
rect 26053 7497 26065 7500
rect 26099 7497 26111 7531
rect 26053 7491 26111 7497
rect 2406 7460 2412 7472
rect 2056 7432 2412 7460
rect 2056 7401 2084 7432
rect 2406 7420 2412 7432
rect 2464 7420 2470 7472
rect 7193 7463 7251 7469
rect 7193 7429 7205 7463
rect 7239 7460 7251 7463
rect 8570 7460 8576 7472
rect 7239 7432 8576 7460
rect 7239 7429 7251 7432
rect 7193 7423 7251 7429
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 10597 7463 10655 7469
rect 10597 7429 10609 7463
rect 10643 7460 10655 7463
rect 10778 7460 10784 7472
rect 10643 7432 10784 7460
rect 10643 7429 10655 7432
rect 10597 7423 10655 7429
rect 10778 7420 10784 7432
rect 10836 7420 10842 7472
rect 16298 7420 16304 7472
rect 16356 7460 16362 7472
rect 20806 7460 20812 7472
rect 16356 7432 20812 7460
rect 16356 7420 16362 7432
rect 20806 7420 20812 7432
rect 20864 7420 20870 7472
rect 21177 7463 21235 7469
rect 21177 7429 21189 7463
rect 21223 7460 21235 7463
rect 24210 7460 24216 7472
rect 21223 7432 24216 7460
rect 21223 7429 21235 7432
rect 21177 7423 21235 7429
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7392 2283 7395
rect 2314 7392 2320 7404
rect 2271 7364 2320 7392
rect 2271 7361 2283 7364
rect 2225 7355 2283 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 3053 7395 3111 7401
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3234 7392 3240 7404
rect 3099 7364 3240 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 3234 7352 3240 7364
rect 3292 7392 3298 7404
rect 3789 7395 3847 7401
rect 3789 7392 3801 7395
rect 3292 7364 3801 7392
rect 3292 7352 3298 7364
rect 3789 7361 3801 7364
rect 3835 7392 3847 7395
rect 4614 7392 4620 7404
rect 3835 7364 4620 7392
rect 3835 7361 3847 7364
rect 3789 7355 3847 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 5261 7395 5319 7401
rect 5261 7392 5273 7395
rect 4764 7364 5273 7392
rect 4764 7352 4770 7364
rect 5261 7361 5273 7364
rect 5307 7361 5319 7395
rect 5261 7355 5319 7361
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8205 7395 8263 7401
rect 8205 7392 8217 7395
rect 8076 7364 8217 7392
rect 8076 7352 8082 7364
rect 8205 7361 8217 7364
rect 8251 7361 8263 7395
rect 8588 7392 8616 7420
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 8588 7364 9873 7392
rect 8205 7355 8263 7361
rect 9861 7361 9873 7364
rect 9907 7392 9919 7395
rect 10134 7392 10140 7404
rect 9907 7364 10140 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 10134 7352 10140 7364
rect 10192 7392 10198 7404
rect 11425 7395 11483 7401
rect 11425 7392 11437 7395
rect 10192 7364 11437 7392
rect 10192 7352 10198 7364
rect 11425 7361 11437 7364
rect 11471 7392 11483 7395
rect 11698 7392 11704 7404
rect 11471 7364 11704 7392
rect 11471 7361 11483 7364
rect 11425 7355 11483 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7392 12955 7395
rect 12943 7364 13492 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 13464 7336 13492 7364
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14826 7392 14832 7404
rect 14424 7364 14832 7392
rect 14424 7352 14430 7364
rect 14826 7352 14832 7364
rect 14884 7352 14890 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16393 7395 16451 7401
rect 16393 7392 16405 7395
rect 15795 7364 16405 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16393 7361 16405 7364
rect 16439 7361 16451 7395
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 16393 7355 16451 7361
rect 3602 7324 3608 7336
rect 3563 7296 3608 7324
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5166 7324 5172 7336
rect 5123 7296 5172 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 8846 7324 8852 7336
rect 5828 7296 8852 7324
rect 1949 7259 2007 7265
rect 1949 7225 1961 7259
rect 1995 7256 2007 7259
rect 2406 7256 2412 7268
rect 1995 7228 2412 7256
rect 1995 7225 2007 7228
rect 1949 7219 2007 7225
rect 2406 7216 2412 7228
rect 2464 7216 2470 7268
rect 3418 7216 3424 7268
rect 3476 7256 3482 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3476 7228 3525 7256
rect 3476 7216 3482 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 3513 7219 3571 7225
rect 4249 7259 4307 7265
rect 4249 7225 4261 7259
rect 4295 7256 4307 7259
rect 4982 7256 4988 7268
rect 4295 7228 4988 7256
rect 4295 7225 4307 7228
rect 4249 7219 4307 7225
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 5040 7228 5212 7256
rect 5040 7216 5046 7228
rect 2590 7188 2596 7200
rect 2551 7160 2596 7188
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 5184 7197 5212 7228
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 5721 7259 5779 7265
rect 5721 7256 5733 7259
rect 5500 7228 5733 7256
rect 5500 7216 5506 7228
rect 5721 7225 5733 7228
rect 5767 7225 5779 7259
rect 5721 7219 5779 7225
rect 5169 7191 5227 7197
rect 5169 7157 5181 7191
rect 5215 7188 5227 7191
rect 5828 7188 5856 7296
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7324 9183 7327
rect 9171 7296 9444 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 9416 7268 9444 7296
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9640 7296 9689 7324
rect 9640 7284 9646 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 10778 7284 10784 7336
rect 10836 7284 10842 7336
rect 11146 7324 11152 7336
rect 11107 7296 11152 7324
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 13127 7296 13369 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 13446 7284 13452 7336
rect 13504 7324 13510 7336
rect 13624 7327 13682 7333
rect 13624 7324 13636 7327
rect 13504 7296 13636 7324
rect 13504 7284 13510 7296
rect 13624 7293 13636 7296
rect 13670 7324 13682 7327
rect 15764 7324 15792 7355
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 19886 7352 19892 7404
rect 19944 7392 19950 7404
rect 20257 7395 20315 7401
rect 20257 7392 20269 7395
rect 19944 7364 20269 7392
rect 19944 7352 19950 7364
rect 20257 7361 20269 7364
rect 20303 7361 20315 7395
rect 20257 7355 20315 7361
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7392 21879 7395
rect 21867 7364 21956 7392
rect 21867 7361 21879 7364
rect 21821 7355 21879 7361
rect 21928 7336 21956 7364
rect 13670 7296 15792 7324
rect 17497 7327 17555 7333
rect 13670 7293 13682 7296
rect 13624 7287 13682 7293
rect 17497 7293 17509 7327
rect 17543 7324 17555 7327
rect 18230 7324 18236 7336
rect 17543 7296 18236 7324
rect 17543 7293 17555 7296
rect 17497 7287 17555 7293
rect 18230 7284 18236 7296
rect 18288 7324 18294 7336
rect 18509 7327 18567 7333
rect 18509 7324 18521 7327
rect 18288 7296 18521 7324
rect 18288 7284 18294 7296
rect 18509 7293 18521 7296
rect 18555 7324 18567 7327
rect 19058 7324 19064 7336
rect 18555 7296 19064 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 19058 7284 19064 7296
rect 19116 7284 19122 7336
rect 20070 7324 20076 7336
rect 20031 7296 20076 7324
rect 20070 7284 20076 7296
rect 20128 7284 20134 7336
rect 21910 7284 21916 7336
rect 21968 7284 21974 7336
rect 23676 7333 23704 7432
rect 24210 7420 24216 7432
rect 24268 7420 24274 7472
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 23842 7284 23848 7336
rect 23900 7324 23906 7336
rect 24762 7324 24768 7336
rect 23900 7296 24768 7324
rect 23900 7284 23906 7296
rect 24762 7284 24768 7296
rect 24820 7284 24826 7336
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 26418 7284 26424 7296
rect 26476 7284 26482 7336
rect 6641 7259 6699 7265
rect 6641 7225 6653 7259
rect 6687 7256 6699 7259
rect 8021 7259 8079 7265
rect 8021 7256 8033 7259
rect 6687 7228 8033 7256
rect 6687 7225 6699 7228
rect 6641 7219 6699 7225
rect 8021 7225 8033 7228
rect 8067 7256 8079 7259
rect 8067 7228 9260 7256
rect 8067 7225 8079 7228
rect 8021 7219 8079 7225
rect 7466 7188 7472 7200
rect 5215 7160 5856 7188
rect 7427 7160 7472 7188
rect 5215 7157 5227 7160
rect 5169 7151 5227 7157
rect 7466 7148 7472 7160
rect 7524 7148 7530 7200
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 9232 7197 9260 7228
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 10796 7256 10824 7284
rect 11241 7259 11299 7265
rect 11241 7256 11253 7259
rect 9456 7228 9628 7256
rect 10796 7228 11253 7256
rect 9456 7216 9462 7228
rect 9600 7197 9628 7228
rect 11241 7225 11253 7228
rect 11287 7225 11299 7259
rect 18874 7256 18880 7268
rect 11241 7219 11299 7225
rect 18616 7228 18880 7256
rect 9217 7191 9275 7197
rect 9217 7157 9229 7191
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 9585 7191 9643 7197
rect 9585 7157 9597 7191
rect 9631 7157 9643 7191
rect 10778 7188 10784 7200
rect 10739 7160 10784 7188
rect 9585 7151 9643 7157
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 14737 7191 14795 7197
rect 14737 7157 14749 7191
rect 14783 7188 14795 7191
rect 14826 7188 14832 7200
rect 14783 7160 14832 7188
rect 14783 7157 14795 7160
rect 14737 7151 14795 7157
rect 14826 7148 14832 7160
rect 14884 7148 14890 7200
rect 16206 7188 16212 7200
rect 16167 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16298 7148 16304 7200
rect 16356 7188 16362 7200
rect 17865 7191 17923 7197
rect 16356 7160 16401 7188
rect 16356 7148 16362 7160
rect 17865 7157 17877 7191
rect 17911 7188 17923 7191
rect 18230 7188 18236 7200
rect 17911 7160 18236 7188
rect 17911 7157 17923 7160
rect 17865 7151 17923 7157
rect 18230 7148 18236 7160
rect 18288 7188 18294 7200
rect 18616 7197 18644 7228
rect 18874 7216 18880 7228
rect 18932 7216 18938 7268
rect 19242 7216 19248 7268
rect 19300 7256 19306 7268
rect 19978 7256 19984 7268
rect 19300 7228 19984 7256
rect 19300 7216 19306 7228
rect 19978 7216 19984 7228
rect 20036 7256 20042 7268
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 20036 7228 20177 7256
rect 20036 7216 20042 7228
rect 20165 7225 20177 7228
rect 20211 7225 20223 7259
rect 21177 7259 21235 7265
rect 21177 7256 21189 7259
rect 20165 7219 20223 7225
rect 20916 7228 21189 7256
rect 18601 7191 18659 7197
rect 18601 7188 18613 7191
rect 18288 7160 18613 7188
rect 18288 7148 18294 7160
rect 18601 7157 18613 7160
rect 18647 7157 18659 7191
rect 18601 7151 18659 7157
rect 18690 7148 18696 7200
rect 18748 7188 18754 7200
rect 19150 7188 19156 7200
rect 18748 7160 19156 7188
rect 18748 7148 18754 7160
rect 19150 7148 19156 7160
rect 19208 7188 19214 7200
rect 20916 7188 20944 7228
rect 21177 7225 21189 7228
rect 21223 7225 21235 7259
rect 21177 7219 21235 7225
rect 21637 7259 21695 7265
rect 21637 7225 21649 7259
rect 21683 7256 21695 7259
rect 21683 7228 21864 7256
rect 21683 7225 21695 7228
rect 21637 7219 21695 7225
rect 19208 7160 20944 7188
rect 20993 7191 21051 7197
rect 19208 7148 19214 7160
rect 20993 7157 21005 7191
rect 21039 7188 21051 7191
rect 21266 7188 21272 7200
rect 21039 7160 21272 7188
rect 21039 7157 21051 7160
rect 20993 7151 21051 7157
rect 21266 7148 21272 7160
rect 21324 7148 21330 7200
rect 21726 7188 21732 7200
rect 21687 7160 21732 7188
rect 21726 7148 21732 7160
rect 21784 7148 21790 7200
rect 21836 7188 21864 7228
rect 22094 7188 22100 7200
rect 21836 7160 22100 7188
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 22557 7191 22615 7197
rect 22557 7157 22569 7191
rect 22603 7188 22615 7191
rect 22738 7188 22744 7200
rect 22603 7160 22744 7188
rect 22603 7157 22615 7160
rect 22557 7151 22615 7157
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 23845 7191 23903 7197
rect 23845 7157 23857 7191
rect 23891 7188 23903 7191
rect 24118 7188 24124 7200
rect 23891 7160 24124 7188
rect 23891 7157 23903 7160
rect 23845 7151 23903 7157
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25958 7188 25964 7200
rect 24995 7160 25964 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25958 7148 25964 7160
rect 26016 7148 26022 7200
rect 1104 7098 26864 7120
rect 1104 7046 10315 7098
rect 10367 7046 10379 7098
rect 10431 7046 10443 7098
rect 10495 7046 10507 7098
rect 10559 7046 19648 7098
rect 19700 7046 19712 7098
rect 19764 7046 19776 7098
rect 19828 7046 19840 7098
rect 19892 7046 26864 7098
rect 1104 7024 26864 7046
rect 2406 6984 2412 6996
rect 2367 6956 2412 6984
rect 2406 6944 2412 6956
rect 2464 6944 2470 6996
rect 2777 6987 2835 6993
rect 2777 6953 2789 6987
rect 2823 6984 2835 6987
rect 3142 6984 3148 6996
rect 2823 6956 3148 6984
rect 2823 6953 2835 6956
rect 2777 6947 2835 6953
rect 3142 6944 3148 6956
rect 3200 6944 3206 6996
rect 4433 6987 4491 6993
rect 4433 6953 4445 6987
rect 4479 6984 4491 6987
rect 4706 6984 4712 6996
rect 4479 6956 4712 6984
rect 4479 6953 4491 6956
rect 4433 6947 4491 6953
rect 4706 6944 4712 6956
rect 4764 6944 4770 6996
rect 6457 6987 6515 6993
rect 6457 6953 6469 6987
rect 6503 6984 6515 6987
rect 6822 6984 6828 6996
rect 6503 6956 6828 6984
rect 6503 6953 6515 6956
rect 6457 6947 6515 6953
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 8570 6944 8576 6996
rect 8628 6984 8634 6996
rect 9217 6987 9275 6993
rect 9217 6984 9229 6987
rect 8628 6956 9229 6984
rect 8628 6944 8634 6956
rect 9217 6953 9229 6956
rect 9263 6953 9275 6987
rect 9950 6984 9956 6996
rect 9911 6956 9956 6984
rect 9217 6947 9275 6953
rect 9950 6944 9956 6956
rect 10008 6944 10014 6996
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 12124 6956 12265 6984
rect 12124 6944 12130 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 13814 6944 13820 6996
rect 13872 6984 13878 6996
rect 15102 6984 15108 6996
rect 13872 6956 15108 6984
rect 13872 6944 13878 6956
rect 15102 6944 15108 6956
rect 15160 6944 15166 6996
rect 15654 6944 15660 6996
rect 15712 6984 15718 6996
rect 18598 6984 18604 6996
rect 15712 6956 16528 6984
rect 18559 6956 18604 6984
rect 15712 6944 15718 6956
rect 1673 6919 1731 6925
rect 1673 6885 1685 6919
rect 1719 6916 1731 6919
rect 2314 6916 2320 6928
rect 1719 6888 2320 6916
rect 1719 6885 1731 6888
rect 1673 6879 1731 6885
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 8386 6916 8392 6928
rect 8299 6888 8392 6916
rect 8386 6876 8392 6888
rect 8444 6916 8450 6928
rect 10778 6916 10784 6928
rect 8444 6888 10784 6916
rect 8444 6876 8450 6888
rect 10778 6876 10784 6888
rect 10836 6876 10842 6928
rect 13173 6919 13231 6925
rect 13173 6916 13185 6919
rect 12268 6888 13185 6916
rect 12268 6860 12296 6888
rect 13173 6885 13185 6888
rect 13219 6885 13231 6919
rect 16298 6916 16304 6928
rect 13173 6879 13231 6885
rect 15120 6888 16304 6916
rect 2869 6851 2927 6857
rect 2869 6817 2881 6851
rect 2915 6848 2927 6851
rect 4062 6848 4068 6860
rect 2915 6820 4068 6848
rect 2915 6817 2927 6820
rect 2869 6811 2927 6817
rect 4062 6808 4068 6820
rect 4120 6808 4126 6860
rect 4522 6848 4528 6860
rect 4483 6820 4528 6848
rect 4522 6808 4528 6820
rect 4580 6808 4586 6860
rect 5810 6848 5816 6860
rect 5771 6820 5816 6848
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7340 6820 7757 6848
rect 7340 6808 7346 6820
rect 7745 6817 7757 6820
rect 7791 6848 7803 6851
rect 8018 6848 8024 6860
rect 7791 6820 8024 6848
rect 7791 6817 7803 6820
rect 7745 6811 7803 6817
rect 8018 6808 8024 6820
rect 8076 6848 8082 6860
rect 10588 6851 10646 6857
rect 8076 6820 8708 6848
rect 8076 6808 8082 6820
rect 8680 6792 8708 6820
rect 10588 6817 10600 6851
rect 10634 6848 10646 6851
rect 11146 6848 11152 6860
rect 10634 6820 11152 6848
rect 10634 6817 10646 6820
rect 10588 6811 10646 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 12250 6808 12256 6860
rect 12308 6808 12314 6860
rect 14734 6808 14740 6860
rect 14792 6848 14798 6860
rect 15013 6851 15071 6857
rect 15013 6848 15025 6851
rect 14792 6820 15025 6848
rect 14792 6808 14798 6820
rect 15013 6817 15025 6820
rect 15059 6848 15071 6851
rect 15120 6848 15148 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 15059 6820 15148 6848
rect 15059 6817 15071 6820
rect 15013 6811 15071 6817
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15252 6820 15577 6848
rect 15252 6808 15258 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 16500 6848 16528 6956
rect 18598 6944 18604 6956
rect 18656 6944 18662 6996
rect 19426 6944 19432 6996
rect 19484 6984 19490 6996
rect 19613 6987 19671 6993
rect 19613 6984 19625 6987
rect 19484 6956 19625 6984
rect 19484 6944 19490 6956
rect 19613 6953 19625 6956
rect 19659 6953 19671 6987
rect 19613 6947 19671 6953
rect 20990 6944 20996 6996
rect 21048 6984 21054 6996
rect 21269 6987 21327 6993
rect 21269 6984 21281 6987
rect 21048 6956 21281 6984
rect 21048 6944 21054 6956
rect 21269 6953 21281 6956
rect 21315 6984 21327 6987
rect 21818 6984 21824 6996
rect 21315 6956 21824 6984
rect 21315 6953 21327 6956
rect 21269 6947 21327 6953
rect 21818 6944 21824 6956
rect 21876 6944 21882 6996
rect 22370 6944 22376 6996
rect 22428 6984 22434 6996
rect 22833 6987 22891 6993
rect 22833 6984 22845 6987
rect 22428 6956 22845 6984
rect 22428 6944 22434 6956
rect 22833 6953 22845 6956
rect 22879 6953 22891 6987
rect 22833 6947 22891 6953
rect 22940 6956 23704 6984
rect 18966 6876 18972 6928
rect 19024 6916 19030 6928
rect 22278 6916 22284 6928
rect 19024 6888 22284 6916
rect 19024 6876 19030 6888
rect 22278 6876 22284 6888
rect 22336 6916 22342 6928
rect 22462 6916 22468 6928
rect 22336 6888 22468 6916
rect 22336 6876 22342 6888
rect 22462 6876 22468 6888
rect 22520 6876 22526 6928
rect 22554 6876 22560 6928
rect 22612 6916 22618 6928
rect 22940 6916 22968 6956
rect 22612 6888 22968 6916
rect 22612 6876 22618 6888
rect 23014 6876 23020 6928
rect 23072 6916 23078 6928
rect 23676 6916 23704 6956
rect 23750 6944 23756 6996
rect 23808 6984 23814 6996
rect 24026 6984 24032 6996
rect 23808 6956 24032 6984
rect 23808 6944 23814 6956
rect 24026 6944 24032 6956
rect 24084 6944 24090 6996
rect 24762 6984 24768 6996
rect 24723 6956 24768 6984
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 23072 6888 23520 6916
rect 23676 6888 23796 6916
rect 23072 6876 23078 6888
rect 16669 6851 16727 6857
rect 16669 6848 16681 6851
rect 16500 6820 16681 6848
rect 15565 6811 15623 6817
rect 16669 6817 16681 6820
rect 16715 6817 16727 6851
rect 16669 6811 16727 6817
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 16925 6851 16983 6857
rect 16925 6848 16937 6851
rect 16816 6820 16937 6848
rect 16816 6808 16822 6820
rect 16925 6817 16937 6820
rect 16971 6817 16983 6851
rect 16925 6811 16983 6817
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6817 19579 6851
rect 19521 6811 19579 6817
rect 2958 6780 2964 6792
rect 2919 6752 2964 6780
rect 2958 6740 2964 6752
rect 3016 6740 3022 6792
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6549 6783 6607 6789
rect 6549 6780 6561 6783
rect 6052 6752 6561 6780
rect 6052 6740 6058 6752
rect 6549 6749 6561 6752
rect 6595 6749 6607 6783
rect 6549 6743 6607 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 3142 6672 3148 6724
rect 3200 6712 3206 6724
rect 3789 6715 3847 6721
rect 3789 6712 3801 6715
rect 3200 6684 3801 6712
rect 3200 6672 3206 6684
rect 3789 6681 3801 6684
rect 3835 6681 3847 6715
rect 3789 6675 3847 6681
rect 5537 6715 5595 6721
rect 5537 6681 5549 6715
rect 5583 6712 5595 6715
rect 5626 6712 5632 6724
rect 5583 6684 5632 6712
rect 5583 6681 5595 6684
rect 5537 6675 5595 6681
rect 5626 6672 5632 6684
rect 5684 6672 5690 6724
rect 6086 6712 6092 6724
rect 6047 6684 6092 6712
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 6362 6672 6368 6724
rect 6420 6712 6426 6724
rect 6656 6712 6684 6743
rect 8294 6740 8300 6792
rect 8352 6780 8358 6792
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 8352 6752 8493 6780
rect 8352 6740 8358 6752
rect 8481 6749 8493 6752
rect 8527 6749 8539 6783
rect 8662 6780 8668 6792
rect 8623 6752 8668 6780
rect 8481 6743 8539 6749
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 9950 6740 9956 6792
rect 10008 6780 10014 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 10008 6752 10333 6780
rect 10008 6740 10014 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 13262 6780 13268 6792
rect 13223 6752 13268 6780
rect 10321 6743 10379 6749
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6749 13415 6783
rect 13357 6743 13415 6749
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14090 6780 14096 6792
rect 13955 6752 14096 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 6420 6684 6684 6712
rect 7377 6715 7435 6721
rect 6420 6672 6426 6684
rect 7377 6681 7389 6715
rect 7423 6712 7435 6715
rect 8202 6712 8208 6724
rect 7423 6684 8208 6712
rect 7423 6681 7435 6684
rect 7377 6675 7435 6681
rect 8202 6672 8208 6684
rect 8260 6672 8266 6724
rect 12802 6712 12808 6724
rect 12763 6684 12808 6712
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 2314 6644 2320 6656
rect 2275 6616 2320 6644
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 2498 6604 2504 6656
rect 2556 6644 2562 6656
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2556 6616 3433 6644
rect 2556 6604 2562 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 4062 6644 4068 6656
rect 4023 6616 4068 6644
rect 3421 6607 3479 6613
rect 4062 6604 4068 6616
rect 4120 6604 4126 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 8018 6644 8024 6656
rect 7979 6616 8024 6644
rect 8018 6604 8024 6616
rect 8076 6604 8082 6656
rect 11698 6644 11704 6656
rect 11611 6616 11704 6644
rect 11698 6604 11704 6616
rect 11756 6644 11762 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 11756 6616 12725 6644
rect 11756 6604 11762 6616
rect 12713 6613 12725 6616
rect 12759 6644 12771 6647
rect 13372 6644 13400 6743
rect 14090 6740 14096 6752
rect 14148 6780 14154 6792
rect 14918 6780 14924 6792
rect 14148 6752 14924 6780
rect 14148 6740 14154 6752
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18012 6752 18981 6780
rect 18012 6740 18018 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6712 14427 6715
rect 15010 6712 15016 6724
rect 14415 6684 15016 6712
rect 14415 6681 14427 6684
rect 14369 6675 14427 6681
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 19536 6656 19564 6811
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21361 6851 21419 6857
rect 21361 6848 21373 6851
rect 20864 6820 21373 6848
rect 20864 6808 20870 6820
rect 21361 6817 21373 6820
rect 21407 6848 21419 6851
rect 21818 6848 21824 6860
rect 21407 6820 21824 6848
rect 21407 6817 21419 6820
rect 21361 6811 21419 6817
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 22373 6851 22431 6857
rect 22373 6817 22385 6851
rect 22419 6848 22431 6851
rect 22925 6851 22983 6857
rect 22925 6848 22937 6851
rect 22419 6820 22937 6848
rect 22419 6817 22431 6820
rect 22373 6811 22431 6817
rect 22925 6817 22937 6820
rect 22971 6848 22983 6851
rect 23382 6848 23388 6860
rect 22971 6820 23388 6848
rect 22971 6817 22983 6820
rect 22925 6811 22983 6817
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 23492 6848 23520 6888
rect 23658 6848 23664 6860
rect 23492 6820 23664 6848
rect 23658 6808 23664 6820
rect 23716 6808 23722 6860
rect 23768 6848 23796 6888
rect 24026 6848 24032 6860
rect 23768 6820 24032 6848
rect 24026 6808 24032 6820
rect 24084 6808 24090 6860
rect 25133 6851 25191 6857
rect 25133 6817 25145 6851
rect 25179 6817 25191 6851
rect 25133 6811 25191 6817
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19668 6752 19717 6780
rect 19668 6740 19674 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 21453 6783 21511 6789
rect 21453 6749 21465 6783
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 20346 6672 20352 6724
rect 20404 6712 20410 6724
rect 20901 6715 20959 6721
rect 20901 6712 20913 6715
rect 20404 6684 20913 6712
rect 20404 6672 20410 6684
rect 20901 6681 20913 6684
rect 20947 6681 20959 6715
rect 20901 6675 20959 6681
rect 21358 6672 21364 6724
rect 21416 6712 21422 6724
rect 21468 6712 21496 6743
rect 21910 6740 21916 6792
rect 21968 6780 21974 6792
rect 23106 6780 23112 6792
rect 21968 6752 23112 6780
rect 21968 6740 21974 6752
rect 23106 6740 23112 6752
rect 23164 6740 23170 6792
rect 25148 6780 25176 6811
rect 25774 6780 25780 6792
rect 23400 6752 25780 6780
rect 23400 6724 23428 6752
rect 25774 6740 25780 6752
rect 25832 6740 25838 6792
rect 21416 6684 21496 6712
rect 21416 6672 21422 6684
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 22465 6715 22523 6721
rect 22465 6712 22477 6715
rect 22152 6684 22477 6712
rect 22152 6672 22158 6684
rect 22465 6681 22477 6684
rect 22511 6712 22523 6715
rect 23290 6712 23296 6724
rect 22511 6684 23296 6712
rect 22511 6681 22523 6684
rect 22465 6675 22523 6681
rect 23290 6672 23296 6684
rect 23348 6672 23354 6724
rect 23382 6672 23388 6724
rect 23440 6672 23446 6724
rect 14734 6644 14740 6656
rect 12759 6616 13400 6644
rect 14695 6616 14740 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16114 6644 16120 6656
rect 16075 6616 16120 6644
rect 16114 6604 16120 6616
rect 16172 6604 16178 6656
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6644 16635 6647
rect 16666 6644 16672 6656
rect 16623 6616 16672 6644
rect 16623 6613 16635 6616
rect 16577 6607 16635 6613
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 17034 6604 17040 6656
rect 17092 6644 17098 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 17092 6616 18061 6644
rect 17092 6604 17098 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 19150 6644 19156 6656
rect 19111 6616 19156 6644
rect 18049 6607 18107 6613
rect 19150 6604 19156 6616
rect 19208 6604 19214 6656
rect 19518 6604 19524 6656
rect 19576 6604 19582 6656
rect 19978 6604 19984 6656
rect 20036 6644 20042 6656
rect 20165 6647 20223 6653
rect 20165 6644 20177 6647
rect 20036 6616 20177 6644
rect 20036 6604 20042 6616
rect 20165 6613 20177 6616
rect 20211 6613 20223 6647
rect 20714 6644 20720 6656
rect 20675 6616 20720 6644
rect 20165 6607 20223 6613
rect 20714 6604 20720 6616
rect 20772 6644 20778 6656
rect 21174 6644 21180 6656
rect 20772 6616 21180 6644
rect 20772 6604 20778 6616
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 22002 6644 22008 6656
rect 21963 6616 22008 6644
rect 22002 6604 22008 6616
rect 22060 6604 22066 6656
rect 23566 6604 23572 6656
rect 23624 6644 23630 6656
rect 24213 6647 24271 6653
rect 24213 6644 24225 6647
rect 23624 6616 24225 6644
rect 23624 6604 23630 6616
rect 24213 6613 24225 6616
rect 24259 6613 24271 6647
rect 24213 6607 24271 6613
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25317 6647 25375 6653
rect 25317 6644 25329 6647
rect 24912 6616 25329 6644
rect 24912 6604 24918 6616
rect 25317 6613 25329 6616
rect 25363 6613 25375 6647
rect 25682 6644 25688 6656
rect 25643 6616 25688 6644
rect 25317 6607 25375 6613
rect 25682 6604 25688 6616
rect 25740 6604 25746 6656
rect 26050 6644 26056 6656
rect 26011 6616 26056 6644
rect 26050 6604 26056 6616
rect 26108 6604 26114 6656
rect 1104 6554 26864 6576
rect 1104 6502 5648 6554
rect 5700 6502 5712 6554
rect 5764 6502 5776 6554
rect 5828 6502 5840 6554
rect 5892 6502 14982 6554
rect 15034 6502 15046 6554
rect 15098 6502 15110 6554
rect 15162 6502 15174 6554
rect 15226 6502 24315 6554
rect 24367 6502 24379 6554
rect 24431 6502 24443 6554
rect 24495 6502 24507 6554
rect 24559 6502 26864 6554
rect 1104 6480 26864 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 3234 6440 3240 6452
rect 3195 6412 3240 6440
rect 3234 6400 3240 6412
rect 3292 6400 3298 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6089 6443 6147 6449
rect 6089 6440 6101 6443
rect 6052 6412 6101 6440
rect 6052 6400 6058 6412
rect 6089 6409 6101 6412
rect 6135 6409 6147 6443
rect 6089 6403 6147 6409
rect 6549 6443 6607 6449
rect 6549 6409 6561 6443
rect 6595 6440 6607 6443
rect 6822 6440 6828 6452
rect 6595 6412 6828 6440
rect 6595 6409 6607 6412
rect 6549 6403 6607 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7282 6440 7288 6452
rect 7243 6412 7288 6440
rect 7282 6400 7288 6412
rect 7340 6400 7346 6452
rect 10410 6440 10416 6452
rect 10371 6412 10416 6440
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6440 11667 6443
rect 11882 6440 11888 6452
rect 11655 6412 11888 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12526 6400 12532 6452
rect 12584 6440 12590 6452
rect 15470 6440 15476 6452
rect 12584 6412 15476 6440
rect 12584 6400 12590 6412
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 16393 6443 16451 6449
rect 16393 6409 16405 6443
rect 16439 6440 16451 6443
rect 16482 6440 16488 6452
rect 16439 6412 16488 6440
rect 16439 6409 16451 6412
rect 16393 6403 16451 6409
rect 16482 6400 16488 6412
rect 16540 6400 16546 6452
rect 18049 6443 18107 6449
rect 18049 6409 18061 6443
rect 18095 6440 18107 6443
rect 19242 6440 19248 6452
rect 18095 6412 19248 6440
rect 18095 6409 18107 6412
rect 18049 6403 18107 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 20990 6440 20996 6452
rect 20951 6412 20996 6440
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 21174 6440 21180 6452
rect 21135 6412 21180 6440
rect 21174 6400 21180 6412
rect 21232 6400 21238 6452
rect 23382 6440 23388 6452
rect 21468 6412 23388 6440
rect 1765 6375 1823 6381
rect 1765 6341 1777 6375
rect 1811 6372 1823 6375
rect 2590 6372 2596 6384
rect 1811 6344 2596 6372
rect 1811 6341 1823 6344
rect 1765 6335 1823 6341
rect 2590 6332 2596 6344
rect 2648 6372 2654 6384
rect 2958 6372 2964 6384
rect 2648 6344 2964 6372
rect 2648 6332 2654 6344
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 5813 6375 5871 6381
rect 5813 6341 5825 6375
rect 5859 6372 5871 6375
rect 5902 6372 5908 6384
rect 5859 6344 5908 6372
rect 5859 6341 5871 6344
rect 5813 6335 5871 6341
rect 5902 6332 5908 6344
rect 5960 6372 5966 6384
rect 6362 6372 6368 6384
rect 5960 6344 6368 6372
rect 5960 6332 5966 6344
rect 6362 6332 6368 6344
rect 6420 6332 6426 6384
rect 10045 6375 10103 6381
rect 10045 6341 10057 6375
rect 10091 6372 10103 6375
rect 10870 6372 10876 6384
rect 10091 6344 10876 6372
rect 10091 6341 10103 6344
rect 10045 6335 10103 6341
rect 10870 6332 10876 6344
rect 10928 6372 10934 6384
rect 10928 6344 11008 6372
rect 10928 6332 10934 6344
rect 2314 6264 2320 6316
rect 2372 6304 2378 6316
rect 10980 6313 11008 6344
rect 14550 6332 14556 6384
rect 14608 6372 14614 6384
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 14608 6344 19073 6372
rect 14608 6332 14614 6344
rect 19061 6341 19073 6344
rect 19107 6372 19119 6375
rect 19702 6372 19708 6384
rect 19107 6344 19708 6372
rect 19107 6341 19119 6344
rect 19061 6335 19119 6341
rect 19702 6332 19708 6344
rect 19760 6372 19766 6384
rect 20254 6372 20260 6384
rect 19760 6344 20260 6372
rect 19760 6332 19766 6344
rect 20254 6332 20260 6344
rect 20312 6332 20318 6384
rect 20622 6332 20628 6384
rect 20680 6372 20686 6384
rect 21468 6372 21496 6412
rect 23382 6400 23388 6412
rect 23440 6400 23446 6452
rect 24026 6400 24032 6452
rect 24084 6440 24090 6452
rect 24673 6443 24731 6449
rect 24673 6440 24685 6443
rect 24084 6412 24685 6440
rect 24084 6400 24090 6412
rect 24673 6409 24685 6412
rect 24719 6409 24731 6443
rect 25130 6440 25136 6452
rect 25091 6412 25136 6440
rect 24673 6403 24731 6409
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 25774 6440 25780 6452
rect 25735 6412 25780 6440
rect 25774 6400 25780 6412
rect 25832 6400 25838 6452
rect 20680 6344 21496 6372
rect 20680 6332 20686 6344
rect 21542 6332 21548 6384
rect 21600 6372 21606 6384
rect 22370 6372 22376 6384
rect 21600 6344 22376 6372
rect 21600 6332 21606 6344
rect 22370 6332 22376 6344
rect 22428 6332 22434 6384
rect 23290 6332 23296 6384
rect 23348 6372 23354 6384
rect 23842 6372 23848 6384
rect 23348 6344 23848 6372
rect 23348 6332 23354 6344
rect 23842 6332 23848 6344
rect 23900 6332 23906 6384
rect 23934 6332 23940 6384
rect 23992 6372 23998 6384
rect 24302 6372 24308 6384
rect 23992 6344 24308 6372
rect 23992 6332 23998 6344
rect 24302 6332 24308 6344
rect 24360 6332 24366 6384
rect 2777 6307 2835 6313
rect 2777 6304 2789 6307
rect 2372 6276 2789 6304
rect 2372 6264 2378 6276
rect 2777 6273 2789 6276
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 7745 6307 7803 6313
rect 7745 6304 7757 6307
rect 7515 6276 7757 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7745 6273 7757 6276
rect 7791 6273 7803 6307
rect 7745 6267 7803 6273
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 11146 6304 11152 6316
rect 11107 6276 11152 6304
rect 10965 6267 11023 6273
rect 11146 6264 11152 6276
rect 11204 6304 11210 6316
rect 11977 6307 12035 6313
rect 11977 6304 11989 6307
rect 11204 6276 11989 6304
rect 11204 6264 11210 6276
rect 11977 6273 11989 6276
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6304 16359 6307
rect 17034 6304 17040 6316
rect 16347 6276 17040 6304
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 18380 6276 18705 6304
rect 18380 6264 18386 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 18874 6304 18880 6316
rect 18739 6276 18880 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 18874 6264 18880 6276
rect 18932 6264 18938 6316
rect 19978 6304 19984 6316
rect 19260 6276 19984 6304
rect 2038 6196 2044 6248
rect 2096 6236 2102 6248
rect 2590 6236 2596 6248
rect 2096 6208 2596 6236
rect 2096 6196 2102 6208
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 3789 6239 3847 6245
rect 3789 6236 3801 6239
rect 3344 6208 3801 6236
rect 3344 6112 3372 6208
rect 3789 6205 3801 6208
rect 3835 6236 3847 6239
rect 3835 6208 4292 6236
rect 3835 6205 3847 6208
rect 3789 6199 3847 6205
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 4034 6171 4092 6177
rect 4034 6168 4046 6171
rect 3476 6140 4046 6168
rect 3476 6128 3482 6140
rect 4034 6137 4046 6140
rect 4080 6137 4092 6171
rect 4264 6168 4292 6208
rect 4338 6196 4344 6248
rect 4396 6236 4402 6248
rect 8938 6236 8944 6248
rect 4396 6208 8944 6236
rect 4396 6196 4402 6208
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 10873 6239 10931 6245
rect 10873 6236 10885 6239
rect 10468 6208 10885 6236
rect 10468 6196 10474 6208
rect 10873 6205 10885 6208
rect 10919 6205 10931 6239
rect 12989 6239 13047 6245
rect 12989 6236 13001 6239
rect 10873 6199 10931 6205
rect 12820 6208 13001 6236
rect 5442 6168 5448 6180
rect 4264 6140 5448 6168
rect 4034 6131 4092 6137
rect 5442 6128 5448 6140
rect 5500 6168 5506 6180
rect 7469 6171 7527 6177
rect 7469 6168 7481 6171
rect 5500 6140 7481 6168
rect 5500 6128 5506 6140
rect 7469 6137 7481 6140
rect 7515 6168 7527 6171
rect 7561 6171 7619 6177
rect 7561 6168 7573 6171
rect 7515 6140 7573 6168
rect 7515 6137 7527 6140
rect 7469 6131 7527 6137
rect 7561 6137 7573 6140
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 8012 6171 8070 6177
rect 8012 6137 8024 6171
rect 8058 6168 8070 6171
rect 8202 6168 8208 6180
rect 8058 6140 8208 6168
rect 8058 6137 8070 6140
rect 8012 6131 8070 6137
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3605 6103 3663 6109
rect 3605 6100 3617 6103
rect 3384 6072 3617 6100
rect 3384 6060 3390 6072
rect 3605 6069 3617 6072
rect 3651 6069 3663 6103
rect 5166 6100 5172 6112
rect 5127 6072 5172 6100
rect 3605 6063 3663 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5258 6060 5264 6112
rect 5316 6100 5322 6112
rect 8754 6100 8760 6112
rect 5316 6072 8760 6100
rect 5316 6060 5322 6072
rect 8754 6060 8760 6072
rect 8812 6060 8818 6112
rect 9125 6103 9183 6109
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 9766 6100 9772 6112
rect 9171 6072 9772 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10505 6103 10563 6109
rect 10505 6069 10517 6103
rect 10551 6100 10563 6103
rect 10778 6100 10784 6112
rect 10551 6072 10784 6100
rect 10551 6069 10563 6072
rect 10505 6063 10563 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11882 6060 11888 6112
rect 11940 6100 11946 6112
rect 12526 6100 12532 6112
rect 11940 6072 12532 6100
rect 11940 6060 11946 6072
rect 12526 6060 12532 6072
rect 12584 6100 12590 6112
rect 12820 6109 12848 6208
rect 12989 6205 13001 6208
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 13256 6239 13314 6245
rect 13256 6205 13268 6239
rect 13302 6236 13314 6239
rect 14090 6236 14096 6248
rect 13302 6208 14096 6236
rect 13302 6205 13314 6208
rect 13256 6199 13314 6205
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 16850 6236 16856 6248
rect 16763 6208 16856 6236
rect 16850 6196 16856 6208
rect 16908 6236 16914 6248
rect 19150 6236 19156 6248
rect 16908 6208 19156 6236
rect 16908 6196 16914 6208
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 15749 6171 15807 6177
rect 15749 6137 15761 6171
rect 15795 6168 15807 6171
rect 16482 6168 16488 6180
rect 15795 6140 16488 6168
rect 15795 6137 15807 6140
rect 15749 6131 15807 6137
rect 16482 6128 16488 6140
rect 16540 6128 16546 6180
rect 16761 6171 16819 6177
rect 16761 6137 16773 6171
rect 16807 6168 16819 6171
rect 17126 6168 17132 6180
rect 16807 6140 17132 6168
rect 16807 6137 16819 6140
rect 16761 6131 16819 6137
rect 17126 6128 17132 6140
rect 17184 6128 17190 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 17773 6171 17831 6177
rect 17773 6168 17785 6171
rect 17368 6140 17785 6168
rect 17368 6128 17374 6140
rect 17773 6137 17785 6140
rect 17819 6168 17831 6171
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 17819 6140 18429 6168
rect 17819 6137 17831 6140
rect 17773 6131 17831 6137
rect 18417 6137 18429 6140
rect 18463 6137 18475 6171
rect 19260 6168 19288 6276
rect 19978 6264 19984 6276
rect 20036 6264 20042 6316
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 20128 6276 20177 6304
rect 20128 6264 20134 6276
rect 20165 6273 20177 6276
rect 20211 6273 20223 6307
rect 20165 6267 20223 6273
rect 21174 6264 21180 6316
rect 21232 6304 21238 6316
rect 21358 6304 21364 6316
rect 21232 6276 21364 6304
rect 21232 6264 21238 6276
rect 21358 6264 21364 6276
rect 21416 6304 21422 6316
rect 21729 6307 21787 6313
rect 21729 6304 21741 6307
rect 21416 6276 21741 6304
rect 21416 6264 21422 6276
rect 21729 6273 21741 6276
rect 21775 6273 21787 6307
rect 21729 6267 21787 6273
rect 23658 6264 23664 6316
rect 23716 6304 23722 6316
rect 24118 6304 24124 6316
rect 23716 6276 24124 6304
rect 23716 6264 23722 6276
rect 24118 6264 24124 6276
rect 24176 6304 24182 6316
rect 24213 6307 24271 6313
rect 24213 6304 24225 6307
rect 24176 6276 24225 6304
rect 24176 6264 24182 6276
rect 24213 6273 24225 6276
rect 24259 6273 24271 6307
rect 24213 6267 24271 6273
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 20714 6236 20720 6248
rect 19392 6208 20720 6236
rect 19392 6196 19398 6208
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 21542 6236 21548 6248
rect 21503 6208 21548 6236
rect 21542 6196 21548 6208
rect 21600 6196 21606 6248
rect 21634 6196 21640 6248
rect 21692 6236 21698 6248
rect 21818 6236 21824 6248
rect 21692 6208 21824 6236
rect 21692 6196 21698 6208
rect 21818 6196 21824 6208
rect 21876 6196 21882 6248
rect 21910 6196 21916 6248
rect 21968 6236 21974 6248
rect 23017 6239 23075 6245
rect 21968 6208 22692 6236
rect 21968 6196 21974 6208
rect 18417 6131 18475 6137
rect 18524 6140 19288 6168
rect 19429 6171 19487 6177
rect 18524 6112 18552 6140
rect 19429 6137 19441 6171
rect 19475 6168 19487 6171
rect 20073 6171 20131 6177
rect 19475 6140 20024 6168
rect 19475 6137 19487 6140
rect 19429 6131 19487 6137
rect 19996 6112 20024 6140
rect 20073 6137 20085 6171
rect 20119 6168 20131 6171
rect 20254 6168 20260 6180
rect 20119 6140 20260 6168
rect 20119 6137 20131 6140
rect 20073 6131 20131 6137
rect 20254 6128 20260 6140
rect 20312 6128 20318 6180
rect 22281 6171 22339 6177
rect 22281 6137 22293 6171
rect 22327 6168 22339 6171
rect 22370 6168 22376 6180
rect 22327 6140 22376 6168
rect 22327 6137 22339 6140
rect 22281 6131 22339 6137
rect 22370 6128 22376 6140
rect 22428 6128 22434 6180
rect 22664 6177 22692 6208
rect 23017 6205 23029 6239
rect 23063 6236 23075 6239
rect 23106 6236 23112 6248
rect 23063 6208 23112 6236
rect 23063 6205 23075 6208
rect 23017 6199 23075 6205
rect 23106 6196 23112 6208
rect 23164 6236 23170 6248
rect 24670 6236 24676 6248
rect 23164 6208 24676 6236
rect 23164 6196 23170 6208
rect 24670 6196 24676 6208
rect 24728 6196 24734 6248
rect 25130 6196 25136 6248
rect 25188 6236 25194 6248
rect 25225 6239 25283 6245
rect 25225 6236 25237 6239
rect 25188 6208 25237 6236
rect 25188 6196 25194 6208
rect 25225 6205 25237 6208
rect 25271 6205 25283 6239
rect 25225 6199 25283 6205
rect 22649 6171 22707 6177
rect 22649 6137 22661 6171
rect 22695 6168 22707 6171
rect 22738 6168 22744 6180
rect 22695 6140 22744 6168
rect 22695 6137 22707 6140
rect 22649 6131 22707 6137
rect 22738 6128 22744 6140
rect 22796 6128 22802 6180
rect 23477 6171 23535 6177
rect 23477 6137 23489 6171
rect 23523 6168 23535 6171
rect 23842 6168 23848 6180
rect 23523 6140 23848 6168
rect 23523 6137 23535 6140
rect 23477 6131 23535 6137
rect 23842 6128 23848 6140
rect 23900 6168 23906 6180
rect 24029 6171 24087 6177
rect 24029 6168 24041 6171
rect 23900 6140 24041 6168
rect 23900 6128 23906 6140
rect 24029 6137 24041 6140
rect 24075 6137 24087 6171
rect 24029 6131 24087 6137
rect 24121 6171 24179 6177
rect 24121 6137 24133 6171
rect 24167 6168 24179 6171
rect 24302 6168 24308 6180
rect 24167 6140 24308 6168
rect 24167 6137 24179 6140
rect 24121 6131 24179 6137
rect 24302 6128 24308 6140
rect 24360 6128 24366 6180
rect 12805 6103 12863 6109
rect 12805 6100 12817 6103
rect 12584 6072 12817 6100
rect 12584 6060 12590 6072
rect 12805 6069 12817 6072
rect 12851 6069 12863 6103
rect 12805 6063 12863 6069
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14369 6103 14427 6109
rect 14369 6100 14381 6103
rect 13780 6072 14381 6100
rect 13780 6060 13786 6072
rect 14369 6069 14381 6072
rect 14415 6100 14427 6103
rect 14458 6100 14464 6112
rect 14415 6072 14464 6100
rect 14415 6069 14427 6072
rect 14369 6063 14427 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 14700 6072 14933 6100
rect 14700 6060 14706 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 15378 6100 15384 6112
rect 15339 6072 15384 6100
rect 14921 6063 14979 6069
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 17405 6103 17463 6109
rect 17405 6100 17417 6103
rect 17000 6072 17417 6100
rect 17000 6060 17006 6072
rect 17405 6069 17417 6072
rect 17451 6069 17463 6103
rect 18506 6100 18512 6112
rect 18467 6072 18512 6100
rect 17405 6063 17463 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 19518 6060 19524 6112
rect 19576 6100 19582 6112
rect 19613 6103 19671 6109
rect 19613 6100 19625 6103
rect 19576 6072 19625 6100
rect 19576 6060 19582 6072
rect 19613 6069 19625 6072
rect 19659 6069 19671 6103
rect 19978 6100 19984 6112
rect 19939 6072 19984 6100
rect 19613 6063 19671 6069
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 21634 6060 21640 6112
rect 21692 6100 21698 6112
rect 23658 6100 23664 6112
rect 21692 6072 21737 6100
rect 23619 6072 23664 6100
rect 21692 6060 21698 6072
rect 23658 6060 23664 6072
rect 23716 6060 23722 6112
rect 25406 6100 25412 6112
rect 25367 6072 25412 6100
rect 25406 6060 25412 6072
rect 25464 6060 25470 6112
rect 26234 6100 26240 6112
rect 26195 6072 26240 6100
rect 26234 6060 26240 6072
rect 26292 6060 26298 6112
rect 1104 6010 26864 6032
rect 1104 5958 10315 6010
rect 10367 5958 10379 6010
rect 10431 5958 10443 6010
rect 10495 5958 10507 6010
rect 10559 5958 19648 6010
rect 19700 5958 19712 6010
rect 19764 5958 19776 6010
rect 19828 5958 19840 6010
rect 19892 5958 26864 6010
rect 1104 5936 26864 5958
rect 1762 5856 1768 5908
rect 1820 5896 1826 5908
rect 2409 5899 2467 5905
rect 2409 5896 2421 5899
rect 1820 5868 2421 5896
rect 1820 5856 1826 5868
rect 2409 5865 2421 5868
rect 2455 5865 2467 5899
rect 2774 5896 2780 5908
rect 2687 5868 2780 5896
rect 2409 5859 2467 5865
rect 2314 5760 2320 5772
rect 2275 5732 2320 5760
rect 2314 5720 2320 5732
rect 2372 5720 2378 5772
rect 1949 5559 2007 5565
rect 1949 5525 1961 5559
rect 1995 5556 2007 5559
rect 2130 5556 2136 5568
rect 1995 5528 2136 5556
rect 1995 5525 2007 5528
rect 1949 5519 2007 5525
rect 2130 5516 2136 5528
rect 2188 5516 2194 5568
rect 2424 5556 2452 5859
rect 2774 5856 2780 5868
rect 2832 5896 2838 5908
rect 4338 5896 4344 5908
rect 2832 5868 4344 5896
rect 2832 5856 2838 5868
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5166 5896 5172 5908
rect 5127 5868 5172 5896
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 6270 5896 6276 5908
rect 5316 5868 5361 5896
rect 6231 5868 6276 5896
rect 5316 5856 5322 5868
rect 6270 5856 6276 5868
rect 6328 5856 6334 5908
rect 6730 5896 6736 5908
rect 6691 5868 6736 5896
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8202 5896 8208 5908
rect 8163 5868 8208 5896
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 8294 5856 8300 5908
rect 8352 5896 8358 5908
rect 8757 5899 8815 5905
rect 8757 5896 8769 5899
rect 8352 5868 8769 5896
rect 8352 5856 8358 5868
rect 8757 5865 8769 5868
rect 8803 5865 8815 5899
rect 12618 5896 12624 5908
rect 12531 5868 12624 5896
rect 8757 5859 8815 5865
rect 12618 5856 12624 5868
rect 12676 5896 12682 5908
rect 13262 5896 13268 5908
rect 12676 5868 13268 5896
rect 12676 5856 12682 5868
rect 13262 5856 13268 5868
rect 13320 5856 13326 5908
rect 14090 5896 14096 5908
rect 14051 5868 14096 5896
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 15286 5896 15292 5908
rect 15247 5868 15292 5896
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15562 5856 15568 5908
rect 15620 5896 15626 5908
rect 15749 5899 15807 5905
rect 15749 5896 15761 5899
rect 15620 5868 15761 5896
rect 15620 5856 15626 5868
rect 15749 5865 15761 5868
rect 15795 5865 15807 5899
rect 15749 5859 15807 5865
rect 16393 5899 16451 5905
rect 16393 5865 16405 5899
rect 16439 5896 16451 5899
rect 16574 5896 16580 5908
rect 16439 5868 16580 5896
rect 16439 5865 16451 5868
rect 16393 5859 16451 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 16758 5896 16764 5908
rect 16719 5868 16764 5896
rect 16758 5856 16764 5868
rect 16816 5896 16822 5908
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 16816 5868 19349 5896
rect 16816 5856 16822 5868
rect 19337 5865 19349 5868
rect 19383 5896 19395 5899
rect 19426 5896 19432 5908
rect 19383 5868 19432 5896
rect 19383 5865 19395 5868
rect 19337 5859 19395 5865
rect 19426 5856 19432 5868
rect 19484 5856 19490 5908
rect 19518 5856 19524 5908
rect 19576 5896 19582 5908
rect 21358 5896 21364 5908
rect 19576 5868 21364 5896
rect 19576 5856 19582 5868
rect 21358 5856 21364 5868
rect 21416 5856 21422 5908
rect 22278 5896 22284 5908
rect 22239 5868 22284 5896
rect 22278 5856 22284 5868
rect 22336 5856 22342 5908
rect 22922 5896 22928 5908
rect 22883 5868 22928 5896
rect 22922 5856 22928 5868
rect 22980 5856 22986 5908
rect 23658 5856 23664 5908
rect 23716 5896 23722 5908
rect 24397 5899 24455 5905
rect 24397 5896 24409 5899
rect 23716 5868 24409 5896
rect 23716 5856 23722 5868
rect 24397 5865 24409 5868
rect 24443 5896 24455 5899
rect 25409 5899 25467 5905
rect 25409 5896 25421 5899
rect 24443 5868 25421 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 25409 5865 25421 5868
rect 25455 5865 25467 5899
rect 25409 5859 25467 5865
rect 6546 5828 6552 5840
rect 5552 5800 6552 5828
rect 2869 5695 2927 5701
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 2958 5692 2964 5704
rect 2915 5664 2964 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2958 5652 2964 5664
rect 3016 5652 3022 5704
rect 3053 5695 3111 5701
rect 3053 5661 3065 5695
rect 3099 5692 3111 5695
rect 3418 5692 3424 5704
rect 3099 5664 3424 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3418 5652 3424 5664
rect 3476 5692 3482 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3476 5664 3801 5692
rect 3476 5652 3482 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 4246 5692 4252 5704
rect 4207 5664 4252 5692
rect 3789 5655 3847 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 5552 5692 5580 5800
rect 6546 5788 6552 5800
rect 6604 5788 6610 5840
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 7282 5828 7288 5840
rect 7064 5800 7288 5828
rect 7064 5788 7070 5800
rect 7282 5788 7288 5800
rect 7340 5788 7346 5840
rect 9493 5831 9551 5837
rect 9493 5797 9505 5831
rect 9539 5828 9551 5831
rect 10870 5828 10876 5840
rect 9539 5800 10876 5828
rect 9539 5797 9551 5800
rect 9493 5791 9551 5797
rect 10870 5788 10876 5800
rect 10928 5788 10934 5840
rect 14550 5788 14556 5840
rect 14608 5828 14614 5840
rect 15580 5828 15608 5856
rect 14608 5800 15608 5828
rect 14608 5788 14614 5800
rect 17034 5788 17040 5840
rect 17092 5828 17098 5840
rect 17190 5831 17248 5837
rect 17190 5828 17202 5831
rect 17092 5800 17202 5828
rect 17092 5788 17098 5800
rect 17190 5797 17202 5800
rect 17236 5797 17248 5831
rect 18874 5828 18880 5840
rect 18835 5800 18880 5828
rect 17190 5791 17248 5797
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 19058 5788 19064 5840
rect 19116 5828 19122 5840
rect 21542 5828 21548 5840
rect 19116 5800 21548 5828
rect 19116 5788 19122 5800
rect 21542 5788 21548 5800
rect 21600 5788 21606 5840
rect 22830 5828 22836 5840
rect 22791 5800 22836 5828
rect 22830 5788 22836 5800
rect 22888 5788 22894 5840
rect 23198 5788 23204 5840
rect 23256 5828 23262 5840
rect 24489 5831 24547 5837
rect 24489 5828 24501 5831
rect 23256 5800 24501 5828
rect 23256 5788 23262 5800
rect 24489 5797 24501 5800
rect 24535 5828 24547 5831
rect 25041 5831 25099 5837
rect 25041 5828 25053 5831
rect 24535 5800 25053 5828
rect 24535 5797 24547 5800
rect 24489 5791 24547 5797
rect 25041 5797 25053 5800
rect 25087 5797 25099 5831
rect 25774 5828 25780 5840
rect 25735 5800 25780 5828
rect 25041 5791 25099 5797
rect 25774 5788 25780 5800
rect 25832 5788 25838 5840
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 6362 5760 6368 5772
rect 5675 5732 6368 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 6362 5720 6368 5732
rect 6420 5760 6426 5772
rect 6638 5760 6644 5772
rect 6420 5732 6644 5760
rect 6420 5720 6426 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 6914 5720 6920 5772
rect 6972 5760 6978 5772
rect 7092 5763 7150 5769
rect 7092 5760 7104 5763
rect 6972 5732 7104 5760
rect 6972 5720 6978 5732
rect 7092 5729 7104 5732
rect 7138 5760 7150 5763
rect 7138 5732 8248 5760
rect 7138 5729 7150 5732
rect 7092 5723 7150 5729
rect 8220 5704 8248 5732
rect 9766 5720 9772 5772
rect 9824 5760 9830 5772
rect 9933 5763 9991 5769
rect 9933 5760 9945 5763
rect 9824 5732 9945 5760
rect 9824 5720 9830 5732
rect 9933 5729 9945 5732
rect 9979 5729 9991 5763
rect 9933 5723 9991 5729
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 12969 5763 13027 5769
rect 12969 5760 12981 5763
rect 12400 5732 12981 5760
rect 12400 5720 12406 5732
rect 12969 5729 12981 5732
rect 13015 5760 13027 5763
rect 13722 5760 13728 5772
rect 13015 5732 13728 5760
rect 13015 5729 13027 5732
rect 12969 5723 13027 5729
rect 13722 5720 13728 5732
rect 13780 5720 13786 5772
rect 15654 5760 15660 5772
rect 15615 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 19426 5760 19432 5772
rect 19387 5732 19432 5760
rect 19426 5720 19432 5732
rect 19484 5720 19490 5772
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 21269 5763 21327 5769
rect 21269 5760 21281 5763
rect 20772 5732 21281 5760
rect 20772 5720 20778 5732
rect 21269 5729 21281 5732
rect 21315 5760 21327 5763
rect 22186 5760 22192 5772
rect 21315 5732 22192 5760
rect 21315 5729 21327 5732
rect 21269 5723 21327 5729
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 23658 5720 23664 5772
rect 23716 5760 23722 5772
rect 26050 5760 26056 5772
rect 23716 5732 26056 5760
rect 23716 5720 23722 5732
rect 26050 5720 26056 5732
rect 26108 5720 26114 5772
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5500 5664 5733 5692
rect 5500 5652 5506 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5902 5692 5908 5704
rect 5863 5664 5908 5692
rect 5721 5655 5779 5661
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6604 5664 6837 5692
rect 6604 5652 6610 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 9677 5695 9735 5701
rect 9677 5661 9689 5695
rect 9723 5661 9735 5695
rect 9677 5655 9735 5661
rect 4801 5627 4859 5633
rect 4801 5593 4813 5627
rect 4847 5624 4859 5627
rect 5920 5624 5948 5652
rect 4847 5596 6868 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 2590 5556 2596 5568
rect 2424 5528 2596 5556
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 2774 5516 2780 5568
rect 2832 5556 2838 5568
rect 3421 5559 3479 5565
rect 3421 5556 3433 5559
rect 2832 5528 3433 5556
rect 2832 5516 2838 5528
rect 3421 5525 3433 5528
rect 3467 5525 3479 5559
rect 6840 5556 6868 5596
rect 7006 5556 7012 5568
rect 6840 5528 7012 5556
rect 3421 5519 3479 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 9692 5556 9720 5655
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11112 5664 12173 5692
rect 11112 5652 11118 5664
rect 12161 5661 12173 5664
rect 12207 5692 12219 5695
rect 12250 5692 12256 5704
rect 12207 5664 12256 5692
rect 12207 5661 12219 5664
rect 12161 5655 12219 5661
rect 12250 5652 12256 5664
rect 12308 5652 12314 5704
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5661 12771 5695
rect 15102 5692 15108 5704
rect 15063 5664 15108 5692
rect 12713 5655 12771 5661
rect 12526 5624 12532 5636
rect 10612 5596 12532 5624
rect 9950 5556 9956 5568
rect 9692 5528 9956 5556
rect 9950 5516 9956 5528
rect 10008 5556 10014 5568
rect 10612 5556 10640 5596
rect 12526 5584 12532 5596
rect 12584 5624 12590 5636
rect 12728 5624 12756 5655
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16114 5692 16120 5704
rect 15887 5664 16120 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 12584 5596 12756 5624
rect 12584 5584 12590 5596
rect 14826 5584 14832 5636
rect 14884 5624 14890 5636
rect 15856 5624 15884 5655
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16942 5692 16948 5704
rect 16903 5664 16948 5692
rect 16942 5652 16948 5664
rect 17000 5652 17006 5704
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 21416 5664 21465 5692
rect 21416 5652 21422 5664
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 23014 5692 23020 5704
rect 22975 5664 23020 5692
rect 21453 5655 21511 5661
rect 23014 5652 23020 5664
rect 23072 5652 23078 5704
rect 24670 5692 24676 5704
rect 24631 5664 24676 5692
rect 24670 5652 24676 5664
rect 24728 5652 24734 5704
rect 18322 5624 18328 5636
rect 14884 5596 15884 5624
rect 18283 5596 18328 5624
rect 14884 5584 14890 5596
rect 18322 5584 18328 5596
rect 18380 5624 18386 5636
rect 20806 5624 20812 5636
rect 18380 5596 20812 5624
rect 18380 5584 18386 5596
rect 20806 5584 20812 5596
rect 20864 5584 20870 5636
rect 20901 5627 20959 5633
rect 20901 5593 20913 5627
rect 20947 5624 20959 5627
rect 21082 5624 21088 5636
rect 20947 5596 21088 5624
rect 20947 5593 20959 5596
rect 20901 5587 20959 5593
rect 21082 5584 21088 5596
rect 21140 5584 21146 5636
rect 21634 5584 21640 5636
rect 21692 5624 21698 5636
rect 22465 5627 22523 5633
rect 22465 5624 22477 5627
rect 21692 5596 22477 5624
rect 21692 5584 21698 5596
rect 22465 5593 22477 5596
rect 22511 5624 22523 5627
rect 23750 5624 23756 5636
rect 22511 5596 23756 5624
rect 22511 5593 22523 5596
rect 22465 5587 22523 5593
rect 23750 5584 23756 5596
rect 23808 5584 23814 5636
rect 24026 5624 24032 5636
rect 23987 5596 24032 5624
rect 24026 5584 24032 5596
rect 24084 5584 24090 5636
rect 24302 5584 24308 5636
rect 24360 5584 24366 5636
rect 10008 5528 10640 5556
rect 10008 5516 10014 5528
rect 10870 5516 10876 5568
rect 10928 5556 10934 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 10928 5528 11069 5556
rect 10928 5516 10934 5528
rect 11057 5525 11069 5528
rect 11103 5556 11115 5559
rect 11146 5556 11152 5568
rect 11103 5528 11152 5556
rect 11103 5525 11115 5528
rect 11057 5519 11115 5525
rect 11146 5516 11152 5528
rect 11204 5516 11210 5568
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 11790 5556 11796 5568
rect 11747 5528 11796 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 14734 5556 14740 5568
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19613 5559 19671 5565
rect 19613 5556 19625 5559
rect 19392 5528 19625 5556
rect 19392 5516 19398 5528
rect 19613 5525 19625 5528
rect 19659 5525 19671 5559
rect 19613 5519 19671 5525
rect 19886 5516 19892 5568
rect 19944 5556 19950 5568
rect 19981 5559 20039 5565
rect 19981 5556 19993 5559
rect 19944 5528 19993 5556
rect 19944 5516 19950 5528
rect 19981 5525 19993 5528
rect 20027 5525 20039 5559
rect 19981 5519 20039 5525
rect 20254 5516 20260 5568
rect 20312 5556 20318 5568
rect 20717 5559 20775 5565
rect 20717 5556 20729 5559
rect 20312 5528 20729 5556
rect 20312 5516 20318 5528
rect 20717 5525 20729 5528
rect 20763 5556 20775 5559
rect 21174 5556 21180 5568
rect 20763 5528 21180 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 21174 5516 21180 5528
rect 21232 5556 21238 5568
rect 21913 5559 21971 5565
rect 21913 5556 21925 5559
rect 21232 5528 21925 5556
rect 21232 5516 21238 5528
rect 21913 5525 21925 5528
rect 21959 5525 21971 5559
rect 21913 5519 21971 5525
rect 23661 5559 23719 5565
rect 23661 5525 23673 5559
rect 23707 5556 23719 5559
rect 24320 5556 24348 5584
rect 23707 5528 24348 5556
rect 26237 5559 26295 5565
rect 23707 5525 23719 5528
rect 23661 5519 23719 5525
rect 26237 5525 26249 5559
rect 26283 5556 26295 5559
rect 26418 5556 26424 5568
rect 26283 5528 26424 5556
rect 26283 5525 26295 5528
rect 26237 5519 26295 5525
rect 26418 5516 26424 5528
rect 26476 5516 26482 5568
rect 1104 5466 26864 5488
rect 1104 5414 5648 5466
rect 5700 5414 5712 5466
rect 5764 5414 5776 5466
rect 5828 5414 5840 5466
rect 5892 5414 14982 5466
rect 15034 5414 15046 5466
rect 15098 5414 15110 5466
rect 15162 5414 15174 5466
rect 15226 5414 24315 5466
rect 24367 5414 24379 5466
rect 24431 5414 24443 5466
rect 24495 5414 24507 5466
rect 24559 5414 26864 5466
rect 1104 5392 26864 5414
rect 3326 5352 3332 5364
rect 2608 5324 3332 5352
rect 2608 5225 2636 5324
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 5132 5324 5181 5352
rect 5132 5312 5138 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 5169 5315 5227 5321
rect 6273 5355 6331 5361
rect 6273 5321 6285 5355
rect 6319 5352 6331 5355
rect 6822 5352 6828 5364
rect 6319 5324 6828 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7285 5355 7343 5361
rect 7285 5321 7297 5355
rect 7331 5352 7343 5355
rect 8294 5352 8300 5364
rect 7331 5324 8300 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 11054 5352 11060 5364
rect 10459 5324 11060 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 13817 5355 13875 5361
rect 13817 5321 13829 5355
rect 13863 5352 13875 5355
rect 14182 5352 14188 5364
rect 13863 5324 14188 5352
rect 13863 5321 13875 5324
rect 13817 5315 13875 5321
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14608 5324 14933 5352
rect 14608 5312 14614 5324
rect 14921 5321 14933 5324
rect 14967 5321 14979 5355
rect 14921 5315 14979 5321
rect 15289 5355 15347 5361
rect 15289 5321 15301 5355
rect 15335 5352 15347 5355
rect 15654 5352 15660 5364
rect 15335 5324 15660 5352
rect 15335 5321 15347 5324
rect 15289 5315 15347 5321
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 17034 5312 17040 5364
rect 17092 5352 17098 5364
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17092 5324 17785 5352
rect 17092 5312 17098 5324
rect 17773 5321 17785 5324
rect 17819 5321 17831 5355
rect 17773 5315 17831 5321
rect 19613 5355 19671 5361
rect 19613 5321 19625 5355
rect 19659 5352 19671 5355
rect 20714 5352 20720 5364
rect 19659 5324 20720 5352
rect 19659 5321 19671 5324
rect 19613 5315 19671 5321
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 22922 5352 22928 5364
rect 22883 5324 22928 5352
rect 22922 5312 22928 5324
rect 22980 5312 22986 5364
rect 23474 5312 23480 5364
rect 23532 5352 23538 5364
rect 23661 5355 23719 5361
rect 23661 5352 23673 5355
rect 23532 5324 23673 5352
rect 23532 5312 23538 5324
rect 23661 5321 23673 5324
rect 23707 5321 23719 5355
rect 24670 5352 24676 5364
rect 24631 5324 24676 5352
rect 23661 5315 23719 5321
rect 24670 5312 24676 5324
rect 24728 5312 24734 5364
rect 25866 5352 25872 5364
rect 25827 5324 25872 5352
rect 25866 5312 25872 5324
rect 25924 5312 25930 5364
rect 10686 5244 10692 5296
rect 10744 5284 10750 5296
rect 11606 5284 11612 5296
rect 10744 5256 11612 5284
rect 10744 5244 10750 5256
rect 11606 5244 11612 5256
rect 11664 5244 11670 5296
rect 13909 5287 13967 5293
rect 13909 5253 13921 5287
rect 13955 5284 13967 5287
rect 15378 5284 15384 5296
rect 13955 5256 15384 5284
rect 13955 5253 13967 5256
rect 13909 5247 13967 5253
rect 15378 5244 15384 5256
rect 15436 5244 15442 5296
rect 20070 5244 20076 5296
rect 20128 5244 20134 5296
rect 22557 5287 22615 5293
rect 22557 5253 22569 5287
rect 22603 5284 22615 5287
rect 22830 5284 22836 5296
rect 22603 5256 22836 5284
rect 22603 5253 22615 5256
rect 22557 5247 22615 5253
rect 22830 5244 22836 5256
rect 22888 5244 22894 5296
rect 23750 5244 23756 5296
rect 23808 5284 23814 5296
rect 25774 5284 25780 5296
rect 23808 5256 25780 5284
rect 23808 5244 23814 5256
rect 25774 5244 25780 5256
rect 25832 5284 25838 5296
rect 26237 5287 26295 5293
rect 26237 5284 26249 5287
rect 25832 5256 26249 5284
rect 25832 5244 25838 5256
rect 26237 5253 26249 5256
rect 26283 5253 26295 5287
rect 26237 5247 26295 5253
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5216 1823 5219
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 1811 5188 2605 5216
rect 1811 5185 1823 5188
rect 1765 5179 1823 5185
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5442 5216 5448 5228
rect 5123 5188 5448 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5216 5871 5219
rect 6270 5216 6276 5228
rect 5859 5188 6276 5216
rect 5859 5185 5871 5188
rect 5813 5179 5871 5185
rect 6270 5176 6276 5188
rect 6328 5216 6334 5228
rect 6914 5216 6920 5228
rect 6328 5188 6920 5216
rect 6328 5176 6334 5188
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 7064 5188 8309 5216
rect 7064 5176 7070 5188
rect 8297 5185 8309 5188
rect 8343 5216 8355 5219
rect 8757 5219 8815 5225
rect 8757 5216 8769 5219
rect 8343 5188 8769 5216
rect 8343 5185 8355 5188
rect 8297 5179 8355 5185
rect 8757 5185 8769 5188
rect 8803 5185 8815 5219
rect 8757 5179 8815 5185
rect 10870 5176 10876 5228
rect 10928 5216 10934 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10928 5188 10977 5216
rect 10928 5176 10934 5188
rect 10965 5185 10977 5188
rect 11011 5216 11023 5219
rect 11425 5219 11483 5225
rect 11425 5216 11437 5219
rect 11011 5188 11437 5216
rect 11011 5185 11023 5188
rect 10965 5179 11023 5185
rect 11425 5185 11437 5188
rect 11471 5185 11483 5219
rect 11425 5179 11483 5185
rect 14553 5219 14611 5225
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 18598 5216 18604 5228
rect 14599 5188 15148 5216
rect 18559 5188 18604 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 3786 5108 3792 5160
rect 3844 5148 3850 5160
rect 4062 5148 4068 5160
rect 3844 5120 4068 5148
rect 3844 5108 3850 5120
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4706 5148 4712 5160
rect 4667 5120 4712 5148
rect 4706 5108 4712 5120
rect 4764 5108 4770 5160
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5148 5687 5151
rect 6086 5148 6092 5160
rect 5675 5120 6092 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 6086 5108 6092 5120
rect 6144 5108 6150 5160
rect 6546 5108 6552 5160
rect 6604 5148 6610 5160
rect 9125 5151 9183 5157
rect 9125 5148 9137 5151
rect 6604 5120 9137 5148
rect 6604 5108 6610 5120
rect 9125 5117 9137 5120
rect 9171 5117 9183 5151
rect 9306 5148 9312 5160
rect 9267 5120 9312 5148
rect 9125 5111 9183 5117
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 10321 5151 10379 5157
rect 10321 5148 10333 5151
rect 10192 5120 10333 5148
rect 10192 5108 10198 5120
rect 10321 5117 10333 5120
rect 10367 5148 10379 5151
rect 10367 5120 10916 5148
rect 10367 5117 10379 5120
rect 10321 5111 10379 5117
rect 750 5040 756 5092
rect 808 5080 814 5092
rect 2133 5083 2191 5089
rect 2133 5080 2145 5083
rect 808 5052 2145 5080
rect 808 5040 814 5052
rect 2133 5049 2145 5052
rect 2179 5080 2191 5083
rect 2682 5080 2688 5092
rect 2179 5052 2688 5080
rect 2179 5049 2191 5052
rect 2133 5043 2191 5049
rect 2682 5040 2688 5052
rect 2740 5040 2746 5092
rect 2860 5083 2918 5089
rect 2860 5049 2872 5083
rect 2906 5080 2918 5083
rect 3234 5080 3240 5092
rect 2906 5052 3240 5080
rect 2906 5049 2918 5052
rect 2860 5043 2918 5049
rect 3234 5040 3240 5052
rect 3292 5040 3298 5092
rect 5537 5083 5595 5089
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 7653 5083 7711 5089
rect 5583 5052 7328 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 2406 5012 2412 5024
rect 2367 4984 2412 5012
rect 2406 4972 2412 4984
rect 2464 5012 2470 5024
rect 2958 5012 2964 5024
rect 2464 4984 2964 5012
rect 2464 4972 2470 4984
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 3786 4972 3792 5024
rect 3844 5012 3850 5024
rect 3973 5015 4031 5021
rect 3973 5012 3985 5015
rect 3844 4984 3985 5012
rect 3844 4972 3850 4984
rect 3973 4981 3985 4984
rect 4019 4981 4031 5015
rect 6546 5012 6552 5024
rect 6507 4984 6552 5012
rect 3973 4975 4031 4981
rect 6546 4972 6552 4984
rect 6604 4972 6610 5024
rect 7300 5012 7328 5052
rect 7653 5049 7665 5083
rect 7699 5080 7711 5083
rect 8110 5080 8116 5092
rect 7699 5052 8116 5080
rect 7699 5049 7711 5052
rect 7653 5043 7711 5049
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 10888 5089 10916 5120
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 11882 5148 11888 5160
rect 11664 5120 11888 5148
rect 11664 5108 11670 5120
rect 11882 5108 11888 5120
rect 11940 5108 11946 5160
rect 12805 5151 12863 5157
rect 12805 5117 12817 5151
rect 12851 5148 12863 5151
rect 13170 5148 13176 5160
rect 12851 5120 13176 5148
rect 12851 5117 12863 5120
rect 12805 5111 12863 5117
rect 13170 5108 13176 5120
rect 13228 5108 13234 5160
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14277 5151 14335 5157
rect 14277 5148 14289 5151
rect 14240 5120 14289 5148
rect 14240 5108 14246 5120
rect 14277 5117 14289 5120
rect 14323 5117 14335 5151
rect 14277 5111 14335 5117
rect 15120 5092 15148 5188
rect 18598 5176 18604 5188
rect 18656 5216 18662 5228
rect 18966 5216 18972 5228
rect 18656 5188 18972 5216
rect 18656 5176 18662 5188
rect 18966 5176 18972 5188
rect 19024 5216 19030 5228
rect 19886 5216 19892 5228
rect 19024 5188 19892 5216
rect 19024 5176 19030 5188
rect 19886 5176 19892 5188
rect 19944 5216 19950 5228
rect 20088 5216 20116 5244
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19944 5188 20177 5216
rect 19944 5176 19950 5188
rect 20165 5185 20177 5188
rect 20211 5216 20223 5219
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20211 5188 20637 5216
rect 20211 5185 20223 5188
rect 20165 5179 20223 5185
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 21729 5219 21787 5225
rect 21729 5216 21741 5219
rect 21048 5188 21741 5216
rect 21048 5176 21054 5188
rect 21729 5185 21741 5188
rect 21775 5185 21787 5219
rect 21729 5179 21787 5185
rect 22462 5176 22468 5228
rect 22520 5216 22526 5228
rect 23198 5216 23204 5228
rect 22520 5188 23204 5216
rect 22520 5176 22526 5188
rect 23198 5176 23204 5188
rect 23256 5176 23262 5228
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24213 5219 24271 5225
rect 24213 5216 24225 5219
rect 24176 5188 24225 5216
rect 24176 5176 24182 5188
rect 24213 5185 24225 5188
rect 24259 5185 24271 5219
rect 24213 5179 24271 5185
rect 15473 5151 15531 5157
rect 15473 5117 15485 5151
rect 15519 5148 15531 5151
rect 15562 5148 15568 5160
rect 15519 5120 15568 5148
rect 15519 5117 15531 5120
rect 15473 5111 15531 5117
rect 15562 5108 15568 5120
rect 15620 5148 15626 5160
rect 16942 5148 16948 5160
rect 15620 5120 16948 5148
rect 15620 5108 15626 5120
rect 16942 5108 16948 5120
rect 17000 5148 17006 5160
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 17000 5120 17417 5148
rect 17000 5108 17006 5120
rect 17405 5117 17417 5120
rect 17451 5117 17463 5151
rect 17405 5111 17463 5117
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 20073 5151 20131 5157
rect 20073 5148 20085 5151
rect 19567 5120 20085 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 20073 5117 20085 5120
rect 20119 5148 20131 5151
rect 20530 5148 20536 5160
rect 20119 5120 20536 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 20530 5108 20536 5120
rect 20588 5108 20594 5160
rect 21082 5108 21088 5160
rect 21140 5148 21146 5160
rect 21545 5151 21603 5157
rect 21545 5148 21557 5151
rect 21140 5120 21557 5148
rect 21140 5108 21146 5120
rect 21545 5117 21557 5120
rect 21591 5117 21603 5151
rect 24026 5148 24032 5160
rect 23987 5120 24032 5148
rect 21545 5111 21603 5117
rect 24026 5108 24032 5120
rect 24084 5108 24090 5160
rect 25225 5151 25283 5157
rect 25225 5117 25237 5151
rect 25271 5148 25283 5151
rect 25866 5148 25872 5160
rect 25271 5120 25872 5148
rect 25271 5117 25283 5120
rect 25225 5111 25283 5117
rect 25866 5108 25872 5120
rect 25924 5108 25930 5160
rect 9953 5083 10011 5089
rect 9953 5049 9965 5083
rect 9999 5080 10011 5083
rect 10873 5083 10931 5089
rect 9999 5052 10824 5080
rect 9999 5049 10011 5052
rect 9953 5043 10011 5049
rect 10796 5024 10824 5052
rect 10873 5049 10885 5083
rect 10919 5080 10931 5083
rect 10962 5080 10968 5092
rect 10919 5052 10968 5080
rect 10919 5049 10931 5052
rect 10873 5043 10931 5049
rect 10962 5040 10968 5052
rect 11020 5040 11026 5092
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 13449 5083 13507 5089
rect 13449 5080 13461 5083
rect 13136 5052 13461 5080
rect 13136 5040 13142 5052
rect 13449 5049 13461 5052
rect 13495 5080 13507 5083
rect 13495 5052 14412 5080
rect 13495 5049 13507 5052
rect 13449 5043 13507 5049
rect 7745 5015 7803 5021
rect 7745 5012 7757 5015
rect 7300 4984 7757 5012
rect 7745 4981 7757 4984
rect 7791 5012 7803 5015
rect 8018 5012 8024 5024
rect 7791 4984 8024 5012
rect 7791 4981 7803 4984
rect 7745 4975 7803 4981
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8205 5015 8263 5021
rect 8205 4981 8217 5015
rect 8251 5012 8263 5015
rect 8294 5012 8300 5024
rect 8251 4984 8300 5012
rect 8251 4981 8263 4984
rect 8205 4975 8263 4981
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 9122 5012 9128 5024
rect 8352 4984 9128 5012
rect 8352 4972 8358 4984
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 10778 5012 10784 5024
rect 10739 4984 10784 5012
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11882 5012 11888 5024
rect 11843 4984 11888 5012
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12584 4984 12633 5012
rect 12584 4972 12590 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13262 5012 13268 5024
rect 13035 4984 13268 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13262 4972 13268 4984
rect 13320 4972 13326 5024
rect 14384 5021 14412 5052
rect 15102 5040 15108 5092
rect 15160 5080 15166 5092
rect 15740 5083 15798 5089
rect 15740 5080 15752 5083
rect 15160 5052 15752 5080
rect 15160 5040 15166 5052
rect 15740 5049 15752 5052
rect 15786 5080 15798 5083
rect 16574 5080 16580 5092
rect 15786 5052 16580 5080
rect 15786 5049 15798 5052
rect 15740 5043 15798 5049
rect 16574 5040 16580 5052
rect 16632 5080 16638 5092
rect 17494 5080 17500 5092
rect 16632 5052 17500 5080
rect 16632 5040 16638 5052
rect 17494 5040 17500 5052
rect 17552 5040 17558 5092
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 21634 5080 21640 5092
rect 20772 5052 21640 5080
rect 20772 5040 20778 5052
rect 21634 5040 21640 5052
rect 21692 5040 21698 5092
rect 22370 5040 22376 5092
rect 22428 5080 22434 5092
rect 26326 5080 26332 5092
rect 22428 5052 26332 5080
rect 22428 5040 22434 5052
rect 26326 5040 26332 5052
rect 26384 5040 26390 5092
rect 14369 5015 14427 5021
rect 14369 4981 14381 5015
rect 14415 5012 14427 5015
rect 14458 5012 14464 5024
rect 14415 4984 14464 5012
rect 14415 4981 14427 4984
rect 14369 4975 14427 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 16853 5015 16911 5021
rect 16853 5012 16865 5015
rect 16816 4984 16865 5012
rect 16816 4972 16822 4984
rect 16853 4981 16865 4984
rect 16899 4981 16911 5015
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 16853 4975 16911 4981
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 18414 5012 18420 5024
rect 18375 4984 18420 5012
rect 18414 4972 18420 4984
rect 18472 4972 18478 5024
rect 18506 4972 18512 5024
rect 18564 5012 18570 5024
rect 19058 5012 19064 5024
rect 18564 4984 18609 5012
rect 19019 4984 19064 5012
rect 18564 4972 18570 4984
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19576 4984 19993 5012
rect 19576 4972 19582 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 20990 5012 20996 5024
rect 20951 4984 20996 5012
rect 19981 4975 20039 4981
rect 20990 4972 20996 4984
rect 21048 4972 21054 5024
rect 21174 5012 21180 5024
rect 21135 4984 21180 5012
rect 21174 4972 21180 4984
rect 21232 4972 21238 5024
rect 22002 4972 22008 5024
rect 22060 5012 22066 5024
rect 23477 5015 23535 5021
rect 23477 5012 23489 5015
rect 22060 4984 23489 5012
rect 22060 4972 22066 4984
rect 23477 4981 23489 4984
rect 23523 5012 23535 5015
rect 24121 5015 24179 5021
rect 24121 5012 24133 5015
rect 23523 4984 24133 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 24121 4981 24133 4984
rect 24167 4981 24179 5015
rect 25038 5012 25044 5024
rect 24999 4984 25044 5012
rect 24121 4975 24179 4981
rect 25038 4972 25044 4984
rect 25096 4972 25102 5024
rect 25130 4972 25136 5024
rect 25188 5012 25194 5024
rect 25409 5015 25467 5021
rect 25409 5012 25421 5015
rect 25188 4984 25421 5012
rect 25188 4972 25194 4984
rect 25409 4981 25421 4984
rect 25455 4981 25467 5015
rect 25409 4975 25467 4981
rect 1104 4922 26864 4944
rect 1104 4870 10315 4922
rect 10367 4870 10379 4922
rect 10431 4870 10443 4922
rect 10495 4870 10507 4922
rect 10559 4870 19648 4922
rect 19700 4870 19712 4922
rect 19764 4870 19776 4922
rect 19828 4870 19840 4922
rect 19892 4870 26864 4922
rect 1104 4848 26864 4870
rect 1946 4808 1952 4820
rect 1907 4780 1952 4808
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2682 4808 2688 4820
rect 2455 4780 2688 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3234 4808 3240 4820
rect 3147 4780 3240 4808
rect 3234 4768 3240 4780
rect 3292 4808 3298 4820
rect 3513 4811 3571 4817
rect 3513 4808 3525 4811
rect 3292 4780 3525 4808
rect 3292 4768 3298 4780
rect 3513 4777 3525 4780
rect 3559 4808 3571 4811
rect 5166 4808 5172 4820
rect 3559 4780 5172 4808
rect 3559 4777 3571 4780
rect 3513 4771 3571 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 8570 4808 8576 4820
rect 8531 4780 8576 4808
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10229 4811 10287 4817
rect 10229 4808 10241 4811
rect 9732 4780 10241 4808
rect 9732 4768 9738 4780
rect 10229 4777 10241 4780
rect 10275 4777 10287 4811
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 10229 4771 10287 4777
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 12342 4768 12348 4820
rect 12400 4808 12406 4820
rect 12618 4808 12624 4820
rect 12400 4780 12624 4808
rect 12400 4768 12406 4780
rect 12618 4768 12624 4780
rect 12676 4768 12682 4820
rect 14093 4811 14151 4817
rect 14093 4777 14105 4811
rect 14139 4808 14151 4811
rect 14274 4808 14280 4820
rect 14139 4780 14280 4808
rect 14139 4777 14151 4780
rect 14093 4771 14151 4777
rect 14274 4768 14280 4780
rect 14332 4768 14338 4820
rect 14826 4768 14832 4820
rect 14884 4808 14890 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 14884 4780 15025 4808
rect 14884 4768 14890 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15013 4771 15071 4777
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 15657 4811 15715 4817
rect 15657 4808 15669 4811
rect 15436 4780 15669 4808
rect 15436 4768 15442 4780
rect 15657 4777 15669 4780
rect 15703 4777 15715 4811
rect 15657 4771 15715 4777
rect 16574 4768 16580 4820
rect 16632 4808 16638 4820
rect 16853 4811 16911 4817
rect 16853 4808 16865 4811
rect 16632 4780 16865 4808
rect 16632 4768 16638 4780
rect 16853 4777 16865 4780
rect 16899 4777 16911 4811
rect 18138 4808 18144 4820
rect 18099 4780 18144 4808
rect 16853 4771 16911 4777
rect 18138 4768 18144 4780
rect 18196 4808 18202 4820
rect 18322 4808 18328 4820
rect 18196 4780 18328 4808
rect 18196 4768 18202 4780
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18417 4811 18475 4817
rect 18417 4777 18429 4811
rect 18463 4777 18475 4811
rect 18417 4771 18475 4777
rect 1397 4675 1455 4681
rect 1397 4641 1409 4675
rect 1443 4672 1455 4675
rect 1964 4672 1992 4768
rect 3786 4700 3792 4752
rect 3844 4740 3850 4752
rect 4310 4743 4368 4749
rect 4310 4740 4322 4743
rect 3844 4712 4322 4740
rect 3844 4700 3850 4712
rect 4310 4709 4322 4712
rect 4356 4709 4368 4743
rect 4310 4703 4368 4709
rect 9766 4700 9772 4752
rect 9824 4740 9830 4752
rect 9950 4740 9956 4752
rect 9824 4712 9956 4740
rect 9824 4700 9830 4712
rect 9950 4700 9956 4712
rect 10008 4700 10014 4752
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 14737 4743 14795 4749
rect 11480 4712 12296 4740
rect 11480 4700 11486 4712
rect 1443 4644 1992 4672
rect 2777 4675 2835 4681
rect 1443 4641 1455 4644
rect 1397 4635 1455 4641
rect 2777 4641 2789 4675
rect 2823 4672 2835 4675
rect 3970 4672 3976 4684
rect 2823 4644 3976 4672
rect 2823 4641 2835 4644
rect 2777 4635 2835 4641
rect 3970 4632 3976 4644
rect 4028 4632 4034 4684
rect 6822 4681 6828 4684
rect 6457 4675 6515 4681
rect 6457 4641 6469 4675
rect 6503 4672 6515 4675
rect 6816 4672 6828 4681
rect 6503 4644 6828 4672
rect 6503 4641 6515 4644
rect 6457 4635 6515 4641
rect 6816 4635 6828 4644
rect 3050 4604 3056 4616
rect 2963 4576 3056 4604
rect 3050 4564 3056 4576
rect 3108 4604 3114 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3108 4576 3249 4604
rect 3108 4564 3114 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 3384 4576 4077 4604
rect 3384 4564 3390 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 1578 4536 1584 4548
rect 1539 4508 1584 4536
rect 1578 4496 1584 4508
rect 1636 4496 1642 4548
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 3418 4468 3424 4480
rect 2363 4440 3424 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 3786 4468 3792 4480
rect 3747 4440 3792 4468
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 4080 4468 4108 4567
rect 5445 4539 5503 4545
rect 5445 4505 5457 4539
rect 5491 4536 5503 4539
rect 6472 4536 6500 4635
rect 6822 4632 6828 4635
rect 6880 4632 6886 4684
rect 10594 4672 10600 4684
rect 10555 4644 10600 4672
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 12268 4681 12296 4712
rect 14737 4709 14749 4743
rect 14783 4740 14795 4743
rect 15102 4740 15108 4752
rect 14783 4712 15108 4740
rect 14783 4709 14795 4712
rect 14737 4703 14795 4709
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11440 4644 12173 4672
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6604 4576 6649 4604
rect 6604 4564 6610 4576
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10134 4604 10140 4616
rect 9824 4576 10140 4604
rect 9824 4564 9830 4576
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10686 4604 10692 4616
rect 10647 4576 10692 4604
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10778 4564 10784 4616
rect 10836 4604 10842 4616
rect 10836 4576 10881 4604
rect 10836 4564 10842 4576
rect 11440 4548 11468 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 12253 4675 12311 4681
rect 12253 4641 12265 4675
rect 12299 4672 12311 4675
rect 12710 4672 12716 4684
rect 12299 4644 12716 4672
rect 12299 4641 12311 4644
rect 12253 4635 12311 4641
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 13998 4672 14004 4684
rect 13959 4644 14004 4672
rect 13998 4632 14004 4644
rect 14056 4632 14062 4684
rect 12342 4604 12348 4616
rect 12303 4576 12348 4604
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 13170 4604 13176 4616
rect 13131 4576 13176 4604
rect 13170 4564 13176 4576
rect 13228 4564 13234 4616
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4604 14335 4607
rect 14752 4604 14780 4703
rect 15102 4700 15108 4712
rect 15160 4700 15166 4752
rect 15286 4700 15292 4752
rect 15344 4740 15350 4752
rect 15749 4743 15807 4749
rect 15749 4740 15761 4743
rect 15344 4712 15761 4740
rect 15344 4700 15350 4712
rect 15749 4709 15761 4712
rect 15795 4740 15807 4743
rect 18432 4740 18460 4771
rect 18690 4768 18696 4820
rect 18748 4808 18754 4820
rect 18785 4811 18843 4817
rect 18785 4808 18797 4811
rect 18748 4780 18797 4808
rect 18748 4768 18754 4780
rect 18785 4777 18797 4780
rect 18831 4777 18843 4811
rect 18785 4771 18843 4777
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 18932 4780 18977 4808
rect 18932 4768 18938 4780
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 19613 4811 19671 4817
rect 19613 4808 19625 4811
rect 19576 4780 19625 4808
rect 19576 4768 19582 4780
rect 19613 4777 19625 4780
rect 19659 4777 19671 4811
rect 20070 4808 20076 4820
rect 20031 4780 20076 4808
rect 19613 4771 19671 4777
rect 20070 4768 20076 4780
rect 20128 4808 20134 4820
rect 20349 4811 20407 4817
rect 20349 4808 20361 4811
rect 20128 4780 20361 4808
rect 20128 4768 20134 4780
rect 20349 4777 20361 4780
rect 20395 4777 20407 4811
rect 20349 4771 20407 4777
rect 22373 4811 22431 4817
rect 22373 4777 22385 4811
rect 22419 4808 22431 4811
rect 23014 4808 23020 4820
rect 22419 4780 23020 4808
rect 22419 4777 22431 4780
rect 22373 4771 22431 4777
rect 23014 4768 23020 4780
rect 23072 4768 23078 4820
rect 23753 4811 23811 4817
rect 23753 4777 23765 4811
rect 23799 4808 23811 4811
rect 24026 4808 24032 4820
rect 23799 4780 24032 4808
rect 23799 4777 23811 4780
rect 23753 4771 23811 4777
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 24118 4768 24124 4820
rect 24176 4808 24182 4820
rect 24176 4780 24221 4808
rect 24176 4768 24182 4780
rect 15795 4712 18460 4740
rect 15795 4709 15807 4712
rect 15749 4703 15807 4709
rect 21358 4700 21364 4752
rect 21416 4740 21422 4752
rect 21821 4743 21879 4749
rect 21821 4740 21833 4743
rect 21416 4712 21833 4740
rect 21416 4700 21422 4712
rect 21821 4709 21833 4712
rect 21867 4740 21879 4743
rect 21913 4743 21971 4749
rect 21913 4740 21925 4743
rect 21867 4712 21925 4740
rect 21867 4709 21879 4712
rect 21821 4703 21879 4709
rect 21913 4709 21925 4712
rect 21959 4709 21971 4743
rect 21913 4703 21971 4709
rect 16758 4672 16764 4684
rect 15948 4644 16764 4672
rect 15948 4613 15976 4644
rect 16758 4632 16764 4644
rect 16816 4632 16822 4684
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17221 4675 17279 4681
rect 17221 4672 17233 4675
rect 17092 4644 17233 4672
rect 17092 4632 17098 4644
rect 17221 4641 17233 4644
rect 17267 4641 17279 4675
rect 17221 4635 17279 4641
rect 21269 4675 21327 4681
rect 21269 4641 21281 4675
rect 21315 4672 21327 4675
rect 22830 4672 22836 4684
rect 21315 4644 21956 4672
rect 22791 4644 22836 4672
rect 21315 4641 21327 4644
rect 21269 4635 21327 4641
rect 21928 4616 21956 4644
rect 22830 4632 22836 4644
rect 22888 4632 22894 4684
rect 22922 4632 22928 4684
rect 22980 4672 22986 4684
rect 24486 4672 24492 4684
rect 22980 4644 23152 4672
rect 24447 4644 24492 4672
rect 22980 4632 22986 4644
rect 14323 4576 14780 4604
rect 15933 4607 15991 4613
rect 14323 4573 14335 4576
rect 14277 4567 14335 4573
rect 15933 4573 15945 4607
rect 15979 4573 15991 4607
rect 15933 4567 15991 4573
rect 5491 4508 6500 4536
rect 5491 4505 5503 4508
rect 5445 4499 5503 4505
rect 11146 4496 11152 4548
rect 11204 4536 11210 4548
rect 11422 4536 11428 4548
rect 11204 4508 11428 4536
rect 11204 4496 11210 4508
rect 11422 4496 11428 4508
rect 11480 4496 11486 4548
rect 12897 4539 12955 4545
rect 12897 4505 12909 4539
rect 12943 4536 12955 4539
rect 13722 4536 13728 4548
rect 12943 4508 13728 4536
rect 12943 4505 12955 4508
rect 12897 4499 12955 4505
rect 13722 4496 13728 4508
rect 13780 4536 13786 4548
rect 14292 4536 14320 4567
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17310 4604 17316 4616
rect 17000 4576 17316 4604
rect 17000 4564 17006 4576
rect 17310 4564 17316 4576
rect 17368 4564 17374 4616
rect 17494 4604 17500 4616
rect 17455 4576 17500 4604
rect 17494 4564 17500 4576
rect 17552 4564 17558 4616
rect 18969 4607 19027 4613
rect 18969 4573 18981 4607
rect 19015 4573 19027 4607
rect 18969 4567 19027 4573
rect 13780 4508 14320 4536
rect 17512 4536 17540 4564
rect 18984 4536 19012 4567
rect 20898 4564 20904 4616
rect 20956 4604 20962 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 20956 4576 21373 4604
rect 20956 4564 20962 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21542 4604 21548 4616
rect 21503 4576 21548 4604
rect 21361 4567 21419 4573
rect 21542 4564 21548 4576
rect 21600 4564 21606 4616
rect 21910 4564 21916 4616
rect 21968 4564 21974 4616
rect 23014 4604 23020 4616
rect 22975 4576 23020 4604
rect 23014 4564 23020 4576
rect 23072 4564 23078 4616
rect 23124 4604 23152 4644
rect 24486 4632 24492 4644
rect 24544 4632 24550 4684
rect 25409 4607 25467 4613
rect 25409 4604 25421 4607
rect 23124 4576 25421 4604
rect 25409 4573 25421 4576
rect 25455 4573 25467 4607
rect 25774 4604 25780 4616
rect 25735 4576 25780 4604
rect 25409 4567 25467 4573
rect 25774 4564 25780 4576
rect 25832 4564 25838 4616
rect 19426 4536 19432 4548
rect 17512 4508 19432 4536
rect 13780 4496 13786 4508
rect 19426 4496 19432 4508
rect 19484 4496 19490 4548
rect 20530 4496 20536 4548
rect 20588 4536 20594 4548
rect 23106 4536 23112 4548
rect 20588 4508 23112 4536
rect 20588 4496 20594 4508
rect 23106 4496 23112 4508
rect 23164 4496 23170 4548
rect 4338 4468 4344 4480
rect 4080 4440 4344 4468
rect 4338 4428 4344 4440
rect 4396 4428 4402 4480
rect 5994 4428 6000 4480
rect 6052 4468 6058 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 6052 4440 6101 4468
rect 6052 4428 6058 4440
rect 6089 4437 6101 4440
rect 6135 4468 6147 4471
rect 6730 4468 6736 4480
rect 6135 4440 6736 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7926 4468 7932 4480
rect 7887 4440 7932 4468
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8938 4468 8944 4480
rect 8899 4440 8944 4468
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9122 4428 9128 4480
rect 9180 4468 9186 4480
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 9180 4440 9321 4468
rect 9180 4428 9186 4440
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 9309 4431 9367 4437
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 11112 4440 11253 4468
rect 11112 4428 11118 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11698 4468 11704 4480
rect 11659 4440 11704 4468
rect 11241 4431 11299 4437
rect 11698 4428 11704 4440
rect 11756 4428 11762 4480
rect 13630 4468 13636 4480
rect 13591 4440 13636 4468
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 15286 4468 15292 4480
rect 15247 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15562 4428 15568 4480
rect 15620 4468 15626 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 15620 4440 16313 4468
rect 15620 4428 15626 4440
rect 16301 4437 16313 4440
rect 16347 4437 16359 4471
rect 16301 4431 16359 4437
rect 20901 4471 20959 4477
rect 20901 4437 20913 4471
rect 20947 4468 20959 4471
rect 20990 4468 20996 4480
rect 20947 4440 20996 4468
rect 20947 4437 20959 4440
rect 20901 4431 20959 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21821 4471 21879 4477
rect 21821 4437 21833 4471
rect 21867 4468 21879 4471
rect 22094 4468 22100 4480
rect 21867 4440 22100 4468
rect 21867 4437 21879 4440
rect 21821 4431 21879 4437
rect 22094 4428 22100 4440
rect 22152 4428 22158 4480
rect 22465 4471 22523 4477
rect 22465 4437 22477 4471
rect 22511 4468 22523 4471
rect 23566 4468 23572 4480
rect 22511 4440 23572 4468
rect 22511 4437 22523 4440
rect 22465 4431 22523 4437
rect 23566 4428 23572 4440
rect 23624 4428 23630 4480
rect 24670 4468 24676 4480
rect 24631 4440 24676 4468
rect 24670 4428 24676 4440
rect 24728 4428 24734 4480
rect 24762 4428 24768 4480
rect 24820 4468 24826 4480
rect 25041 4471 25099 4477
rect 25041 4468 25053 4471
rect 24820 4440 25053 4468
rect 24820 4428 24826 4440
rect 25041 4437 25053 4440
rect 25087 4437 25099 4471
rect 26234 4468 26240 4480
rect 26195 4440 26240 4468
rect 25041 4431 25099 4437
rect 26234 4428 26240 4440
rect 26292 4428 26298 4480
rect 1104 4378 26864 4400
rect 1104 4326 5648 4378
rect 5700 4326 5712 4378
rect 5764 4326 5776 4378
rect 5828 4326 5840 4378
rect 5892 4326 14982 4378
rect 15034 4326 15046 4378
rect 15098 4326 15110 4378
rect 15162 4326 15174 4378
rect 15226 4326 24315 4378
rect 24367 4326 24379 4378
rect 24431 4326 24443 4378
rect 24495 4326 24507 4378
rect 24559 4326 26864 4378
rect 1104 4304 26864 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 3329 4267 3387 4273
rect 3329 4264 3341 4267
rect 2924 4236 3341 4264
rect 2924 4224 2930 4236
rect 3329 4233 3341 4236
rect 3375 4233 3387 4267
rect 3329 4227 3387 4233
rect 4062 4224 4068 4276
rect 4120 4224 4126 4276
rect 4338 4264 4344 4276
rect 4299 4236 4344 4264
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 10686 4264 10692 4276
rect 10647 4236 10692 4264
rect 10686 4224 10692 4236
rect 10744 4224 10750 4276
rect 11241 4267 11299 4273
rect 11241 4233 11253 4267
rect 11287 4264 11299 4267
rect 11422 4264 11428 4276
rect 11287 4236 11428 4264
rect 11287 4233 11299 4236
rect 11241 4227 11299 4233
rect 11422 4224 11428 4236
rect 11480 4264 11486 4276
rect 11480 4236 11928 4264
rect 11480 4224 11486 4236
rect 3786 4196 3792 4208
rect 2424 4168 3792 4196
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2424 4137 2452 4168
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 2409 4131 2467 4137
rect 2409 4128 2421 4131
rect 2372 4100 2421 4128
rect 2372 4088 2378 4100
rect 2409 4097 2421 4100
rect 2455 4097 2467 4131
rect 2409 4091 2467 4097
rect 3418 4088 3424 4140
rect 3476 4128 3482 4140
rect 3881 4131 3939 4137
rect 3881 4128 3893 4131
rect 3476 4100 3893 4128
rect 3476 4088 3482 4100
rect 3881 4097 3893 4100
rect 3927 4097 3939 4131
rect 4080 4128 4108 4224
rect 11900 4208 11928 4236
rect 12342 4224 12348 4276
rect 12400 4264 12406 4276
rect 18506 4264 18512 4276
rect 12400 4236 18512 4264
rect 12400 4224 12406 4236
rect 18506 4224 18512 4236
rect 18564 4224 18570 4276
rect 18690 4224 18696 4276
rect 18748 4264 18754 4276
rect 19061 4267 19119 4273
rect 19061 4264 19073 4267
rect 18748 4236 19073 4264
rect 18748 4224 18754 4236
rect 19061 4233 19073 4236
rect 19107 4233 19119 4267
rect 19061 4227 19119 4233
rect 20990 4224 20996 4276
rect 21048 4264 21054 4276
rect 22922 4264 22928 4276
rect 21048 4236 22928 4264
rect 21048 4224 21054 4236
rect 22922 4224 22928 4236
rect 22980 4224 22986 4276
rect 24118 4224 24124 4276
rect 24176 4264 24182 4276
rect 24673 4267 24731 4273
rect 24673 4264 24685 4267
rect 24176 4236 24685 4264
rect 24176 4224 24182 4236
rect 24673 4233 24685 4236
rect 24719 4233 24731 4267
rect 24673 4227 24731 4233
rect 4617 4199 4675 4205
rect 4617 4165 4629 4199
rect 4663 4196 4675 4199
rect 4893 4199 4951 4205
rect 4893 4196 4905 4199
rect 4663 4168 4905 4196
rect 4663 4165 4675 4168
rect 4617 4159 4675 4165
rect 4893 4165 4905 4168
rect 4939 4165 4951 4199
rect 5994 4196 6000 4208
rect 4893 4159 4951 4165
rect 5460 4168 6000 4196
rect 5460 4140 5488 4168
rect 5994 4156 6000 4168
rect 6052 4156 6058 4208
rect 9122 4156 9128 4208
rect 9180 4196 9186 4208
rect 9180 4168 9904 4196
rect 9180 4156 9186 4168
rect 5166 4128 5172 4140
rect 4080 4100 5172 4128
rect 3881 4091 3939 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5442 4128 5448 4140
rect 5355 4100 5448 4128
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 8662 4088 8668 4140
rect 8720 4128 8726 4140
rect 9876 4137 9904 4168
rect 11882 4156 11888 4208
rect 11940 4156 11946 4208
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 14182 4196 14188 4208
rect 13688 4168 13768 4196
rect 14143 4168 14188 4196
rect 13688 4156 13694 4168
rect 9769 4131 9827 4137
rect 9769 4128 9781 4131
rect 8720 4100 9781 4128
rect 8720 4088 8726 4100
rect 9769 4097 9781 4100
rect 9815 4097 9827 4131
rect 9769 4091 9827 4097
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 11296 4100 12265 4128
rect 11296 4088 11302 4100
rect 12253 4097 12265 4100
rect 12299 4128 12311 4131
rect 13357 4131 13415 4137
rect 12299 4100 13124 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 13096 4072 13124 4100
rect 13357 4097 13369 4131
rect 13403 4097 13415 4131
rect 13740 4128 13768 4168
rect 14182 4156 14188 4168
rect 14240 4156 14246 4208
rect 15841 4199 15899 4205
rect 15841 4165 15853 4199
rect 15887 4196 15899 4199
rect 15930 4196 15936 4208
rect 15887 4168 15936 4196
rect 15887 4165 15899 4168
rect 15841 4159 15899 4165
rect 15930 4156 15936 4168
rect 15988 4196 15994 4208
rect 16298 4196 16304 4208
rect 15988 4168 16304 4196
rect 15988 4156 15994 4168
rect 16298 4156 16304 4168
rect 16356 4156 16362 4208
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 21358 4196 21364 4208
rect 18104 4168 19288 4196
rect 18104 4156 18110 4168
rect 14734 4128 14740 4140
rect 13740 4100 14740 4128
rect 13357 4091 13415 4097
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4060 2283 4063
rect 2682 4060 2688 4072
rect 2271 4032 2688 4060
rect 2271 4029 2283 4032
rect 2225 4023 2283 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 2832 4032 3249 4060
rect 2832 4020 2838 4032
rect 3237 4029 3249 4032
rect 3283 4060 3295 4063
rect 3789 4063 3847 4069
rect 3789 4060 3801 4063
rect 3283 4032 3801 4060
rect 3283 4029 3295 4032
rect 3237 4023 3295 4029
rect 3789 4029 3801 4032
rect 3835 4060 3847 4063
rect 4062 4060 4068 4072
rect 3835 4032 4068 4060
rect 3835 4029 3847 4032
rect 3789 4023 3847 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4246 4020 4252 4072
rect 4304 4060 4310 4072
rect 5074 4060 5080 4072
rect 4304 4032 5080 4060
rect 4304 4020 4310 4032
rect 5074 4020 5080 4032
rect 5132 4060 5138 4072
rect 5261 4063 5319 4069
rect 5261 4060 5273 4063
rect 5132 4032 5273 4060
rect 5132 4020 5138 4032
rect 5261 4029 5273 4032
rect 5307 4029 5319 4063
rect 6546 4060 6552 4072
rect 6459 4032 6552 4060
rect 5261 4023 5319 4029
rect 6546 4020 6552 4032
rect 6604 4060 6610 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6604 4032 6837 4060
rect 6604 4020 6610 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9677 4063 9735 4069
rect 9677 4060 9689 4063
rect 9263 4032 9689 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9677 4029 9689 4032
rect 9723 4060 9735 4063
rect 10962 4060 10968 4072
rect 9723 4032 10968 4060
rect 9723 4029 9735 4032
rect 9677 4023 9735 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11333 4063 11391 4069
rect 11333 4029 11345 4063
rect 11379 4060 11391 4063
rect 12618 4060 12624 4072
rect 11379 4032 12624 4060
rect 11379 4029 11391 4032
rect 11333 4023 11391 4029
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 13078 4060 13084 4072
rect 12991 4032 13084 4060
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13372 4060 13400 4091
rect 14734 4088 14740 4100
rect 14792 4088 14798 4140
rect 14918 4128 14924 4140
rect 14879 4100 14924 4128
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 16577 4131 16635 4137
rect 16577 4097 16589 4131
rect 16623 4128 16635 4131
rect 16758 4128 16764 4140
rect 16623 4100 16764 4128
rect 16623 4097 16635 4100
rect 16577 4091 16635 4097
rect 16758 4088 16764 4100
rect 16816 4088 16822 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18138 4128 18144 4140
rect 17911 4100 18144 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 18138 4088 18144 4100
rect 18196 4128 18202 4140
rect 18598 4128 18604 4140
rect 18196 4100 18460 4128
rect 18559 4100 18604 4128
rect 18196 4088 18202 4100
rect 13722 4060 13728 4072
rect 13372 4032 13728 4060
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14642 4060 14648 4072
rect 14603 4032 14648 4060
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 16301 4063 16359 4069
rect 16301 4060 16313 4063
rect 15519 4032 16313 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 16301 4029 16313 4032
rect 16347 4060 16359 4063
rect 16390 4060 16396 4072
rect 16347 4032 16396 4060
rect 16347 4029 16359 4032
rect 16301 4023 16359 4029
rect 16390 4020 16396 4032
rect 16448 4020 16454 4072
rect 18432 4069 18460 4100
rect 18598 4088 18604 4100
rect 18656 4088 18662 4140
rect 19260 4128 19288 4168
rect 20272 4168 21364 4196
rect 20070 4128 20076 4140
rect 19260 4100 20076 4128
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20272 4137 20300 4168
rect 21358 4156 21364 4168
rect 21416 4156 21422 4208
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4097 20315 4131
rect 21726 4128 21732 4140
rect 21687 4100 21732 4128
rect 20257 4091 20315 4097
rect 21726 4088 21732 4100
rect 21784 4128 21790 4140
rect 22189 4131 22247 4137
rect 22189 4128 22201 4131
rect 21784 4100 22201 4128
rect 21784 4088 21790 4100
rect 22189 4097 22201 4100
rect 22235 4097 22247 4131
rect 22189 4091 22247 4097
rect 23474 4088 23480 4140
rect 23532 4128 23538 4140
rect 24213 4131 24271 4137
rect 24213 4128 24225 4131
rect 23532 4100 24225 4128
rect 23532 4088 23538 4100
rect 24213 4097 24225 4100
rect 24259 4097 24271 4131
rect 24213 4091 24271 4097
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4029 18475 4063
rect 19426 4060 19432 4072
rect 19387 4032 19432 4060
rect 18417 4023 18475 4029
rect 19426 4020 19432 4032
rect 19484 4020 19490 4072
rect 20714 4060 20720 4072
rect 19628 4032 20720 4060
rect 1670 3992 1676 4004
rect 1631 3964 1676 3992
rect 1670 3952 1676 3964
rect 1728 3952 1734 4004
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 2498 3992 2504 4004
rect 2179 3964 2504 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2498 3952 2504 3964
rect 2556 3952 2562 4004
rect 3878 3952 3884 4004
rect 3936 3992 3942 4004
rect 4617 3995 4675 4001
rect 4617 3992 4629 3995
rect 3936 3964 4629 3992
rect 3936 3952 3942 3964
rect 4617 3961 4629 3964
rect 4663 3961 4675 3995
rect 4798 3992 4804 4004
rect 4711 3964 4804 3992
rect 4617 3955 4675 3961
rect 4798 3952 4804 3964
rect 4856 3992 4862 4004
rect 5353 3995 5411 4001
rect 5353 3992 5365 3995
rect 4856 3964 5365 3992
rect 4856 3952 4862 3964
rect 5353 3961 5365 3964
rect 5399 3961 5411 3995
rect 5353 3955 5411 3961
rect 1762 3924 1768 3936
rect 1723 3896 1768 3924
rect 1762 3884 1768 3896
rect 1820 3884 1826 3936
rect 2682 3884 2688 3936
rect 2740 3924 2746 3936
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 2740 3896 2789 3924
rect 2740 3884 2746 3896
rect 2777 3893 2789 3896
rect 2823 3924 2835 3927
rect 3697 3927 3755 3933
rect 3697 3924 3709 3927
rect 2823 3896 3709 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 3697 3893 3709 3896
rect 3743 3893 3755 3927
rect 3697 3887 3755 3893
rect 5994 3884 6000 3936
rect 6052 3924 6058 3936
rect 6564 3933 6592 4020
rect 7092 3995 7150 4001
rect 7092 3961 7104 3995
rect 7138 3992 7150 3995
rect 7926 3992 7932 4004
rect 7138 3964 7932 3992
rect 7138 3961 7150 3964
rect 7092 3955 7150 3961
rect 7926 3952 7932 3964
rect 7984 3992 7990 4004
rect 7984 3964 8892 3992
rect 7984 3952 7990 3964
rect 8864 3936 8892 3964
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 10870 3992 10876 4004
rect 10652 3964 10876 3992
rect 10652 3952 10658 3964
rect 10870 3952 10876 3964
rect 10928 3952 10934 4004
rect 14660 3992 14688 4020
rect 17862 3992 17868 4004
rect 12728 3964 14688 3992
rect 15948 3964 17868 3992
rect 6181 3927 6239 3933
rect 6181 3924 6193 3927
rect 6052 3896 6193 3924
rect 6052 3884 6058 3896
rect 6181 3893 6193 3896
rect 6227 3924 6239 3927
rect 6549 3927 6607 3933
rect 6549 3924 6561 3927
rect 6227 3896 6561 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6549 3893 6561 3896
rect 6595 3893 6607 3927
rect 8202 3924 8208 3936
rect 8163 3896 8208 3924
rect 6549 3887 6607 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8846 3924 8852 3936
rect 8807 3896 8852 3924
rect 8846 3884 8852 3896
rect 8904 3884 8910 3936
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 9272 3896 9321 3924
rect 9272 3884 9278 3896
rect 9309 3893 9321 3896
rect 9355 3893 9367 3927
rect 9309 3887 9367 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10321 3927 10379 3933
rect 10321 3924 10333 3927
rect 10008 3896 10333 3924
rect 10008 3884 10014 3896
rect 10321 3893 10333 3896
rect 10367 3924 10379 3927
rect 10612 3924 10640 3952
rect 10367 3896 10640 3924
rect 11885 3927 11943 3933
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 11885 3893 11897 3927
rect 11931 3924 11943 3927
rect 12618 3924 12624 3936
rect 11931 3896 12624 3924
rect 11931 3893 11943 3896
rect 11885 3887 11943 3893
rect 12618 3884 12624 3896
rect 12676 3884 12682 3936
rect 12728 3933 12756 3964
rect 12713 3927 12771 3933
rect 12713 3893 12725 3927
rect 12759 3893 12771 3927
rect 12713 3887 12771 3893
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 13817 3927 13875 3933
rect 13228 3896 13273 3924
rect 13228 3884 13234 3896
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13998 3924 14004 3936
rect 13863 3896 14004 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13998 3884 14004 3896
rect 14056 3884 14062 3936
rect 14274 3924 14280 3936
rect 14235 3896 14280 3924
rect 14274 3884 14280 3896
rect 14332 3884 14338 3936
rect 15948 3933 15976 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 19242 3992 19248 4004
rect 18064 3964 19248 3992
rect 15933 3927 15991 3933
rect 15933 3893 15945 3927
rect 15979 3893 15991 3927
rect 15933 3887 15991 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16393 3927 16451 3933
rect 16393 3924 16405 3927
rect 16356 3896 16405 3924
rect 16356 3884 16362 3896
rect 16393 3893 16405 3896
rect 16439 3893 16451 3927
rect 16942 3924 16948 3936
rect 16903 3896 16948 3924
rect 16393 3887 16451 3893
rect 16942 3884 16948 3896
rect 17000 3884 17006 3936
rect 17034 3884 17040 3936
rect 17092 3924 17098 3936
rect 18064 3933 18092 3964
rect 19242 3952 19248 3964
rect 19300 3952 19306 4004
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 17092 3896 17325 3924
rect 17092 3884 17098 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 19628 3933 19656 4032
rect 20714 4020 20720 4032
rect 20772 4020 20778 4072
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 21637 4063 21695 4069
rect 21637 4060 21649 4063
rect 20864 4032 21649 4060
rect 20864 4020 20870 4032
rect 21637 4029 21649 4032
rect 21683 4060 21695 4063
rect 22002 4060 22008 4072
rect 21683 4032 22008 4060
rect 21683 4029 21695 4032
rect 21637 4023 21695 4029
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 22554 4020 22560 4072
rect 22612 4060 22618 4072
rect 22925 4063 22983 4069
rect 22925 4060 22937 4063
rect 22612 4032 22937 4060
rect 22612 4020 22618 4032
rect 22925 4029 22937 4032
rect 22971 4060 22983 4063
rect 23014 4060 23020 4072
rect 22971 4032 23020 4060
rect 22971 4029 22983 4032
rect 22925 4023 22983 4029
rect 23014 4020 23020 4032
rect 23072 4020 23078 4072
rect 23566 4020 23572 4072
rect 23624 4060 23630 4072
rect 24121 4063 24179 4069
rect 24121 4060 24133 4063
rect 23624 4032 24133 4060
rect 23624 4020 23630 4032
rect 24121 4029 24133 4032
rect 24167 4029 24179 4063
rect 25222 4060 25228 4072
rect 25135 4032 25228 4060
rect 24121 4023 24179 4029
rect 19981 3995 20039 4001
rect 19981 3961 19993 3995
rect 20027 3992 20039 3995
rect 20162 3992 20168 4004
rect 20027 3964 20168 3992
rect 20027 3961 20039 3964
rect 19981 3955 20039 3961
rect 20162 3952 20168 3964
rect 20220 3952 20226 4004
rect 21545 3995 21603 4001
rect 21545 3992 21557 3995
rect 20732 3964 21557 3992
rect 20732 3936 20760 3964
rect 21545 3961 21557 3964
rect 21591 3961 21603 3995
rect 21545 3955 21603 3961
rect 23750 3952 23756 4004
rect 23808 3992 23814 4004
rect 23934 3992 23940 4004
rect 23808 3964 23940 3992
rect 23808 3952 23814 3964
rect 23934 3952 23940 3964
rect 23992 3952 23998 4004
rect 24136 3992 24164 4023
rect 25222 4020 25228 4032
rect 25280 4060 25286 4072
rect 25777 4063 25835 4069
rect 25777 4060 25789 4063
rect 25280 4032 25789 4060
rect 25280 4020 25286 4032
rect 25777 4029 25789 4032
rect 25823 4029 25835 4063
rect 25777 4023 25835 4029
rect 26237 3995 26295 4001
rect 26237 3992 26249 3995
rect 24136 3964 26249 3992
rect 26237 3961 26249 3964
rect 26283 3961 26295 3995
rect 26237 3955 26295 3961
rect 18509 3927 18567 3933
rect 18509 3924 18521 3927
rect 18380 3896 18521 3924
rect 18380 3884 18386 3896
rect 18509 3893 18521 3896
rect 18555 3893 18567 3927
rect 18509 3887 18567 3893
rect 19613 3927 19671 3933
rect 19613 3893 19625 3927
rect 19659 3893 19671 3927
rect 20714 3924 20720 3936
rect 20675 3896 20720 3924
rect 19613 3887 19671 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 20806 3884 20812 3936
rect 20864 3924 20870 3936
rect 20993 3927 21051 3933
rect 20993 3924 21005 3927
rect 20864 3896 21005 3924
rect 20864 3884 20870 3896
rect 20993 3893 21005 3896
rect 21039 3893 21051 3927
rect 21174 3924 21180 3936
rect 21135 3896 21180 3924
rect 20993 3887 21051 3893
rect 21174 3884 21180 3896
rect 21232 3884 21238 3936
rect 22649 3927 22707 3933
rect 22649 3893 22661 3927
rect 22695 3924 22707 3927
rect 23014 3924 23020 3936
rect 22695 3896 23020 3924
rect 22695 3893 22707 3896
rect 22649 3887 22707 3893
rect 23014 3884 23020 3896
rect 23072 3884 23078 3936
rect 23474 3924 23480 3936
rect 23435 3896 23480 3924
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 23658 3924 23664 3936
rect 23619 3896 23664 3924
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 24029 3927 24087 3933
rect 24029 3893 24041 3927
rect 24075 3924 24087 3927
rect 24118 3924 24124 3936
rect 24075 3896 24124 3924
rect 24075 3893 24087 3896
rect 24029 3887 24087 3893
rect 24118 3884 24124 3896
rect 24176 3924 24182 3936
rect 24762 3924 24768 3936
rect 24176 3896 24768 3924
rect 24176 3884 24182 3896
rect 24762 3884 24768 3896
rect 24820 3884 24826 3936
rect 25038 3924 25044 3936
rect 24999 3896 25044 3924
rect 25038 3884 25044 3896
rect 25096 3884 25102 3936
rect 25406 3924 25412 3936
rect 25367 3896 25412 3924
rect 25406 3884 25412 3896
rect 25464 3884 25470 3936
rect 1104 3834 26864 3856
rect 1104 3782 10315 3834
rect 10367 3782 10379 3834
rect 10431 3782 10443 3834
rect 10495 3782 10507 3834
rect 10559 3782 19648 3834
rect 19700 3782 19712 3834
rect 19764 3782 19776 3834
rect 19828 3782 19840 3834
rect 19892 3782 26864 3834
rect 1104 3760 26864 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 1949 3723 2007 3729
rect 1949 3689 1961 3723
rect 1995 3720 2007 3723
rect 2314 3720 2320 3732
rect 1995 3692 2320 3720
rect 1995 3689 2007 3692
rect 1949 3683 2007 3689
rect 2314 3680 2320 3692
rect 2372 3680 2378 3732
rect 2409 3723 2467 3729
rect 2409 3689 2421 3723
rect 2455 3720 2467 3723
rect 2498 3720 2504 3732
rect 2455 3692 2504 3720
rect 2455 3689 2467 3692
rect 2409 3683 2467 3689
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2869 3723 2927 3729
rect 2869 3720 2881 3723
rect 2648 3692 2881 3720
rect 2648 3680 2654 3692
rect 2869 3689 2881 3692
rect 2915 3689 2927 3723
rect 2869 3683 2927 3689
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 4065 3723 4123 3729
rect 4065 3720 4077 3723
rect 4028 3692 4077 3720
rect 4028 3680 4034 3692
rect 4065 3689 4077 3692
rect 4111 3689 4123 3723
rect 5074 3720 5080 3732
rect 5035 3692 5080 3720
rect 4065 3683 4123 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 6972 3692 7205 3720
rect 6972 3680 6978 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 9674 3720 9680 3732
rect 9635 3692 9680 3720
rect 7193 3683 7251 3689
rect 2777 3655 2835 3661
rect 2777 3621 2789 3655
rect 2823 3652 2835 3655
rect 3878 3652 3884 3664
rect 2823 3624 3884 3652
rect 2823 3621 2835 3624
rect 2777 3615 2835 3621
rect 3878 3612 3884 3624
rect 3936 3612 3942 3664
rect 4433 3655 4491 3661
rect 4433 3652 4445 3655
rect 3988 3624 4445 3652
rect 3988 3596 4016 3624
rect 4433 3621 4445 3624
rect 4479 3652 4491 3655
rect 4982 3652 4988 3664
rect 4479 3624 4988 3652
rect 4479 3621 4491 3624
rect 4433 3615 4491 3621
rect 4982 3612 4988 3624
rect 5040 3612 5046 3664
rect 5721 3655 5779 3661
rect 5721 3621 5733 3655
rect 5767 3652 5779 3655
rect 7208 3652 7236 3683
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9916 3692 10057 3720
rect 9916 3680 9922 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10045 3683 10103 3689
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 12158 3720 12164 3732
rect 10888 3692 12164 3720
rect 10686 3652 10692 3664
rect 5767 3624 6123 3652
rect 7208 3624 10692 3652
rect 5767 3621 5779 3624
rect 5721 3615 5779 3621
rect 1394 3584 1400 3596
rect 1355 3556 1400 3584
rect 1394 3544 1400 3556
rect 1452 3544 1458 3596
rect 3970 3544 3976 3596
rect 4028 3544 4034 3596
rect 4522 3584 4528 3596
rect 4483 3556 4528 3584
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 5813 3587 5871 3593
rect 5813 3553 5825 3587
rect 5859 3584 5871 3587
rect 5902 3584 5908 3596
rect 5859 3556 5908 3584
rect 5859 3553 5871 3556
rect 5813 3547 5871 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6095 3593 6123 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 6080 3587 6138 3593
rect 6080 3553 6092 3587
rect 6126 3584 6138 3587
rect 8294 3584 8300 3596
rect 6126 3556 8300 3584
rect 6126 3553 6138 3556
rect 6080 3547 6138 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9493 3587 9551 3593
rect 9493 3584 9505 3587
rect 8904 3556 9505 3584
rect 8904 3544 8910 3556
rect 9493 3553 9505 3556
rect 9539 3584 9551 3587
rect 9539 3556 10364 3584
rect 9539 3553 9551 3556
rect 9493 3547 9551 3553
rect 3050 3516 3056 3528
rect 3011 3488 3056 3516
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 3513 3519 3571 3525
rect 3513 3516 3525 3519
rect 3476 3488 3525 3516
rect 3476 3476 3482 3488
rect 3513 3485 3525 3488
rect 3559 3516 3571 3519
rect 3881 3519 3939 3525
rect 3881 3516 3893 3519
rect 3559 3488 3893 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3881 3485 3893 3488
rect 3927 3516 3939 3519
rect 4062 3516 4068 3528
rect 3927 3488 4068 3516
rect 3927 3485 3939 3488
rect 3881 3479 3939 3485
rect 4062 3476 4068 3488
rect 4120 3516 4126 3528
rect 4709 3519 4767 3525
rect 4709 3516 4721 3519
rect 4120 3488 4721 3516
rect 4120 3476 4126 3488
rect 4709 3485 4721 3488
rect 4755 3516 4767 3519
rect 5442 3516 5448 3528
rect 4755 3488 5448 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 8573 3519 8631 3525
rect 7064 3488 8340 3516
rect 7064 3476 7070 3488
rect 7834 3448 7840 3460
rect 7795 3420 7840 3448
rect 7834 3408 7840 3420
rect 7892 3408 7898 3460
rect 8312 3448 8340 3488
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 9582 3516 9588 3528
rect 8619 3488 9588 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 10336 3525 10364 3556
rect 10321 3519 10379 3525
rect 10321 3485 10333 3519
rect 10367 3516 10379 3519
rect 10888 3516 10916 3692
rect 12158 3680 12164 3692
rect 12216 3720 12222 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 12216 3692 12265 3720
rect 12216 3680 12222 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12768 3692 12817 3720
rect 12768 3680 12774 3692
rect 12805 3689 12817 3692
rect 12851 3720 12863 3723
rect 13170 3720 13176 3732
rect 12851 3692 13176 3720
rect 12851 3689 12863 3692
rect 12805 3683 12863 3689
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13722 3720 13728 3732
rect 13587 3692 13728 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14001 3723 14059 3729
rect 14001 3689 14013 3723
rect 14047 3720 14059 3723
rect 14274 3720 14280 3732
rect 14047 3692 14280 3720
rect 14047 3689 14059 3692
rect 14001 3683 14059 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 16025 3723 16083 3729
rect 16025 3720 16037 3723
rect 15896 3692 16037 3720
rect 15896 3680 15902 3692
rect 16025 3689 16037 3692
rect 16071 3689 16083 3723
rect 16025 3683 16083 3689
rect 16117 3723 16175 3729
rect 16117 3689 16129 3723
rect 16163 3720 16175 3723
rect 16482 3720 16488 3732
rect 16163 3692 16488 3720
rect 16163 3689 16175 3692
rect 16117 3683 16175 3689
rect 16482 3680 16488 3692
rect 16540 3680 16546 3732
rect 16945 3723 17003 3729
rect 16945 3689 16957 3723
rect 16991 3720 17003 3723
rect 17402 3720 17408 3732
rect 16991 3692 17408 3720
rect 16991 3689 17003 3692
rect 16945 3683 17003 3689
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 17862 3720 17868 3732
rect 17635 3692 17868 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 20162 3720 20168 3732
rect 18831 3692 20168 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 20162 3680 20168 3692
rect 20220 3680 20226 3732
rect 20901 3723 20959 3729
rect 20901 3689 20913 3723
rect 20947 3720 20959 3723
rect 21910 3720 21916 3732
rect 20947 3692 21916 3720
rect 20947 3689 20959 3692
rect 20901 3683 20959 3689
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22094 3680 22100 3732
rect 22152 3720 22158 3732
rect 22281 3723 22339 3729
rect 22281 3720 22293 3723
rect 22152 3692 22293 3720
rect 22152 3680 22158 3692
rect 22281 3689 22293 3692
rect 22327 3689 22339 3723
rect 22281 3683 22339 3689
rect 22465 3723 22523 3729
rect 22465 3689 22477 3723
rect 22511 3720 22523 3723
rect 22830 3720 22836 3732
rect 22511 3692 22836 3720
rect 22511 3689 22523 3692
rect 22465 3683 22523 3689
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 24486 3720 24492 3732
rect 24447 3692 24492 3720
rect 24486 3680 24492 3692
rect 24544 3720 24550 3732
rect 25222 3720 25228 3732
rect 24544 3692 25228 3720
rect 24544 3680 24550 3692
rect 25222 3680 25228 3692
rect 25280 3680 25286 3732
rect 11514 3612 11520 3664
rect 11572 3652 11578 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11572 3624 11621 3652
rect 11572 3612 11578 3624
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 14090 3652 14096 3664
rect 14003 3624 14096 3652
rect 11609 3615 11667 3621
rect 14090 3612 14096 3624
rect 14148 3652 14154 3664
rect 15102 3652 15108 3664
rect 14148 3624 15108 3652
rect 14148 3612 14154 3624
rect 15102 3612 15108 3624
rect 15160 3612 15166 3664
rect 18509 3655 18567 3661
rect 18509 3621 18521 3655
rect 18555 3652 18567 3655
rect 18874 3652 18880 3664
rect 18555 3624 18880 3652
rect 18555 3621 18567 3624
rect 18509 3615 18567 3621
rect 18874 3612 18880 3624
rect 18932 3612 18938 3664
rect 19242 3652 19248 3664
rect 19203 3624 19248 3652
rect 19242 3612 19248 3624
rect 19300 3612 19306 3664
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 19797 3655 19855 3661
rect 19797 3652 19809 3655
rect 19484 3624 19809 3652
rect 19484 3612 19490 3624
rect 19797 3621 19809 3624
rect 19843 3652 19855 3655
rect 20530 3652 20536 3664
rect 19843 3624 20536 3652
rect 19843 3621 19855 3624
rect 19797 3615 19855 3621
rect 20530 3612 20536 3624
rect 20588 3652 20594 3664
rect 20625 3655 20683 3661
rect 20625 3652 20637 3655
rect 20588 3624 20637 3652
rect 20588 3612 20594 3624
rect 20625 3621 20637 3624
rect 20671 3652 20683 3655
rect 20671 3624 21404 3652
rect 20671 3621 20683 3624
rect 20625 3615 20683 3621
rect 11146 3584 11152 3596
rect 11059 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3584 11210 3596
rect 14737 3587 14795 3593
rect 11204 3556 11836 3584
rect 11204 3544 11210 3556
rect 11698 3516 11704 3528
rect 10367 3488 10916 3516
rect 11659 3488 11704 3516
rect 10367 3485 10379 3488
rect 10321 3479 10379 3485
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 11808 3525 11836 3556
rect 14737 3553 14749 3587
rect 14783 3584 14795 3587
rect 14918 3584 14924 3596
rect 14783 3556 14924 3584
rect 14783 3553 14795 3556
rect 14737 3547 14795 3553
rect 14918 3544 14924 3556
rect 14976 3584 14982 3596
rect 14976 3556 15148 3584
rect 14976 3544 14982 3556
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14826 3516 14832 3528
rect 14323 3488 14832 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 9033 3451 9091 3457
rect 9033 3448 9045 3451
rect 8312 3420 9045 3448
rect 9033 3417 9045 3420
rect 9079 3448 9091 3451
rect 9122 3448 9128 3460
rect 9079 3420 9128 3448
rect 9079 3417 9091 3420
rect 9033 3411 9091 3417
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 13173 3451 13231 3457
rect 13173 3417 13185 3451
rect 13219 3448 13231 3451
rect 14292 3448 14320 3479
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 15120 3525 15148 3556
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 17586 3584 17592 3596
rect 16632 3556 17592 3584
rect 16632 3544 16638 3556
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 18046 3544 18052 3596
rect 18104 3584 18110 3596
rect 19058 3584 19064 3596
rect 18104 3556 19064 3584
rect 18104 3544 18110 3556
rect 19058 3544 19064 3556
rect 19116 3584 19122 3596
rect 19153 3587 19211 3593
rect 19153 3584 19165 3587
rect 19116 3556 19165 3584
rect 19116 3544 19122 3556
rect 19153 3553 19165 3556
rect 19199 3553 19211 3587
rect 21266 3584 21272 3596
rect 21227 3556 21272 3584
rect 19153 3547 19211 3553
rect 21266 3544 21272 3556
rect 21324 3544 21330 3596
rect 21376 3584 21404 3624
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 25409 3655 25467 3661
rect 25409 3652 25421 3655
rect 24360 3624 25421 3652
rect 24360 3612 24366 3624
rect 25409 3621 25421 3624
rect 25455 3621 25467 3655
rect 26234 3652 26240 3664
rect 26195 3624 26240 3652
rect 25409 3615 25467 3621
rect 26234 3612 26240 3624
rect 26292 3612 26298 3664
rect 22830 3584 22836 3596
rect 21376 3556 21496 3584
rect 22791 3556 22836 3584
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15378 3516 15384 3528
rect 15151 3488 15384 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15378 3476 15384 3488
rect 15436 3516 15442 3528
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 15436 3488 15577 3516
rect 15436 3476 15442 3488
rect 15565 3485 15577 3488
rect 15611 3516 15623 3519
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 15611 3488 16313 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 16301 3485 16313 3488
rect 16347 3516 16359 3519
rect 16758 3516 16764 3528
rect 16347 3488 16764 3516
rect 16347 3485 16359 3488
rect 16301 3479 16359 3485
rect 16758 3476 16764 3488
rect 16816 3476 16822 3528
rect 17681 3519 17739 3525
rect 17681 3485 17693 3519
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 13219 3420 14320 3448
rect 13219 3417 13231 3420
rect 13173 3411 13231 3417
rect 14550 3408 14556 3460
rect 14608 3448 14614 3460
rect 15010 3448 15016 3460
rect 14608 3420 15016 3448
rect 14608 3408 14614 3420
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 16666 3448 16672 3460
rect 15703 3420 16672 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 16666 3408 16672 3420
rect 16724 3448 16730 3460
rect 17696 3448 17724 3479
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 17828 3488 17873 3516
rect 17828 3476 17834 3488
rect 18966 3476 18972 3528
rect 19024 3516 19030 3528
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 19024 3488 19349 3516
rect 19024 3476 19030 3488
rect 19337 3485 19349 3488
rect 19383 3485 19395 3519
rect 19337 3479 19395 3485
rect 20990 3476 20996 3528
rect 21048 3516 21054 3528
rect 21358 3516 21364 3528
rect 21048 3488 21364 3516
rect 21048 3476 21054 3488
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 21468 3525 21496 3556
rect 22830 3544 22836 3556
rect 22888 3544 22894 3596
rect 22922 3544 22928 3596
rect 22980 3584 22986 3596
rect 24397 3587 24455 3593
rect 22980 3556 23025 3584
rect 22980 3544 22986 3556
rect 24397 3553 24409 3587
rect 24443 3584 24455 3587
rect 24946 3584 24952 3596
rect 24443 3556 24952 3584
rect 24443 3553 24455 3556
rect 24397 3547 24455 3553
rect 24946 3544 24952 3556
rect 25004 3544 25010 3596
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 21634 3516 21640 3528
rect 21499 3488 21640 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 21634 3476 21640 3488
rect 21692 3516 21698 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 21692 3488 21925 3516
rect 21692 3476 21698 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 21913 3479 21971 3485
rect 23014 3476 23020 3488
rect 23072 3516 23078 3528
rect 23566 3516 23572 3528
rect 23072 3488 23572 3516
rect 23072 3476 23078 3488
rect 23566 3476 23572 3488
rect 23624 3516 23630 3528
rect 23845 3519 23903 3525
rect 23845 3516 23857 3519
rect 23624 3488 23857 3516
rect 23624 3476 23630 3488
rect 23845 3485 23857 3488
rect 23891 3516 23903 3519
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23891 3488 24593 3516
rect 23891 3485 23903 3488
rect 23845 3479 23903 3485
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 16724 3420 17724 3448
rect 16724 3408 16730 3420
rect 23934 3408 23940 3460
rect 23992 3448 23998 3460
rect 25777 3451 25835 3457
rect 25777 3448 25789 3451
rect 23992 3420 25789 3448
rect 23992 3408 23998 3420
rect 25777 3417 25789 3420
rect 25823 3417 25835 3451
rect 25777 3411 25835 3417
rect 8481 3383 8539 3389
rect 8481 3349 8493 3383
rect 8527 3380 8539 3383
rect 8662 3380 8668 3392
rect 8527 3352 8668 3380
rect 8527 3349 8539 3352
rect 8481 3343 8539 3349
rect 8662 3340 8668 3352
rect 8720 3340 8726 3392
rect 11238 3380 11244 3392
rect 11199 3352 11244 3380
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 13630 3380 13636 3392
rect 13591 3352 13636 3380
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 17126 3380 17132 3392
rect 13780 3352 17132 3380
rect 13780 3340 13786 3352
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 18322 3380 18328 3392
rect 17267 3352 18328 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 20165 3383 20223 3389
rect 20165 3380 20177 3383
rect 19484 3352 20177 3380
rect 19484 3340 19490 3352
rect 20165 3349 20177 3352
rect 20211 3380 20223 3383
rect 20254 3380 20260 3392
rect 20211 3352 20260 3380
rect 20211 3349 20223 3352
rect 20165 3343 20223 3349
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 23474 3380 23480 3392
rect 23435 3352 23480 3380
rect 23474 3340 23480 3352
rect 23532 3340 23538 3392
rect 24026 3380 24032 3392
rect 23987 3352 24032 3380
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 25038 3380 25044 3392
rect 24999 3352 25044 3380
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 1104 3290 26864 3312
rect 1104 3238 5648 3290
rect 5700 3238 5712 3290
rect 5764 3238 5776 3290
rect 5828 3238 5840 3290
rect 5892 3238 14982 3290
rect 15034 3238 15046 3290
rect 15098 3238 15110 3290
rect 15162 3238 15174 3290
rect 15226 3238 24315 3290
rect 24367 3238 24379 3290
rect 24431 3238 24443 3290
rect 24495 3238 24507 3290
rect 24559 3238 26864 3290
rect 1104 3216 26864 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 1857 3179 1915 3185
rect 1857 3176 1869 3179
rect 1728 3148 1869 3176
rect 1728 3136 1734 3148
rect 1857 3145 1869 3148
rect 1903 3176 1915 3179
rect 3050 3176 3056 3188
rect 1903 3148 3056 3176
rect 1903 3145 1915 3148
rect 1857 3139 1915 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3510 3176 3516 3188
rect 3471 3148 3516 3176
rect 3510 3136 3516 3148
rect 3568 3176 3574 3188
rect 3786 3176 3792 3188
rect 3568 3148 3792 3176
rect 3568 3136 3574 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 6638 3136 6644 3188
rect 6696 3176 6702 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 6696 3148 6837 3176
rect 6696 3136 6702 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 6825 3139 6883 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10689 3179 10747 3185
rect 10689 3176 10701 3179
rect 10192 3148 10701 3176
rect 10192 3136 10198 3148
rect 10689 3145 10701 3148
rect 10735 3176 10747 3179
rect 13722 3176 13728 3188
rect 10735 3148 13728 3176
rect 10735 3145 10747 3148
rect 10689 3139 10747 3145
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 15470 3176 15476 3188
rect 13872 3148 15476 3176
rect 13872 3136 13878 3148
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16482 3176 16488 3188
rect 16395 3148 16488 3176
rect 16482 3136 16488 3148
rect 16540 3176 16546 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 16540 3148 17509 3176
rect 16540 3136 16546 3148
rect 17497 3145 17509 3148
rect 17543 3176 17555 3179
rect 17770 3176 17776 3188
rect 17543 3148 17776 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3176 18107 3179
rect 18782 3176 18788 3188
rect 18095 3148 18788 3176
rect 18095 3145 18107 3148
rect 18049 3139 18107 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19613 3179 19671 3185
rect 19613 3145 19625 3179
rect 19659 3176 19671 3179
rect 20898 3176 20904 3188
rect 19659 3148 20904 3176
rect 19659 3145 19671 3148
rect 19613 3139 19671 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21266 3176 21272 3188
rect 21008 3148 21272 3176
rect 4522 3108 4528 3120
rect 4483 3080 4528 3108
rect 4522 3068 4528 3080
rect 4580 3068 4586 3120
rect 4982 3108 4988 3120
rect 4943 3080 4988 3108
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 5077 3111 5135 3117
rect 5077 3077 5089 3111
rect 5123 3108 5135 3111
rect 5166 3108 5172 3120
rect 5123 3080 5172 3108
rect 5123 3077 5135 3080
rect 5077 3071 5135 3077
rect 5166 3068 5172 3080
rect 5224 3068 5230 3120
rect 6549 3111 6607 3117
rect 6549 3077 6561 3111
rect 6595 3108 6607 3111
rect 7282 3108 7288 3120
rect 6595 3080 7288 3108
rect 6595 3077 6607 3080
rect 6549 3071 6607 3077
rect 7282 3068 7288 3080
rect 7340 3068 7346 3120
rect 9858 3068 9864 3120
rect 9916 3108 9922 3120
rect 10321 3111 10379 3117
rect 10321 3108 10333 3111
rect 9916 3080 10333 3108
rect 9916 3068 9922 3080
rect 10321 3077 10333 3080
rect 10367 3077 10379 3111
rect 11425 3111 11483 3117
rect 10321 3071 10379 3077
rect 10888 3080 11376 3108
rect 2314 3000 2320 3052
rect 2372 3040 2378 3052
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2372 3012 2513 3040
rect 2372 3000 2378 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3053 3043 3111 3049
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 4062 3040 4068 3052
rect 3099 3012 4068 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5629 3043 5687 3049
rect 5629 3040 5641 3043
rect 5316 3012 5641 3040
rect 5316 3000 5322 3012
rect 5629 3009 5641 3012
rect 5675 3009 5687 3043
rect 5629 3003 5687 3009
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6638 3040 6644 3052
rect 6512 3012 6644 3040
rect 6512 3000 6518 3012
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7377 3043 7435 3049
rect 7377 3040 7389 3043
rect 7064 3012 7389 3040
rect 7064 3000 7070 3012
rect 7377 3009 7389 3012
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 10888 3040 10916 3080
rect 9456 3012 10916 3040
rect 9456 3000 9462 3012
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11348 3040 11376 3080
rect 11425 3077 11437 3111
rect 11471 3108 11483 3111
rect 12434 3108 12440 3120
rect 11471 3080 12440 3108
rect 11471 3077 11483 3080
rect 11425 3071 11483 3077
rect 12434 3068 12440 3080
rect 12492 3068 12498 3120
rect 16758 3068 16764 3120
rect 16816 3108 16822 3120
rect 17037 3111 17095 3117
rect 17037 3108 17049 3111
rect 16816 3080 17049 3108
rect 16816 3068 16822 3080
rect 17037 3077 17049 3080
rect 17083 3077 17095 3111
rect 17037 3071 17095 3077
rect 19521 3111 19579 3117
rect 19521 3077 19533 3111
rect 19567 3108 19579 3111
rect 20622 3108 20628 3120
rect 19567 3080 20628 3108
rect 19567 3077 19579 3080
rect 19521 3071 19579 3077
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 11112 3012 11284 3040
rect 11348 3012 12572 3040
rect 11112 3000 11118 3012
rect 2409 2975 2467 2981
rect 2409 2941 2421 2975
rect 2455 2972 2467 2975
rect 2866 2972 2872 2984
rect 2455 2944 2872 2972
rect 2455 2941 2467 2944
rect 2409 2935 2467 2941
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 5350 2932 5356 2984
rect 5408 2972 5414 2984
rect 5445 2975 5503 2981
rect 5445 2972 5457 2975
rect 5408 2944 5457 2972
rect 5408 2932 5414 2944
rect 5445 2941 5457 2944
rect 5491 2941 5503 2975
rect 5445 2935 5503 2941
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 6086 2972 6092 2984
rect 5583 2944 6092 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 6086 2932 6092 2944
rect 6144 2932 6150 2984
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2972 7254 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7248 2944 7849 2972
rect 7248 2932 7254 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 7837 2935 7895 2941
rect 8220 2944 8401 2972
rect 2130 2864 2136 2916
rect 2188 2904 2194 2916
rect 2317 2907 2375 2913
rect 2317 2904 2329 2907
rect 2188 2876 2329 2904
rect 2188 2864 2194 2876
rect 2317 2873 2329 2876
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 3421 2907 3479 2913
rect 3421 2873 3433 2907
rect 3467 2904 3479 2907
rect 7282 2904 7288 2916
rect 3467 2876 4016 2904
rect 7243 2876 7288 2904
rect 3467 2873 3479 2876
rect 3421 2867 3479 2873
rect 1946 2836 1952 2848
rect 1907 2808 1952 2836
rect 1946 2796 1952 2808
rect 2004 2796 2010 2848
rect 2406 2796 2412 2848
rect 2464 2836 2470 2848
rect 2774 2836 2780 2848
rect 2464 2808 2780 2836
rect 2464 2796 2470 2808
rect 2774 2796 2780 2808
rect 2832 2796 2838 2848
rect 3878 2836 3884 2848
rect 3839 2808 3884 2836
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 3988 2845 4016 2876
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 3973 2839 4031 2845
rect 3973 2805 3985 2839
rect 4019 2836 4031 2839
rect 4062 2836 4068 2848
rect 4019 2808 4068 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4430 2796 4436 2848
rect 4488 2836 4494 2848
rect 5994 2836 6000 2848
rect 4488 2808 6000 2836
rect 4488 2796 4494 2808
rect 5994 2796 6000 2808
rect 6052 2836 6058 2848
rect 6089 2839 6147 2845
rect 6089 2836 6101 2839
rect 6052 2808 6101 2836
rect 6052 2796 6058 2808
rect 6089 2805 6101 2808
rect 6135 2836 6147 2839
rect 6546 2836 6552 2848
rect 6135 2808 6552 2836
rect 6135 2805 6147 2808
rect 6089 2799 6147 2805
rect 6546 2796 6552 2808
rect 6604 2836 6610 2848
rect 8220 2845 8248 2944
rect 8389 2941 8401 2944
rect 8435 2972 8447 2975
rect 8478 2972 8484 2984
rect 8435 2944 8484 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 8662 2981 8668 2984
rect 8656 2972 8668 2981
rect 8623 2944 8668 2972
rect 8656 2935 8668 2944
rect 8662 2932 8668 2935
rect 8720 2932 8726 2984
rect 9490 2932 9496 2984
rect 9548 2932 9554 2984
rect 11256 2981 11284 3012
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2941 11299 2975
rect 12437 2975 12495 2981
rect 12437 2972 12449 2975
rect 11241 2935 11299 2941
rect 11808 2944 12449 2972
rect 9508 2904 9536 2932
rect 8404 2876 9536 2904
rect 8404 2848 8432 2876
rect 10778 2864 10784 2916
rect 10836 2904 10842 2916
rect 11808 2904 11836 2944
rect 12437 2941 12449 2944
rect 12483 2941 12495 2975
rect 12544 2972 12572 3012
rect 13832 3012 14841 3040
rect 13832 2972 13860 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17644 3012 17877 3040
rect 17644 3000 17650 3012
rect 17865 3009 17877 3012
rect 17911 3040 17923 3043
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 17911 3012 18613 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 12544 2944 13860 2972
rect 12437 2935 12495 2941
rect 14642 2932 14648 2984
rect 14700 2932 14706 2984
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 15378 2981 15384 2984
rect 15372 2972 15384 2981
rect 15339 2944 15384 2972
rect 15372 2935 15384 2944
rect 15378 2932 15384 2935
rect 15436 2932 15442 2984
rect 18414 2972 18420 2984
rect 18375 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 18506 2932 18512 2984
rect 18564 2972 18570 2984
rect 19996 2981 20024 3080
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 20717 3111 20775 3117
rect 20717 3077 20729 3111
rect 20763 3108 20775 3111
rect 21008 3108 21036 3148
rect 21266 3136 21272 3148
rect 21324 3136 21330 3188
rect 21818 3136 21824 3188
rect 21876 3176 21882 3188
rect 22189 3179 22247 3185
rect 22189 3176 22201 3179
rect 21876 3148 22201 3176
rect 21876 3136 21882 3148
rect 22189 3145 22201 3148
rect 22235 3145 22247 3179
rect 23474 3176 23480 3188
rect 23435 3148 23480 3176
rect 22189 3139 22247 3145
rect 23474 3136 23480 3148
rect 23532 3136 23538 3188
rect 24670 3136 24676 3188
rect 24728 3176 24734 3188
rect 24946 3176 24952 3188
rect 24728 3148 24952 3176
rect 24728 3136 24734 3148
rect 24946 3136 24952 3148
rect 25004 3176 25010 3188
rect 25041 3179 25099 3185
rect 25041 3176 25053 3179
rect 25004 3148 25053 3176
rect 25004 3136 25010 3148
rect 25041 3145 25053 3148
rect 25087 3145 25099 3179
rect 25041 3139 25099 3145
rect 20763 3080 21036 3108
rect 21177 3111 21235 3117
rect 20763 3077 20775 3080
rect 20717 3071 20775 3077
rect 21177 3077 21189 3111
rect 21223 3077 21235 3111
rect 21177 3071 21235 3077
rect 20257 3043 20315 3049
rect 20257 3009 20269 3043
rect 20303 3040 20315 3043
rect 20530 3040 20536 3052
rect 20303 3012 20536 3040
rect 20303 3009 20315 3012
rect 20257 3003 20315 3009
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 19981 2975 20039 2981
rect 18564 2944 18609 2972
rect 18564 2932 18570 2944
rect 19981 2941 19993 2975
rect 20027 2941 20039 2975
rect 19981 2935 20039 2941
rect 20073 2975 20131 2981
rect 20073 2941 20085 2975
rect 20119 2972 20131 2975
rect 20346 2972 20352 2984
rect 20119 2944 20352 2972
rect 20119 2941 20131 2944
rect 20073 2935 20131 2941
rect 20346 2932 20352 2944
rect 20404 2932 20410 2984
rect 21192 2972 21220 3071
rect 22094 3068 22100 3120
rect 22152 3108 22158 3120
rect 22925 3111 22983 3117
rect 22925 3108 22937 3111
rect 22152 3080 22937 3108
rect 22152 3068 22158 3080
rect 22925 3077 22937 3080
rect 22971 3108 22983 3111
rect 23014 3108 23020 3120
rect 22971 3080 23020 3108
rect 22971 3077 22983 3080
rect 22925 3071 22983 3077
rect 23014 3068 23020 3080
rect 23072 3068 23078 3120
rect 23106 3068 23112 3120
rect 23164 3108 23170 3120
rect 24578 3108 24584 3120
rect 23164 3080 24584 3108
rect 23164 3068 23170 3080
rect 24578 3068 24584 3080
rect 24636 3068 24642 3120
rect 24765 3111 24823 3117
rect 24765 3077 24777 3111
rect 24811 3108 24823 3111
rect 25222 3108 25228 3120
rect 24811 3080 25228 3108
rect 24811 3077 24823 3080
rect 24765 3071 24823 3077
rect 25222 3068 25228 3080
rect 25280 3068 25286 3120
rect 21634 3000 21640 3052
rect 21692 3040 21698 3052
rect 21729 3043 21787 3049
rect 21729 3040 21741 3043
rect 21692 3012 21741 3040
rect 21692 3000 21698 3012
rect 21729 3009 21741 3012
rect 21775 3009 21787 3043
rect 21729 3003 21787 3009
rect 22370 3000 22376 3052
rect 22428 3040 22434 3052
rect 23842 3040 23848 3052
rect 22428 3012 23848 3040
rect 22428 3000 22434 3012
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 23934 3000 23940 3052
rect 23992 3040 23998 3052
rect 24121 3043 24179 3049
rect 24121 3040 24133 3043
rect 23992 3012 24133 3040
rect 23992 3000 23998 3012
rect 24121 3009 24133 3012
rect 24167 3009 24179 3043
rect 24121 3003 24179 3009
rect 24213 3043 24271 3049
rect 24213 3009 24225 3043
rect 24259 3009 24271 3043
rect 24213 3003 24271 3009
rect 22922 2972 22928 2984
rect 21192 2944 22928 2972
rect 22922 2932 22928 2944
rect 22980 2932 22986 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 24228 2972 24256 3003
rect 25222 2972 25228 2984
rect 23624 2944 24256 2972
rect 25135 2944 25228 2972
rect 23624 2932 23630 2944
rect 25222 2932 25228 2944
rect 25280 2972 25286 2984
rect 25777 2975 25835 2981
rect 25777 2972 25789 2975
rect 25280 2944 25789 2972
rect 25280 2932 25286 2944
rect 25777 2941 25789 2944
rect 25823 2941 25835 2975
rect 25777 2935 25835 2941
rect 10836 2876 11836 2904
rect 10836 2864 10842 2876
rect 8205 2839 8263 2845
rect 8205 2836 8217 2839
rect 6604 2808 8217 2836
rect 6604 2796 6610 2808
rect 8205 2805 8217 2808
rect 8251 2805 8263 2839
rect 8205 2799 8263 2805
rect 8386 2796 8392 2848
rect 8444 2796 8450 2848
rect 8662 2796 8668 2848
rect 8720 2836 8726 2848
rect 9490 2836 9496 2848
rect 8720 2808 9496 2836
rect 8720 2796 8726 2808
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2836 11207 2839
rect 11330 2836 11336 2848
rect 11195 2808 11336 2836
rect 11195 2805 11207 2808
rect 11149 2799 11207 2805
rect 11330 2796 11336 2808
rect 11388 2796 11394 2848
rect 11808 2836 11836 2876
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12704 2907 12762 2913
rect 12704 2904 12716 2907
rect 11931 2876 12716 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 12704 2873 12716 2876
rect 12750 2904 12762 2907
rect 13722 2904 13728 2916
rect 12750 2876 13728 2904
rect 12750 2873 12762 2876
rect 12704 2867 12762 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 14660 2904 14688 2932
rect 15654 2904 15660 2916
rect 14660 2876 15660 2904
rect 15654 2864 15660 2876
rect 15712 2864 15718 2916
rect 21358 2864 21364 2916
rect 21416 2904 21422 2916
rect 22557 2907 22615 2913
rect 22557 2904 22569 2907
rect 21416 2876 22569 2904
rect 21416 2864 21422 2876
rect 22557 2873 22569 2876
rect 22603 2904 22615 2907
rect 22738 2904 22744 2916
rect 22603 2876 22744 2904
rect 22603 2873 22615 2876
rect 22557 2867 22615 2873
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 23474 2864 23480 2916
rect 23532 2904 23538 2916
rect 24029 2907 24087 2913
rect 24029 2904 24041 2907
rect 23532 2876 24041 2904
rect 23532 2864 23538 2876
rect 24029 2873 24041 2876
rect 24075 2873 24087 2907
rect 24029 2867 24087 2873
rect 12161 2839 12219 2845
rect 12161 2836 12173 2839
rect 11808 2808 12173 2836
rect 12161 2805 12173 2808
rect 12207 2836 12219 2839
rect 12526 2836 12532 2848
rect 12207 2808 12532 2836
rect 12207 2805 12219 2808
rect 12161 2799 12219 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 14642 2836 14648 2848
rect 14603 2808 14648 2836
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 14829 2839 14887 2845
rect 14829 2805 14841 2839
rect 14875 2836 14887 2839
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 14875 2808 15025 2836
rect 14875 2805 14887 2808
rect 14829 2799 14887 2805
rect 15013 2805 15025 2808
rect 15059 2836 15071 2839
rect 15838 2836 15844 2848
rect 15059 2808 15844 2836
rect 15059 2805 15071 2808
rect 15013 2799 15071 2805
rect 15838 2796 15844 2808
rect 15896 2796 15902 2848
rect 20990 2796 20996 2848
rect 21048 2836 21054 2848
rect 21085 2839 21143 2845
rect 21085 2836 21097 2839
rect 21048 2808 21097 2836
rect 21048 2796 21054 2808
rect 21085 2805 21097 2808
rect 21131 2836 21143 2839
rect 21545 2839 21603 2845
rect 21545 2836 21557 2839
rect 21131 2808 21557 2836
rect 21131 2805 21143 2808
rect 21085 2799 21143 2805
rect 21545 2805 21557 2808
rect 21591 2805 21603 2839
rect 21545 2799 21603 2805
rect 21637 2839 21695 2845
rect 21637 2805 21649 2839
rect 21683 2836 21695 2839
rect 21818 2836 21824 2848
rect 21683 2808 21824 2836
rect 21683 2805 21695 2808
rect 21637 2799 21695 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 23658 2836 23664 2848
rect 23619 2808 23664 2836
rect 23658 2796 23664 2808
rect 23716 2796 23722 2848
rect 25130 2796 25136 2848
rect 25188 2836 25194 2848
rect 25409 2839 25467 2845
rect 25409 2836 25421 2839
rect 25188 2808 25421 2836
rect 25188 2796 25194 2808
rect 25409 2805 25421 2808
rect 25455 2805 25467 2839
rect 26234 2836 26240 2848
rect 26195 2808 26240 2836
rect 25409 2799 25467 2805
rect 26234 2796 26240 2808
rect 26292 2796 26298 2848
rect 1104 2746 26864 2768
rect 1104 2694 10315 2746
rect 10367 2694 10379 2746
rect 10431 2694 10443 2746
rect 10495 2694 10507 2746
rect 10559 2694 19648 2746
rect 19700 2694 19712 2746
rect 19764 2694 19776 2746
rect 19828 2694 19840 2746
rect 19892 2694 26864 2746
rect 1104 2672 26864 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2409 2635 2467 2641
rect 2409 2632 2421 2635
rect 2188 2604 2421 2632
rect 2188 2592 2194 2604
rect 2409 2601 2421 2604
rect 2455 2601 2467 2635
rect 2409 2595 2467 2601
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 3786 2632 3792 2644
rect 2823 2604 3792 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 4798 2632 4804 2644
rect 3936 2604 4804 2632
rect 3936 2592 3942 2604
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 5721 2635 5779 2641
rect 5721 2601 5733 2635
rect 5767 2632 5779 2635
rect 6178 2632 6184 2644
rect 5767 2604 6184 2632
rect 5767 2601 5779 2604
rect 5721 2595 5779 2601
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 6604 2604 6653 2632
rect 6604 2592 6610 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 2869 2567 2927 2573
rect 2869 2533 2881 2567
rect 2915 2564 2927 2567
rect 3142 2564 3148 2576
rect 2915 2536 3148 2564
rect 2915 2533 2927 2536
rect 2869 2527 2927 2533
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 3605 2567 3663 2573
rect 3605 2533 3617 2567
rect 3651 2564 3663 2567
rect 3896 2564 3924 2592
rect 3651 2536 3924 2564
rect 3651 2533 3663 2536
rect 3605 2527 3663 2533
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1946 2496 1952 2508
rect 1443 2468 1952 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2428 2375 2431
rect 3050 2428 3056 2440
rect 2363 2400 3056 2428
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 1762 2320 1768 2372
rect 1820 2360 1826 2372
rect 3620 2360 3648 2527
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4430 2496 4436 2508
rect 4387 2468 4436 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 4608 2499 4666 2505
rect 4608 2465 4620 2499
rect 4654 2496 4666 2499
rect 5074 2496 5080 2508
rect 4654 2468 5080 2496
rect 4654 2465 4666 2468
rect 4608 2459 4666 2465
rect 5074 2456 5080 2468
rect 5132 2496 5138 2508
rect 6273 2499 6331 2505
rect 6273 2496 6285 2499
rect 5132 2468 6285 2496
rect 5132 2456 5138 2468
rect 6273 2465 6285 2468
rect 6319 2465 6331 2499
rect 6656 2496 6684 2595
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7834 2632 7840 2644
rect 7432 2604 7840 2632
rect 7432 2592 7438 2604
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 12250 2632 12256 2644
rect 10192 2604 12256 2632
rect 10192 2592 10198 2604
rect 12250 2592 12256 2604
rect 12308 2592 12314 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12526 2632 12532 2644
rect 12483 2604 12532 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12526 2592 12532 2604
rect 12584 2632 12590 2644
rect 13446 2632 13452 2644
rect 12584 2604 13452 2632
rect 12584 2592 12590 2604
rect 7184 2567 7242 2573
rect 7184 2533 7196 2567
rect 7230 2564 7242 2567
rect 7926 2564 7932 2576
rect 7230 2536 7932 2564
rect 7230 2533 7242 2536
rect 7184 2527 7242 2533
rect 7926 2524 7932 2536
rect 7984 2524 7990 2576
rect 8478 2524 8484 2576
rect 8536 2564 8542 2576
rect 8849 2567 8907 2573
rect 8849 2564 8861 2567
rect 8536 2536 8861 2564
rect 8536 2524 8542 2536
rect 8849 2533 8861 2536
rect 8895 2564 8907 2567
rect 9493 2567 9551 2573
rect 9493 2564 9505 2567
rect 8895 2536 9505 2564
rect 8895 2533 8907 2536
rect 8849 2527 8907 2533
rect 9493 2533 9505 2536
rect 9539 2533 9551 2567
rect 9493 2527 9551 2533
rect 10036 2567 10094 2573
rect 10036 2533 10048 2567
rect 10082 2564 10094 2567
rect 11330 2564 11336 2576
rect 10082 2536 11336 2564
rect 10082 2533 10094 2536
rect 10036 2527 10094 2533
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6656 2468 6929 2496
rect 6273 2459 6331 2465
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 9508 2496 9536 2527
rect 11330 2524 11336 2536
rect 11388 2524 11394 2576
rect 13170 2573 13176 2576
rect 12069 2567 12127 2573
rect 12069 2533 12081 2567
rect 12115 2564 12127 2567
rect 13164 2564 13176 2573
rect 12115 2536 13176 2564
rect 12115 2533 12127 2536
rect 12069 2527 12127 2533
rect 13164 2527 13176 2536
rect 13170 2524 13176 2527
rect 13228 2524 13234 2576
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9508 2468 9781 2496
rect 6917 2459 6975 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 10778 2496 10784 2508
rect 9815 2468 10784 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 12897 2499 12955 2505
rect 12897 2465 12909 2499
rect 12943 2496 12955 2499
rect 13280 2496 13308 2604
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14277 2635 14335 2641
rect 14277 2632 14289 2635
rect 13872 2604 14289 2632
rect 13872 2592 13878 2604
rect 14277 2601 14289 2604
rect 14323 2632 14335 2635
rect 14550 2632 14556 2644
rect 14323 2604 14556 2632
rect 14323 2601 14335 2604
rect 14277 2595 14335 2601
rect 14550 2592 14556 2604
rect 14608 2592 14614 2644
rect 16850 2632 16856 2644
rect 16763 2604 16856 2632
rect 16850 2592 16856 2604
rect 16908 2632 16914 2644
rect 17586 2632 17592 2644
rect 16908 2604 17592 2632
rect 16908 2592 16914 2604
rect 17586 2592 17592 2604
rect 17644 2592 17650 2644
rect 18046 2632 18052 2644
rect 18007 2604 18052 2632
rect 18046 2592 18052 2604
rect 18104 2632 18110 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18104 2604 18797 2632
rect 18104 2592 18110 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 21174 2632 21180 2644
rect 21135 2604 21180 2632
rect 18785 2595 18843 2601
rect 21174 2592 21180 2604
rect 21232 2592 21238 2644
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 21818 2632 21824 2644
rect 21692 2604 21824 2632
rect 21692 2592 21698 2604
rect 21818 2592 21824 2604
rect 21876 2592 21882 2644
rect 23198 2592 23204 2644
rect 23256 2632 23262 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 23256 2604 23305 2632
rect 23256 2592 23262 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 23566 2592 23572 2644
rect 23624 2632 23630 2644
rect 23661 2635 23719 2641
rect 23661 2632 23673 2635
rect 23624 2604 23673 2632
rect 23624 2592 23630 2604
rect 23661 2601 23673 2604
rect 23707 2601 23719 2635
rect 23661 2595 23719 2601
rect 24029 2635 24087 2641
rect 24029 2601 24041 2635
rect 24075 2632 24087 2635
rect 24118 2632 24124 2644
rect 24075 2604 24124 2632
rect 24075 2601 24087 2604
rect 24029 2595 24087 2601
rect 24118 2592 24124 2604
rect 24176 2592 24182 2644
rect 24946 2592 24952 2644
rect 25004 2632 25010 2644
rect 25409 2635 25467 2641
rect 25409 2632 25421 2635
rect 25004 2604 25421 2632
rect 25004 2592 25010 2604
rect 25409 2601 25421 2604
rect 25455 2601 25467 2635
rect 25409 2595 25467 2601
rect 25777 2635 25835 2641
rect 25777 2601 25789 2635
rect 25823 2632 25835 2635
rect 25866 2632 25872 2644
rect 25823 2604 25872 2632
rect 25823 2601 25835 2604
rect 25777 2595 25835 2601
rect 25866 2592 25872 2604
rect 25924 2592 25930 2644
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 14921 2567 14979 2573
rect 14921 2564 14933 2567
rect 14884 2536 14933 2564
rect 14884 2524 14890 2536
rect 14921 2533 14933 2536
rect 14967 2564 14979 2567
rect 15740 2567 15798 2573
rect 15740 2564 15752 2567
rect 14967 2536 15752 2564
rect 14967 2533 14979 2536
rect 14921 2527 14979 2533
rect 15740 2533 15752 2536
rect 15786 2564 15798 2567
rect 16482 2564 16488 2576
rect 15786 2536 16488 2564
rect 15786 2533 15798 2536
rect 15740 2527 15798 2533
rect 16482 2524 16488 2536
rect 16540 2524 16546 2576
rect 19705 2567 19763 2573
rect 19705 2533 19717 2567
rect 19751 2564 19763 2567
rect 20346 2564 20352 2576
rect 19751 2536 20352 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 12943 2468 13308 2496
rect 12943 2465 12955 2468
rect 12897 2459 12955 2465
rect 15194 2456 15200 2508
rect 15252 2496 15258 2508
rect 15289 2499 15347 2505
rect 15289 2496 15301 2499
rect 15252 2468 15301 2496
rect 15252 2456 15258 2468
rect 15289 2465 15301 2468
rect 15335 2496 15347 2499
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15335 2468 15485 2496
rect 15335 2465 15347 2468
rect 15289 2459 15347 2465
rect 15473 2465 15485 2468
rect 15519 2496 15531 2499
rect 15562 2496 15568 2508
rect 15519 2468 15568 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 18690 2496 18696 2508
rect 17696 2468 18696 2496
rect 1820 2332 3648 2360
rect 1820 2320 1826 2332
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 1946 2292 1952 2304
rect 1907 2264 1952 2292
rect 1946 2252 1952 2264
rect 2004 2252 2010 2304
rect 2866 2252 2872 2304
rect 2924 2292 2930 2304
rect 6270 2292 6276 2304
rect 2924 2264 6276 2292
rect 2924 2252 2930 2264
rect 6270 2252 6276 2264
rect 6328 2252 6334 2304
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11238 2292 11244 2304
rect 11195 2264 11244 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 14458 2252 14464 2304
rect 14516 2292 14522 2304
rect 17696 2301 17724 2468
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19904 2505 19932 2536
rect 20346 2524 20352 2536
rect 20404 2564 20410 2576
rect 22189 2567 22247 2573
rect 22189 2564 22201 2567
rect 20404 2536 22201 2564
rect 20404 2524 20410 2536
rect 22189 2533 22201 2536
rect 22235 2533 22247 2567
rect 22189 2527 22247 2533
rect 19889 2499 19947 2505
rect 19889 2465 19901 2499
rect 19935 2465 19947 2499
rect 19889 2459 19947 2465
rect 21545 2499 21603 2505
rect 21545 2465 21557 2499
rect 21591 2465 21603 2499
rect 21545 2459 21603 2465
rect 18782 2388 18788 2440
rect 18840 2428 18846 2440
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18840 2400 18889 2428
rect 18840 2388 18846 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19794 2320 19800 2372
rect 19852 2360 19858 2372
rect 20533 2363 20591 2369
rect 20533 2360 20545 2363
rect 19852 2332 20545 2360
rect 19852 2320 19858 2332
rect 20533 2329 20545 2332
rect 20579 2360 20591 2363
rect 21560 2360 21588 2459
rect 21634 2456 21640 2508
rect 21692 2496 21698 2508
rect 22370 2496 22376 2508
rect 21692 2468 22376 2496
rect 21692 2456 21698 2468
rect 22370 2456 22376 2468
rect 22428 2456 22434 2508
rect 22741 2499 22799 2505
rect 22741 2465 22753 2499
rect 22787 2496 22799 2499
rect 23216 2496 23244 2592
rect 24397 2567 24455 2573
rect 24397 2564 24409 2567
rect 24044 2536 24409 2564
rect 24044 2508 24072 2536
rect 24397 2533 24409 2536
rect 24443 2564 24455 2567
rect 26421 2567 26479 2573
rect 26421 2564 26433 2567
rect 24443 2536 26433 2564
rect 24443 2533 24455 2536
rect 24397 2527 24455 2533
rect 26421 2533 26433 2536
rect 26467 2533 26479 2567
rect 26421 2527 26479 2533
rect 22787 2468 23244 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 24026 2456 24032 2508
rect 24084 2456 24090 2508
rect 24118 2456 24124 2508
rect 24176 2496 24182 2508
rect 24762 2496 24768 2508
rect 24176 2468 24768 2496
rect 24176 2456 24182 2468
rect 24762 2456 24768 2468
rect 24820 2456 24826 2508
rect 25593 2499 25651 2505
rect 25593 2465 25605 2499
rect 25639 2496 25651 2499
rect 26050 2496 26056 2508
rect 25639 2468 26056 2496
rect 25639 2465 25651 2468
rect 25593 2459 25651 2465
rect 26050 2456 26056 2468
rect 26108 2456 26114 2508
rect 21818 2428 21824 2440
rect 21779 2400 21824 2428
rect 21818 2388 21824 2400
rect 21876 2428 21882 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 21876 2400 22569 2428
rect 21876 2388 21882 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 23658 2388 23664 2440
rect 23716 2428 23722 2440
rect 24489 2431 24547 2437
rect 24489 2428 24501 2431
rect 23716 2400 24501 2428
rect 23716 2388 23722 2400
rect 24489 2397 24501 2400
rect 24535 2397 24547 2431
rect 24489 2391 24547 2397
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 24857 2431 24915 2437
rect 24857 2428 24869 2431
rect 24719 2400 24869 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 24857 2397 24869 2400
rect 24903 2397 24915 2431
rect 24857 2391 24915 2397
rect 20579 2332 21588 2360
rect 24504 2360 24532 2391
rect 26053 2363 26111 2369
rect 26053 2360 26065 2363
rect 24504 2332 26065 2360
rect 20579 2329 20591 2332
rect 20533 2323 20591 2329
rect 26053 2329 26065 2332
rect 26099 2329 26111 2363
rect 26053 2323 26111 2329
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 14516 2264 17693 2292
rect 14516 2252 14522 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 18322 2292 18328 2304
rect 18283 2264 18328 2292
rect 17681 2255 17739 2261
rect 18322 2252 18328 2264
rect 18380 2252 18386 2304
rect 19886 2252 19892 2304
rect 19944 2292 19950 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 19944 2264 20085 2292
rect 19944 2252 19950 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20898 2292 20904 2304
rect 20859 2264 20904 2292
rect 20073 2255 20131 2261
rect 20898 2252 20904 2264
rect 20956 2292 20962 2304
rect 21634 2292 21640 2304
rect 20956 2264 21640 2292
rect 20956 2252 20962 2264
rect 21634 2252 21640 2264
rect 21692 2252 21698 2304
rect 22922 2292 22928 2304
rect 22883 2264 22928 2292
rect 22922 2252 22928 2264
rect 22980 2252 22986 2304
rect 23842 2252 23848 2304
rect 23900 2292 23906 2304
rect 24857 2295 24915 2301
rect 24857 2292 24869 2295
rect 23900 2264 24869 2292
rect 23900 2252 23906 2264
rect 24857 2261 24869 2264
rect 24903 2292 24915 2295
rect 25041 2295 25099 2301
rect 25041 2292 25053 2295
rect 24903 2264 25053 2292
rect 24903 2261 24915 2264
rect 24857 2255 24915 2261
rect 25041 2261 25053 2264
rect 25087 2261 25099 2295
rect 25041 2255 25099 2261
rect 1104 2202 26864 2224
rect 1104 2150 5648 2202
rect 5700 2150 5712 2202
rect 5764 2150 5776 2202
rect 5828 2150 5840 2202
rect 5892 2150 14982 2202
rect 15034 2150 15046 2202
rect 15098 2150 15110 2202
rect 15162 2150 15174 2202
rect 15226 2150 24315 2202
rect 24367 2150 24379 2202
rect 24431 2150 24443 2202
rect 24495 2150 24507 2202
rect 24559 2150 26864 2202
rect 1104 2128 26864 2150
rect 12894 2048 12900 2100
rect 12952 2088 12958 2100
rect 15378 2088 15384 2100
rect 12952 2060 15384 2088
rect 12952 2048 12958 2060
rect 15378 2048 15384 2060
rect 15436 2048 15442 2100
rect 13262 1980 13268 2032
rect 13320 2020 13326 2032
rect 17126 2020 17132 2032
rect 13320 1992 17132 2020
rect 13320 1980 13326 1992
rect 17126 1980 17132 1992
rect 17184 1980 17190 2032
rect 12066 1572 12072 1624
rect 12124 1612 12130 1624
rect 12526 1612 12532 1624
rect 12124 1584 12532 1612
rect 12124 1572 12130 1584
rect 12526 1572 12532 1584
rect 12584 1572 12590 1624
rect 6546 1504 6552 1556
rect 6604 1544 6610 1556
rect 9214 1544 9220 1556
rect 6604 1516 9220 1544
rect 6604 1504 6610 1516
rect 9214 1504 9220 1516
rect 9272 1504 9278 1556
rect 3418 1436 3424 1488
rect 3476 1476 3482 1488
rect 4522 1476 4528 1488
rect 3476 1448 4528 1476
rect 3476 1436 3482 1448
rect 4522 1436 4528 1448
rect 4580 1436 4586 1488
<< via1 >>
rect 18236 26664 18288 26716
rect 24768 26664 24820 26716
rect 22008 26392 22060 26444
rect 24768 26392 24820 26444
rect 10048 26188 10100 26240
rect 16580 26188 16632 26240
rect 6368 26120 6420 26172
rect 17408 26120 17460 26172
rect 9128 26052 9180 26104
rect 23480 26052 23532 26104
rect 11244 25984 11296 26036
rect 20352 25984 20404 26036
rect 6920 25916 6972 25968
rect 9496 25916 9548 25968
rect 12164 25916 12216 25968
rect 19432 25916 19484 25968
rect 1768 25848 1820 25900
rect 11980 25848 12032 25900
rect 13452 25848 13504 25900
rect 18972 25848 19024 25900
rect 6092 25780 6144 25832
rect 9496 25780 9548 25832
rect 10968 25780 11020 25832
rect 21364 25780 21416 25832
rect 10784 25712 10836 25764
rect 19340 25712 19392 25764
rect 4896 25644 4948 25696
rect 14004 25644 14056 25696
rect 15476 25644 15528 25696
rect 24676 25644 24728 25696
rect 10315 25542 10367 25594
rect 10379 25542 10431 25594
rect 10443 25542 10495 25594
rect 10507 25542 10559 25594
rect 19648 25542 19700 25594
rect 19712 25542 19764 25594
rect 19776 25542 19828 25594
rect 19840 25542 19892 25594
rect 3240 25440 3292 25492
rect 7840 25440 7892 25492
rect 10968 25483 11020 25492
rect 6276 25372 6328 25424
rect 2136 25304 2188 25356
rect 3424 25304 3476 25356
rect 4160 25304 4212 25356
rect 5172 25279 5224 25288
rect 5172 25245 5181 25279
rect 5181 25245 5215 25279
rect 5215 25245 5224 25279
rect 5172 25236 5224 25245
rect 3056 25168 3108 25220
rect 5080 25168 5132 25220
rect 5264 25168 5316 25220
rect 8116 25279 8168 25288
rect 8116 25245 8125 25279
rect 8125 25245 8159 25279
rect 8159 25245 8168 25279
rect 8116 25236 8168 25245
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 10968 25449 10977 25483
rect 10977 25449 11011 25483
rect 11011 25449 11020 25483
rect 10968 25440 11020 25449
rect 11060 25440 11112 25492
rect 12440 25372 12492 25424
rect 18328 25440 18380 25492
rect 22376 25440 22428 25492
rect 11244 25304 11296 25356
rect 10968 25236 11020 25288
rect 11060 25236 11112 25288
rect 13084 25279 13136 25288
rect 8024 25168 8076 25220
rect 8300 25168 8352 25220
rect 10048 25211 10100 25220
rect 10048 25177 10057 25211
rect 10057 25177 10091 25211
rect 10091 25177 10100 25211
rect 10048 25168 10100 25177
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 15292 25304 15344 25356
rect 15384 25236 15436 25288
rect 11796 25168 11848 25220
rect 17868 25372 17920 25424
rect 24860 25372 24912 25424
rect 17132 25304 17184 25356
rect 21088 25304 21140 25356
rect 16948 25279 17000 25288
rect 16948 25245 16957 25279
rect 16957 25245 16991 25279
rect 16991 25245 17000 25279
rect 16948 25236 17000 25245
rect 17224 25236 17276 25288
rect 19064 25279 19116 25288
rect 19064 25245 19073 25279
rect 19073 25245 19107 25279
rect 19107 25245 19116 25279
rect 19064 25236 19116 25245
rect 19156 25279 19208 25288
rect 19156 25245 19165 25279
rect 19165 25245 19199 25279
rect 19199 25245 19208 25279
rect 19156 25236 19208 25245
rect 19340 25236 19392 25288
rect 22836 25236 22888 25288
rect 25780 25168 25832 25220
rect 1400 25100 1452 25152
rect 2044 25143 2096 25152
rect 2044 25109 2053 25143
rect 2053 25109 2087 25143
rect 2087 25109 2096 25143
rect 2044 25100 2096 25109
rect 3516 25100 3568 25152
rect 3700 25143 3752 25152
rect 3700 25109 3709 25143
rect 3709 25109 3743 25143
rect 3743 25109 3752 25143
rect 3700 25100 3752 25109
rect 3976 25100 4028 25152
rect 4988 25143 5040 25152
rect 4988 25109 4997 25143
rect 4997 25109 5031 25143
rect 5031 25109 5040 25143
rect 4988 25100 5040 25109
rect 5356 25100 5408 25152
rect 7104 25100 7156 25152
rect 7932 25100 7984 25152
rect 8944 25100 8996 25152
rect 12256 25100 12308 25152
rect 14372 25100 14424 25152
rect 14740 25100 14792 25152
rect 15844 25143 15896 25152
rect 15844 25109 15853 25143
rect 15853 25109 15887 25143
rect 15887 25109 15896 25143
rect 15844 25100 15896 25109
rect 16120 25100 16172 25152
rect 16764 25100 16816 25152
rect 18236 25100 18288 25152
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 19708 25143 19760 25152
rect 19708 25109 19717 25143
rect 19717 25109 19751 25143
rect 19751 25109 19760 25143
rect 19708 25100 19760 25109
rect 5648 24998 5700 25050
rect 5712 24998 5764 25050
rect 5776 24998 5828 25050
rect 5840 24998 5892 25050
rect 14982 24998 15034 25050
rect 15046 24998 15098 25050
rect 15110 24998 15162 25050
rect 15174 24998 15226 25050
rect 24315 24998 24367 25050
rect 24379 24998 24431 25050
rect 24443 24998 24495 25050
rect 24507 24998 24559 25050
rect 3056 24896 3108 24948
rect 6644 24939 6696 24948
rect 6644 24905 6653 24939
rect 6653 24905 6687 24939
rect 6687 24905 6696 24939
rect 6644 24896 6696 24905
rect 8024 24896 8076 24948
rect 1768 24828 1820 24880
rect 4436 24828 4488 24880
rect 1584 24692 1636 24744
rect 2504 24735 2556 24744
rect 2504 24701 2513 24735
rect 2513 24701 2547 24735
rect 2547 24701 2556 24735
rect 3424 24803 3476 24812
rect 3424 24769 3433 24803
rect 3433 24769 3467 24803
rect 3467 24769 3476 24803
rect 3424 24760 3476 24769
rect 4160 24803 4212 24812
rect 4160 24769 4169 24803
rect 4169 24769 4203 24803
rect 4203 24769 4212 24803
rect 4160 24760 4212 24769
rect 4896 24760 4948 24812
rect 8116 24828 8168 24880
rect 2504 24692 2556 24701
rect 2780 24692 2832 24744
rect 4988 24735 5040 24744
rect 2964 24624 3016 24676
rect 4988 24701 4997 24735
rect 4997 24701 5031 24735
rect 5031 24701 5040 24735
rect 4988 24692 5040 24701
rect 7104 24735 7156 24744
rect 7104 24701 7113 24735
rect 7113 24701 7147 24735
rect 7147 24701 7156 24735
rect 7104 24692 7156 24701
rect 8392 24692 8444 24744
rect 8944 24692 8996 24744
rect 12072 24896 12124 24948
rect 19064 24896 19116 24948
rect 24768 24896 24820 24948
rect 9864 24828 9916 24880
rect 15016 24828 15068 24880
rect 15292 24828 15344 24880
rect 16396 24828 16448 24880
rect 9956 24760 10008 24812
rect 11980 24760 12032 24812
rect 12256 24760 12308 24812
rect 12624 24760 12676 24812
rect 13636 24760 13688 24812
rect 14372 24760 14424 24812
rect 15752 24760 15804 24812
rect 9864 24692 9916 24744
rect 12348 24692 12400 24744
rect 12532 24692 12584 24744
rect 7840 24624 7892 24676
rect 2136 24556 2188 24608
rect 2688 24599 2740 24608
rect 2688 24565 2697 24599
rect 2697 24565 2731 24599
rect 2731 24565 2740 24599
rect 2688 24556 2740 24565
rect 4436 24599 4488 24608
rect 4436 24565 4445 24599
rect 4445 24565 4479 24599
rect 4479 24565 4488 24599
rect 4436 24556 4488 24565
rect 5080 24599 5132 24608
rect 5080 24565 5089 24599
rect 5089 24565 5123 24599
rect 5123 24565 5132 24599
rect 5080 24556 5132 24565
rect 6000 24599 6052 24608
rect 6000 24565 6009 24599
rect 6009 24565 6043 24599
rect 6043 24565 6052 24599
rect 6000 24556 6052 24565
rect 7288 24599 7340 24608
rect 7288 24565 7297 24599
rect 7297 24565 7331 24599
rect 7331 24565 7340 24599
rect 7288 24556 7340 24565
rect 8116 24599 8168 24608
rect 8116 24565 8125 24599
rect 8125 24565 8159 24599
rect 8159 24565 8168 24599
rect 8116 24556 8168 24565
rect 11980 24624 12032 24676
rect 13176 24624 13228 24676
rect 14004 24667 14056 24676
rect 14004 24633 14013 24667
rect 14013 24633 14047 24667
rect 14047 24633 14056 24667
rect 15844 24692 15896 24744
rect 19708 24828 19760 24880
rect 20996 24828 21048 24880
rect 24216 24828 24268 24880
rect 17868 24803 17920 24812
rect 17868 24769 17877 24803
rect 17877 24769 17911 24803
rect 17911 24769 17920 24803
rect 17868 24760 17920 24769
rect 17132 24735 17184 24744
rect 17132 24701 17141 24735
rect 17141 24701 17175 24735
rect 17175 24701 17184 24735
rect 17132 24692 17184 24701
rect 17224 24692 17276 24744
rect 19156 24760 19208 24812
rect 20444 24760 20496 24812
rect 18052 24692 18104 24744
rect 18512 24692 18564 24744
rect 14004 24624 14056 24633
rect 8300 24556 8352 24608
rect 9772 24599 9824 24608
rect 9772 24565 9781 24599
rect 9781 24565 9815 24599
rect 9815 24565 9824 24599
rect 9772 24556 9824 24565
rect 11060 24599 11112 24608
rect 11060 24565 11069 24599
rect 11069 24565 11103 24599
rect 11103 24565 11112 24599
rect 11060 24556 11112 24565
rect 12716 24556 12768 24608
rect 13728 24556 13780 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 14464 24599 14516 24608
rect 14464 24565 14473 24599
rect 14473 24565 14507 24599
rect 14507 24565 14516 24599
rect 14464 24556 14516 24565
rect 14648 24556 14700 24608
rect 15660 24556 15712 24608
rect 17316 24624 17368 24676
rect 19708 24624 19760 24676
rect 20168 24624 20220 24676
rect 21180 24692 21232 24744
rect 23940 24735 23992 24744
rect 23940 24701 23949 24735
rect 23949 24701 23983 24735
rect 23983 24701 23992 24735
rect 23940 24692 23992 24701
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 17868 24556 17920 24608
rect 18236 24556 18288 24608
rect 19524 24556 19576 24608
rect 20260 24556 20312 24608
rect 27252 24624 27304 24676
rect 20628 24599 20680 24608
rect 20628 24565 20637 24599
rect 20637 24565 20671 24599
rect 20671 24565 20680 24599
rect 20628 24556 20680 24565
rect 21088 24556 21140 24608
rect 21824 24599 21876 24608
rect 21824 24565 21833 24599
rect 21833 24565 21867 24599
rect 21867 24565 21876 24599
rect 21824 24556 21876 24565
rect 24216 24556 24268 24608
rect 10315 24454 10367 24506
rect 10379 24454 10431 24506
rect 10443 24454 10495 24506
rect 10507 24454 10559 24506
rect 19648 24454 19700 24506
rect 19712 24454 19764 24506
rect 19776 24454 19828 24506
rect 19840 24454 19892 24506
rect 2412 24352 2464 24404
rect 4988 24352 5040 24404
rect 9680 24352 9732 24404
rect 1952 24284 2004 24336
rect 5356 24284 5408 24336
rect 9956 24284 10008 24336
rect 13084 24352 13136 24404
rect 13452 24395 13504 24404
rect 13452 24361 13461 24395
rect 13461 24361 13495 24395
rect 13495 24361 13504 24395
rect 13452 24352 13504 24361
rect 15476 24395 15528 24404
rect 15476 24361 15485 24395
rect 15485 24361 15519 24395
rect 15519 24361 15528 24395
rect 15476 24352 15528 24361
rect 18604 24395 18656 24404
rect 18604 24361 18613 24395
rect 18613 24361 18647 24395
rect 18647 24361 18656 24395
rect 18604 24352 18656 24361
rect 19984 24352 20036 24404
rect 21364 24395 21416 24404
rect 21364 24361 21373 24395
rect 21373 24361 21407 24395
rect 21407 24361 21416 24395
rect 21364 24352 21416 24361
rect 24124 24352 24176 24404
rect 24676 24395 24728 24404
rect 24676 24361 24685 24395
rect 24685 24361 24719 24395
rect 24719 24361 24728 24395
rect 24676 24352 24728 24361
rect 11336 24284 11388 24336
rect 14464 24284 14516 24336
rect 15108 24327 15160 24336
rect 15108 24293 15117 24327
rect 15117 24293 15151 24327
rect 15151 24293 15160 24327
rect 15108 24284 15160 24293
rect 15200 24284 15252 24336
rect 16212 24284 16264 24336
rect 16948 24327 17000 24336
rect 16948 24293 16957 24327
rect 16957 24293 16991 24327
rect 16991 24293 17000 24327
rect 16948 24284 17000 24293
rect 20628 24284 20680 24336
rect 5172 24216 5224 24268
rect 6184 24216 6236 24268
rect 7196 24216 7248 24268
rect 13360 24259 13412 24268
rect 13360 24225 13369 24259
rect 13369 24225 13403 24259
rect 13403 24225 13412 24259
rect 13360 24216 13412 24225
rect 13912 24216 13964 24268
rect 14372 24216 14424 24268
rect 14832 24216 14884 24268
rect 15292 24259 15344 24268
rect 15292 24225 15301 24259
rect 15301 24225 15335 24259
rect 15335 24225 15344 24259
rect 15292 24216 15344 24225
rect 19156 24259 19208 24268
rect 2504 24148 2556 24200
rect 3332 24148 3384 24200
rect 3424 24148 3476 24200
rect 4068 24080 4120 24132
rect 4252 24148 4304 24200
rect 5908 24191 5960 24200
rect 1768 24012 1820 24064
rect 3148 24055 3200 24064
rect 3148 24021 3157 24055
rect 3157 24021 3191 24055
rect 3191 24021 3200 24055
rect 3148 24012 3200 24021
rect 4160 24012 4212 24064
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 6552 24148 6604 24200
rect 10508 24191 10560 24200
rect 10508 24157 10517 24191
rect 10517 24157 10551 24191
rect 10551 24157 10560 24191
rect 10508 24148 10560 24157
rect 11520 24148 11572 24200
rect 12256 24148 12308 24200
rect 13452 24148 13504 24200
rect 13636 24191 13688 24200
rect 13636 24157 13645 24191
rect 13645 24157 13679 24191
rect 13679 24157 13688 24191
rect 13636 24148 13688 24157
rect 13268 24080 13320 24132
rect 14832 24080 14884 24132
rect 16948 24080 17000 24132
rect 17500 24148 17552 24200
rect 19156 24225 19165 24259
rect 19165 24225 19199 24259
rect 19199 24225 19208 24259
rect 19156 24216 19208 24225
rect 19708 24259 19760 24268
rect 19708 24225 19717 24259
rect 19717 24225 19751 24259
rect 19751 24225 19760 24259
rect 19708 24216 19760 24225
rect 21548 24216 21600 24268
rect 22652 24216 22704 24268
rect 24676 24216 24728 24268
rect 20168 24148 20220 24200
rect 20352 24148 20404 24200
rect 17684 24123 17736 24132
rect 17684 24089 17693 24123
rect 17693 24089 17727 24123
rect 17727 24089 17736 24123
rect 17684 24080 17736 24089
rect 18052 24123 18104 24132
rect 18052 24089 18061 24123
rect 18061 24089 18095 24123
rect 18095 24089 18104 24123
rect 18052 24080 18104 24089
rect 19340 24080 19392 24132
rect 19984 24080 20036 24132
rect 20444 24080 20496 24132
rect 20904 24123 20956 24132
rect 20904 24089 20913 24123
rect 20913 24089 20947 24123
rect 20947 24089 20956 24123
rect 20904 24080 20956 24089
rect 6000 24012 6052 24064
rect 7288 24012 7340 24064
rect 7564 24012 7616 24064
rect 9312 24012 9364 24064
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 9956 24055 10008 24064
rect 9956 24021 9965 24055
rect 9965 24021 9999 24055
rect 9999 24021 10008 24055
rect 9956 24012 10008 24021
rect 11244 24012 11296 24064
rect 11428 24012 11480 24064
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 14464 24012 14516 24064
rect 15752 24012 15804 24064
rect 16580 24055 16632 24064
rect 16580 24021 16589 24055
rect 16589 24021 16623 24055
rect 16623 24021 16632 24055
rect 16580 24012 16632 24021
rect 17224 24012 17276 24064
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 5648 23910 5700 23962
rect 5712 23910 5764 23962
rect 5776 23910 5828 23962
rect 5840 23910 5892 23962
rect 14982 23910 15034 23962
rect 15046 23910 15098 23962
rect 15110 23910 15162 23962
rect 15174 23910 15226 23962
rect 24315 23910 24367 23962
rect 24379 23910 24431 23962
rect 24443 23910 24495 23962
rect 24507 23910 24559 23962
rect 3516 23808 3568 23860
rect 6184 23851 6236 23860
rect 6184 23817 6193 23851
rect 6193 23817 6227 23851
rect 6227 23817 6236 23851
rect 6184 23808 6236 23817
rect 6552 23851 6604 23860
rect 6552 23817 6561 23851
rect 6561 23817 6595 23851
rect 6595 23817 6604 23851
rect 6552 23808 6604 23817
rect 2044 23672 2096 23724
rect 2504 23672 2556 23724
rect 3148 23672 3200 23724
rect 4436 23672 4488 23724
rect 5540 23672 5592 23724
rect 6000 23672 6052 23724
rect 7472 23715 7524 23724
rect 7472 23681 7481 23715
rect 7481 23681 7515 23715
rect 7515 23681 7524 23715
rect 7472 23672 7524 23681
rect 9956 23808 10008 23860
rect 12256 23851 12308 23860
rect 12256 23817 12265 23851
rect 12265 23817 12299 23851
rect 12299 23817 12308 23851
rect 12256 23808 12308 23817
rect 10968 23740 11020 23792
rect 11796 23740 11848 23792
rect 11244 23715 11296 23724
rect 11244 23681 11253 23715
rect 11253 23681 11287 23715
rect 11287 23681 11296 23715
rect 11244 23672 11296 23681
rect 11428 23715 11480 23724
rect 11428 23681 11437 23715
rect 11437 23681 11471 23715
rect 11471 23681 11480 23715
rect 11428 23672 11480 23681
rect 13636 23808 13688 23860
rect 14004 23808 14056 23860
rect 14464 23808 14516 23860
rect 20260 23808 20312 23860
rect 20628 23808 20680 23860
rect 21548 23851 21600 23860
rect 21548 23817 21557 23851
rect 21557 23817 21591 23851
rect 21591 23817 21600 23851
rect 21548 23808 21600 23817
rect 21916 23808 21968 23860
rect 24768 23851 24820 23860
rect 24768 23817 24777 23851
rect 24777 23817 24811 23851
rect 24811 23817 24820 23851
rect 24768 23808 24820 23817
rect 15200 23783 15252 23792
rect 15200 23749 15209 23783
rect 15209 23749 15243 23783
rect 15243 23749 15252 23783
rect 15200 23740 15252 23749
rect 16304 23740 16356 23792
rect 16488 23740 16540 23792
rect 8300 23604 8352 23656
rect 10508 23604 10560 23656
rect 10784 23604 10836 23656
rect 12348 23604 12400 23656
rect 12532 23604 12584 23656
rect 20444 23672 20496 23724
rect 24308 23672 24360 23724
rect 24676 23672 24728 23724
rect 15568 23647 15620 23656
rect 15568 23613 15591 23647
rect 15591 23613 15620 23647
rect 15568 23604 15620 23613
rect 16488 23604 16540 23656
rect 18696 23604 18748 23656
rect 2228 23536 2280 23588
rect 6092 23536 6144 23588
rect 9312 23536 9364 23588
rect 12624 23536 12676 23588
rect 18604 23536 18656 23588
rect 1492 23468 1544 23520
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 2780 23468 2832 23477
rect 3332 23468 3384 23520
rect 3700 23468 3752 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 8576 23468 8628 23520
rect 9680 23468 9732 23520
rect 11152 23511 11204 23520
rect 11152 23477 11161 23511
rect 11161 23477 11195 23511
rect 11195 23477 11204 23511
rect 11152 23468 11204 23477
rect 13820 23511 13872 23520
rect 13820 23477 13829 23511
rect 13829 23477 13863 23511
rect 13863 23477 13872 23511
rect 13820 23468 13872 23477
rect 16948 23468 17000 23520
rect 17500 23511 17552 23520
rect 17500 23477 17509 23511
rect 17509 23477 17543 23511
rect 17543 23477 17552 23511
rect 17500 23468 17552 23477
rect 19524 23468 19576 23520
rect 19708 23536 19760 23588
rect 20628 23536 20680 23588
rect 20720 23536 20772 23588
rect 22008 23536 22060 23588
rect 20996 23511 21048 23520
rect 20996 23477 21005 23511
rect 21005 23477 21039 23511
rect 21039 23477 21048 23511
rect 20996 23468 21048 23477
rect 21916 23511 21968 23520
rect 21916 23477 21925 23511
rect 21925 23477 21959 23511
rect 21959 23477 21968 23511
rect 22652 23511 22704 23520
rect 21916 23468 21968 23477
rect 22652 23477 22661 23511
rect 22661 23477 22695 23511
rect 22695 23477 22704 23511
rect 22652 23468 22704 23477
rect 24492 23511 24544 23520
rect 24492 23477 24501 23511
rect 24501 23477 24535 23511
rect 24535 23477 24544 23511
rect 24492 23468 24544 23477
rect 10315 23366 10367 23418
rect 10379 23366 10431 23418
rect 10443 23366 10495 23418
rect 10507 23366 10559 23418
rect 19648 23366 19700 23418
rect 19712 23366 19764 23418
rect 19776 23366 19828 23418
rect 19840 23366 19892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 1676 23264 1728 23316
rect 1952 23264 2004 23316
rect 2412 23307 2464 23316
rect 2412 23273 2421 23307
rect 2421 23273 2455 23307
rect 2455 23273 2464 23307
rect 2412 23264 2464 23273
rect 2872 23264 2924 23316
rect 3332 23307 3384 23316
rect 3332 23273 3341 23307
rect 3341 23273 3375 23307
rect 3375 23273 3384 23307
rect 3332 23264 3384 23273
rect 4252 23264 4304 23316
rect 4528 23307 4580 23316
rect 4528 23273 4537 23307
rect 4537 23273 4571 23307
rect 4571 23273 4580 23307
rect 4528 23264 4580 23273
rect 7196 23307 7248 23316
rect 7196 23273 7205 23307
rect 7205 23273 7239 23307
rect 7239 23273 7248 23307
rect 7196 23264 7248 23273
rect 3608 23196 3660 23248
rect 3424 23128 3476 23180
rect 5448 23196 5500 23248
rect 9772 23264 9824 23316
rect 10140 23307 10192 23316
rect 10140 23273 10149 23307
rect 10149 23273 10183 23307
rect 10183 23273 10192 23307
rect 10140 23264 10192 23273
rect 12808 23307 12860 23316
rect 12808 23273 12817 23307
rect 12817 23273 12851 23307
rect 12851 23273 12860 23307
rect 12808 23264 12860 23273
rect 13084 23264 13136 23316
rect 15568 23264 15620 23316
rect 16672 23264 16724 23316
rect 18144 23264 18196 23316
rect 20444 23264 20496 23316
rect 20720 23264 20772 23316
rect 22008 23307 22060 23316
rect 22008 23273 22017 23307
rect 22017 23273 22051 23307
rect 22051 23273 22060 23307
rect 22008 23264 22060 23273
rect 22836 23264 22888 23316
rect 24768 23307 24820 23316
rect 24768 23273 24777 23307
rect 24777 23273 24811 23307
rect 24811 23273 24820 23307
rect 24768 23264 24820 23273
rect 8576 23196 8628 23248
rect 6000 23128 6052 23180
rect 2412 23060 2464 23112
rect 2412 22924 2464 22976
rect 2780 22924 2832 22976
rect 3608 22992 3660 23044
rect 8024 23035 8076 23044
rect 8024 23001 8033 23035
rect 8033 23001 8067 23035
rect 8067 23001 8076 23035
rect 8024 22992 8076 23001
rect 8484 23103 8536 23112
rect 8484 23069 8493 23103
rect 8493 23069 8527 23103
rect 8527 23069 8536 23103
rect 8484 23060 8536 23069
rect 9496 23171 9548 23180
rect 9496 23137 9505 23171
rect 9505 23137 9539 23171
rect 9539 23137 9548 23171
rect 9496 23128 9548 23137
rect 9312 23060 9364 23112
rect 10968 23196 11020 23248
rect 11796 23196 11848 23248
rect 13912 23239 13964 23248
rect 13912 23205 13921 23239
rect 13921 23205 13955 23239
rect 13955 23205 13964 23239
rect 13912 23196 13964 23205
rect 16948 23196 17000 23248
rect 23480 23239 23532 23248
rect 23480 23205 23489 23239
rect 23489 23205 23523 23239
rect 23523 23205 23532 23239
rect 23480 23196 23532 23205
rect 11060 23128 11112 23180
rect 13544 23128 13596 23180
rect 15384 23128 15436 23180
rect 19340 23128 19392 23180
rect 20168 23128 20220 23180
rect 20444 23128 20496 23180
rect 21640 23128 21692 23180
rect 22836 23171 22888 23180
rect 22836 23137 22845 23171
rect 22845 23137 22879 23171
rect 22879 23137 22888 23171
rect 22836 23128 22888 23137
rect 24676 23128 24728 23180
rect 11152 23060 11204 23112
rect 12164 23060 12216 23112
rect 13728 23060 13780 23112
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 16488 23060 16540 23069
rect 19524 23103 19576 23112
rect 19524 23069 19533 23103
rect 19533 23069 19567 23103
rect 19567 23069 19576 23103
rect 19524 23060 19576 23069
rect 20904 23060 20956 23112
rect 21456 23103 21508 23112
rect 21456 23069 21465 23103
rect 21465 23069 21499 23103
rect 21499 23069 21508 23103
rect 23020 23103 23072 23112
rect 21456 23060 21508 23069
rect 23020 23069 23029 23103
rect 23029 23069 23063 23103
rect 23063 23069 23072 23103
rect 23020 23060 23072 23069
rect 9036 22992 9088 23044
rect 15936 22992 15988 23044
rect 19248 22992 19300 23044
rect 21824 22992 21876 23044
rect 3056 22924 3108 22976
rect 3424 22924 3476 22976
rect 4436 22924 4488 22976
rect 7196 22924 7248 22976
rect 10784 22924 10836 22976
rect 12532 22924 12584 22976
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 16304 22967 16356 22976
rect 16304 22933 16313 22967
rect 16313 22933 16347 22967
rect 16347 22933 16356 22967
rect 16304 22924 16356 22933
rect 17500 22924 17552 22976
rect 18880 22924 18932 22976
rect 20720 22924 20772 22976
rect 22100 22924 22152 22976
rect 23480 22924 23532 22976
rect 5648 22822 5700 22874
rect 5712 22822 5764 22874
rect 5776 22822 5828 22874
rect 5840 22822 5892 22874
rect 14982 22822 15034 22874
rect 15046 22822 15098 22874
rect 15110 22822 15162 22874
rect 15174 22822 15226 22874
rect 24315 22822 24367 22874
rect 24379 22822 24431 22874
rect 24443 22822 24495 22874
rect 24507 22822 24559 22874
rect 1492 22720 1544 22772
rect 1860 22720 1912 22772
rect 2596 22720 2648 22772
rect 2872 22720 2924 22772
rect 3700 22763 3752 22772
rect 3700 22729 3709 22763
rect 3709 22729 3743 22763
rect 3743 22729 3752 22763
rect 3700 22720 3752 22729
rect 5540 22720 5592 22772
rect 8300 22720 8352 22772
rect 2780 22652 2832 22704
rect 1676 22516 1728 22568
rect 2320 22516 2372 22568
rect 3516 22516 3568 22568
rect 1860 22448 1912 22500
rect 2228 22448 2280 22500
rect 3148 22380 3200 22432
rect 6000 22584 6052 22636
rect 7564 22584 7616 22636
rect 9956 22720 10008 22772
rect 11152 22720 11204 22772
rect 11428 22763 11480 22772
rect 11428 22729 11437 22763
rect 11437 22729 11471 22763
rect 11471 22729 11480 22763
rect 11428 22720 11480 22729
rect 12164 22763 12216 22772
rect 12164 22729 12173 22763
rect 12173 22729 12207 22763
rect 12207 22729 12216 22763
rect 12164 22720 12216 22729
rect 12440 22763 12492 22772
rect 12440 22729 12449 22763
rect 12449 22729 12483 22763
rect 12483 22729 12492 22763
rect 12440 22720 12492 22729
rect 13084 22720 13136 22772
rect 15568 22720 15620 22772
rect 17040 22763 17092 22772
rect 17040 22729 17049 22763
rect 17049 22729 17083 22763
rect 17083 22729 17092 22763
rect 17040 22720 17092 22729
rect 18696 22763 18748 22772
rect 18696 22729 18705 22763
rect 18705 22729 18739 22763
rect 18739 22729 18748 22763
rect 18696 22720 18748 22729
rect 22836 22763 22888 22772
rect 11060 22695 11112 22704
rect 11060 22661 11069 22695
rect 11069 22661 11103 22695
rect 11103 22661 11112 22695
rect 11060 22652 11112 22661
rect 11244 22652 11296 22704
rect 13912 22652 13964 22704
rect 17224 22652 17276 22704
rect 20904 22695 20956 22704
rect 20904 22661 20913 22695
rect 20913 22661 20947 22695
rect 20947 22661 20956 22695
rect 20904 22652 20956 22661
rect 20996 22652 21048 22704
rect 12164 22584 12216 22636
rect 12900 22584 12952 22636
rect 15568 22584 15620 22636
rect 15752 22584 15804 22636
rect 18328 22584 18380 22636
rect 5448 22516 5500 22568
rect 11244 22559 11296 22568
rect 11244 22525 11253 22559
rect 11253 22525 11287 22559
rect 11287 22525 11296 22559
rect 11244 22516 11296 22525
rect 12716 22516 12768 22568
rect 13360 22516 13412 22568
rect 14464 22516 14516 22568
rect 14648 22559 14700 22568
rect 14648 22525 14671 22559
rect 14671 22525 14700 22559
rect 16856 22559 16908 22568
rect 14648 22516 14700 22525
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 18696 22516 18748 22568
rect 19156 22559 19208 22568
rect 19156 22525 19190 22559
rect 19190 22525 19208 22559
rect 4436 22448 4488 22500
rect 6736 22448 6788 22500
rect 8116 22491 8168 22500
rect 8116 22457 8125 22491
rect 8125 22457 8159 22491
rect 8159 22457 8168 22491
rect 8852 22491 8904 22500
rect 8116 22448 8168 22457
rect 8852 22457 8886 22491
rect 8886 22457 8904 22491
rect 8852 22448 8904 22457
rect 12992 22448 13044 22500
rect 19156 22516 19208 22525
rect 19524 22516 19576 22568
rect 19984 22516 20036 22568
rect 20904 22516 20956 22568
rect 19064 22448 19116 22500
rect 21456 22584 21508 22636
rect 21732 22516 21784 22568
rect 22008 22516 22060 22568
rect 22836 22729 22845 22763
rect 22845 22729 22879 22763
rect 22879 22729 22888 22763
rect 22836 22720 22888 22729
rect 24124 22720 24176 22772
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 22744 22584 22796 22636
rect 23848 22584 23900 22636
rect 24676 22584 24728 22636
rect 23664 22559 23716 22568
rect 23664 22525 23673 22559
rect 23673 22525 23707 22559
rect 23707 22525 23716 22559
rect 23664 22516 23716 22525
rect 6000 22380 6052 22432
rect 7196 22423 7248 22432
rect 7196 22389 7205 22423
rect 7205 22389 7239 22423
rect 7239 22389 7248 22423
rect 7196 22380 7248 22389
rect 9956 22423 10008 22432
rect 9956 22389 9965 22423
rect 9965 22389 9999 22423
rect 9999 22389 10008 22423
rect 9956 22380 10008 22389
rect 11796 22423 11848 22432
rect 11796 22389 11805 22423
rect 11805 22389 11839 22423
rect 11839 22389 11848 22423
rect 11796 22380 11848 22389
rect 11980 22380 12032 22432
rect 13084 22380 13136 22432
rect 13268 22380 13320 22432
rect 13452 22380 13504 22432
rect 15292 22380 15344 22432
rect 16488 22423 16540 22432
rect 16488 22389 16497 22423
rect 16497 22389 16531 22423
rect 16531 22389 16540 22423
rect 16488 22380 16540 22389
rect 17776 22423 17828 22432
rect 17776 22389 17785 22423
rect 17785 22389 17819 22423
rect 17819 22389 17828 22423
rect 17776 22380 17828 22389
rect 19340 22380 19392 22432
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 23756 22448 23808 22500
rect 23020 22380 23072 22432
rect 24952 22423 25004 22432
rect 24952 22389 24961 22423
rect 24961 22389 24995 22423
rect 24995 22389 25004 22423
rect 24952 22380 25004 22389
rect 10315 22278 10367 22330
rect 10379 22278 10431 22330
rect 10443 22278 10495 22330
rect 10507 22278 10559 22330
rect 19648 22278 19700 22330
rect 19712 22278 19764 22330
rect 19776 22278 19828 22330
rect 19840 22278 19892 22330
rect 2044 22176 2096 22228
rect 5908 22176 5960 22228
rect 6644 22176 6696 22228
rect 9312 22176 9364 22228
rect 2412 22108 2464 22160
rect 4068 22108 4120 22160
rect 7104 22108 7156 22160
rect 8300 22108 8352 22160
rect 8576 22108 8628 22160
rect 10140 22176 10192 22228
rect 10692 22176 10744 22228
rect 12256 22176 12308 22228
rect 12440 22176 12492 22228
rect 12624 22176 12676 22228
rect 12716 22176 12768 22228
rect 12900 22219 12952 22228
rect 12900 22185 12909 22219
rect 12909 22185 12943 22219
rect 12943 22185 12952 22219
rect 12900 22176 12952 22185
rect 13544 22176 13596 22228
rect 17776 22219 17828 22228
rect 2320 22083 2372 22092
rect 2320 22049 2329 22083
rect 2329 22049 2363 22083
rect 2363 22049 2372 22083
rect 2320 22040 2372 22049
rect 4160 22040 4212 22092
rect 5080 22040 5132 22092
rect 6368 22083 6420 22092
rect 6368 22049 6377 22083
rect 6377 22049 6411 22083
rect 6411 22049 6420 22083
rect 6368 22040 6420 22049
rect 6736 22040 6788 22092
rect 7012 22040 7064 22092
rect 7564 22040 7616 22092
rect 9956 22108 10008 22160
rect 13820 22151 13872 22160
rect 9772 22040 9824 22092
rect 9864 22040 9916 22092
rect 11520 22040 11572 22092
rect 13820 22117 13829 22151
rect 13829 22117 13863 22151
rect 13863 22117 13872 22151
rect 13820 22108 13872 22117
rect 14556 22108 14608 22160
rect 15752 22108 15804 22160
rect 17776 22185 17785 22219
rect 17785 22185 17819 22219
rect 17819 22185 17828 22219
rect 17776 22176 17828 22185
rect 19156 22176 19208 22228
rect 21456 22176 21508 22228
rect 19616 22108 19668 22160
rect 20076 22108 20128 22160
rect 15936 22040 15988 22092
rect 16948 22040 17000 22092
rect 18144 22083 18196 22092
rect 18144 22049 18153 22083
rect 18153 22049 18187 22083
rect 18187 22049 18196 22083
rect 18144 22040 18196 22049
rect 19524 22040 19576 22092
rect 20352 22040 20404 22092
rect 23204 22219 23256 22228
rect 23204 22185 23213 22219
rect 23213 22185 23247 22219
rect 23247 22185 23256 22219
rect 23204 22176 23256 22185
rect 24676 22108 24728 22160
rect 22192 22040 22244 22092
rect 23940 22083 23992 22092
rect 2412 22015 2464 22024
rect 2412 21981 2421 22015
rect 2421 21981 2455 22015
rect 2455 21981 2464 22015
rect 2412 21972 2464 21981
rect 2596 22015 2648 22024
rect 2596 21981 2605 22015
rect 2605 21981 2639 22015
rect 2639 21981 2648 22015
rect 2596 21972 2648 21981
rect 4068 21972 4120 22024
rect 4620 21972 4672 22024
rect 6552 21972 6604 22024
rect 8484 22015 8536 22024
rect 8484 21981 8493 22015
rect 8493 21981 8527 22015
rect 8527 21981 8536 22015
rect 8484 21972 8536 21981
rect 3056 21947 3108 21956
rect 3056 21913 3065 21947
rect 3065 21913 3099 21947
rect 3099 21913 3108 21947
rect 3056 21904 3108 21913
rect 1216 21836 1268 21888
rect 2320 21836 2372 21888
rect 3608 21879 3660 21888
rect 3608 21845 3617 21879
rect 3617 21845 3651 21879
rect 3651 21845 3660 21879
rect 3608 21836 3660 21845
rect 3884 21836 3936 21888
rect 5448 21904 5500 21956
rect 8208 21904 8260 21956
rect 8300 21904 8352 21956
rect 9588 21972 9640 22024
rect 10784 21972 10836 22024
rect 10968 22015 11020 22024
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 14004 22015 14056 22024
rect 14004 21981 14013 22015
rect 14013 21981 14047 22015
rect 14047 21981 14056 22015
rect 14004 21972 14056 21981
rect 15292 22015 15344 22024
rect 15292 21981 15301 22015
rect 15301 21981 15335 22015
rect 15335 21981 15344 22015
rect 15292 21972 15344 21981
rect 17500 21972 17552 22024
rect 18328 22015 18380 22024
rect 18328 21981 18337 22015
rect 18337 21981 18371 22015
rect 18371 21981 18380 22015
rect 18328 21972 18380 21981
rect 9680 21904 9732 21956
rect 16672 21947 16724 21956
rect 16672 21913 16681 21947
rect 16681 21913 16715 21947
rect 16715 21913 16724 21947
rect 16672 21904 16724 21913
rect 18880 21904 18932 21956
rect 20536 21972 20588 22024
rect 20720 21972 20772 22024
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 23296 22015 23348 22024
rect 21824 21972 21876 21981
rect 23296 21981 23305 22015
rect 23305 21981 23339 22015
rect 23339 21981 23348 22015
rect 23296 21972 23348 21981
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 25320 22040 25372 22092
rect 21272 21947 21324 21956
rect 21272 21913 21281 21947
rect 21281 21913 21315 21947
rect 21315 21913 21324 21947
rect 21272 21904 21324 21913
rect 22468 21904 22520 21956
rect 25780 21904 25832 21956
rect 6828 21836 6880 21888
rect 7564 21836 7616 21888
rect 9496 21836 9548 21888
rect 10784 21836 10836 21888
rect 13360 21879 13412 21888
rect 13360 21845 13369 21879
rect 13369 21845 13403 21879
rect 13403 21845 13412 21879
rect 13360 21836 13412 21845
rect 14832 21879 14884 21888
rect 14832 21845 14841 21879
rect 14841 21845 14875 21879
rect 14875 21845 14884 21879
rect 14832 21836 14884 21845
rect 20536 21836 20588 21888
rect 21088 21879 21140 21888
rect 21088 21845 21097 21879
rect 21097 21845 21131 21879
rect 21131 21845 21140 21879
rect 21088 21836 21140 21845
rect 21640 21836 21692 21888
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 26148 21836 26200 21888
rect 5648 21734 5700 21786
rect 5712 21734 5764 21786
rect 5776 21734 5828 21786
rect 5840 21734 5892 21786
rect 14982 21734 15034 21786
rect 15046 21734 15098 21786
rect 15110 21734 15162 21786
rect 15174 21734 15226 21786
rect 24315 21734 24367 21786
rect 24379 21734 24431 21786
rect 24443 21734 24495 21786
rect 24507 21734 24559 21786
rect 1308 21632 1360 21684
rect 2504 21632 2556 21684
rect 3516 21675 3568 21684
rect 3516 21641 3525 21675
rect 3525 21641 3559 21675
rect 3559 21641 3568 21675
rect 3516 21632 3568 21641
rect 5080 21675 5132 21684
rect 5080 21641 5089 21675
rect 5089 21641 5123 21675
rect 5123 21641 5132 21675
rect 5080 21632 5132 21641
rect 5356 21632 5408 21684
rect 2596 21539 2648 21548
rect 2596 21505 2605 21539
rect 2605 21505 2639 21539
rect 2639 21505 2648 21539
rect 2596 21496 2648 21505
rect 756 21428 808 21480
rect 3516 21428 3568 21480
rect 3608 21428 3660 21480
rect 6552 21632 6604 21684
rect 7656 21632 7708 21684
rect 8852 21632 8904 21684
rect 11520 21675 11572 21684
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 12440 21632 12492 21684
rect 12900 21632 12952 21684
rect 14372 21632 14424 21684
rect 16304 21675 16356 21684
rect 16304 21641 16313 21675
rect 16313 21641 16347 21675
rect 16347 21641 16356 21675
rect 16304 21632 16356 21641
rect 17500 21675 17552 21684
rect 17500 21641 17509 21675
rect 17509 21641 17543 21675
rect 17543 21641 17552 21675
rect 17500 21632 17552 21641
rect 18328 21632 18380 21684
rect 21456 21675 21508 21684
rect 21456 21641 21465 21675
rect 21465 21641 21499 21675
rect 21499 21641 21508 21675
rect 21456 21632 21508 21641
rect 23204 21675 23256 21684
rect 23204 21641 23213 21675
rect 23213 21641 23247 21675
rect 23247 21641 23256 21675
rect 23204 21632 23256 21641
rect 25412 21675 25464 21684
rect 25412 21641 25421 21675
rect 25421 21641 25455 21675
rect 25455 21641 25464 21675
rect 25412 21632 25464 21641
rect 11060 21564 11112 21616
rect 10692 21496 10744 21548
rect 11888 21496 11940 21548
rect 15384 21496 15436 21548
rect 15844 21496 15896 21548
rect 24860 21564 24912 21616
rect 25320 21564 25372 21616
rect 17500 21496 17552 21548
rect 18880 21496 18932 21548
rect 19248 21496 19300 21548
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 21272 21496 21324 21548
rect 22284 21539 22336 21548
rect 22284 21505 22293 21539
rect 22293 21505 22327 21539
rect 22327 21505 22336 21539
rect 22284 21496 22336 21505
rect 24124 21539 24176 21548
rect 24124 21505 24133 21539
rect 24133 21505 24167 21539
rect 24167 21505 24176 21539
rect 24124 21496 24176 21505
rect 20 21360 72 21412
rect 848 21360 900 21412
rect 7104 21428 7156 21480
rect 7564 21428 7616 21480
rect 10048 21428 10100 21480
rect 10968 21428 11020 21480
rect 13360 21428 13412 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 16764 21471 16816 21480
rect 16764 21437 16773 21471
rect 16773 21437 16807 21471
rect 16807 21437 16816 21471
rect 16764 21428 16816 21437
rect 17776 21428 17828 21480
rect 19616 21428 19668 21480
rect 20076 21428 20128 21480
rect 20628 21428 20680 21480
rect 23940 21428 23992 21480
rect 8300 21360 8352 21412
rect 9772 21403 9824 21412
rect 9772 21369 9781 21403
rect 9781 21369 9815 21403
rect 9815 21369 9824 21403
rect 9772 21360 9824 21369
rect 3608 21292 3660 21344
rect 4620 21335 4672 21344
rect 4620 21301 4629 21335
rect 4629 21301 4663 21335
rect 4663 21301 4672 21335
rect 4620 21292 4672 21301
rect 5540 21335 5592 21344
rect 5540 21301 5549 21335
rect 5549 21301 5583 21335
rect 5583 21301 5592 21335
rect 6368 21335 6420 21344
rect 5540 21292 5592 21301
rect 6368 21301 6377 21335
rect 6377 21301 6411 21335
rect 6411 21301 6420 21335
rect 6368 21292 6420 21301
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 10784 21292 10836 21344
rect 10968 21292 11020 21344
rect 11888 21335 11940 21344
rect 11888 21301 11897 21335
rect 11897 21301 11931 21335
rect 11931 21301 11940 21335
rect 11888 21292 11940 21301
rect 13636 21360 13688 21412
rect 14188 21360 14240 21412
rect 16304 21360 16356 21412
rect 16856 21403 16908 21412
rect 16856 21369 16865 21403
rect 16865 21369 16899 21403
rect 16899 21369 16908 21403
rect 16856 21360 16908 21369
rect 17868 21360 17920 21412
rect 19708 21403 19760 21412
rect 19708 21369 19717 21403
rect 19717 21369 19751 21403
rect 19751 21369 19760 21403
rect 19708 21360 19760 21369
rect 21824 21360 21876 21412
rect 23020 21360 23072 21412
rect 23204 21360 23256 21412
rect 25136 21428 25188 21480
rect 14464 21292 14516 21344
rect 15200 21292 15252 21344
rect 15936 21292 15988 21344
rect 18420 21292 18472 21344
rect 18788 21292 18840 21344
rect 19524 21292 19576 21344
rect 19984 21292 20036 21344
rect 21640 21335 21692 21344
rect 21640 21301 21649 21335
rect 21649 21301 21683 21335
rect 21683 21301 21692 21335
rect 21640 21292 21692 21301
rect 21916 21292 21968 21344
rect 23388 21292 23440 21344
rect 23664 21335 23716 21344
rect 23664 21301 23673 21335
rect 23673 21301 23707 21335
rect 23707 21301 23716 21335
rect 23664 21292 23716 21301
rect 10315 21190 10367 21242
rect 10379 21190 10431 21242
rect 10443 21190 10495 21242
rect 10507 21190 10559 21242
rect 19648 21190 19700 21242
rect 19712 21190 19764 21242
rect 19776 21190 19828 21242
rect 19840 21190 19892 21242
rect 1860 21088 1912 21140
rect 2320 21131 2372 21140
rect 2320 21097 2329 21131
rect 2329 21097 2363 21131
rect 2363 21097 2372 21131
rect 2320 21088 2372 21097
rect 3148 21088 3200 21140
rect 4068 21131 4120 21140
rect 4068 21097 4077 21131
rect 4077 21097 4111 21131
rect 4111 21097 4120 21131
rect 4068 21088 4120 21097
rect 4528 21131 4580 21140
rect 4528 21097 4537 21131
rect 4537 21097 4571 21131
rect 4571 21097 4580 21131
rect 4528 21088 4580 21097
rect 4804 21088 4856 21140
rect 7288 21088 7340 21140
rect 8024 21088 8076 21140
rect 9036 21131 9088 21140
rect 9036 21097 9045 21131
rect 9045 21097 9079 21131
rect 9079 21097 9088 21131
rect 9036 21088 9088 21097
rect 2412 21020 2464 21072
rect 6368 21020 6420 21072
rect 9680 21020 9732 21072
rect 12072 21088 12124 21140
rect 13728 21088 13780 21140
rect 14280 21131 14332 21140
rect 14280 21097 14289 21131
rect 14289 21097 14323 21131
rect 14323 21097 14332 21131
rect 14280 21088 14332 21097
rect 14464 21088 14516 21140
rect 14832 21088 14884 21140
rect 16856 21131 16908 21140
rect 16856 21097 16865 21131
rect 16865 21097 16899 21131
rect 16899 21097 16908 21131
rect 16856 21088 16908 21097
rect 18144 21088 18196 21140
rect 18972 21131 19024 21140
rect 18972 21097 18981 21131
rect 18981 21097 19015 21131
rect 19015 21097 19024 21131
rect 18972 21088 19024 21097
rect 19064 21088 19116 21140
rect 20352 21131 20404 21140
rect 3976 20952 4028 21004
rect 6276 20952 6328 21004
rect 8300 20995 8352 21004
rect 8300 20961 8309 20995
rect 8309 20961 8343 20995
rect 8343 20961 8352 20995
rect 12716 21020 12768 21072
rect 13636 21020 13688 21072
rect 16580 21020 16632 21072
rect 17868 21020 17920 21072
rect 19248 21020 19300 21072
rect 19524 21020 19576 21072
rect 8300 20952 8352 20961
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 12624 20995 12676 21004
rect 12624 20961 12633 20995
rect 12633 20961 12667 20995
rect 12667 20961 12676 20995
rect 12624 20952 12676 20961
rect 14740 20952 14792 21004
rect 2596 20927 2648 20936
rect 2596 20893 2605 20927
rect 2605 20893 2639 20927
rect 2639 20893 2648 20927
rect 2596 20884 2648 20893
rect 5356 20884 5408 20936
rect 6460 20884 6512 20936
rect 7656 20927 7708 20936
rect 7656 20893 7665 20927
rect 7665 20893 7699 20927
rect 7699 20893 7708 20927
rect 7656 20884 7708 20893
rect 7748 20927 7800 20936
rect 7748 20893 7757 20927
rect 7757 20893 7791 20927
rect 7791 20893 7800 20927
rect 7748 20884 7800 20893
rect 11612 20927 11664 20936
rect 2872 20816 2924 20868
rect 3884 20816 3936 20868
rect 5540 20816 5592 20868
rect 8484 20816 8536 20868
rect 9588 20816 9640 20868
rect 3608 20791 3660 20800
rect 3608 20757 3617 20791
rect 3617 20757 3651 20791
rect 3651 20757 3660 20791
rect 3608 20748 3660 20757
rect 7196 20791 7248 20800
rect 7196 20757 7205 20791
rect 7205 20757 7239 20791
rect 7239 20757 7248 20791
rect 7196 20748 7248 20757
rect 9404 20791 9456 20800
rect 9404 20757 9413 20791
rect 9413 20757 9447 20791
rect 9447 20757 9456 20791
rect 9404 20748 9456 20757
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 12716 20927 12768 20936
rect 12716 20893 12725 20927
rect 12725 20893 12759 20927
rect 12759 20893 12768 20927
rect 12716 20884 12768 20893
rect 10048 20748 10100 20800
rect 14648 20791 14700 20800
rect 14648 20757 14657 20791
rect 14657 20757 14691 20791
rect 14691 20757 14700 20791
rect 14648 20748 14700 20757
rect 14832 20748 14884 20800
rect 16948 20952 17000 21004
rect 17592 20952 17644 21004
rect 18144 20952 18196 21004
rect 18512 20952 18564 21004
rect 18880 20995 18932 21004
rect 18880 20961 18889 20995
rect 18889 20961 18923 20995
rect 18923 20961 18932 20995
rect 18880 20952 18932 20961
rect 15752 20927 15804 20936
rect 15752 20893 15761 20927
rect 15761 20893 15795 20927
rect 15795 20893 15804 20927
rect 15936 20927 15988 20936
rect 15752 20884 15804 20893
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 16212 20884 16264 20936
rect 17500 20927 17552 20936
rect 17500 20893 17509 20927
rect 17509 20893 17543 20927
rect 17543 20893 17552 20927
rect 17500 20884 17552 20893
rect 19064 20927 19116 20936
rect 19064 20893 19073 20927
rect 19073 20893 19107 20927
rect 19107 20893 19116 20927
rect 19064 20884 19116 20893
rect 20352 21097 20361 21131
rect 20361 21097 20395 21131
rect 20395 21097 20404 21131
rect 20352 21088 20404 21097
rect 20720 21131 20772 21140
rect 20720 21097 20729 21131
rect 20729 21097 20763 21131
rect 20763 21097 20772 21131
rect 20720 21088 20772 21097
rect 21732 21131 21784 21140
rect 21732 21097 21741 21131
rect 21741 21097 21775 21131
rect 21775 21097 21784 21131
rect 21732 21088 21784 21097
rect 23664 21088 23716 21140
rect 20628 21020 20680 21072
rect 22192 21063 22244 21072
rect 22192 21029 22226 21063
rect 22226 21029 22244 21063
rect 22192 21020 22244 21029
rect 22468 21020 22520 21072
rect 24124 21020 24176 21072
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 20812 20816 20864 20868
rect 23480 20884 23532 20936
rect 25044 20927 25096 20936
rect 25044 20893 25053 20927
rect 25053 20893 25087 20927
rect 25087 20893 25096 20927
rect 25044 20884 25096 20893
rect 26240 20816 26292 20868
rect 15936 20748 15988 20800
rect 16212 20748 16264 20800
rect 16488 20748 16540 20800
rect 18512 20791 18564 20800
rect 18512 20757 18521 20791
rect 18521 20757 18555 20791
rect 18555 20757 18564 20791
rect 18512 20748 18564 20757
rect 19156 20748 19208 20800
rect 19432 20748 19484 20800
rect 21824 20748 21876 20800
rect 23572 20748 23624 20800
rect 24124 20748 24176 20800
rect 5648 20646 5700 20698
rect 5712 20646 5764 20698
rect 5776 20646 5828 20698
rect 5840 20646 5892 20698
rect 14982 20646 15034 20698
rect 15046 20646 15098 20698
rect 15110 20646 15162 20698
rect 15174 20646 15226 20698
rect 24315 20646 24367 20698
rect 24379 20646 24431 20698
rect 24443 20646 24495 20698
rect 24507 20646 24559 20698
rect 940 20544 992 20596
rect 2136 20544 2188 20596
rect 2872 20544 2924 20596
rect 3700 20544 3752 20596
rect 6276 20544 6328 20596
rect 6460 20587 6512 20596
rect 6460 20553 6469 20587
rect 6469 20553 6503 20587
rect 6503 20553 6512 20587
rect 6460 20544 6512 20553
rect 6920 20544 6972 20596
rect 7748 20544 7800 20596
rect 9588 20544 9640 20596
rect 10876 20544 10928 20596
rect 12532 20544 12584 20596
rect 12808 20544 12860 20596
rect 14372 20544 14424 20596
rect 3148 20476 3200 20528
rect 3516 20476 3568 20528
rect 2412 20451 2464 20460
rect 2412 20417 2421 20451
rect 2421 20417 2455 20451
rect 2455 20417 2464 20451
rect 2412 20408 2464 20417
rect 2596 20451 2648 20460
rect 2596 20417 2605 20451
rect 2605 20417 2639 20451
rect 2639 20417 2648 20451
rect 2596 20408 2648 20417
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 7748 20408 7800 20460
rect 10968 20476 11020 20528
rect 12624 20476 12676 20528
rect 14924 20476 14976 20528
rect 15476 20476 15528 20528
rect 3792 20383 3844 20392
rect 3792 20349 3801 20383
rect 3801 20349 3835 20383
rect 3835 20349 3844 20383
rect 3792 20340 3844 20349
rect 4620 20340 4672 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 6368 20340 6420 20392
rect 9680 20408 9732 20460
rect 11888 20408 11940 20460
rect 14556 20451 14608 20460
rect 14556 20417 14565 20451
rect 14565 20417 14599 20451
rect 14599 20417 14608 20451
rect 14556 20408 14608 20417
rect 8576 20340 8628 20392
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 11520 20272 11572 20324
rect 12624 20340 12676 20392
rect 12900 20383 12952 20392
rect 12900 20349 12909 20383
rect 12909 20349 12943 20383
rect 12943 20349 12952 20383
rect 12900 20340 12952 20349
rect 13452 20340 13504 20392
rect 15752 20340 15804 20392
rect 14556 20272 14608 20324
rect 16488 20544 16540 20596
rect 17500 20587 17552 20596
rect 17500 20553 17509 20587
rect 17509 20553 17543 20587
rect 17543 20553 17552 20587
rect 17500 20544 17552 20553
rect 18972 20587 19024 20596
rect 18972 20553 18981 20587
rect 18981 20553 19015 20587
rect 19015 20553 19024 20587
rect 18972 20544 19024 20553
rect 21456 20544 21508 20596
rect 22192 20544 22244 20596
rect 23480 20587 23532 20596
rect 23480 20553 23489 20587
rect 23489 20553 23523 20587
rect 23523 20553 23532 20587
rect 23480 20544 23532 20553
rect 19156 20476 19208 20528
rect 20812 20476 20864 20528
rect 22652 20476 22704 20528
rect 22836 20476 22888 20528
rect 16948 20451 17000 20460
rect 16948 20417 16957 20451
rect 16957 20417 16991 20451
rect 16991 20417 17000 20451
rect 16948 20408 17000 20417
rect 20536 20408 20588 20460
rect 22284 20451 22336 20460
rect 22284 20417 22293 20451
rect 22293 20417 22327 20451
rect 22327 20417 22336 20451
rect 22284 20408 22336 20417
rect 24860 20544 24912 20596
rect 26240 20587 26292 20596
rect 26240 20553 26249 20587
rect 26249 20553 26283 20587
rect 26283 20553 26292 20587
rect 26240 20544 26292 20553
rect 24308 20451 24360 20460
rect 16764 20383 16816 20392
rect 16764 20349 16773 20383
rect 16773 20349 16807 20383
rect 16807 20349 16816 20383
rect 16764 20340 16816 20349
rect 18052 20383 18104 20392
rect 18052 20349 18061 20383
rect 18061 20349 18095 20383
rect 18095 20349 18104 20383
rect 18052 20340 18104 20349
rect 19248 20340 19300 20392
rect 21640 20340 21692 20392
rect 21732 20340 21784 20392
rect 22468 20340 22520 20392
rect 24308 20417 24317 20451
rect 24317 20417 24351 20451
rect 24351 20417 24360 20451
rect 24308 20408 24360 20417
rect 16856 20315 16908 20324
rect 16856 20281 16865 20315
rect 16865 20281 16899 20315
rect 16899 20281 16908 20315
rect 16856 20272 16908 20281
rect 17776 20315 17828 20324
rect 17776 20281 17785 20315
rect 17785 20281 17819 20315
rect 17819 20281 17828 20315
rect 17776 20272 17828 20281
rect 19524 20272 19576 20324
rect 24216 20272 24268 20324
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 4528 20204 4580 20256
rect 7656 20247 7708 20256
rect 7656 20213 7665 20247
rect 7665 20213 7699 20247
rect 7699 20213 7708 20247
rect 7656 20204 7708 20213
rect 8300 20204 8352 20256
rect 10048 20204 10100 20256
rect 10692 20247 10744 20256
rect 10692 20213 10701 20247
rect 10701 20213 10735 20247
rect 10735 20213 10744 20247
rect 10692 20204 10744 20213
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 12624 20204 12676 20256
rect 13176 20204 13228 20256
rect 14004 20247 14056 20256
rect 14004 20213 14013 20247
rect 14013 20213 14047 20247
rect 14047 20213 14056 20247
rect 14004 20204 14056 20213
rect 14372 20247 14424 20256
rect 14372 20213 14381 20247
rect 14381 20213 14415 20247
rect 14415 20213 14424 20247
rect 14372 20204 14424 20213
rect 15200 20204 15252 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 22652 20247 22704 20256
rect 22652 20213 22661 20247
rect 22661 20213 22695 20247
rect 22695 20213 22704 20247
rect 22652 20204 22704 20213
rect 25044 20247 25096 20256
rect 25044 20213 25053 20247
rect 25053 20213 25087 20247
rect 25087 20213 25096 20247
rect 25044 20204 25096 20213
rect 10315 20102 10367 20154
rect 10379 20102 10431 20154
rect 10443 20102 10495 20154
rect 10507 20102 10559 20154
rect 19648 20102 19700 20154
rect 19712 20102 19764 20154
rect 19776 20102 19828 20154
rect 19840 20102 19892 20154
rect 1124 20000 1176 20052
rect 2320 20000 2372 20052
rect 4620 20000 4672 20052
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 7748 20000 7800 20052
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9864 20000 9916 20052
rect 11060 20000 11112 20052
rect 11336 20000 11388 20052
rect 11612 20000 11664 20052
rect 12900 20000 12952 20052
rect 13636 20000 13688 20052
rect 14556 20000 14608 20052
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 16028 20000 16080 20052
rect 16764 20000 16816 20052
rect 18328 20000 18380 20052
rect 18604 20000 18656 20052
rect 19340 20000 19392 20052
rect 19524 20000 19576 20052
rect 2872 19975 2924 19984
rect 2872 19941 2881 19975
rect 2881 19941 2915 19975
rect 2915 19941 2924 19975
rect 2872 19932 2924 19941
rect 3976 19932 4028 19984
rect 4804 19932 4856 19984
rect 5540 19932 5592 19984
rect 6460 19932 6512 19984
rect 9404 19932 9456 19984
rect 12624 19932 12676 19984
rect 3884 19864 3936 19916
rect 4068 19907 4120 19916
rect 4068 19873 4077 19907
rect 4077 19873 4111 19907
rect 4111 19873 4120 19907
rect 4068 19864 4120 19873
rect 2596 19796 2648 19848
rect 4528 19796 4580 19848
rect 6276 19864 6328 19916
rect 6552 19864 6604 19916
rect 8760 19864 8812 19916
rect 9680 19864 9732 19916
rect 10232 19864 10284 19916
rect 12256 19864 12308 19916
rect 12808 19864 12860 19916
rect 15936 19864 15988 19916
rect 17408 19907 17460 19916
rect 17408 19873 17417 19907
rect 17417 19873 17451 19907
rect 17451 19873 17460 19907
rect 17408 19864 17460 19873
rect 17684 19864 17736 19916
rect 18420 19864 18472 19916
rect 6828 19796 6880 19848
rect 7104 19796 7156 19848
rect 8024 19796 8076 19848
rect 11336 19839 11388 19848
rect 3884 19728 3936 19780
rect 8300 19728 8352 19780
rect 11336 19805 11345 19839
rect 11345 19805 11379 19839
rect 11379 19805 11388 19839
rect 11336 19796 11388 19805
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 13820 19728 13872 19780
rect 14372 19728 14424 19780
rect 16856 19728 16908 19780
rect 19156 19796 19208 19848
rect 20536 20000 20588 20052
rect 22284 20000 22336 20052
rect 23572 19932 23624 19984
rect 24308 19932 24360 19984
rect 20812 19864 20864 19916
rect 21456 19864 21508 19916
rect 23388 19839 23440 19848
rect 23388 19805 23397 19839
rect 23397 19805 23431 19839
rect 23431 19805 23440 19839
rect 23388 19796 23440 19805
rect 18788 19728 18840 19780
rect 22192 19728 22244 19780
rect 22376 19728 22428 19780
rect 2320 19660 2372 19712
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 4252 19703 4304 19712
rect 4252 19669 4261 19703
rect 4261 19669 4295 19703
rect 4295 19669 4304 19703
rect 4252 19660 4304 19669
rect 5448 19703 5500 19712
rect 5448 19669 5457 19703
rect 5457 19669 5491 19703
rect 5491 19669 5500 19703
rect 5448 19660 5500 19669
rect 9128 19703 9180 19712
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 9496 19703 9548 19712
rect 9496 19669 9505 19703
rect 9505 19669 9539 19703
rect 9539 19669 9548 19703
rect 9496 19660 9548 19669
rect 9680 19660 9732 19712
rect 9772 19660 9824 19712
rect 10600 19660 10652 19712
rect 11796 19660 11848 19712
rect 13084 19660 13136 19712
rect 14464 19660 14516 19712
rect 16948 19703 17000 19712
rect 16948 19669 16957 19703
rect 16957 19669 16991 19703
rect 16991 19669 17000 19703
rect 16948 19660 17000 19669
rect 17592 19660 17644 19712
rect 19248 19660 19300 19712
rect 22008 19660 22060 19712
rect 23296 19703 23348 19712
rect 23296 19669 23305 19703
rect 23305 19669 23339 19703
rect 23339 19669 23348 19703
rect 23296 19660 23348 19669
rect 5648 19558 5700 19610
rect 5712 19558 5764 19610
rect 5776 19558 5828 19610
rect 5840 19558 5892 19610
rect 14982 19558 15034 19610
rect 15046 19558 15098 19610
rect 15110 19558 15162 19610
rect 15174 19558 15226 19610
rect 24315 19558 24367 19610
rect 24379 19558 24431 19610
rect 24443 19558 24495 19610
rect 24507 19558 24559 19610
rect 1584 19388 1636 19440
rect 2044 19388 2096 19440
rect 2688 19320 2740 19372
rect 2872 19456 2924 19508
rect 4068 19499 4120 19508
rect 4068 19465 4077 19499
rect 4077 19465 4111 19499
rect 4111 19465 4120 19499
rect 4068 19456 4120 19465
rect 6460 19456 6512 19508
rect 9496 19456 9548 19508
rect 10692 19456 10744 19508
rect 10968 19456 11020 19508
rect 11152 19456 11204 19508
rect 11428 19456 11480 19508
rect 12256 19456 12308 19508
rect 1860 19252 1912 19304
rect 2136 19252 2188 19304
rect 2412 19252 2464 19304
rect 3792 19388 3844 19440
rect 3884 19320 3936 19372
rect 3056 19295 3108 19304
rect 3056 19261 3065 19295
rect 3065 19261 3099 19295
rect 3099 19261 3108 19295
rect 3056 19252 3108 19261
rect 4528 19295 4580 19304
rect 4528 19261 4562 19295
rect 4562 19261 4580 19295
rect 3792 19227 3844 19236
rect 3792 19193 3801 19227
rect 3801 19193 3835 19227
rect 3835 19193 3844 19227
rect 4528 19252 4580 19261
rect 6276 19320 6328 19372
rect 7656 19320 7708 19372
rect 9404 19320 9456 19372
rect 7012 19252 7064 19304
rect 11612 19388 11664 19440
rect 11336 19363 11388 19372
rect 11336 19329 11345 19363
rect 11345 19329 11379 19363
rect 11379 19329 11388 19363
rect 11336 19320 11388 19329
rect 12624 19456 12676 19508
rect 14556 19499 14608 19508
rect 14556 19465 14565 19499
rect 14565 19465 14599 19499
rect 14599 19465 14608 19499
rect 14556 19456 14608 19465
rect 16856 19499 16908 19508
rect 12440 19388 12492 19440
rect 12900 19388 12952 19440
rect 13084 19388 13136 19440
rect 12808 19363 12860 19372
rect 12808 19329 12817 19363
rect 12817 19329 12851 19363
rect 12851 19329 12860 19363
rect 12808 19320 12860 19329
rect 13268 19320 13320 19372
rect 11244 19295 11296 19304
rect 3792 19184 3844 19193
rect 1584 19159 1636 19168
rect 1584 19125 1593 19159
rect 1593 19125 1627 19159
rect 1627 19125 1636 19159
rect 1584 19116 1636 19125
rect 2688 19159 2740 19168
rect 2688 19125 2697 19159
rect 2697 19125 2731 19159
rect 2731 19125 2740 19159
rect 2688 19116 2740 19125
rect 3332 19116 3384 19168
rect 5632 19159 5684 19168
rect 5632 19125 5641 19159
rect 5641 19125 5675 19159
rect 5675 19125 5684 19159
rect 5632 19116 5684 19125
rect 8116 19184 8168 19236
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12532 19252 12584 19304
rect 14464 19320 14516 19372
rect 14924 19320 14976 19372
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 20720 19456 20772 19508
rect 21456 19456 21508 19508
rect 24216 19456 24268 19508
rect 20812 19388 20864 19440
rect 24308 19388 24360 19440
rect 15844 19320 15896 19372
rect 14280 19295 14332 19304
rect 14280 19261 14289 19295
rect 14289 19261 14323 19295
rect 14323 19261 14332 19295
rect 14280 19252 14332 19261
rect 15568 19295 15620 19304
rect 15568 19261 15577 19295
rect 15577 19261 15611 19295
rect 15611 19261 15620 19295
rect 15568 19252 15620 19261
rect 16948 19295 17000 19304
rect 16948 19261 16957 19295
rect 16957 19261 16991 19295
rect 16991 19261 17000 19295
rect 16948 19252 17000 19261
rect 6276 19159 6328 19168
rect 6276 19125 6285 19159
rect 6285 19125 6319 19159
rect 6319 19125 6328 19159
rect 6276 19116 6328 19125
rect 7012 19159 7064 19168
rect 7012 19125 7021 19159
rect 7021 19125 7055 19159
rect 7055 19125 7064 19159
rect 7012 19116 7064 19125
rect 7472 19159 7524 19168
rect 7472 19125 7481 19159
rect 7481 19125 7515 19159
rect 7515 19125 7524 19159
rect 7472 19116 7524 19125
rect 11520 19116 11572 19168
rect 13728 19184 13780 19236
rect 14832 19184 14884 19236
rect 13544 19159 13596 19168
rect 13544 19125 13553 19159
rect 13553 19125 13587 19159
rect 13587 19125 13596 19159
rect 13544 19116 13596 19125
rect 15292 19184 15344 19236
rect 17040 19184 17092 19236
rect 17408 19227 17460 19236
rect 17408 19193 17417 19227
rect 17417 19193 17451 19227
rect 17451 19193 17460 19227
rect 17408 19184 17460 19193
rect 20536 19320 20588 19372
rect 22376 19320 22428 19372
rect 22652 19320 22704 19372
rect 23388 19363 23440 19372
rect 23388 19329 23397 19363
rect 23397 19329 23431 19363
rect 23431 19329 23440 19363
rect 23388 19320 23440 19329
rect 24216 19363 24268 19372
rect 24216 19329 24225 19363
rect 24225 19329 24259 19363
rect 24259 19329 24268 19363
rect 24216 19320 24268 19329
rect 19340 19252 19392 19304
rect 19984 19252 20036 19304
rect 23296 19252 23348 19304
rect 23940 19252 23992 19304
rect 25320 19252 25372 19304
rect 15936 19116 15988 19168
rect 17316 19116 17368 19168
rect 17684 19116 17736 19168
rect 18420 19159 18472 19168
rect 18420 19125 18429 19159
rect 18429 19125 18463 19159
rect 18463 19125 18472 19159
rect 18420 19116 18472 19125
rect 18604 19159 18656 19168
rect 18604 19125 18613 19159
rect 18613 19125 18647 19159
rect 18647 19125 18656 19159
rect 18604 19116 18656 19125
rect 18972 19159 19024 19168
rect 18972 19125 18981 19159
rect 18981 19125 19015 19159
rect 19015 19125 19024 19159
rect 18972 19116 19024 19125
rect 19248 19116 19300 19168
rect 19340 19116 19392 19168
rect 20260 19116 20312 19168
rect 20628 19159 20680 19168
rect 20628 19125 20637 19159
rect 20637 19125 20671 19159
rect 20671 19125 20680 19159
rect 20628 19116 20680 19125
rect 22100 19116 22152 19168
rect 22836 19116 22888 19168
rect 23020 19159 23072 19168
rect 23020 19125 23029 19159
rect 23029 19125 23063 19159
rect 23063 19125 23072 19159
rect 23020 19116 23072 19125
rect 23664 19159 23716 19168
rect 23664 19125 23673 19159
rect 23673 19125 23707 19159
rect 23707 19125 23716 19159
rect 23664 19116 23716 19125
rect 25504 19116 25556 19168
rect 25596 19116 25648 19168
rect 26332 19116 26384 19168
rect 10315 19014 10367 19066
rect 10379 19014 10431 19066
rect 10443 19014 10495 19066
rect 10507 19014 10559 19066
rect 19648 19014 19700 19066
rect 19712 19014 19764 19066
rect 19776 19014 19828 19066
rect 19840 19014 19892 19066
rect 2596 18912 2648 18964
rect 3148 18912 3200 18964
rect 3884 18955 3936 18964
rect 3884 18921 3893 18955
rect 3893 18921 3927 18955
rect 3927 18921 3936 18955
rect 3884 18912 3936 18921
rect 4528 18912 4580 18964
rect 5540 18912 5592 18964
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 9404 18912 9456 18964
rect 9588 18912 9640 18964
rect 9864 18955 9916 18964
rect 9864 18921 9873 18955
rect 9873 18921 9907 18955
rect 9907 18921 9916 18955
rect 9864 18912 9916 18921
rect 11336 18912 11388 18964
rect 12532 18912 12584 18964
rect 13268 18955 13320 18964
rect 13268 18921 13277 18955
rect 13277 18921 13311 18955
rect 13311 18921 13320 18955
rect 13268 18912 13320 18921
rect 15568 18912 15620 18964
rect 16028 18912 16080 18964
rect 17500 18912 17552 18964
rect 18512 18912 18564 18964
rect 19984 18912 20036 18964
rect 21364 18912 21416 18964
rect 22376 18912 22428 18964
rect 23020 18912 23072 18964
rect 24216 18912 24268 18964
rect 24860 18912 24912 18964
rect 5632 18887 5684 18896
rect 2136 18776 2188 18828
rect 3884 18776 3936 18828
rect 5632 18853 5666 18887
rect 5666 18853 5684 18887
rect 5632 18844 5684 18853
rect 6276 18844 6328 18896
rect 6460 18844 6512 18896
rect 4528 18776 4580 18828
rect 2228 18708 2280 18760
rect 2412 18708 2464 18760
rect 3240 18708 3292 18760
rect 4160 18708 4212 18760
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 7932 18844 7984 18896
rect 11152 18844 11204 18896
rect 12900 18844 12952 18896
rect 20812 18844 20864 18896
rect 21272 18844 21324 18896
rect 7656 18776 7708 18828
rect 9864 18776 9916 18828
rect 10048 18776 10100 18828
rect 11520 18776 11572 18828
rect 12808 18776 12860 18828
rect 13084 18776 13136 18828
rect 15292 18819 15344 18828
rect 15292 18785 15301 18819
rect 15301 18785 15335 18819
rect 15335 18785 15344 18819
rect 15292 18776 15344 18785
rect 15476 18776 15528 18828
rect 17408 18776 17460 18828
rect 20260 18776 20312 18828
rect 22652 18776 22704 18828
rect 23940 18776 23992 18828
rect 24952 18776 25004 18828
rect 8300 18708 8352 18760
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 13636 18708 13688 18760
rect 14556 18708 14608 18760
rect 17868 18708 17920 18760
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 21088 18708 21140 18760
rect 21824 18708 21876 18760
rect 2964 18640 3016 18692
rect 16120 18640 16172 18692
rect 3332 18572 3384 18624
rect 4068 18572 4120 18624
rect 8116 18572 8168 18624
rect 13544 18572 13596 18624
rect 13728 18572 13780 18624
rect 14372 18615 14424 18624
rect 14372 18581 14381 18615
rect 14381 18581 14415 18615
rect 14415 18581 14424 18615
rect 14372 18572 14424 18581
rect 15844 18615 15896 18624
rect 15844 18581 15853 18615
rect 15853 18581 15887 18615
rect 15887 18581 15896 18615
rect 15844 18572 15896 18581
rect 18512 18572 18564 18624
rect 18972 18640 19024 18692
rect 21916 18640 21968 18692
rect 19156 18572 19208 18624
rect 19524 18572 19576 18624
rect 21732 18572 21784 18624
rect 22192 18572 22244 18624
rect 5648 18470 5700 18522
rect 5712 18470 5764 18522
rect 5776 18470 5828 18522
rect 5840 18470 5892 18522
rect 14982 18470 15034 18522
rect 15046 18470 15098 18522
rect 15110 18470 15162 18522
rect 15174 18470 15226 18522
rect 24315 18470 24367 18522
rect 24379 18470 24431 18522
rect 24443 18470 24495 18522
rect 24507 18470 24559 18522
rect 3148 18368 3200 18420
rect 3424 18368 3476 18420
rect 4528 18411 4580 18420
rect 4528 18377 4537 18411
rect 4537 18377 4571 18411
rect 4571 18377 4580 18411
rect 4528 18368 4580 18377
rect 2136 18343 2188 18352
rect 2136 18309 2145 18343
rect 2145 18309 2179 18343
rect 2179 18309 2188 18343
rect 2136 18300 2188 18309
rect 3240 18300 3292 18352
rect 5540 18368 5592 18420
rect 6276 18368 6328 18420
rect 8576 18368 8628 18420
rect 9220 18411 9272 18420
rect 9220 18377 9229 18411
rect 9229 18377 9263 18411
rect 9263 18377 9272 18411
rect 9220 18368 9272 18377
rect 9588 18368 9640 18420
rect 11520 18368 11572 18420
rect 11888 18368 11940 18420
rect 13084 18411 13136 18420
rect 8392 18300 8444 18352
rect 2228 18275 2280 18284
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 5172 18232 5224 18284
rect 6276 18232 6328 18284
rect 7840 18232 7892 18284
rect 8208 18275 8260 18284
rect 8208 18241 8217 18275
rect 8217 18241 8251 18275
rect 8251 18241 8260 18275
rect 8208 18232 8260 18241
rect 8484 18232 8536 18284
rect 9404 18232 9456 18284
rect 11152 18300 11204 18352
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 13452 18368 13504 18420
rect 14556 18411 14608 18420
rect 14556 18377 14565 18411
rect 14565 18377 14599 18411
rect 14599 18377 14608 18411
rect 14556 18368 14608 18377
rect 17408 18411 17460 18420
rect 17408 18377 17417 18411
rect 17417 18377 17451 18411
rect 17451 18377 17460 18411
rect 17408 18368 17460 18377
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 18788 18368 18840 18420
rect 19340 18368 19392 18420
rect 19708 18368 19760 18420
rect 20812 18368 20864 18420
rect 21364 18411 21416 18420
rect 21364 18377 21373 18411
rect 21373 18377 21407 18411
rect 21407 18377 21416 18411
rect 21364 18368 21416 18377
rect 23296 18368 23348 18420
rect 24216 18368 24268 18420
rect 24952 18368 25004 18420
rect 25412 18411 25464 18420
rect 25412 18377 25421 18411
rect 25421 18377 25455 18411
rect 25455 18377 25464 18411
rect 25412 18368 25464 18377
rect 12900 18232 12952 18284
rect 13084 18232 13136 18284
rect 14004 18232 14056 18284
rect 16120 18300 16172 18352
rect 16488 18343 16540 18352
rect 16488 18309 16497 18343
rect 16497 18309 16531 18343
rect 16531 18309 16540 18343
rect 16488 18300 16540 18309
rect 2872 18164 2924 18216
rect 7656 18164 7708 18216
rect 7932 18207 7984 18216
rect 7932 18173 7941 18207
rect 7941 18173 7975 18207
rect 7975 18173 7984 18207
rect 7932 18164 7984 18173
rect 9128 18164 9180 18216
rect 9588 18207 9640 18216
rect 9588 18173 9597 18207
rect 9597 18173 9631 18207
rect 9631 18173 9640 18207
rect 9588 18164 9640 18173
rect 9864 18164 9916 18216
rect 10968 18164 11020 18216
rect 11520 18164 11572 18216
rect 13360 18164 13412 18216
rect 14280 18164 14332 18216
rect 15108 18207 15160 18216
rect 5540 18139 5592 18148
rect 5540 18105 5549 18139
rect 5549 18105 5583 18139
rect 5583 18105 5592 18139
rect 5540 18096 5592 18105
rect 10876 18096 10928 18148
rect 12808 18096 12860 18148
rect 5172 18071 5224 18080
rect 5172 18037 5181 18071
rect 5181 18037 5215 18071
rect 5215 18037 5224 18071
rect 5172 18028 5224 18037
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 6644 18028 6696 18080
rect 7472 18028 7524 18080
rect 11060 18028 11112 18080
rect 11244 18071 11296 18080
rect 11244 18037 11253 18071
rect 11253 18037 11287 18071
rect 11287 18037 11296 18071
rect 11244 18028 11296 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 13636 18028 13688 18080
rect 14096 18096 14148 18148
rect 15108 18173 15117 18207
rect 15117 18173 15151 18207
rect 15151 18173 15160 18207
rect 15108 18164 15160 18173
rect 15844 18164 15896 18216
rect 15476 18028 15528 18080
rect 18236 18232 18288 18284
rect 18420 18232 18472 18284
rect 23572 18300 23624 18352
rect 22192 18275 22244 18284
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 23848 18232 23900 18284
rect 18972 18096 19024 18148
rect 18052 18028 18104 18080
rect 18236 18071 18288 18080
rect 18236 18037 18245 18071
rect 18245 18037 18279 18071
rect 18279 18037 18288 18071
rect 18236 18028 18288 18037
rect 19340 18028 19392 18080
rect 19708 18164 19760 18216
rect 21364 18164 21416 18216
rect 23572 18164 23624 18216
rect 25228 18207 25280 18216
rect 25228 18173 25237 18207
rect 25237 18173 25271 18207
rect 25271 18173 25280 18207
rect 25228 18164 25280 18173
rect 19616 18096 19668 18148
rect 21272 18096 21324 18148
rect 21824 18096 21876 18148
rect 25320 18096 25372 18148
rect 19524 18028 19576 18080
rect 20812 18028 20864 18080
rect 21548 18071 21600 18080
rect 21548 18037 21557 18071
rect 21557 18037 21591 18071
rect 21591 18037 21600 18071
rect 21548 18028 21600 18037
rect 21640 18028 21692 18080
rect 22008 18071 22060 18080
rect 22008 18037 22017 18071
rect 22017 18037 22051 18071
rect 22051 18037 22060 18071
rect 22008 18028 22060 18037
rect 22744 18028 22796 18080
rect 10315 17926 10367 17978
rect 10379 17926 10431 17978
rect 10443 17926 10495 17978
rect 10507 17926 10559 17978
rect 19648 17926 19700 17978
rect 19712 17926 19764 17978
rect 19776 17926 19828 17978
rect 19840 17926 19892 17978
rect 2964 17824 3016 17876
rect 3884 17867 3936 17876
rect 3884 17833 3893 17867
rect 3893 17833 3927 17867
rect 3927 17833 3936 17867
rect 3884 17824 3936 17833
rect 5448 17824 5500 17876
rect 6276 17867 6328 17876
rect 6276 17833 6285 17867
rect 6285 17833 6319 17867
rect 6319 17833 6328 17867
rect 6276 17824 6328 17833
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 11428 17824 11480 17876
rect 2228 17688 2280 17740
rect 2872 17756 2924 17808
rect 5356 17756 5408 17808
rect 6552 17756 6604 17808
rect 8760 17756 8812 17808
rect 9036 17756 9088 17808
rect 12532 17756 12584 17808
rect 13820 17824 13872 17876
rect 17592 17867 17644 17876
rect 17592 17833 17601 17867
rect 17601 17833 17635 17867
rect 17635 17833 17644 17867
rect 17592 17824 17644 17833
rect 17960 17867 18012 17876
rect 17960 17833 17969 17867
rect 17969 17833 18003 17867
rect 18003 17833 18012 17867
rect 17960 17824 18012 17833
rect 20260 17867 20312 17876
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 8300 17688 8352 17740
rect 9680 17688 9732 17740
rect 12808 17688 12860 17740
rect 14004 17756 14056 17808
rect 14096 17756 14148 17808
rect 15568 17799 15620 17808
rect 15568 17765 15602 17799
rect 15602 17765 15620 17799
rect 15568 17756 15620 17765
rect 16028 17756 16080 17808
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 21088 17824 21140 17876
rect 22376 17824 22428 17876
rect 24860 17824 24912 17876
rect 3424 17620 3476 17672
rect 5080 17620 5132 17672
rect 6552 17620 6604 17672
rect 6920 17663 6972 17672
rect 6920 17629 6929 17663
rect 6929 17629 6963 17663
rect 6963 17629 6972 17663
rect 6920 17620 6972 17629
rect 8668 17663 8720 17672
rect 5540 17552 5592 17604
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 9036 17620 9088 17672
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 13268 17663 13320 17672
rect 13268 17629 13277 17663
rect 13277 17629 13311 17663
rect 13311 17629 13320 17663
rect 13268 17620 13320 17629
rect 13636 17620 13688 17672
rect 14004 17620 14056 17672
rect 15108 17620 15160 17672
rect 8392 17552 8444 17604
rect 11704 17552 11756 17604
rect 12072 17552 12124 17604
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 6644 17484 6696 17536
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 11244 17527 11296 17536
rect 11244 17493 11253 17527
rect 11253 17493 11287 17527
rect 11287 17493 11296 17527
rect 11244 17484 11296 17493
rect 12532 17484 12584 17536
rect 14096 17484 14148 17536
rect 17868 17688 17920 17740
rect 20628 17756 20680 17808
rect 21272 17799 21324 17808
rect 21272 17765 21281 17799
rect 21281 17765 21315 17799
rect 21315 17765 21324 17799
rect 21272 17756 21324 17765
rect 22836 17756 22888 17808
rect 23204 17756 23256 17808
rect 23388 17756 23440 17808
rect 25044 17799 25096 17808
rect 25044 17765 25053 17799
rect 25053 17765 25087 17799
rect 25087 17765 25096 17799
rect 25044 17756 25096 17765
rect 20720 17688 20772 17740
rect 20904 17688 20956 17740
rect 21088 17688 21140 17740
rect 22652 17688 22704 17740
rect 23020 17731 23072 17740
rect 23020 17697 23043 17731
rect 23043 17697 23072 17731
rect 23020 17688 23072 17697
rect 25136 17688 25188 17740
rect 25780 17688 25832 17740
rect 18052 17620 18104 17672
rect 20260 17620 20312 17672
rect 22744 17663 22796 17672
rect 20720 17552 20772 17604
rect 22744 17629 22753 17663
rect 22753 17629 22787 17663
rect 22787 17629 22796 17663
rect 22744 17620 22796 17629
rect 23756 17552 23808 17604
rect 15476 17484 15528 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 17592 17484 17644 17536
rect 20904 17527 20956 17536
rect 20904 17493 20913 17527
rect 20913 17493 20947 17527
rect 20947 17493 20956 17527
rect 20904 17484 20956 17493
rect 21548 17484 21600 17536
rect 22008 17484 22060 17536
rect 22192 17484 22244 17536
rect 25780 17484 25832 17536
rect 25964 17484 26016 17536
rect 5648 17382 5700 17434
rect 5712 17382 5764 17434
rect 5776 17382 5828 17434
rect 5840 17382 5892 17434
rect 14982 17382 15034 17434
rect 15046 17382 15098 17434
rect 15110 17382 15162 17434
rect 15174 17382 15226 17434
rect 24315 17382 24367 17434
rect 24379 17382 24431 17434
rect 24443 17382 24495 17434
rect 24507 17382 24559 17434
rect 2136 17280 2188 17332
rect 3516 17280 3568 17332
rect 5080 17280 5132 17332
rect 5448 17280 5500 17332
rect 8668 17280 8720 17332
rect 10232 17280 10284 17332
rect 11888 17280 11940 17332
rect 3700 17212 3752 17264
rect 9680 17255 9732 17264
rect 2872 17008 2924 17060
rect 3792 17008 3844 17060
rect 9680 17221 9689 17255
rect 9689 17221 9723 17255
rect 9723 17221 9732 17255
rect 9680 17212 9732 17221
rect 5540 17144 5592 17196
rect 16120 17280 16172 17332
rect 17500 17323 17552 17332
rect 15568 17212 15620 17264
rect 5632 17119 5684 17128
rect 5632 17085 5641 17119
rect 5641 17085 5675 17119
rect 5675 17085 5684 17119
rect 5632 17076 5684 17085
rect 6644 17076 6696 17128
rect 9956 17076 10008 17128
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 17500 17289 17509 17323
rect 17509 17289 17543 17323
rect 17543 17289 17552 17323
rect 17500 17280 17552 17289
rect 17868 17323 17920 17332
rect 17868 17289 17877 17323
rect 17877 17289 17911 17323
rect 17911 17289 17920 17323
rect 17868 17280 17920 17289
rect 20628 17280 20680 17332
rect 23572 17280 23624 17332
rect 24676 17280 24728 17332
rect 25688 17280 25740 17332
rect 26056 17280 26108 17332
rect 18052 17212 18104 17264
rect 17592 17144 17644 17196
rect 17500 17076 17552 17128
rect 19340 17119 19392 17128
rect 19340 17085 19374 17119
rect 19374 17085 19392 17119
rect 23020 17212 23072 17264
rect 22100 17187 22152 17196
rect 22100 17153 22109 17187
rect 22109 17153 22143 17187
rect 22143 17153 22152 17187
rect 22100 17144 22152 17153
rect 19340 17076 19392 17085
rect 22468 17076 22520 17128
rect 23388 17076 23440 17128
rect 24768 17076 24820 17128
rect 25228 17119 25280 17128
rect 25228 17085 25237 17119
rect 25237 17085 25271 17119
rect 25271 17085 25280 17119
rect 25228 17076 25280 17085
rect 6276 17008 6328 17060
rect 7932 17008 7984 17060
rect 9404 17008 9456 17060
rect 11704 17008 11756 17060
rect 12624 17008 12676 17060
rect 13636 17008 13688 17060
rect 19984 17008 20036 17060
rect 2136 16940 2188 16992
rect 3424 16940 3476 16992
rect 6552 16983 6604 16992
rect 6552 16949 6561 16983
rect 6561 16949 6595 16983
rect 6595 16949 6604 16983
rect 6552 16940 6604 16949
rect 8208 16983 8260 16992
rect 8208 16949 8217 16983
rect 8217 16949 8251 16983
rect 8251 16949 8260 16983
rect 8208 16940 8260 16949
rect 11152 16940 11204 16992
rect 13820 16983 13872 16992
rect 13820 16949 13829 16983
rect 13829 16949 13863 16983
rect 13863 16949 13872 16983
rect 13820 16940 13872 16949
rect 15108 16940 15160 16992
rect 15476 16940 15528 16992
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 16948 16940 17000 16992
rect 17684 16940 17736 16992
rect 18052 16983 18104 16992
rect 18052 16949 18061 16983
rect 18061 16949 18095 16983
rect 18095 16949 18104 16983
rect 18052 16940 18104 16949
rect 20904 16940 20956 16992
rect 22192 17008 22244 17060
rect 21456 16940 21508 16992
rect 22744 16983 22796 16992
rect 22744 16949 22753 16983
rect 22753 16949 22787 16983
rect 22787 16949 22796 16983
rect 22744 16940 22796 16949
rect 23664 16983 23716 16992
rect 23664 16949 23673 16983
rect 23673 16949 23707 16983
rect 23707 16949 23716 16983
rect 23664 16940 23716 16949
rect 25136 16983 25188 16992
rect 25136 16949 25145 16983
rect 25145 16949 25179 16983
rect 25179 16949 25188 16983
rect 25136 16940 25188 16949
rect 10315 16838 10367 16890
rect 10379 16838 10431 16890
rect 10443 16838 10495 16890
rect 10507 16838 10559 16890
rect 19648 16838 19700 16890
rect 19712 16838 19764 16890
rect 19776 16838 19828 16890
rect 19840 16838 19892 16890
rect 2596 16736 2648 16788
rect 2780 16736 2832 16788
rect 3516 16779 3568 16788
rect 3516 16745 3525 16779
rect 3525 16745 3559 16779
rect 3559 16745 3568 16779
rect 3516 16736 3568 16745
rect 3792 16779 3844 16788
rect 3792 16745 3801 16779
rect 3801 16745 3835 16779
rect 3835 16745 3844 16779
rect 3792 16736 3844 16745
rect 5540 16736 5592 16788
rect 7932 16779 7984 16788
rect 2504 16668 2556 16720
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 2044 16600 2096 16652
rect 3056 16600 3108 16652
rect 1952 16532 2004 16584
rect 2412 16532 2464 16584
rect 2964 16575 3016 16584
rect 2964 16541 2973 16575
rect 2973 16541 3007 16575
rect 3007 16541 3016 16575
rect 2964 16532 3016 16541
rect 3424 16668 3476 16720
rect 7932 16745 7941 16779
rect 7941 16745 7975 16779
rect 7975 16745 7984 16779
rect 7932 16736 7984 16745
rect 8024 16736 8076 16788
rect 8576 16736 8628 16788
rect 8668 16736 8720 16788
rect 9404 16779 9456 16788
rect 9404 16745 9413 16779
rect 9413 16745 9447 16779
rect 9447 16745 9456 16779
rect 9404 16736 9456 16745
rect 9956 16779 10008 16788
rect 9956 16745 9965 16779
rect 9965 16745 9999 16779
rect 9999 16745 10008 16779
rect 9956 16736 10008 16745
rect 11704 16779 11756 16788
rect 11704 16745 11713 16779
rect 11713 16745 11747 16779
rect 11747 16745 11756 16779
rect 11704 16736 11756 16745
rect 12808 16779 12860 16788
rect 12808 16745 12817 16779
rect 12817 16745 12851 16779
rect 12851 16745 12860 16779
rect 12808 16736 12860 16745
rect 14188 16779 14240 16788
rect 14188 16745 14197 16779
rect 14197 16745 14231 16779
rect 14231 16745 14240 16779
rect 14188 16736 14240 16745
rect 14556 16779 14608 16788
rect 14556 16745 14565 16779
rect 14565 16745 14599 16779
rect 14599 16745 14608 16779
rect 14556 16736 14608 16745
rect 14832 16736 14884 16788
rect 16028 16736 16080 16788
rect 16580 16736 16632 16788
rect 17408 16736 17460 16788
rect 17868 16736 17920 16788
rect 18328 16736 18380 16788
rect 19248 16736 19300 16788
rect 20260 16779 20312 16788
rect 20260 16745 20269 16779
rect 20269 16745 20303 16779
rect 20303 16745 20312 16779
rect 20260 16736 20312 16745
rect 20628 16779 20680 16788
rect 20628 16745 20637 16779
rect 20637 16745 20671 16779
rect 20671 16745 20680 16779
rect 20628 16736 20680 16745
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 22652 16779 22704 16788
rect 7012 16668 7064 16720
rect 4620 16600 4672 16652
rect 6368 16600 6420 16652
rect 6460 16600 6512 16652
rect 8484 16600 8536 16652
rect 9036 16643 9088 16652
rect 9036 16609 9045 16643
rect 9045 16609 9079 16643
rect 9079 16609 9088 16643
rect 9036 16600 9088 16609
rect 10140 16668 10192 16720
rect 13452 16668 13504 16720
rect 14924 16711 14976 16720
rect 14924 16677 14933 16711
rect 14933 16677 14967 16711
rect 14967 16677 14976 16711
rect 14924 16668 14976 16677
rect 10324 16643 10376 16652
rect 10324 16609 10333 16643
rect 10333 16609 10367 16643
rect 10367 16609 10376 16643
rect 10324 16600 10376 16609
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 15752 16643 15804 16652
rect 15752 16609 15761 16643
rect 15761 16609 15795 16643
rect 15795 16609 15804 16643
rect 15752 16600 15804 16609
rect 3608 16532 3660 16584
rect 6276 16532 6328 16584
rect 13268 16575 13320 16584
rect 13268 16541 13277 16575
rect 13277 16541 13311 16575
rect 13311 16541 13320 16575
rect 13268 16532 13320 16541
rect 13728 16532 13780 16584
rect 15936 16532 15988 16584
rect 2412 16439 2464 16448
rect 2412 16405 2421 16439
rect 2421 16405 2455 16439
rect 2455 16405 2464 16439
rect 2412 16396 2464 16405
rect 2688 16396 2740 16448
rect 4988 16396 5040 16448
rect 5448 16439 5500 16448
rect 5448 16405 5457 16439
rect 5457 16405 5491 16439
rect 5491 16405 5500 16439
rect 5448 16396 5500 16405
rect 11428 16464 11480 16516
rect 11704 16464 11756 16516
rect 16304 16464 16356 16516
rect 16856 16464 16908 16516
rect 18144 16668 18196 16720
rect 18972 16668 19024 16720
rect 19984 16668 20036 16720
rect 19340 16600 19392 16652
rect 20812 16668 20864 16720
rect 21364 16711 21416 16720
rect 21364 16677 21373 16711
rect 21373 16677 21407 16711
rect 21407 16677 21416 16711
rect 21364 16668 21416 16677
rect 21272 16643 21324 16652
rect 17684 16532 17736 16584
rect 19156 16532 19208 16584
rect 21272 16609 21281 16643
rect 21281 16609 21315 16643
rect 21315 16609 21324 16643
rect 21272 16600 21324 16609
rect 22652 16745 22661 16779
rect 22661 16745 22695 16779
rect 22695 16745 22704 16779
rect 22652 16736 22704 16745
rect 22836 16736 22888 16788
rect 25596 16736 25648 16788
rect 22284 16668 22336 16720
rect 24860 16668 24912 16720
rect 20812 16532 20864 16584
rect 22652 16532 22704 16584
rect 17960 16464 18012 16516
rect 19984 16464 20036 16516
rect 22100 16464 22152 16516
rect 25044 16532 25096 16584
rect 26056 16464 26108 16516
rect 7196 16396 7248 16448
rect 12624 16396 12676 16448
rect 16764 16439 16816 16448
rect 16764 16405 16773 16439
rect 16773 16405 16807 16439
rect 16807 16405 16816 16439
rect 16764 16396 16816 16405
rect 18052 16439 18104 16448
rect 18052 16405 18061 16439
rect 18061 16405 18095 16439
rect 18095 16405 18104 16439
rect 18052 16396 18104 16405
rect 18328 16439 18380 16448
rect 18328 16405 18337 16439
rect 18337 16405 18371 16439
rect 18371 16405 18380 16439
rect 18328 16396 18380 16405
rect 23756 16396 23808 16448
rect 23940 16396 23992 16448
rect 24676 16396 24728 16448
rect 5648 16294 5700 16346
rect 5712 16294 5764 16346
rect 5776 16294 5828 16346
rect 5840 16294 5892 16346
rect 14982 16294 15034 16346
rect 15046 16294 15098 16346
rect 15110 16294 15162 16346
rect 15174 16294 15226 16346
rect 24315 16294 24367 16346
rect 24379 16294 24431 16346
rect 24443 16294 24495 16346
rect 24507 16294 24559 16346
rect 2964 16192 3016 16244
rect 5540 16192 5592 16244
rect 2504 16056 2556 16108
rect 3056 16056 3108 16108
rect 5632 16124 5684 16176
rect 6276 16192 6328 16244
rect 8668 16099 8720 16108
rect 1860 15988 1912 16040
rect 2228 15920 2280 15972
rect 2044 15895 2096 15904
rect 2044 15861 2053 15895
rect 2053 15861 2087 15895
rect 2087 15861 2096 15895
rect 2044 15852 2096 15861
rect 3700 15988 3752 16040
rect 3976 15988 4028 16040
rect 8668 16065 8677 16099
rect 8677 16065 8711 16099
rect 8711 16065 8720 16099
rect 8668 16056 8720 16065
rect 10324 16192 10376 16244
rect 10784 16235 10836 16244
rect 10784 16201 10793 16235
rect 10793 16201 10827 16235
rect 10827 16201 10836 16235
rect 10784 16192 10836 16201
rect 12532 16235 12584 16244
rect 12532 16201 12541 16235
rect 12541 16201 12575 16235
rect 12575 16201 12584 16235
rect 12532 16192 12584 16201
rect 9220 16056 9272 16108
rect 10140 16056 10192 16108
rect 12992 16099 13044 16108
rect 12992 16065 13001 16099
rect 13001 16065 13035 16099
rect 13035 16065 13044 16099
rect 12992 16056 13044 16065
rect 13728 16192 13780 16244
rect 15936 16235 15988 16244
rect 15936 16201 15945 16235
rect 15945 16201 15979 16235
rect 15979 16201 15988 16235
rect 15936 16192 15988 16201
rect 16396 16235 16448 16244
rect 16396 16201 16405 16235
rect 16405 16201 16439 16235
rect 16439 16201 16448 16235
rect 16396 16192 16448 16201
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 18972 16192 19024 16244
rect 19524 16192 19576 16244
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 22284 16192 22336 16244
rect 22652 16192 22704 16244
rect 23388 16235 23440 16244
rect 23388 16201 23397 16235
rect 23397 16201 23431 16235
rect 23431 16201 23440 16235
rect 23388 16192 23440 16201
rect 23848 16192 23900 16244
rect 24124 16192 24176 16244
rect 25412 16235 25464 16244
rect 25412 16201 25421 16235
rect 25421 16201 25455 16235
rect 25455 16201 25464 16235
rect 25412 16192 25464 16201
rect 17408 16167 17460 16176
rect 8392 15988 8444 16040
rect 8576 16031 8628 16040
rect 8576 15997 8585 16031
rect 8585 15997 8619 16031
rect 8619 15997 8628 16031
rect 8576 15988 8628 15997
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 12072 15988 12124 16040
rect 17408 16133 17417 16167
rect 17417 16133 17451 16167
rect 17451 16133 17460 16167
rect 17408 16124 17460 16133
rect 21272 16124 21324 16176
rect 14004 16056 14056 16108
rect 16304 16056 16356 16108
rect 17684 16056 17736 16108
rect 18052 16056 18104 16108
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19432 16056 19484 16108
rect 20536 16056 20588 16108
rect 21916 16056 21968 16108
rect 22100 16056 22152 16108
rect 14464 15988 14516 16040
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 19984 16031 20036 16040
rect 19984 15997 19993 16031
rect 19993 15997 20027 16031
rect 20027 15997 20036 16031
rect 19984 15988 20036 15997
rect 20720 15988 20772 16040
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 25228 16031 25280 16040
rect 25228 15997 25237 16031
rect 25237 15997 25271 16031
rect 25271 15997 25280 16031
rect 25228 15988 25280 15997
rect 8024 15920 8076 15972
rect 14004 15963 14056 15972
rect 14004 15929 14013 15963
rect 14013 15929 14047 15963
rect 14047 15929 14056 15963
rect 14004 15920 14056 15929
rect 15292 15963 15344 15972
rect 15292 15929 15301 15963
rect 15301 15929 15335 15963
rect 15335 15929 15344 15963
rect 15292 15920 15344 15929
rect 2688 15852 2740 15904
rect 3424 15895 3476 15904
rect 3424 15861 3433 15895
rect 3433 15861 3467 15895
rect 3467 15861 3476 15895
rect 3424 15852 3476 15861
rect 3608 15895 3660 15904
rect 3608 15861 3617 15895
rect 3617 15861 3651 15895
rect 3651 15861 3660 15895
rect 3608 15852 3660 15861
rect 3884 15852 3936 15904
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 5540 15895 5592 15904
rect 5540 15861 5549 15895
rect 5549 15861 5583 15895
rect 5583 15861 5592 15895
rect 5540 15852 5592 15861
rect 6368 15852 6420 15904
rect 6552 15895 6604 15904
rect 6552 15861 6561 15895
rect 6561 15861 6595 15895
rect 6595 15861 6604 15895
rect 6552 15852 6604 15861
rect 7012 15895 7064 15904
rect 7012 15861 7021 15895
rect 7021 15861 7055 15895
rect 7055 15861 7064 15895
rect 7012 15852 7064 15861
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 9680 15852 9732 15904
rect 13820 15852 13872 15904
rect 15016 15852 15068 15904
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 16212 15852 16264 15904
rect 16672 15852 16724 15904
rect 16856 15895 16908 15904
rect 16856 15861 16865 15895
rect 16865 15861 16899 15895
rect 16899 15861 16908 15895
rect 16856 15852 16908 15861
rect 17592 15852 17644 15904
rect 20628 15920 20680 15972
rect 21088 15920 21140 15972
rect 23296 15920 23348 15972
rect 25320 15920 25372 15972
rect 19156 15852 19208 15904
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 20904 15852 20956 15904
rect 24032 15895 24084 15904
rect 24032 15861 24041 15895
rect 24041 15861 24075 15895
rect 24075 15861 24084 15895
rect 24032 15852 24084 15861
rect 25044 15895 25096 15904
rect 25044 15861 25053 15895
rect 25053 15861 25087 15895
rect 25087 15861 25096 15895
rect 25044 15852 25096 15861
rect 10315 15750 10367 15802
rect 10379 15750 10431 15802
rect 10443 15750 10495 15802
rect 10507 15750 10559 15802
rect 19648 15750 19700 15802
rect 19712 15750 19764 15802
rect 19776 15750 19828 15802
rect 19840 15750 19892 15802
rect 3700 15691 3752 15700
rect 3700 15657 3709 15691
rect 3709 15657 3743 15691
rect 3743 15657 3752 15691
rect 3700 15648 3752 15657
rect 6276 15691 6328 15700
rect 6276 15657 6285 15691
rect 6285 15657 6319 15691
rect 6319 15657 6328 15691
rect 6276 15648 6328 15657
rect 7196 15691 7248 15700
rect 7196 15657 7205 15691
rect 7205 15657 7239 15691
rect 7239 15657 7248 15691
rect 7196 15648 7248 15657
rect 8116 15648 8168 15700
rect 8852 15648 8904 15700
rect 9404 15691 9456 15700
rect 9404 15657 9413 15691
rect 9413 15657 9447 15691
rect 9447 15657 9456 15691
rect 9404 15648 9456 15657
rect 9496 15648 9548 15700
rect 10140 15691 10192 15700
rect 10140 15657 10149 15691
rect 10149 15657 10183 15691
rect 10183 15657 10192 15691
rect 10140 15648 10192 15657
rect 12440 15648 12492 15700
rect 13544 15648 13596 15700
rect 14372 15691 14424 15700
rect 14372 15657 14381 15691
rect 14381 15657 14415 15691
rect 14415 15657 14424 15691
rect 14372 15648 14424 15657
rect 14740 15691 14792 15700
rect 14740 15657 14749 15691
rect 14749 15657 14783 15691
rect 14783 15657 14792 15691
rect 14740 15648 14792 15657
rect 15568 15691 15620 15700
rect 15568 15657 15577 15691
rect 15577 15657 15611 15691
rect 15611 15657 15620 15691
rect 15568 15648 15620 15657
rect 17316 15648 17368 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 17960 15648 18012 15700
rect 18328 15648 18380 15700
rect 20168 15648 20220 15700
rect 21548 15648 21600 15700
rect 3792 15580 3844 15632
rect 5448 15580 5500 15632
rect 8668 15580 8720 15632
rect 11060 15580 11112 15632
rect 13268 15580 13320 15632
rect 13728 15623 13780 15632
rect 13728 15589 13737 15623
rect 13737 15589 13771 15623
rect 13771 15589 13780 15623
rect 13728 15580 13780 15589
rect 18420 15580 18472 15632
rect 20536 15580 20588 15632
rect 20720 15580 20772 15632
rect 22100 15648 22152 15700
rect 24492 15691 24544 15700
rect 24492 15657 24501 15691
rect 24501 15657 24535 15691
rect 24535 15657 24544 15691
rect 24492 15648 24544 15657
rect 24860 15648 24912 15700
rect 22652 15580 22704 15632
rect 24032 15580 24084 15632
rect 2412 15512 2464 15564
rect 2964 15512 3016 15564
rect 4620 15512 4672 15564
rect 6552 15512 6604 15564
rect 8484 15512 8536 15564
rect 10784 15512 10836 15564
rect 15568 15512 15620 15564
rect 16304 15512 16356 15564
rect 17684 15512 17736 15564
rect 19984 15512 20036 15564
rect 20996 15512 21048 15564
rect 21732 15512 21784 15564
rect 22008 15555 22060 15564
rect 22008 15521 22017 15555
rect 22017 15521 22051 15555
rect 22051 15521 22060 15555
rect 22008 15512 22060 15521
rect 22836 15512 22888 15564
rect 24952 15580 25004 15632
rect 3056 15487 3108 15496
rect 3056 15453 3065 15487
rect 3065 15453 3099 15487
rect 3099 15453 3108 15487
rect 3056 15444 3108 15453
rect 4068 15444 4120 15496
rect 4712 15444 4764 15496
rect 14004 15487 14056 15496
rect 1860 15376 1912 15428
rect 8024 15419 8076 15428
rect 8024 15385 8033 15419
rect 8033 15385 8067 15419
rect 8067 15385 8076 15419
rect 8024 15376 8076 15385
rect 8300 15376 8352 15428
rect 14004 15453 14013 15487
rect 14013 15453 14047 15487
rect 14047 15453 14056 15487
rect 14004 15444 14056 15453
rect 13452 15376 13504 15428
rect 18696 15444 18748 15496
rect 20812 15444 20864 15496
rect 24952 15487 25004 15496
rect 24952 15453 24961 15487
rect 24961 15453 24995 15487
rect 24995 15453 25004 15487
rect 24952 15444 25004 15453
rect 18144 15376 18196 15428
rect 19524 15376 19576 15428
rect 21916 15376 21968 15428
rect 24768 15376 24820 15428
rect 25964 15376 26016 15428
rect 2228 15308 2280 15360
rect 2596 15308 2648 15360
rect 8576 15308 8628 15360
rect 10508 15351 10560 15360
rect 10508 15317 10517 15351
rect 10517 15317 10551 15351
rect 10551 15317 10560 15351
rect 10508 15308 10560 15317
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 13360 15351 13412 15360
rect 13360 15317 13369 15351
rect 13369 15317 13403 15351
rect 13403 15317 13412 15351
rect 13360 15308 13412 15317
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 20352 15351 20404 15360
rect 20352 15317 20361 15351
rect 20361 15317 20395 15351
rect 20395 15317 20404 15351
rect 20352 15308 20404 15317
rect 20628 15308 20680 15360
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 24124 15308 24176 15360
rect 5648 15206 5700 15258
rect 5712 15206 5764 15258
rect 5776 15206 5828 15258
rect 5840 15206 5892 15258
rect 14982 15206 15034 15258
rect 15046 15206 15098 15258
rect 15110 15206 15162 15258
rect 15174 15206 15226 15258
rect 24315 15206 24367 15258
rect 24379 15206 24431 15258
rect 24443 15206 24495 15258
rect 24507 15206 24559 15258
rect 2872 15104 2924 15156
rect 1584 15079 1636 15088
rect 1584 15045 1593 15079
rect 1593 15045 1627 15079
rect 1627 15045 1636 15079
rect 1584 15036 1636 15045
rect 6276 15104 6328 15156
rect 6920 15104 6972 15156
rect 8484 15104 8536 15156
rect 8852 15104 8904 15156
rect 10784 15104 10836 15156
rect 11152 15104 11204 15156
rect 11428 15104 11480 15156
rect 13544 15147 13596 15156
rect 13544 15113 13553 15147
rect 13553 15113 13587 15147
rect 13587 15113 13596 15147
rect 13544 15104 13596 15113
rect 13912 15104 13964 15156
rect 16764 15104 16816 15156
rect 17684 15104 17736 15156
rect 17868 15147 17920 15156
rect 17868 15113 17877 15147
rect 17877 15113 17911 15147
rect 17911 15113 17920 15147
rect 17868 15104 17920 15113
rect 22468 15104 22520 15156
rect 22836 15104 22888 15156
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 24216 15104 24268 15156
rect 25964 15104 26016 15156
rect 3792 15036 3844 15088
rect 4068 15036 4120 15088
rect 14004 15036 14056 15088
rect 22008 15036 22060 15088
rect 22284 15036 22336 15088
rect 22652 15036 22704 15088
rect 3516 14968 3568 15020
rect 7472 14968 7524 15020
rect 8300 14968 8352 15020
rect 11060 14968 11112 15020
rect 13452 14968 13504 15020
rect 13820 14968 13872 15020
rect 20720 14968 20772 15020
rect 24860 15036 24912 15088
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 3056 14832 3108 14884
rect 4712 14900 4764 14952
rect 7196 14900 7248 14952
rect 8024 14900 8076 14952
rect 14188 14900 14240 14952
rect 14464 14900 14516 14952
rect 15568 14900 15620 14952
rect 18236 14900 18288 14952
rect 19340 14943 19392 14952
rect 19340 14909 19349 14943
rect 19349 14909 19383 14943
rect 19383 14909 19392 14943
rect 19340 14900 19392 14909
rect 19524 14900 19576 14952
rect 22100 14900 22152 14952
rect 4528 14832 4580 14884
rect 7380 14832 7432 14884
rect 7748 14832 7800 14884
rect 8576 14832 8628 14884
rect 9036 14832 9088 14884
rect 10784 14832 10836 14884
rect 13360 14832 13412 14884
rect 13728 14832 13780 14884
rect 16488 14832 16540 14884
rect 18052 14832 18104 14884
rect 18880 14875 18932 14884
rect 18880 14841 18889 14875
rect 18889 14841 18923 14875
rect 18923 14841 18932 14875
rect 18880 14832 18932 14841
rect 20352 14832 20404 14884
rect 23940 14900 23992 14952
rect 24952 14900 25004 14952
rect 24032 14875 24084 14884
rect 24032 14841 24041 14875
rect 24041 14841 24075 14875
rect 24075 14841 24084 14875
rect 24032 14832 24084 14841
rect 2044 14807 2096 14816
rect 2044 14773 2053 14807
rect 2053 14773 2087 14807
rect 2087 14773 2096 14807
rect 2044 14764 2096 14773
rect 2872 14764 2924 14816
rect 5540 14807 5592 14816
rect 5540 14773 5549 14807
rect 5549 14773 5583 14807
rect 5583 14773 5592 14807
rect 5540 14764 5592 14773
rect 6552 14764 6604 14816
rect 9496 14764 9548 14816
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 11152 14764 11204 14773
rect 12532 14807 12584 14816
rect 12532 14773 12541 14807
rect 12541 14773 12575 14807
rect 12575 14773 12584 14807
rect 12532 14764 12584 14773
rect 13084 14764 13136 14816
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 18512 14807 18564 14816
rect 18512 14773 18521 14807
rect 18521 14773 18555 14807
rect 18555 14773 18564 14807
rect 18512 14764 18564 14773
rect 21916 14807 21968 14816
rect 21916 14773 21925 14807
rect 21925 14773 21959 14807
rect 21959 14773 21968 14807
rect 21916 14764 21968 14773
rect 22284 14807 22336 14816
rect 22284 14773 22293 14807
rect 22293 14773 22327 14807
rect 22327 14773 22336 14807
rect 22284 14764 22336 14773
rect 23664 14807 23716 14816
rect 23664 14773 23673 14807
rect 23673 14773 23707 14807
rect 23707 14773 23716 14807
rect 23664 14764 23716 14773
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 10315 14662 10367 14714
rect 10379 14662 10431 14714
rect 10443 14662 10495 14714
rect 10507 14662 10559 14714
rect 19648 14662 19700 14714
rect 19712 14662 19764 14714
rect 19776 14662 19828 14714
rect 19840 14662 19892 14714
rect 2320 14560 2372 14612
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 3332 14560 3384 14612
rect 4528 14560 4580 14612
rect 6276 14603 6328 14612
rect 6276 14569 6285 14603
rect 6285 14569 6319 14603
rect 6319 14569 6328 14603
rect 6276 14560 6328 14569
rect 7472 14603 7524 14612
rect 7472 14569 7481 14603
rect 7481 14569 7515 14603
rect 7515 14569 7524 14603
rect 7472 14560 7524 14569
rect 11060 14603 11112 14612
rect 2872 14535 2924 14544
rect 2872 14501 2881 14535
rect 2881 14501 2915 14535
rect 2915 14501 2924 14535
rect 2872 14492 2924 14501
rect 3516 14535 3568 14544
rect 3516 14501 3525 14535
rect 3525 14501 3559 14535
rect 3559 14501 3568 14535
rect 3516 14492 3568 14501
rect 2780 14467 2832 14476
rect 2780 14433 2789 14467
rect 2789 14433 2823 14467
rect 2823 14433 2832 14467
rect 2780 14424 2832 14433
rect 4712 14492 4764 14544
rect 5540 14492 5592 14544
rect 11060 14569 11069 14603
rect 11069 14569 11103 14603
rect 11103 14569 11112 14603
rect 11060 14560 11112 14569
rect 11336 14603 11388 14612
rect 11336 14569 11345 14603
rect 11345 14569 11379 14603
rect 11379 14569 11388 14603
rect 11336 14560 11388 14569
rect 12992 14560 13044 14612
rect 13360 14560 13412 14612
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14832 14603 14884 14612
rect 14832 14569 14841 14603
rect 14841 14569 14875 14603
rect 14875 14569 14884 14603
rect 14832 14560 14884 14569
rect 16304 14603 16356 14612
rect 16304 14569 16313 14603
rect 16313 14569 16347 14603
rect 16347 14569 16356 14603
rect 16304 14560 16356 14569
rect 16856 14560 16908 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21824 14560 21876 14612
rect 22284 14560 22336 14612
rect 22836 14560 22888 14612
rect 23112 14560 23164 14612
rect 24952 14603 25004 14612
rect 24952 14569 24961 14603
rect 24961 14569 24995 14603
rect 24995 14569 25004 14603
rect 24952 14560 25004 14569
rect 5632 14424 5684 14476
rect 6828 14467 6880 14476
rect 6828 14433 6837 14467
rect 6837 14433 6871 14467
rect 6871 14433 6880 14467
rect 6828 14424 6880 14433
rect 8392 14467 8444 14476
rect 8392 14433 8401 14467
rect 8401 14433 8435 14467
rect 8435 14433 8444 14467
rect 8392 14424 8444 14433
rect 12256 14492 12308 14544
rect 12440 14535 12492 14544
rect 12440 14501 12474 14535
rect 12474 14501 12492 14535
rect 14556 14535 14608 14544
rect 12440 14492 12492 14501
rect 14556 14501 14565 14535
rect 14565 14501 14599 14535
rect 14599 14501 14608 14535
rect 14556 14492 14608 14501
rect 15108 14492 15160 14544
rect 17776 14492 17828 14544
rect 2136 14356 2188 14408
rect 10784 14424 10836 14476
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 15568 14424 15620 14476
rect 16396 14424 16448 14476
rect 18880 14492 18932 14544
rect 7012 14331 7064 14340
rect 7012 14297 7021 14331
rect 7021 14297 7055 14331
rect 7055 14297 7064 14331
rect 7012 14288 7064 14297
rect 7840 14288 7892 14340
rect 8760 14356 8812 14408
rect 10048 14356 10100 14408
rect 11060 14356 11112 14408
rect 12164 14399 12216 14408
rect 12164 14365 12173 14399
rect 12173 14365 12207 14399
rect 12207 14365 12216 14399
rect 12164 14356 12216 14365
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 17592 14356 17644 14408
rect 18788 14356 18840 14408
rect 19248 14356 19300 14408
rect 20996 14492 21048 14544
rect 22468 14492 22520 14544
rect 19616 14424 19668 14476
rect 20260 14356 20312 14408
rect 20444 14356 20496 14408
rect 21088 14424 21140 14476
rect 22008 14467 22060 14476
rect 22008 14433 22017 14467
rect 22017 14433 22051 14467
rect 22051 14433 22060 14467
rect 22008 14424 22060 14433
rect 24216 14424 24268 14476
rect 24860 14467 24912 14476
rect 24860 14433 24869 14467
rect 24869 14433 24903 14467
rect 24903 14433 24912 14467
rect 24860 14424 24912 14433
rect 25228 14424 25280 14476
rect 24676 14356 24728 14408
rect 9220 14288 9272 14340
rect 14280 14288 14332 14340
rect 15844 14331 15896 14340
rect 15844 14297 15853 14331
rect 15853 14297 15887 14331
rect 15887 14297 15896 14331
rect 15844 14288 15896 14297
rect 22008 14288 22060 14340
rect 23480 14288 23532 14340
rect 24032 14288 24084 14340
rect 1860 14220 1912 14272
rect 4160 14220 4212 14272
rect 5540 14220 5592 14272
rect 6276 14220 6328 14272
rect 9036 14263 9088 14272
rect 9036 14229 9045 14263
rect 9045 14229 9079 14263
rect 9079 14229 9088 14263
rect 9036 14220 9088 14229
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 9956 14263 10008 14272
rect 9956 14229 9965 14263
rect 9965 14229 9999 14263
rect 9999 14229 10008 14263
rect 9956 14220 10008 14229
rect 17868 14263 17920 14272
rect 17868 14229 17877 14263
rect 17877 14229 17911 14263
rect 17911 14229 17920 14263
rect 17868 14220 17920 14229
rect 19524 14220 19576 14272
rect 20076 14220 20128 14272
rect 20444 14220 20496 14272
rect 20536 14220 20588 14272
rect 24952 14288 25004 14340
rect 24676 14220 24728 14272
rect 25228 14220 25280 14272
rect 5648 14118 5700 14170
rect 5712 14118 5764 14170
rect 5776 14118 5828 14170
rect 5840 14118 5892 14170
rect 14982 14118 15034 14170
rect 15046 14118 15098 14170
rect 15110 14118 15162 14170
rect 15174 14118 15226 14170
rect 24315 14118 24367 14170
rect 24379 14118 24431 14170
rect 24443 14118 24495 14170
rect 24507 14118 24559 14170
rect 2780 14016 2832 14068
rect 3240 14016 3292 14068
rect 3700 14016 3752 14068
rect 5172 14016 5224 14068
rect 9220 14059 9272 14068
rect 9220 14025 9229 14059
rect 9229 14025 9263 14059
rect 9263 14025 9272 14059
rect 9220 14016 9272 14025
rect 2228 13948 2280 14000
rect 3516 13948 3568 14000
rect 4988 13991 5040 14000
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 1952 13812 2004 13864
rect 4988 13957 4997 13991
rect 4997 13957 5031 13991
rect 5031 13957 5040 13991
rect 4988 13948 5040 13957
rect 8576 13991 8628 14000
rect 8576 13957 8585 13991
rect 8585 13957 8619 13991
rect 8619 13957 8628 13991
rect 8576 13948 8628 13957
rect 11060 14016 11112 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 12900 14016 12952 14068
rect 13452 14059 13504 14068
rect 13452 14025 13461 14059
rect 13461 14025 13495 14059
rect 13495 14025 13504 14059
rect 13452 14016 13504 14025
rect 16212 14016 16264 14068
rect 16396 14016 16448 14068
rect 4160 13880 4212 13932
rect 9036 13880 9088 13932
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 6276 13812 6328 13864
rect 7840 13812 7892 13864
rect 4620 13744 4672 13796
rect 5356 13787 5408 13796
rect 5356 13753 5365 13787
rect 5365 13753 5399 13787
rect 5399 13753 5408 13787
rect 5356 13744 5408 13753
rect 6460 13744 6512 13796
rect 12440 13880 12492 13932
rect 12992 13880 13044 13932
rect 13452 13880 13504 13932
rect 17776 14016 17828 14068
rect 19248 14016 19300 14068
rect 20536 14016 20588 14068
rect 20628 14016 20680 14068
rect 21088 14016 21140 14068
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 22100 14016 22152 14068
rect 23296 14016 23348 14068
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 12900 13812 12952 13821
rect 13820 13812 13872 13864
rect 14924 13812 14976 13864
rect 15844 13812 15896 13864
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 16488 13812 16540 13864
rect 17868 13812 17920 13864
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 20720 13880 20772 13932
rect 22100 13812 22152 13864
rect 22836 13812 22888 13864
rect 24032 14016 24084 14068
rect 24860 14016 24912 14068
rect 24952 14016 25004 14068
rect 25504 14016 25556 14068
rect 23480 13948 23532 14000
rect 24216 13923 24268 13932
rect 24216 13889 24225 13923
rect 24225 13889 24259 13923
rect 24259 13889 24268 13923
rect 24216 13880 24268 13889
rect 24860 13812 24912 13864
rect 26240 13855 26292 13864
rect 26240 13821 26249 13855
rect 26249 13821 26283 13855
rect 26283 13821 26292 13855
rect 26240 13812 26292 13821
rect 9496 13744 9548 13796
rect 10600 13744 10652 13796
rect 11060 13744 11112 13796
rect 12532 13744 12584 13796
rect 13728 13744 13780 13796
rect 16028 13744 16080 13796
rect 17960 13744 18012 13796
rect 19524 13744 19576 13796
rect 22376 13744 22428 13796
rect 23020 13744 23072 13796
rect 1768 13676 1820 13728
rect 2320 13676 2372 13728
rect 2596 13676 2648 13728
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 6552 13719 6604 13728
rect 6552 13685 6561 13719
rect 6561 13685 6595 13719
rect 6595 13685 6604 13719
rect 6552 13676 6604 13685
rect 13268 13676 13320 13728
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 14188 13676 14240 13728
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 18328 13719 18380 13728
rect 18328 13685 18337 13719
rect 18337 13685 18371 13719
rect 18371 13685 18380 13719
rect 18328 13676 18380 13685
rect 19156 13676 19208 13728
rect 21916 13676 21968 13728
rect 22100 13676 22152 13728
rect 22468 13676 22520 13728
rect 23572 13676 23624 13728
rect 25228 13676 25280 13728
rect 10315 13574 10367 13626
rect 10379 13574 10431 13626
rect 10443 13574 10495 13626
rect 10507 13574 10559 13626
rect 19648 13574 19700 13626
rect 19712 13574 19764 13626
rect 19776 13574 19828 13626
rect 19840 13574 19892 13626
rect 2136 13472 2188 13524
rect 2412 13472 2464 13524
rect 3240 13515 3292 13524
rect 3240 13481 3249 13515
rect 3249 13481 3283 13515
rect 3283 13481 3292 13515
rect 3240 13472 3292 13481
rect 4712 13515 4764 13524
rect 4712 13481 4721 13515
rect 4721 13481 4755 13515
rect 4755 13481 4764 13515
rect 4712 13472 4764 13481
rect 4896 13515 4948 13524
rect 4896 13481 4905 13515
rect 4905 13481 4939 13515
rect 4939 13481 4948 13515
rect 4896 13472 4948 13481
rect 7840 13515 7892 13524
rect 7840 13481 7849 13515
rect 7849 13481 7883 13515
rect 7883 13481 7892 13515
rect 7840 13472 7892 13481
rect 8760 13515 8812 13524
rect 8760 13481 8769 13515
rect 8769 13481 8803 13515
rect 8803 13481 8812 13515
rect 8760 13472 8812 13481
rect 9496 13515 9548 13524
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 9956 13472 10008 13524
rect 11336 13472 11388 13524
rect 2688 13404 2740 13456
rect 4988 13404 5040 13456
rect 6552 13404 6604 13456
rect 2228 13379 2280 13388
rect 2228 13345 2237 13379
rect 2237 13345 2271 13379
rect 2271 13345 2280 13379
rect 2228 13336 2280 13345
rect 3608 13336 3660 13388
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 3056 13268 3108 13320
rect 3424 13268 3476 13320
rect 4160 13268 4212 13320
rect 4528 13268 4580 13320
rect 4712 13268 4764 13320
rect 6000 13336 6052 13388
rect 9772 13336 9824 13388
rect 5448 13311 5500 13320
rect 5448 13277 5457 13311
rect 5457 13277 5491 13311
rect 5491 13277 5500 13311
rect 6460 13311 6512 13320
rect 5448 13268 5500 13277
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 9588 13268 9640 13320
rect 10600 13336 10652 13388
rect 1400 13200 1452 13252
rect 1952 13200 2004 13252
rect 8392 13200 8444 13252
rect 9036 13200 9088 13252
rect 11244 13243 11296 13252
rect 11244 13209 11253 13243
rect 11253 13209 11287 13243
rect 11287 13209 11296 13243
rect 11244 13200 11296 13209
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 13636 13472 13688 13524
rect 14096 13472 14148 13524
rect 14556 13515 14608 13524
rect 14556 13481 14565 13515
rect 14565 13481 14599 13515
rect 14599 13481 14608 13515
rect 14556 13472 14608 13481
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 18236 13515 18288 13524
rect 18236 13481 18245 13515
rect 18245 13481 18279 13515
rect 18279 13481 18288 13515
rect 18236 13472 18288 13481
rect 20904 13515 20956 13524
rect 20904 13481 20913 13515
rect 20913 13481 20947 13515
rect 20947 13481 20956 13515
rect 20904 13472 20956 13481
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 12992 13404 13044 13456
rect 21548 13472 21600 13524
rect 23388 13472 23440 13524
rect 23756 13472 23808 13524
rect 23020 13447 23072 13456
rect 23020 13413 23029 13447
rect 23029 13413 23063 13447
rect 23063 13413 23072 13447
rect 23020 13404 23072 13413
rect 23572 13404 23624 13456
rect 12440 13336 12492 13388
rect 12808 13336 12860 13388
rect 14096 13336 14148 13388
rect 14556 13336 14608 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 18420 13336 18472 13388
rect 20628 13336 20680 13388
rect 21272 13336 21324 13388
rect 21548 13336 21600 13388
rect 22192 13336 22244 13388
rect 22376 13379 22428 13388
rect 22376 13345 22385 13379
rect 22385 13345 22419 13379
rect 22419 13345 22428 13379
rect 22376 13336 22428 13345
rect 22836 13336 22888 13388
rect 23480 13336 23532 13388
rect 24768 13336 24820 13388
rect 12624 13268 12676 13320
rect 12992 13268 13044 13320
rect 13268 13311 13320 13320
rect 13268 13277 13277 13311
rect 13277 13277 13311 13311
rect 13311 13277 13320 13311
rect 13268 13268 13320 13277
rect 13452 13311 13504 13320
rect 13452 13277 13461 13311
rect 13461 13277 13495 13311
rect 13495 13277 13504 13311
rect 13452 13268 13504 13277
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 18052 13268 18104 13320
rect 20812 13268 20864 13320
rect 22652 13268 22704 13320
rect 23112 13311 23164 13320
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 24216 13268 24268 13320
rect 12348 13200 12400 13252
rect 6000 13175 6052 13184
rect 6000 13141 6009 13175
rect 6009 13141 6043 13175
rect 6043 13141 6052 13175
rect 6000 13132 6052 13141
rect 10784 13132 10836 13184
rect 14832 13200 14884 13252
rect 15936 13243 15988 13252
rect 15936 13209 15945 13243
rect 15945 13209 15979 13243
rect 15979 13209 15988 13243
rect 15936 13200 15988 13209
rect 23020 13200 23072 13252
rect 14648 13132 14700 13184
rect 17040 13175 17092 13184
rect 17040 13141 17049 13175
rect 17049 13141 17083 13175
rect 17083 13141 17092 13175
rect 17040 13132 17092 13141
rect 19524 13132 19576 13184
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 19708 13132 19760 13141
rect 20720 13175 20772 13184
rect 20720 13141 20729 13175
rect 20729 13141 20763 13175
rect 20763 13141 20772 13175
rect 20720 13132 20772 13141
rect 22100 13175 22152 13184
rect 22100 13141 22109 13175
rect 22109 13141 22143 13175
rect 22143 13141 22152 13175
rect 22100 13132 22152 13141
rect 22652 13132 22704 13184
rect 25044 13132 25096 13184
rect 25596 13268 25648 13320
rect 25504 13175 25556 13184
rect 25504 13141 25513 13175
rect 25513 13141 25547 13175
rect 25547 13141 25556 13175
rect 25504 13132 25556 13141
rect 25596 13132 25648 13184
rect 26240 13175 26292 13184
rect 26240 13141 26249 13175
rect 26249 13141 26283 13175
rect 26283 13141 26292 13175
rect 26240 13132 26292 13141
rect 5648 13030 5700 13082
rect 5712 13030 5764 13082
rect 5776 13030 5828 13082
rect 5840 13030 5892 13082
rect 14982 13030 15034 13082
rect 15046 13030 15098 13082
rect 15110 13030 15162 13082
rect 15174 13030 15226 13082
rect 24315 13030 24367 13082
rect 24379 13030 24431 13082
rect 24443 13030 24495 13082
rect 24507 13030 24559 13082
rect 296 12928 348 12980
rect 2044 12971 2096 12980
rect 2044 12937 2053 12971
rect 2053 12937 2087 12971
rect 2087 12937 2096 12971
rect 2044 12928 2096 12937
rect 2780 12928 2832 12980
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 3608 12971 3660 12980
rect 3608 12937 3617 12971
rect 3617 12937 3651 12971
rect 3651 12937 3660 12971
rect 3608 12928 3660 12937
rect 8392 12971 8444 12980
rect 8392 12937 8401 12971
rect 8401 12937 8435 12971
rect 8435 12937 8444 12971
rect 8392 12928 8444 12937
rect 8484 12928 8536 12980
rect 8852 12928 8904 12980
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 11428 12928 11480 12980
rect 11704 12928 11756 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13268 12928 13320 12980
rect 5448 12860 5500 12912
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 3976 12792 4028 12844
rect 3884 12724 3936 12776
rect 4252 12792 4304 12844
rect 4988 12792 5040 12844
rect 5172 12792 5224 12844
rect 6184 12860 6236 12912
rect 6460 12860 6512 12912
rect 7196 12860 7248 12912
rect 9588 12860 9640 12912
rect 13820 12928 13872 12980
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 15292 12928 15344 12980
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 16028 12971 16080 12980
rect 16028 12937 16037 12971
rect 16037 12937 16071 12971
rect 16071 12937 16080 12971
rect 16028 12928 16080 12937
rect 16304 12928 16356 12980
rect 18604 12928 18656 12980
rect 19984 12928 20036 12980
rect 20812 12928 20864 12980
rect 21732 12971 21784 12980
rect 21732 12937 21741 12971
rect 21741 12937 21775 12971
rect 21775 12937 21784 12971
rect 21732 12928 21784 12937
rect 13452 12860 13504 12912
rect 6000 12792 6052 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 10600 12835 10652 12844
rect 2136 12656 2188 12708
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 3976 12631 4028 12640
rect 3976 12597 3985 12631
rect 3985 12597 4019 12631
rect 4019 12597 4028 12631
rect 3976 12588 4028 12597
rect 4896 12588 4948 12640
rect 5448 12656 5500 12708
rect 9956 12724 10008 12776
rect 10232 12724 10284 12776
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 11336 12792 11388 12844
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 14648 12792 14700 12844
rect 17224 12860 17276 12912
rect 17592 12860 17644 12912
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 10508 12724 10560 12776
rect 10876 12724 10928 12776
rect 12256 12724 12308 12776
rect 14832 12724 14884 12776
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 18052 12724 18104 12776
rect 5356 12588 5408 12640
rect 5816 12656 5868 12708
rect 9496 12656 9548 12708
rect 6000 12588 6052 12640
rect 6552 12631 6604 12640
rect 6552 12597 6561 12631
rect 6561 12597 6595 12631
rect 6595 12597 6604 12631
rect 6552 12588 6604 12597
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 7288 12631 7340 12640
rect 7288 12597 7297 12631
rect 7297 12597 7331 12631
rect 7331 12597 7340 12631
rect 7288 12588 7340 12597
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 9220 12588 9272 12640
rect 10692 12656 10744 12708
rect 10968 12656 11020 12708
rect 11704 12656 11756 12708
rect 9864 12588 9916 12640
rect 10876 12588 10928 12640
rect 11152 12588 11204 12640
rect 11336 12588 11388 12640
rect 11520 12588 11572 12640
rect 11612 12588 11664 12640
rect 14188 12656 14240 12708
rect 16672 12656 16724 12708
rect 18604 12656 18656 12708
rect 20076 12792 20128 12844
rect 20996 12792 21048 12844
rect 23112 12928 23164 12980
rect 23480 12971 23532 12980
rect 23480 12937 23489 12971
rect 23489 12937 23523 12971
rect 23523 12937 23532 12971
rect 23480 12928 23532 12937
rect 23940 12928 23992 12980
rect 24216 12928 24268 12980
rect 25412 12971 25464 12980
rect 25412 12937 25421 12971
rect 25421 12937 25455 12971
rect 25455 12937 25464 12971
rect 25412 12928 25464 12937
rect 26332 12928 26384 12980
rect 23756 12860 23808 12912
rect 24308 12860 24360 12912
rect 19432 12724 19484 12776
rect 20812 12724 20864 12776
rect 22744 12724 22796 12776
rect 23112 12724 23164 12776
rect 23480 12724 23532 12776
rect 24768 12724 24820 12776
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 25228 12724 25280 12733
rect 25412 12724 25464 12776
rect 19340 12656 19392 12708
rect 22652 12656 22704 12708
rect 24308 12656 24360 12708
rect 13176 12588 13228 12640
rect 13452 12631 13504 12640
rect 13452 12597 13461 12631
rect 13461 12597 13495 12631
rect 13495 12597 13504 12631
rect 13452 12588 13504 12597
rect 14372 12588 14424 12640
rect 15016 12631 15068 12640
rect 15016 12597 15025 12631
rect 15025 12597 15059 12631
rect 15059 12597 15068 12631
rect 15016 12588 15068 12597
rect 16396 12631 16448 12640
rect 16396 12597 16405 12631
rect 16405 12597 16439 12631
rect 16439 12597 16448 12631
rect 16396 12588 16448 12597
rect 18052 12588 18104 12640
rect 18420 12588 18472 12640
rect 20812 12588 20864 12640
rect 22008 12588 22060 12640
rect 23940 12588 23992 12640
rect 25596 12656 25648 12708
rect 10315 12486 10367 12538
rect 10379 12486 10431 12538
rect 10443 12486 10495 12538
rect 10507 12486 10559 12538
rect 19648 12486 19700 12538
rect 19712 12486 19764 12538
rect 19776 12486 19828 12538
rect 19840 12486 19892 12538
rect 1676 12384 1728 12436
rect 2780 12384 2832 12436
rect 4160 12384 4212 12436
rect 4896 12384 4948 12436
rect 7012 12384 7064 12436
rect 7288 12384 7340 12436
rect 8116 12384 8168 12436
rect 8576 12384 8628 12436
rect 20 12316 72 12368
rect 2412 12316 2464 12368
rect 2504 12316 2556 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 3148 12248 3200 12300
rect 4712 12316 4764 12368
rect 5448 12316 5500 12368
rect 2412 12180 2464 12232
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 5632 12248 5684 12300
rect 3516 12180 3568 12189
rect 5540 12180 5592 12232
rect 6644 12316 6696 12368
rect 6828 12248 6880 12300
rect 2320 12112 2372 12164
rect 4160 12112 4212 12164
rect 5816 12112 5868 12164
rect 6276 12180 6328 12232
rect 6644 12180 6696 12232
rect 7104 12180 7156 12232
rect 7656 12316 7708 12368
rect 8300 12316 8352 12368
rect 7288 12248 7340 12300
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 7748 12248 7800 12300
rect 7656 12223 7708 12232
rect 7656 12189 7665 12223
rect 7665 12189 7699 12223
rect 7699 12189 7708 12223
rect 7656 12180 7708 12189
rect 8944 12180 8996 12232
rect 6736 12112 6788 12164
rect 9772 12384 9824 12436
rect 9864 12384 9916 12436
rect 14648 12427 14700 12436
rect 14648 12393 14657 12427
rect 14657 12393 14691 12427
rect 14691 12393 14700 12427
rect 14648 12384 14700 12393
rect 14832 12384 14884 12436
rect 15752 12384 15804 12436
rect 16488 12384 16540 12436
rect 16672 12427 16724 12436
rect 16672 12393 16681 12427
rect 16681 12393 16715 12427
rect 16715 12393 16724 12427
rect 16672 12384 16724 12393
rect 17684 12384 17736 12436
rect 18420 12427 18472 12436
rect 18420 12393 18429 12427
rect 18429 12393 18463 12427
rect 18463 12393 18472 12427
rect 18420 12384 18472 12393
rect 20352 12427 20404 12436
rect 20352 12393 20361 12427
rect 20361 12393 20395 12427
rect 20395 12393 20404 12427
rect 20352 12384 20404 12393
rect 20720 12384 20772 12436
rect 22008 12384 22060 12436
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 23020 12427 23072 12436
rect 23020 12393 23029 12427
rect 23029 12393 23063 12427
rect 23063 12393 23072 12427
rect 23020 12384 23072 12393
rect 23388 12384 23440 12436
rect 24216 12384 24268 12436
rect 11888 12316 11940 12368
rect 13728 12316 13780 12368
rect 16396 12316 16448 12368
rect 20628 12316 20680 12368
rect 22100 12316 22152 12368
rect 9588 12248 9640 12300
rect 9772 12248 9824 12300
rect 9864 12248 9916 12300
rect 11060 12248 11112 12300
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 17224 12291 17276 12300
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 12164 12180 12216 12232
rect 13176 12180 13228 12232
rect 13636 12223 13688 12232
rect 13636 12189 13645 12223
rect 13645 12189 13679 12223
rect 13679 12189 13688 12223
rect 13636 12180 13688 12189
rect 14096 12112 14148 12164
rect 17224 12257 17233 12291
rect 17233 12257 17267 12291
rect 17267 12257 17276 12291
rect 17224 12248 17276 12257
rect 18972 12248 19024 12300
rect 20076 12248 20128 12300
rect 21732 12248 21784 12300
rect 17408 12180 17460 12232
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 21640 12180 21692 12232
rect 22468 12316 22520 12368
rect 23112 12248 23164 12300
rect 23480 12291 23532 12300
rect 23480 12257 23489 12291
rect 23489 12257 23523 12291
rect 23523 12257 23532 12291
rect 23480 12248 23532 12257
rect 23848 12316 23900 12368
rect 24308 12248 24360 12300
rect 24952 12248 25004 12300
rect 25596 12248 25648 12300
rect 17500 12112 17552 12164
rect 18972 12112 19024 12164
rect 19708 12112 19760 12164
rect 23020 12112 23072 12164
rect 23296 12112 23348 12164
rect 23848 12112 23900 12164
rect 24584 12112 24636 12164
rect 24768 12112 24820 12164
rect 25228 12223 25280 12232
rect 25228 12189 25237 12223
rect 25237 12189 25271 12223
rect 25271 12189 25280 12223
rect 25228 12180 25280 12189
rect 2688 12044 2740 12096
rect 3148 12044 3200 12096
rect 5356 12044 5408 12096
rect 6644 12044 6696 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 12440 12044 12492 12096
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 14280 12044 14332 12096
rect 15660 12044 15712 12096
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 16580 12044 16632 12096
rect 17224 12044 17276 12096
rect 18052 12044 18104 12096
rect 18880 12087 18932 12096
rect 18880 12053 18889 12087
rect 18889 12053 18923 12087
rect 18923 12053 18932 12087
rect 18880 12044 18932 12053
rect 20076 12044 20128 12096
rect 22744 12044 22796 12096
rect 24860 12044 24912 12096
rect 5648 11942 5700 11994
rect 5712 11942 5764 11994
rect 5776 11942 5828 11994
rect 5840 11942 5892 11994
rect 14982 11942 15034 11994
rect 15046 11942 15098 11994
rect 15110 11942 15162 11994
rect 15174 11942 15226 11994
rect 24315 11942 24367 11994
rect 24379 11942 24431 11994
rect 24443 11942 24495 11994
rect 24507 11942 24559 11994
rect 1400 11840 1452 11892
rect 3148 11840 3200 11892
rect 6276 11883 6328 11892
rect 6276 11849 6285 11883
rect 6285 11849 6319 11883
rect 6319 11849 6328 11883
rect 6276 11840 6328 11849
rect 8760 11883 8812 11892
rect 8760 11849 8769 11883
rect 8769 11849 8803 11883
rect 8803 11849 8812 11883
rect 8760 11840 8812 11849
rect 4620 11772 4672 11824
rect 4896 11772 4948 11824
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 10416 11840 10468 11892
rect 13544 11840 13596 11892
rect 12072 11772 12124 11824
rect 14188 11772 14240 11824
rect 16856 11840 16908 11892
rect 20076 11883 20128 11892
rect 20076 11849 20085 11883
rect 20085 11849 20119 11883
rect 20119 11849 20128 11883
rect 20076 11840 20128 11849
rect 21364 11840 21416 11892
rect 21640 11883 21692 11892
rect 21640 11849 21649 11883
rect 21649 11849 21683 11883
rect 21683 11849 21692 11883
rect 21640 11840 21692 11849
rect 23480 11840 23532 11892
rect 25320 11840 25372 11892
rect 26240 11883 26292 11892
rect 26240 11849 26249 11883
rect 26249 11849 26283 11883
rect 26283 11849 26292 11883
rect 26240 11840 26292 11849
rect 19432 11815 19484 11824
rect 19432 11781 19441 11815
rect 19441 11781 19475 11815
rect 19475 11781 19484 11815
rect 19432 11772 19484 11781
rect 19984 11772 20036 11824
rect 24584 11772 24636 11824
rect 17132 11704 17184 11756
rect 17684 11704 17736 11756
rect 2136 11679 2188 11688
rect 2136 11645 2145 11679
rect 2145 11645 2179 11679
rect 2179 11645 2188 11679
rect 2136 11636 2188 11645
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 5632 11636 5684 11688
rect 6552 11636 6604 11688
rect 3976 11568 4028 11620
rect 7196 11568 7248 11620
rect 15568 11636 15620 11688
rect 16764 11636 16816 11688
rect 18052 11679 18104 11688
rect 18052 11645 18061 11679
rect 18061 11645 18095 11679
rect 18095 11645 18104 11679
rect 18052 11636 18104 11645
rect 19708 11636 19760 11688
rect 9588 11568 9640 11620
rect 12532 11568 12584 11620
rect 13636 11568 13688 11620
rect 15660 11568 15712 11620
rect 22468 11704 22520 11756
rect 23020 11747 23072 11756
rect 23020 11713 23029 11747
rect 23029 11713 23063 11747
rect 23063 11713 23072 11747
rect 23020 11704 23072 11713
rect 23112 11704 23164 11756
rect 25136 11704 25188 11756
rect 20628 11679 20680 11688
rect 20628 11645 20637 11679
rect 20637 11645 20671 11679
rect 20671 11645 20680 11679
rect 20628 11636 20680 11645
rect 20720 11636 20772 11688
rect 21548 11636 21600 11688
rect 24952 11636 25004 11688
rect 20812 11568 20864 11620
rect 21456 11611 21508 11620
rect 21456 11577 21465 11611
rect 21465 11577 21499 11611
rect 21499 11577 21508 11611
rect 21456 11568 21508 11577
rect 1768 11543 1820 11552
rect 1768 11509 1777 11543
rect 1777 11509 1811 11543
rect 1811 11509 1820 11543
rect 1768 11500 1820 11509
rect 4620 11500 4672 11552
rect 7656 11500 7708 11552
rect 8576 11500 8628 11552
rect 10876 11500 10928 11552
rect 11060 11500 11112 11552
rect 12072 11500 12124 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 19340 11500 19392 11552
rect 20444 11500 20496 11552
rect 21732 11500 21784 11552
rect 21916 11500 21968 11552
rect 23480 11543 23532 11552
rect 23480 11509 23489 11543
rect 23489 11509 23523 11543
rect 23523 11509 23532 11543
rect 23480 11500 23532 11509
rect 24216 11500 24268 11552
rect 25596 11500 25648 11552
rect 10315 11398 10367 11450
rect 10379 11398 10431 11450
rect 10443 11398 10495 11450
rect 10507 11398 10559 11450
rect 19648 11398 19700 11450
rect 19712 11398 19764 11450
rect 19776 11398 19828 11450
rect 19840 11398 19892 11450
rect 2136 11296 2188 11348
rect 2780 11339 2832 11348
rect 2780 11305 2789 11339
rect 2789 11305 2823 11339
rect 2823 11305 2832 11339
rect 2780 11296 2832 11305
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 3516 11339 3568 11348
rect 2872 11296 2924 11305
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 4436 11296 4488 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 6552 11296 6604 11348
rect 7288 11339 7340 11348
rect 7288 11305 7297 11339
rect 7297 11305 7331 11339
rect 7331 11305 7340 11339
rect 7288 11296 7340 11305
rect 8208 11296 8260 11348
rect 9680 11296 9732 11348
rect 11520 11339 11572 11348
rect 11520 11305 11529 11339
rect 11529 11305 11563 11339
rect 11563 11305 11572 11339
rect 11520 11296 11572 11305
rect 11888 11339 11940 11348
rect 11888 11305 11897 11339
rect 11897 11305 11931 11339
rect 11931 11305 11940 11339
rect 11888 11296 11940 11305
rect 14096 11339 14148 11348
rect 14096 11305 14105 11339
rect 14105 11305 14139 11339
rect 14139 11305 14148 11339
rect 14096 11296 14148 11305
rect 14740 11296 14792 11348
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 17408 11296 17460 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 19432 11296 19484 11348
rect 20076 11296 20128 11348
rect 21088 11296 21140 11348
rect 21548 11296 21600 11348
rect 21916 11339 21968 11348
rect 21916 11305 21925 11339
rect 21925 11305 21959 11339
rect 21959 11305 21968 11339
rect 21916 11296 21968 11305
rect 22376 11296 22428 11348
rect 22928 11339 22980 11348
rect 22928 11305 22937 11339
rect 22937 11305 22971 11339
rect 22971 11305 22980 11339
rect 22928 11296 22980 11305
rect 23020 11296 23072 11348
rect 23296 11296 23348 11348
rect 23940 11296 23992 11348
rect 24124 11296 24176 11348
rect 2504 11228 2556 11280
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 4436 11160 4488 11212
rect 5632 11228 5684 11280
rect 7196 11228 7248 11280
rect 7932 11228 7984 11280
rect 10784 11228 10836 11280
rect 12072 11228 12124 11280
rect 4620 11160 4672 11212
rect 5356 11160 5408 11212
rect 7564 11160 7616 11212
rect 8116 11160 8168 11212
rect 9588 11160 9640 11212
rect 9680 11160 9732 11212
rect 12532 11160 12584 11212
rect 13084 11228 13136 11280
rect 13820 11228 13872 11280
rect 14648 11271 14700 11280
rect 14648 11237 14657 11271
rect 14657 11237 14691 11271
rect 14691 11237 14700 11271
rect 14648 11228 14700 11237
rect 15568 11228 15620 11280
rect 13544 11160 13596 11212
rect 14740 11160 14792 11212
rect 15292 11203 15344 11212
rect 15292 11169 15301 11203
rect 15301 11169 15335 11203
rect 15335 11169 15344 11203
rect 15292 11160 15344 11169
rect 3516 11092 3568 11144
rect 4068 11092 4120 11144
rect 7288 11092 7340 11144
rect 8392 11135 8444 11144
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 1860 11024 1912 11076
rect 2136 11024 2188 11076
rect 6368 11024 6420 11076
rect 7840 11067 7892 11076
rect 7840 11033 7849 11067
rect 7849 11033 7883 11067
rect 7883 11033 7892 11067
rect 7840 11024 7892 11033
rect 3976 10956 4028 11008
rect 5448 10956 5500 11008
rect 6276 10956 6328 11008
rect 7564 10956 7616 11008
rect 8208 10956 8260 11008
rect 9680 10956 9732 11008
rect 10784 11092 10836 11144
rect 11244 11092 11296 11144
rect 12440 11135 12492 11144
rect 12440 11101 12449 11135
rect 12449 11101 12483 11135
rect 12483 11101 12492 11135
rect 12440 11092 12492 11101
rect 16764 11228 16816 11280
rect 16856 11203 16908 11212
rect 16856 11169 16890 11203
rect 16890 11169 16908 11203
rect 16856 11160 16908 11169
rect 10508 11067 10560 11076
rect 10508 11033 10517 11067
rect 10517 11033 10551 11067
rect 10551 11033 10560 11067
rect 10508 11024 10560 11033
rect 13728 11024 13780 11076
rect 11520 10956 11572 11008
rect 13820 10956 13872 11008
rect 14372 10956 14424 11008
rect 19432 11203 19484 11212
rect 19432 11169 19441 11203
rect 19441 11169 19475 11203
rect 19475 11169 19484 11203
rect 19432 11160 19484 11169
rect 20996 11228 21048 11280
rect 22100 11228 22152 11280
rect 24768 11296 24820 11348
rect 25136 11339 25188 11348
rect 25136 11305 25145 11339
rect 25145 11305 25179 11339
rect 25179 11305 25188 11339
rect 25136 11296 25188 11305
rect 25780 11339 25832 11348
rect 25780 11305 25789 11339
rect 25789 11305 25823 11339
rect 25823 11305 25832 11339
rect 25780 11296 25832 11305
rect 22468 11160 22520 11212
rect 22836 11203 22888 11212
rect 22836 11169 22845 11203
rect 22845 11169 22879 11203
rect 22879 11169 22888 11203
rect 22836 11160 22888 11169
rect 25228 11228 25280 11280
rect 25412 11271 25464 11280
rect 25412 11237 25421 11271
rect 25421 11237 25455 11271
rect 25455 11237 25464 11271
rect 25412 11228 25464 11237
rect 25596 11160 25648 11212
rect 25780 11160 25832 11212
rect 18696 11092 18748 11144
rect 20720 11092 20772 11144
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 24124 11092 24176 11144
rect 25320 11092 25372 11144
rect 18880 11067 18932 11076
rect 18880 11033 18889 11067
rect 18889 11033 18923 11067
rect 18923 11033 18932 11067
rect 18880 11024 18932 11033
rect 19156 11024 19208 11076
rect 19984 11024 20036 11076
rect 18420 10956 18472 11008
rect 20260 10956 20312 11008
rect 20812 10956 20864 11008
rect 21640 10956 21692 11008
rect 24216 10956 24268 11008
rect 25320 10956 25372 11008
rect 5648 10854 5700 10906
rect 5712 10854 5764 10906
rect 5776 10854 5828 10906
rect 5840 10854 5892 10906
rect 14982 10854 15034 10906
rect 15046 10854 15098 10906
rect 15110 10854 15162 10906
rect 15174 10854 15226 10906
rect 24315 10854 24367 10906
rect 24379 10854 24431 10906
rect 24443 10854 24495 10906
rect 24507 10854 24559 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 4528 10752 4580 10804
rect 4436 10684 4488 10736
rect 5264 10752 5316 10804
rect 5356 10752 5408 10804
rect 6552 10795 6604 10804
rect 6552 10761 6561 10795
rect 6561 10761 6595 10795
rect 6595 10761 6604 10795
rect 6552 10752 6604 10761
rect 11152 10752 11204 10804
rect 12624 10752 12676 10804
rect 16764 10752 16816 10804
rect 18328 10752 18380 10804
rect 5724 10616 5776 10668
rect 6276 10616 6328 10668
rect 7472 10684 7524 10736
rect 8208 10684 8260 10736
rect 11704 10684 11756 10736
rect 13820 10684 13872 10736
rect 15660 10727 15712 10736
rect 15660 10693 15669 10727
rect 15669 10693 15703 10727
rect 15703 10693 15712 10727
rect 15660 10684 15712 10693
rect 3332 10548 3384 10600
rect 4804 10548 4856 10600
rect 2964 10523 3016 10532
rect 2964 10489 2998 10523
rect 2998 10489 3016 10523
rect 2964 10480 3016 10489
rect 6276 10480 6328 10532
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 11244 10659 11296 10668
rect 11244 10625 11253 10659
rect 11253 10625 11287 10659
rect 11287 10625 11296 10659
rect 11244 10616 11296 10625
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 7932 10548 7984 10600
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 11152 10591 11204 10600
rect 11152 10557 11161 10591
rect 11161 10557 11195 10591
rect 11195 10557 11204 10591
rect 11152 10548 11204 10557
rect 13728 10548 13780 10600
rect 14096 10616 14148 10668
rect 19432 10684 19484 10736
rect 20076 10684 20128 10736
rect 20996 10752 21048 10804
rect 22100 10752 22152 10804
rect 22928 10752 22980 10804
rect 23112 10752 23164 10804
rect 23480 10752 23532 10804
rect 25228 10752 25280 10804
rect 21916 10684 21968 10736
rect 24032 10684 24084 10736
rect 18512 10659 18564 10668
rect 18512 10625 18521 10659
rect 18521 10625 18555 10659
rect 18555 10625 18564 10659
rect 18512 10616 18564 10625
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19524 10659 19576 10668
rect 19524 10625 19533 10659
rect 19533 10625 19567 10659
rect 19567 10625 19576 10659
rect 20260 10659 20312 10668
rect 19524 10616 19576 10625
rect 14556 10591 14608 10600
rect 14556 10557 14579 10591
rect 14579 10557 14608 10591
rect 7840 10480 7892 10532
rect 8116 10480 8168 10532
rect 9036 10480 9088 10532
rect 9312 10480 9364 10532
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 3976 10412 4028 10464
rect 4252 10412 4304 10464
rect 7564 10412 7616 10464
rect 8852 10412 8904 10464
rect 14556 10548 14608 10557
rect 16580 10548 16632 10600
rect 17040 10548 17092 10600
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 21640 10616 21692 10668
rect 23112 10616 23164 10668
rect 23296 10616 23348 10668
rect 21548 10591 21600 10600
rect 21548 10557 21557 10591
rect 21557 10557 21591 10591
rect 21591 10557 21600 10591
rect 21548 10548 21600 10557
rect 23940 10548 23992 10600
rect 15568 10480 15620 10532
rect 16028 10480 16080 10532
rect 17960 10480 18012 10532
rect 20904 10480 20956 10532
rect 21088 10523 21140 10532
rect 21088 10489 21097 10523
rect 21097 10489 21131 10523
rect 21131 10489 21140 10523
rect 21088 10480 21140 10489
rect 21732 10480 21784 10532
rect 22008 10480 22060 10532
rect 24124 10480 24176 10532
rect 11060 10455 11112 10464
rect 11060 10421 11069 10455
rect 11069 10421 11103 10455
rect 11103 10421 11112 10455
rect 11060 10412 11112 10421
rect 13728 10412 13780 10464
rect 16212 10455 16264 10464
rect 16212 10421 16221 10455
rect 16221 10421 16255 10455
rect 16255 10421 16264 10455
rect 16212 10412 16264 10421
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 18236 10412 18288 10464
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 21180 10455 21232 10464
rect 21180 10421 21189 10455
rect 21189 10421 21223 10455
rect 21223 10421 21232 10455
rect 21180 10412 21232 10421
rect 22836 10412 22888 10464
rect 23940 10412 23992 10464
rect 25412 10412 25464 10464
rect 26332 10455 26384 10464
rect 26332 10421 26341 10455
rect 26341 10421 26375 10455
rect 26375 10421 26384 10455
rect 26332 10412 26384 10421
rect 10315 10310 10367 10362
rect 10379 10310 10431 10362
rect 10443 10310 10495 10362
rect 10507 10310 10559 10362
rect 19648 10310 19700 10362
rect 19712 10310 19764 10362
rect 19776 10310 19828 10362
rect 19840 10310 19892 10362
rect 2504 10208 2556 10260
rect 2596 10208 2648 10260
rect 2872 10208 2924 10260
rect 3148 10208 3200 10260
rect 3700 10208 3752 10260
rect 4344 10208 4396 10260
rect 4712 10208 4764 10260
rect 4804 10208 4856 10260
rect 5724 10208 5776 10260
rect 5908 10251 5960 10260
rect 5908 10217 5917 10251
rect 5917 10217 5951 10251
rect 5951 10217 5960 10251
rect 5908 10208 5960 10217
rect 7748 10251 7800 10260
rect 7748 10217 7757 10251
rect 7757 10217 7791 10251
rect 7791 10217 7800 10251
rect 7748 10208 7800 10217
rect 7932 10208 7984 10260
rect 8116 10251 8168 10260
rect 8116 10217 8125 10251
rect 8125 10217 8159 10251
rect 8159 10217 8168 10251
rect 8116 10208 8168 10217
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 9956 10208 10008 10260
rect 10140 10251 10192 10260
rect 10140 10217 10149 10251
rect 10149 10217 10183 10251
rect 10183 10217 10192 10251
rect 10140 10208 10192 10217
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 12532 10208 12584 10260
rect 14556 10208 14608 10260
rect 15200 10208 15252 10260
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 17776 10208 17828 10260
rect 18420 10208 18472 10260
rect 18696 10208 18748 10260
rect 19432 10251 19484 10260
rect 19432 10217 19441 10251
rect 19441 10217 19475 10251
rect 19475 10217 19484 10251
rect 19432 10208 19484 10217
rect 21364 10208 21416 10260
rect 21548 10208 21600 10260
rect 22284 10251 22336 10260
rect 22284 10217 22293 10251
rect 22293 10217 22327 10251
rect 22327 10217 22336 10251
rect 22284 10208 22336 10217
rect 23020 10251 23072 10260
rect 23020 10217 23029 10251
rect 23029 10217 23063 10251
rect 23063 10217 23072 10251
rect 23020 10208 23072 10217
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 23572 10208 23624 10260
rect 24768 10208 24820 10260
rect 25136 10208 25188 10260
rect 25688 10208 25740 10260
rect 26332 10251 26384 10260
rect 26332 10217 26341 10251
rect 26341 10217 26375 10251
rect 26375 10217 26384 10251
rect 26332 10208 26384 10217
rect 3884 10140 3936 10192
rect 6184 10140 6236 10192
rect 3056 10072 3108 10124
rect 6552 10115 6604 10124
rect 6552 10081 6561 10115
rect 6561 10081 6595 10115
rect 6595 10081 6604 10115
rect 6552 10072 6604 10081
rect 7288 10140 7340 10192
rect 7840 10140 7892 10192
rect 9588 10140 9640 10192
rect 10876 10140 10928 10192
rect 9680 10115 9732 10124
rect 2964 10047 3016 10056
rect 2964 10013 2973 10047
rect 2973 10013 3007 10047
rect 3007 10013 3016 10047
rect 2964 10004 3016 10013
rect 2412 9979 2464 9988
rect 2412 9945 2421 9979
rect 2421 9945 2455 9979
rect 2455 9945 2464 9979
rect 2412 9936 2464 9945
rect 4160 10004 4212 10056
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 9680 10081 9689 10115
rect 9689 10081 9723 10115
rect 9723 10081 9732 10115
rect 9680 10072 9732 10081
rect 11244 10115 11296 10124
rect 11244 10081 11253 10115
rect 11253 10081 11287 10115
rect 11287 10081 11296 10115
rect 11244 10072 11296 10081
rect 11888 10115 11940 10124
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9312 10004 9364 10056
rect 11152 10004 11204 10056
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 12532 10072 12584 10124
rect 12808 10115 12860 10124
rect 12808 10081 12817 10115
rect 12817 10081 12851 10115
rect 12851 10081 12860 10115
rect 12808 10072 12860 10081
rect 16212 10140 16264 10192
rect 16856 10140 16908 10192
rect 24032 10183 24084 10192
rect 16304 10115 16356 10124
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 17868 10115 17920 10124
rect 17868 10081 17877 10115
rect 17877 10081 17911 10115
rect 17911 10081 17920 10115
rect 17868 10072 17920 10081
rect 12440 10004 12492 10056
rect 13084 10047 13136 10056
rect 13084 10013 13093 10047
rect 13093 10013 13127 10047
rect 13127 10013 13136 10047
rect 13084 10004 13136 10013
rect 14464 10004 14516 10056
rect 15752 10004 15804 10056
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 17040 10004 17092 10056
rect 5816 9936 5868 9988
rect 8116 9936 8168 9988
rect 11060 9936 11112 9988
rect 24032 10149 24041 10183
rect 24041 10149 24075 10183
rect 24075 10149 24084 10183
rect 24032 10140 24084 10149
rect 20904 10072 20956 10124
rect 22008 10072 22060 10124
rect 22192 10072 22244 10124
rect 22928 10072 22980 10124
rect 23664 10072 23716 10124
rect 23756 10072 23808 10124
rect 24124 10072 24176 10124
rect 24952 10072 25004 10124
rect 19616 10004 19668 10056
rect 20260 10004 20312 10056
rect 21640 10004 21692 10056
rect 22652 10004 22704 10056
rect 20444 9936 20496 9988
rect 21732 9936 21784 9988
rect 23388 9936 23440 9988
rect 25964 9936 26016 9988
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 3056 9868 3108 9920
rect 3608 9868 3660 9920
rect 8392 9868 8444 9920
rect 8852 9868 8904 9920
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 13636 9868 13688 9920
rect 18788 9868 18840 9920
rect 19064 9911 19116 9920
rect 19064 9877 19073 9911
rect 19073 9877 19107 9911
rect 19107 9877 19116 9911
rect 19064 9868 19116 9877
rect 20076 9911 20128 9920
rect 20076 9877 20085 9911
rect 20085 9877 20119 9911
rect 20119 9877 20128 9911
rect 20076 9868 20128 9877
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 21640 9868 21692 9920
rect 22284 9868 22336 9920
rect 22836 9868 22888 9920
rect 5648 9766 5700 9818
rect 5712 9766 5764 9818
rect 5776 9766 5828 9818
rect 5840 9766 5892 9818
rect 14982 9766 15034 9818
rect 15046 9766 15098 9818
rect 15110 9766 15162 9818
rect 15174 9766 15226 9818
rect 24315 9766 24367 9818
rect 24379 9766 24431 9818
rect 24443 9766 24495 9818
rect 24507 9766 24559 9818
rect 6184 9664 6236 9716
rect 6460 9664 6512 9716
rect 6920 9664 6972 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 11152 9664 11204 9716
rect 11244 9664 11296 9716
rect 8024 9596 8076 9648
rect 2228 9528 2280 9580
rect 3056 9528 3108 9580
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 7196 9528 7248 9580
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 7932 9528 7984 9580
rect 8852 9528 8904 9580
rect 2136 9460 2188 9512
rect 1768 9367 1820 9376
rect 1768 9333 1777 9367
rect 1777 9333 1811 9367
rect 1811 9333 1820 9367
rect 1768 9324 1820 9333
rect 3148 9460 3200 9512
rect 8668 9460 8720 9512
rect 2504 9392 2556 9444
rect 2964 9392 3016 9444
rect 4160 9392 4212 9444
rect 3056 9324 3108 9376
rect 4712 9367 4764 9376
rect 4712 9333 4721 9367
rect 4721 9333 4755 9367
rect 4755 9333 4764 9367
rect 4712 9324 4764 9333
rect 5908 9324 5960 9376
rect 7656 9324 7708 9376
rect 8576 9324 8628 9376
rect 9588 9460 9640 9512
rect 12348 9664 12400 9716
rect 12440 9707 12492 9716
rect 12440 9673 12449 9707
rect 12449 9673 12483 9707
rect 12483 9673 12492 9707
rect 12440 9664 12492 9673
rect 13084 9664 13136 9716
rect 15292 9664 15344 9716
rect 15660 9664 15712 9716
rect 16304 9664 16356 9716
rect 15936 9596 15988 9648
rect 18512 9664 18564 9716
rect 18972 9596 19024 9648
rect 19616 9664 19668 9716
rect 20628 9664 20680 9716
rect 20904 9707 20956 9716
rect 20904 9673 20913 9707
rect 20913 9673 20947 9707
rect 20947 9673 20956 9707
rect 20904 9664 20956 9673
rect 22652 9707 22704 9716
rect 22652 9673 22661 9707
rect 22661 9673 22695 9707
rect 22695 9673 22704 9707
rect 22652 9664 22704 9673
rect 22928 9707 22980 9716
rect 22928 9673 22937 9707
rect 22937 9673 22971 9707
rect 22971 9673 22980 9707
rect 22928 9664 22980 9673
rect 23664 9664 23716 9716
rect 24124 9664 24176 9716
rect 19432 9639 19484 9648
rect 19432 9605 19441 9639
rect 19441 9605 19475 9639
rect 19475 9605 19484 9639
rect 19432 9596 19484 9605
rect 19524 9596 19576 9648
rect 12532 9528 12584 9580
rect 12624 9528 12676 9580
rect 13728 9528 13780 9580
rect 16212 9528 16264 9580
rect 16304 9528 16356 9580
rect 16396 9571 16448 9580
rect 16396 9537 16405 9571
rect 16405 9537 16439 9571
rect 16439 9537 16448 9571
rect 16396 9528 16448 9537
rect 18420 9528 18472 9580
rect 19616 9528 19668 9580
rect 19892 9528 19944 9580
rect 20260 9571 20312 9580
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 21272 9596 21324 9648
rect 24676 9596 24728 9648
rect 25596 9596 25648 9648
rect 26332 9639 26384 9648
rect 26332 9605 26341 9639
rect 26341 9605 26375 9639
rect 26375 9605 26384 9639
rect 26332 9596 26384 9605
rect 20628 9528 20680 9580
rect 21640 9571 21692 9580
rect 21640 9537 21649 9571
rect 21649 9537 21683 9571
rect 21683 9537 21692 9571
rect 21640 9528 21692 9537
rect 22192 9571 22244 9580
rect 9404 9392 9456 9444
rect 9588 9324 9640 9376
rect 11520 9324 11572 9376
rect 11612 9324 11664 9376
rect 15384 9460 15436 9512
rect 20076 9460 20128 9512
rect 21180 9460 21232 9512
rect 22192 9537 22201 9571
rect 22201 9537 22235 9571
rect 22235 9537 22244 9571
rect 22192 9528 22244 9537
rect 21916 9460 21968 9512
rect 23388 9460 23440 9512
rect 24860 9460 24912 9512
rect 12808 9367 12860 9376
rect 12808 9333 12817 9367
rect 12817 9333 12851 9367
rect 12851 9333 12860 9367
rect 12808 9324 12860 9333
rect 13268 9324 13320 9376
rect 16488 9392 16540 9444
rect 19432 9392 19484 9444
rect 15660 9367 15712 9376
rect 15660 9333 15669 9367
rect 15669 9333 15703 9367
rect 15703 9333 15712 9367
rect 15660 9324 15712 9333
rect 15844 9324 15896 9376
rect 17408 9367 17460 9376
rect 17408 9333 17417 9367
rect 17417 9333 17451 9367
rect 17451 9333 17460 9367
rect 18420 9367 18472 9376
rect 17408 9324 17460 9333
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 19064 9324 19116 9376
rect 19984 9324 20036 9376
rect 23296 9367 23348 9376
rect 23296 9333 23305 9367
rect 23305 9333 23339 9367
rect 23339 9333 23348 9367
rect 23296 9324 23348 9333
rect 10315 9222 10367 9274
rect 10379 9222 10431 9274
rect 10443 9222 10495 9274
rect 10507 9222 10559 9274
rect 19648 9222 19700 9274
rect 19712 9222 19764 9274
rect 19776 9222 19828 9274
rect 19840 9222 19892 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 2688 9120 2740 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 4620 9163 4672 9172
rect 4620 9129 4629 9163
rect 4629 9129 4663 9163
rect 4663 9129 4672 9163
rect 4620 9120 4672 9129
rect 5080 9120 5132 9172
rect 8116 9120 8168 9172
rect 9312 9120 9364 9172
rect 10784 9120 10836 9172
rect 13176 9120 13228 9172
rect 14004 9120 14056 9172
rect 15292 9120 15344 9172
rect 20720 9163 20772 9172
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 21180 9120 21232 9172
rect 21364 9163 21416 9172
rect 21364 9129 21373 9163
rect 21373 9129 21407 9163
rect 21407 9129 21416 9163
rect 21364 9120 21416 9129
rect 21916 9163 21968 9172
rect 21916 9129 21925 9163
rect 21925 9129 21959 9163
rect 21959 9129 21968 9163
rect 21916 9120 21968 9129
rect 22652 9120 22704 9172
rect 24400 9163 24452 9172
rect 24400 9129 24409 9163
rect 24409 9129 24443 9163
rect 24443 9129 24452 9163
rect 24400 9120 24452 9129
rect 24768 9163 24820 9172
rect 24768 9129 24777 9163
rect 24777 9129 24811 9163
rect 24811 9129 24820 9163
rect 24768 9120 24820 9129
rect 25872 9163 25924 9172
rect 25872 9129 25881 9163
rect 25881 9129 25915 9163
rect 25915 9129 25924 9163
rect 25872 9120 25924 9129
rect 2596 9052 2648 9104
rect 4804 9052 4856 9104
rect 5264 9095 5316 9104
rect 5264 9061 5273 9095
rect 5273 9061 5307 9095
rect 5307 9061 5316 9095
rect 5264 9052 5316 9061
rect 8300 9052 8352 9104
rect 10232 9052 10284 9104
rect 2504 8984 2556 9036
rect 4252 8984 4304 9036
rect 6552 8984 6604 9036
rect 6736 9027 6788 9036
rect 6736 8993 6770 9027
rect 6770 8993 6788 9027
rect 6736 8984 6788 8993
rect 10140 8984 10192 9036
rect 13544 9095 13596 9104
rect 13544 9061 13553 9095
rect 13553 9061 13587 9095
rect 13587 9061 13596 9095
rect 13544 9052 13596 9061
rect 13820 9052 13872 9104
rect 15476 9052 15528 9104
rect 11244 8984 11296 9036
rect 14648 8984 14700 9036
rect 17960 9052 18012 9104
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 20076 8984 20128 9036
rect 20812 9052 20864 9104
rect 21548 9052 21600 9104
rect 22008 8984 22060 9036
rect 23020 8984 23072 9036
rect 23848 9052 23900 9104
rect 2044 8916 2096 8968
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3516 8916 3568 8968
rect 9680 8959 9732 8968
rect 1676 8848 1728 8900
rect 5908 8848 5960 8900
rect 9680 8925 9689 8959
rect 9689 8925 9723 8959
rect 9723 8925 9732 8959
rect 9680 8916 9732 8925
rect 12440 8916 12492 8968
rect 12808 8916 12860 8968
rect 13728 8959 13780 8968
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 1768 8780 1820 8832
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 5264 8780 5316 8832
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 12348 8848 12400 8900
rect 7748 8780 7800 8832
rect 10876 8780 10928 8832
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 13728 8780 13780 8832
rect 17776 8916 17828 8968
rect 18328 8959 18380 8968
rect 18328 8925 18337 8959
rect 18337 8925 18371 8959
rect 18371 8925 18380 8959
rect 18328 8916 18380 8925
rect 20260 8959 20312 8968
rect 20260 8925 20269 8959
rect 20269 8925 20303 8959
rect 20303 8925 20312 8959
rect 20260 8916 20312 8925
rect 22928 8959 22980 8968
rect 19248 8848 19300 8900
rect 22928 8925 22937 8959
rect 22937 8925 22971 8959
rect 22971 8925 22980 8959
rect 22928 8916 22980 8925
rect 21548 8848 21600 8900
rect 23388 8848 23440 8900
rect 24124 8984 24176 9036
rect 24860 8984 24912 9036
rect 25964 8916 26016 8968
rect 26148 8916 26200 8968
rect 15568 8780 15620 8832
rect 16764 8780 16816 8832
rect 17868 8780 17920 8832
rect 19064 8823 19116 8832
rect 19064 8789 19073 8823
rect 19073 8789 19107 8823
rect 19107 8789 19116 8823
rect 19064 8780 19116 8789
rect 19892 8823 19944 8832
rect 19892 8789 19901 8823
rect 19901 8789 19935 8823
rect 19935 8789 19944 8823
rect 19892 8780 19944 8789
rect 22192 8780 22244 8832
rect 25596 8823 25648 8832
rect 25596 8789 25605 8823
rect 25605 8789 25639 8823
rect 25639 8789 25648 8823
rect 25596 8780 25648 8789
rect 26148 8780 26200 8832
rect 5648 8678 5700 8730
rect 5712 8678 5764 8730
rect 5776 8678 5828 8730
rect 5840 8678 5892 8730
rect 14982 8678 15034 8730
rect 15046 8678 15098 8730
rect 15110 8678 15162 8730
rect 15174 8678 15226 8730
rect 24315 8678 24367 8730
rect 24379 8678 24431 8730
rect 24443 8678 24495 8730
rect 24507 8678 24559 8730
rect 1492 8576 1544 8628
rect 3240 8576 3292 8628
rect 3424 8576 3476 8628
rect 4160 8576 4212 8628
rect 7196 8619 7248 8628
rect 572 8508 624 8560
rect 2596 8508 2648 8560
rect 4528 8508 4580 8560
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2044 8372 2096 8424
rect 7196 8585 7205 8619
rect 7205 8585 7239 8619
rect 7239 8585 7248 8619
rect 7196 8576 7248 8585
rect 9312 8576 9364 8628
rect 9956 8576 10008 8628
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 11520 8576 11572 8628
rect 12624 8576 12676 8628
rect 13176 8576 13228 8628
rect 13544 8576 13596 8628
rect 14464 8576 14516 8628
rect 15292 8576 15344 8628
rect 15752 8619 15804 8628
rect 15752 8585 15761 8619
rect 15761 8585 15795 8619
rect 15795 8585 15804 8619
rect 15752 8576 15804 8585
rect 15844 8576 15896 8628
rect 16396 8576 16448 8628
rect 20076 8619 20128 8628
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 20260 8576 20312 8628
rect 21548 8619 21600 8628
rect 21548 8585 21557 8619
rect 21557 8585 21591 8619
rect 21591 8585 21600 8619
rect 21548 8576 21600 8585
rect 24124 8576 24176 8628
rect 25504 8619 25556 8628
rect 25504 8585 25513 8619
rect 25513 8585 25547 8619
rect 25547 8585 25556 8619
rect 25504 8576 25556 8585
rect 26056 8576 26108 8628
rect 26332 8619 26384 8628
rect 26332 8585 26341 8619
rect 26341 8585 26375 8619
rect 26375 8585 26384 8619
rect 26332 8576 26384 8585
rect 4712 8440 4764 8492
rect 3148 8304 3200 8356
rect 4896 8415 4948 8424
rect 4896 8381 4905 8415
rect 4905 8381 4939 8415
rect 4939 8381 4948 8415
rect 4896 8372 4948 8381
rect 5356 8372 5408 8424
rect 6552 8440 6604 8492
rect 7656 8483 7708 8492
rect 7656 8449 7665 8483
rect 7665 8449 7699 8483
rect 7699 8449 7708 8483
rect 7656 8440 7708 8449
rect 9772 8440 9824 8492
rect 9956 8440 10008 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 15568 8508 15620 8560
rect 19340 8508 19392 8560
rect 20720 8440 20772 8492
rect 22652 8508 22704 8560
rect 24860 8551 24912 8560
rect 24860 8517 24869 8551
rect 24869 8517 24903 8551
rect 24903 8517 24912 8551
rect 24860 8508 24912 8517
rect 23572 8440 23624 8492
rect 10968 8372 11020 8424
rect 16120 8415 16172 8424
rect 4252 8304 4304 8356
rect 5448 8304 5500 8356
rect 6736 8304 6788 8356
rect 7748 8304 7800 8356
rect 9772 8304 9824 8356
rect 13728 8304 13780 8356
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 19984 8372 20036 8424
rect 23020 8415 23072 8424
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 6276 8236 6328 8288
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 10784 8236 10836 8288
rect 11152 8236 11204 8288
rect 13452 8236 13504 8288
rect 13636 8236 13688 8288
rect 15568 8347 15620 8356
rect 15568 8313 15577 8347
rect 15577 8313 15611 8347
rect 15611 8313 15620 8347
rect 15568 8304 15620 8313
rect 16672 8304 16724 8356
rect 18328 8347 18380 8356
rect 18328 8313 18362 8347
rect 18362 8313 18380 8347
rect 18328 8304 18380 8313
rect 21732 8304 21784 8356
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 23664 8415 23716 8424
rect 23664 8381 23673 8415
rect 23673 8381 23707 8415
rect 23707 8381 23716 8415
rect 23664 8372 23716 8381
rect 18604 8236 18656 8288
rect 19156 8236 19208 8288
rect 20720 8236 20772 8288
rect 21824 8236 21876 8288
rect 23204 8304 23256 8356
rect 23480 8304 23532 8356
rect 23848 8279 23900 8288
rect 23848 8245 23857 8279
rect 23857 8245 23891 8279
rect 23891 8245 23900 8279
rect 23848 8236 23900 8245
rect 10315 8134 10367 8186
rect 10379 8134 10431 8186
rect 10443 8134 10495 8186
rect 10507 8134 10559 8186
rect 19648 8134 19700 8186
rect 19712 8134 19764 8186
rect 19776 8134 19828 8186
rect 19840 8134 19892 8186
rect 1952 8032 2004 8084
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 3240 8032 3292 8084
rect 3792 8032 3844 8084
rect 4896 8032 4948 8084
rect 7196 8032 7248 8084
rect 7564 8032 7616 8084
rect 9588 8032 9640 8084
rect 9772 8075 9824 8084
rect 9772 8041 9781 8075
rect 9781 8041 9815 8075
rect 9815 8041 9824 8075
rect 9772 8032 9824 8041
rect 9956 8032 10008 8084
rect 10692 8032 10744 8084
rect 11060 8032 11112 8084
rect 12348 8032 12400 8084
rect 13452 8032 13504 8084
rect 13912 8032 13964 8084
rect 15108 8075 15160 8084
rect 15108 8041 15117 8075
rect 15117 8041 15151 8075
rect 15151 8041 15160 8075
rect 15108 8032 15160 8041
rect 15568 8032 15620 8084
rect 16212 8032 16264 8084
rect 16672 8075 16724 8084
rect 16672 8041 16681 8075
rect 16681 8041 16715 8075
rect 16715 8041 16724 8075
rect 16672 8032 16724 8041
rect 17776 8075 17828 8084
rect 17776 8041 17785 8075
rect 17785 8041 17819 8075
rect 17819 8041 17828 8075
rect 17776 8032 17828 8041
rect 18144 8032 18196 8084
rect 19432 8032 19484 8084
rect 22560 8032 22612 8084
rect 2964 7964 3016 8016
rect 3516 7964 3568 8016
rect 6368 7964 6420 8016
rect 7748 8007 7800 8016
rect 7748 7973 7757 8007
rect 7757 7973 7791 8007
rect 7791 7973 7800 8007
rect 7748 7964 7800 7973
rect 4068 7939 4120 7948
rect 4068 7905 4077 7939
rect 4077 7905 4111 7939
rect 4111 7905 4120 7939
rect 4068 7896 4120 7905
rect 4712 7896 4764 7948
rect 5356 7896 5408 7948
rect 8668 7896 8720 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2596 7760 2648 7812
rect 3976 7828 4028 7880
rect 7472 7828 7524 7880
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 9680 7964 9732 8016
rect 11152 7964 11204 8016
rect 12072 7964 12124 8016
rect 11244 7896 11296 7948
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 15660 7964 15712 8016
rect 18696 7964 18748 8016
rect 18972 7964 19024 8016
rect 16120 7896 16172 7948
rect 8576 7828 8628 7837
rect 8116 7760 8168 7812
rect 8392 7760 8444 7812
rect 9588 7760 9640 7812
rect 14188 7760 14240 7812
rect 14372 7760 14424 7812
rect 17684 7896 17736 7948
rect 18604 7896 18656 7948
rect 20352 7964 20404 8016
rect 19524 7896 19576 7948
rect 19892 7939 19944 7948
rect 19892 7905 19901 7939
rect 19901 7905 19935 7939
rect 19935 7905 19944 7939
rect 19892 7896 19944 7905
rect 19984 7896 20036 7948
rect 20444 7896 20496 7948
rect 20720 7828 20772 7880
rect 18696 7760 18748 7812
rect 20076 7760 20128 7812
rect 22468 7964 22520 8016
rect 21180 7896 21232 7948
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 22744 7896 22796 7948
rect 23296 7896 23348 7948
rect 24768 7896 24820 7948
rect 25044 7896 25096 7948
rect 21088 7828 21140 7880
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 21548 7871 21600 7880
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 23020 7871 23072 7880
rect 21548 7828 21600 7837
rect 23020 7837 23029 7871
rect 23029 7837 23063 7871
rect 23063 7837 23072 7871
rect 23020 7828 23072 7837
rect 22836 7760 22888 7812
rect 23480 7828 23532 7880
rect 25504 7760 25556 7812
rect 1492 7692 1544 7744
rect 3516 7692 3568 7744
rect 6276 7692 6328 7744
rect 8208 7692 8260 7744
rect 11704 7692 11756 7744
rect 13452 7692 13504 7744
rect 13820 7692 13872 7744
rect 16212 7692 16264 7744
rect 20444 7692 20496 7744
rect 20720 7735 20772 7744
rect 20720 7701 20729 7735
rect 20729 7701 20763 7735
rect 20763 7701 20772 7735
rect 20720 7692 20772 7701
rect 21548 7692 21600 7744
rect 21732 7692 21784 7744
rect 23204 7692 23256 7744
rect 23296 7692 23348 7744
rect 24032 7692 24084 7744
rect 24952 7735 25004 7744
rect 24952 7701 24961 7735
rect 24961 7701 24995 7735
rect 24995 7701 25004 7735
rect 24952 7692 25004 7701
rect 25320 7735 25372 7744
rect 25320 7701 25329 7735
rect 25329 7701 25363 7735
rect 25363 7701 25372 7735
rect 25320 7692 25372 7701
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 26056 7735 26108 7744
rect 26056 7701 26065 7735
rect 26065 7701 26099 7735
rect 26099 7701 26108 7735
rect 26056 7692 26108 7701
rect 5648 7590 5700 7642
rect 5712 7590 5764 7642
rect 5776 7590 5828 7642
rect 5840 7590 5892 7642
rect 14982 7590 15034 7642
rect 15046 7590 15098 7642
rect 15110 7590 15162 7642
rect 15174 7590 15226 7642
rect 24315 7590 24367 7642
rect 24379 7590 24431 7642
rect 24443 7590 24495 7642
rect 24507 7590 24559 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 5172 7488 5224 7540
rect 6368 7488 6420 7540
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 8668 7531 8720 7540
rect 8668 7497 8677 7531
rect 8677 7497 8711 7531
rect 8711 7497 8720 7531
rect 8668 7488 8720 7497
rect 10692 7488 10744 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 13544 7488 13596 7540
rect 15660 7488 15712 7540
rect 15844 7531 15896 7540
rect 15844 7497 15853 7531
rect 15853 7497 15887 7531
rect 15887 7497 15896 7531
rect 15844 7488 15896 7497
rect 17684 7488 17736 7540
rect 18144 7531 18196 7540
rect 18144 7497 18153 7531
rect 18153 7497 18187 7531
rect 18187 7497 18196 7531
rect 18144 7488 18196 7497
rect 19524 7488 19576 7540
rect 20628 7488 20680 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 22560 7488 22612 7540
rect 23020 7488 23072 7540
rect 24768 7488 24820 7540
rect 25044 7488 25096 7540
rect 25780 7531 25832 7540
rect 25780 7497 25789 7531
rect 25789 7497 25823 7531
rect 25823 7497 25832 7531
rect 25780 7488 25832 7497
rect 25872 7488 25924 7540
rect 2412 7420 2464 7472
rect 8576 7420 8628 7472
rect 10784 7420 10836 7472
rect 16304 7420 16356 7472
rect 20812 7420 20864 7472
rect 24216 7463 24268 7472
rect 2320 7352 2372 7404
rect 3240 7352 3292 7404
rect 4620 7352 4672 7404
rect 4712 7352 4764 7404
rect 8024 7352 8076 7404
rect 10140 7352 10192 7404
rect 11704 7352 11756 7404
rect 14372 7352 14424 7404
rect 14832 7352 14884 7404
rect 18696 7395 18748 7404
rect 3608 7327 3660 7336
rect 3608 7293 3617 7327
rect 3617 7293 3651 7327
rect 3651 7293 3660 7327
rect 3608 7284 3660 7293
rect 5172 7284 5224 7336
rect 2412 7216 2464 7268
rect 3424 7216 3476 7268
rect 4988 7216 5040 7268
rect 2596 7191 2648 7200
rect 2596 7157 2605 7191
rect 2605 7157 2639 7191
rect 2639 7157 2648 7191
rect 2596 7148 2648 7157
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 5448 7216 5500 7268
rect 8852 7284 8904 7336
rect 9588 7284 9640 7336
rect 10784 7284 10836 7336
rect 11152 7327 11204 7336
rect 11152 7293 11161 7327
rect 11161 7293 11195 7327
rect 11195 7293 11204 7327
rect 11152 7284 11204 7293
rect 13452 7284 13504 7336
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 19892 7352 19944 7404
rect 18236 7284 18288 7336
rect 19064 7284 19116 7336
rect 20076 7327 20128 7336
rect 20076 7293 20085 7327
rect 20085 7293 20119 7327
rect 20119 7293 20128 7327
rect 20076 7284 20128 7293
rect 21916 7284 21968 7336
rect 24216 7429 24225 7463
rect 24225 7429 24259 7463
rect 24259 7429 24268 7463
rect 24216 7420 24268 7429
rect 23848 7284 23900 7336
rect 24768 7327 24820 7336
rect 24768 7293 24777 7327
rect 24777 7293 24811 7327
rect 24811 7293 24820 7327
rect 24768 7284 24820 7293
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 9404 7216 9456 7268
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 14832 7148 14884 7200
rect 16212 7191 16264 7200
rect 16212 7157 16221 7191
rect 16221 7157 16255 7191
rect 16255 7157 16264 7191
rect 16212 7148 16264 7157
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 18236 7148 18288 7200
rect 18880 7216 18932 7268
rect 19248 7216 19300 7268
rect 19984 7216 20036 7268
rect 18696 7148 18748 7200
rect 19156 7148 19208 7200
rect 21272 7148 21324 7200
rect 21732 7191 21784 7200
rect 21732 7157 21741 7191
rect 21741 7157 21775 7191
rect 21775 7157 21784 7191
rect 21732 7148 21784 7157
rect 22100 7148 22152 7200
rect 22744 7148 22796 7200
rect 24124 7148 24176 7200
rect 25964 7148 26016 7200
rect 10315 7046 10367 7098
rect 10379 7046 10431 7098
rect 10443 7046 10495 7098
rect 10507 7046 10559 7098
rect 19648 7046 19700 7098
rect 19712 7046 19764 7098
rect 19776 7046 19828 7098
rect 19840 7046 19892 7098
rect 2412 6987 2464 6996
rect 2412 6953 2421 6987
rect 2421 6953 2455 6987
rect 2455 6953 2464 6987
rect 2412 6944 2464 6953
rect 3148 6944 3200 6996
rect 4712 6944 4764 6996
rect 6828 6944 6880 6996
rect 8576 6944 8628 6996
rect 9956 6987 10008 6996
rect 9956 6953 9965 6987
rect 9965 6953 9999 6987
rect 9999 6953 10008 6987
rect 9956 6944 10008 6953
rect 12072 6944 12124 6996
rect 13820 6944 13872 6996
rect 15108 6944 15160 6996
rect 15660 6944 15712 6996
rect 18604 6987 18656 6996
rect 2320 6876 2372 6928
rect 8392 6919 8444 6928
rect 8392 6885 8401 6919
rect 8401 6885 8435 6919
rect 8435 6885 8444 6919
rect 8392 6876 8444 6885
rect 10784 6876 10836 6928
rect 4068 6808 4120 6860
rect 4528 6851 4580 6860
rect 4528 6817 4537 6851
rect 4537 6817 4571 6851
rect 4571 6817 4580 6851
rect 4528 6808 4580 6817
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 7288 6808 7340 6860
rect 8024 6808 8076 6860
rect 11152 6808 11204 6860
rect 12256 6808 12308 6860
rect 14740 6808 14792 6860
rect 16304 6876 16356 6928
rect 15200 6808 15252 6860
rect 18604 6953 18613 6987
rect 18613 6953 18647 6987
rect 18647 6953 18656 6987
rect 18604 6944 18656 6953
rect 19432 6944 19484 6996
rect 20996 6944 21048 6996
rect 21824 6944 21876 6996
rect 22376 6944 22428 6996
rect 18972 6876 19024 6928
rect 22284 6876 22336 6928
rect 22468 6876 22520 6928
rect 22560 6876 22612 6928
rect 23020 6876 23072 6928
rect 23756 6944 23808 6996
rect 24032 6944 24084 6996
rect 24768 6987 24820 6996
rect 24768 6953 24777 6987
rect 24777 6953 24811 6987
rect 24811 6953 24820 6987
rect 24768 6944 24820 6953
rect 16764 6808 16816 6860
rect 2964 6783 3016 6792
rect 2964 6749 2973 6783
rect 2973 6749 3007 6783
rect 3007 6749 3016 6783
rect 2964 6740 3016 6749
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 6000 6740 6052 6792
rect 3148 6672 3200 6724
rect 5632 6672 5684 6724
rect 6092 6715 6144 6724
rect 6092 6681 6101 6715
rect 6101 6681 6135 6715
rect 6135 6681 6144 6715
rect 6092 6672 6144 6681
rect 6368 6672 6420 6724
rect 8300 6740 8352 6792
rect 8668 6783 8720 6792
rect 8668 6749 8677 6783
rect 8677 6749 8711 6783
rect 8711 6749 8720 6783
rect 8668 6740 8720 6749
rect 9956 6740 10008 6792
rect 13268 6783 13320 6792
rect 13268 6749 13277 6783
rect 13277 6749 13311 6783
rect 13311 6749 13320 6783
rect 13268 6740 13320 6749
rect 8208 6672 8260 6724
rect 12808 6715 12860 6724
rect 12808 6681 12817 6715
rect 12817 6681 12851 6715
rect 12851 6681 12860 6715
rect 12808 6672 12860 6681
rect 2320 6647 2372 6656
rect 2320 6613 2329 6647
rect 2329 6613 2363 6647
rect 2363 6613 2372 6647
rect 2320 6604 2372 6613
rect 2504 6604 2556 6656
rect 4068 6647 4120 6656
rect 4068 6613 4077 6647
rect 4077 6613 4111 6647
rect 4111 6613 4120 6647
rect 4068 6604 4120 6613
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 8024 6647 8076 6656
rect 8024 6613 8033 6647
rect 8033 6613 8067 6647
rect 8067 6613 8076 6647
rect 8024 6604 8076 6613
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 14096 6740 14148 6792
rect 14924 6740 14976 6792
rect 17960 6740 18012 6792
rect 15016 6672 15068 6724
rect 20812 6808 20864 6860
rect 21824 6808 21876 6860
rect 23388 6808 23440 6860
rect 23664 6851 23716 6860
rect 23664 6817 23673 6851
rect 23673 6817 23707 6851
rect 23707 6817 23716 6851
rect 23664 6808 23716 6817
rect 24032 6851 24084 6860
rect 24032 6817 24041 6851
rect 24041 6817 24075 6851
rect 24075 6817 24084 6851
rect 24032 6808 24084 6817
rect 19616 6740 19668 6792
rect 20352 6672 20404 6724
rect 21364 6672 21416 6724
rect 21916 6740 21968 6792
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 25780 6740 25832 6792
rect 22100 6672 22152 6724
rect 23296 6672 23348 6724
rect 23388 6672 23440 6724
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16120 6647 16172 6656
rect 16120 6613 16129 6647
rect 16129 6613 16163 6647
rect 16163 6613 16172 6647
rect 16120 6604 16172 6613
rect 16672 6604 16724 6656
rect 17040 6604 17092 6656
rect 19156 6647 19208 6656
rect 19156 6613 19165 6647
rect 19165 6613 19199 6647
rect 19199 6613 19208 6647
rect 19156 6604 19208 6613
rect 19524 6604 19576 6656
rect 19984 6604 20036 6656
rect 20720 6647 20772 6656
rect 20720 6613 20729 6647
rect 20729 6613 20763 6647
rect 20763 6613 20772 6647
rect 20720 6604 20772 6613
rect 21180 6604 21232 6656
rect 22008 6647 22060 6656
rect 22008 6613 22017 6647
rect 22017 6613 22051 6647
rect 22051 6613 22060 6647
rect 22008 6604 22060 6613
rect 23572 6604 23624 6656
rect 24860 6604 24912 6656
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 26056 6647 26108 6656
rect 26056 6613 26065 6647
rect 26065 6613 26099 6647
rect 26099 6613 26108 6647
rect 26056 6604 26108 6613
rect 5648 6502 5700 6554
rect 5712 6502 5764 6554
rect 5776 6502 5828 6554
rect 5840 6502 5892 6554
rect 14982 6502 15034 6554
rect 15046 6502 15098 6554
rect 15110 6502 15162 6554
rect 15174 6502 15226 6554
rect 24315 6502 24367 6554
rect 24379 6502 24431 6554
rect 24443 6502 24495 6554
rect 24507 6502 24559 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 3240 6443 3292 6452
rect 3240 6409 3249 6443
rect 3249 6409 3283 6443
rect 3283 6409 3292 6443
rect 3240 6400 3292 6409
rect 6000 6400 6052 6452
rect 6828 6400 6880 6452
rect 7288 6443 7340 6452
rect 7288 6409 7297 6443
rect 7297 6409 7331 6443
rect 7331 6409 7340 6443
rect 7288 6400 7340 6409
rect 10416 6443 10468 6452
rect 10416 6409 10425 6443
rect 10425 6409 10459 6443
rect 10459 6409 10468 6443
rect 10416 6400 10468 6409
rect 11888 6400 11940 6452
rect 12532 6400 12584 6452
rect 15476 6400 15528 6452
rect 16488 6400 16540 6452
rect 19248 6400 19300 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 21180 6443 21232 6452
rect 21180 6409 21189 6443
rect 21189 6409 21223 6443
rect 21223 6409 21232 6443
rect 21180 6400 21232 6409
rect 2596 6332 2648 6384
rect 2964 6332 3016 6384
rect 5908 6332 5960 6384
rect 6368 6332 6420 6384
rect 10876 6332 10928 6384
rect 2320 6264 2372 6316
rect 14556 6332 14608 6384
rect 19708 6332 19760 6384
rect 20260 6332 20312 6384
rect 20628 6332 20680 6384
rect 23388 6400 23440 6452
rect 24032 6400 24084 6452
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 25780 6443 25832 6452
rect 25780 6409 25789 6443
rect 25789 6409 25823 6443
rect 25823 6409 25832 6443
rect 25780 6400 25832 6409
rect 21548 6332 21600 6384
rect 22376 6332 22428 6384
rect 23296 6332 23348 6384
rect 23848 6332 23900 6384
rect 23940 6332 23992 6384
rect 24308 6332 24360 6384
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 18328 6264 18380 6316
rect 18880 6264 18932 6316
rect 2044 6196 2096 6248
rect 2596 6239 2648 6248
rect 2596 6205 2605 6239
rect 2605 6205 2639 6239
rect 2639 6205 2648 6239
rect 2596 6196 2648 6205
rect 3424 6128 3476 6180
rect 4344 6196 4396 6248
rect 8944 6196 8996 6248
rect 10416 6196 10468 6248
rect 5448 6128 5500 6180
rect 8208 6128 8260 6180
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3332 6060 3384 6112
rect 5172 6103 5224 6112
rect 5172 6069 5181 6103
rect 5181 6069 5215 6103
rect 5215 6069 5224 6103
rect 5172 6060 5224 6069
rect 5264 6060 5316 6112
rect 8760 6060 8812 6112
rect 9772 6060 9824 6112
rect 10784 6060 10836 6112
rect 11888 6060 11940 6112
rect 12532 6060 12584 6112
rect 14096 6196 14148 6248
rect 16856 6239 16908 6248
rect 16856 6205 16865 6239
rect 16865 6205 16899 6239
rect 16899 6205 16908 6239
rect 16856 6196 16908 6205
rect 19156 6196 19208 6248
rect 16488 6128 16540 6180
rect 17132 6128 17184 6180
rect 17316 6128 17368 6180
rect 19984 6264 20036 6316
rect 20076 6264 20128 6316
rect 21180 6264 21232 6316
rect 21364 6264 21416 6316
rect 23664 6264 23716 6316
rect 24124 6264 24176 6316
rect 19340 6196 19392 6248
rect 20720 6196 20772 6248
rect 21548 6239 21600 6248
rect 21548 6205 21557 6239
rect 21557 6205 21591 6239
rect 21591 6205 21600 6239
rect 21548 6196 21600 6205
rect 21640 6196 21692 6248
rect 21824 6196 21876 6248
rect 21916 6196 21968 6248
rect 20260 6128 20312 6180
rect 22376 6128 22428 6180
rect 23112 6196 23164 6248
rect 24676 6196 24728 6248
rect 25136 6196 25188 6248
rect 22744 6128 22796 6180
rect 23848 6128 23900 6180
rect 24308 6128 24360 6180
rect 13728 6060 13780 6112
rect 14464 6060 14516 6112
rect 14648 6060 14700 6112
rect 15384 6103 15436 6112
rect 15384 6069 15393 6103
rect 15393 6069 15427 6103
rect 15427 6069 15436 6103
rect 15384 6060 15436 6069
rect 16948 6060 17000 6112
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 19524 6060 19576 6112
rect 19984 6103 20036 6112
rect 19984 6069 19993 6103
rect 19993 6069 20027 6103
rect 20027 6069 20036 6103
rect 19984 6060 20036 6069
rect 21640 6103 21692 6112
rect 21640 6069 21649 6103
rect 21649 6069 21683 6103
rect 21683 6069 21692 6103
rect 23664 6103 23716 6112
rect 21640 6060 21692 6069
rect 23664 6069 23673 6103
rect 23673 6069 23707 6103
rect 23707 6069 23716 6103
rect 23664 6060 23716 6069
rect 25412 6103 25464 6112
rect 25412 6069 25421 6103
rect 25421 6069 25455 6103
rect 25455 6069 25464 6103
rect 25412 6060 25464 6069
rect 26240 6103 26292 6112
rect 26240 6069 26249 6103
rect 26249 6069 26283 6103
rect 26283 6069 26292 6103
rect 26240 6060 26292 6069
rect 10315 5958 10367 6010
rect 10379 5958 10431 6010
rect 10443 5958 10495 6010
rect 10507 5958 10559 6010
rect 19648 5958 19700 6010
rect 19712 5958 19764 6010
rect 19776 5958 19828 6010
rect 19840 5958 19892 6010
rect 1768 5856 1820 5908
rect 2780 5899 2832 5908
rect 2320 5763 2372 5772
rect 2320 5729 2329 5763
rect 2329 5729 2363 5763
rect 2363 5729 2372 5763
rect 2320 5720 2372 5729
rect 2136 5516 2188 5568
rect 2780 5865 2789 5899
rect 2789 5865 2823 5899
rect 2823 5865 2832 5899
rect 2780 5856 2832 5865
rect 4344 5856 4396 5908
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 5264 5899 5316 5908
rect 5264 5865 5273 5899
rect 5273 5865 5307 5899
rect 5307 5865 5316 5899
rect 6276 5899 6328 5908
rect 5264 5856 5316 5865
rect 6276 5865 6285 5899
rect 6285 5865 6319 5899
rect 6319 5865 6328 5899
rect 6276 5856 6328 5865
rect 6736 5899 6788 5908
rect 6736 5865 6745 5899
rect 6745 5865 6779 5899
rect 6779 5865 6788 5899
rect 6736 5856 6788 5865
rect 8208 5899 8260 5908
rect 8208 5865 8217 5899
rect 8217 5865 8251 5899
rect 8251 5865 8260 5899
rect 8208 5856 8260 5865
rect 8300 5856 8352 5908
rect 12624 5899 12676 5908
rect 12624 5865 12633 5899
rect 12633 5865 12667 5899
rect 12667 5865 12676 5899
rect 12624 5856 12676 5865
rect 13268 5856 13320 5908
rect 14096 5899 14148 5908
rect 14096 5865 14105 5899
rect 14105 5865 14139 5899
rect 14139 5865 14148 5899
rect 14096 5856 14148 5865
rect 15292 5899 15344 5908
rect 15292 5865 15301 5899
rect 15301 5865 15335 5899
rect 15335 5865 15344 5899
rect 15292 5856 15344 5865
rect 15568 5856 15620 5908
rect 16580 5856 16632 5908
rect 16764 5899 16816 5908
rect 16764 5865 16773 5899
rect 16773 5865 16807 5899
rect 16807 5865 16816 5899
rect 16764 5856 16816 5865
rect 19432 5856 19484 5908
rect 19524 5856 19576 5908
rect 21364 5899 21416 5908
rect 21364 5865 21373 5899
rect 21373 5865 21407 5899
rect 21407 5865 21416 5899
rect 21364 5856 21416 5865
rect 22284 5899 22336 5908
rect 22284 5865 22293 5899
rect 22293 5865 22327 5899
rect 22327 5865 22336 5899
rect 22284 5856 22336 5865
rect 22928 5899 22980 5908
rect 22928 5865 22937 5899
rect 22937 5865 22971 5899
rect 22971 5865 22980 5899
rect 22928 5856 22980 5865
rect 23664 5856 23716 5908
rect 2964 5652 3016 5704
rect 3424 5652 3476 5704
rect 4252 5695 4304 5704
rect 4252 5661 4261 5695
rect 4261 5661 4295 5695
rect 4295 5661 4304 5695
rect 4252 5652 4304 5661
rect 5448 5652 5500 5704
rect 6552 5788 6604 5840
rect 7012 5788 7064 5840
rect 7288 5788 7340 5840
rect 10876 5788 10928 5840
rect 14556 5788 14608 5840
rect 17040 5788 17092 5840
rect 18880 5831 18932 5840
rect 18880 5797 18889 5831
rect 18889 5797 18923 5831
rect 18923 5797 18932 5831
rect 18880 5788 18932 5797
rect 19064 5788 19116 5840
rect 21548 5788 21600 5840
rect 22836 5831 22888 5840
rect 22836 5797 22845 5831
rect 22845 5797 22879 5831
rect 22879 5797 22888 5831
rect 22836 5788 22888 5797
rect 23204 5788 23256 5840
rect 25780 5831 25832 5840
rect 25780 5797 25789 5831
rect 25789 5797 25823 5831
rect 25823 5797 25832 5831
rect 25780 5788 25832 5797
rect 6368 5720 6420 5772
rect 6644 5720 6696 5772
rect 6920 5720 6972 5772
rect 9772 5720 9824 5772
rect 12348 5720 12400 5772
rect 13728 5720 13780 5772
rect 15660 5763 15712 5772
rect 15660 5729 15669 5763
rect 15669 5729 15703 5763
rect 15703 5729 15712 5763
rect 15660 5720 15712 5729
rect 19432 5763 19484 5772
rect 19432 5729 19441 5763
rect 19441 5729 19475 5763
rect 19475 5729 19484 5763
rect 19432 5720 19484 5729
rect 20720 5720 20772 5772
rect 22192 5720 22244 5772
rect 23664 5720 23716 5772
rect 26056 5720 26108 5772
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6552 5652 6604 5704
rect 8208 5652 8260 5704
rect 2596 5516 2648 5568
rect 2780 5516 2832 5568
rect 7012 5516 7064 5568
rect 11060 5652 11112 5704
rect 12256 5652 12308 5704
rect 15108 5695 15160 5704
rect 9956 5516 10008 5568
rect 12532 5584 12584 5636
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 14832 5584 14884 5636
rect 16120 5652 16172 5704
rect 16948 5695 17000 5704
rect 16948 5661 16957 5695
rect 16957 5661 16991 5695
rect 16991 5661 17000 5695
rect 16948 5652 17000 5661
rect 21364 5652 21416 5704
rect 23020 5695 23072 5704
rect 23020 5661 23029 5695
rect 23029 5661 23063 5695
rect 23063 5661 23072 5695
rect 23020 5652 23072 5661
rect 24676 5695 24728 5704
rect 24676 5661 24685 5695
rect 24685 5661 24719 5695
rect 24719 5661 24728 5695
rect 24676 5652 24728 5661
rect 18328 5627 18380 5636
rect 18328 5593 18337 5627
rect 18337 5593 18371 5627
rect 18371 5593 18380 5627
rect 18328 5584 18380 5593
rect 20812 5584 20864 5636
rect 21088 5584 21140 5636
rect 21640 5584 21692 5636
rect 23756 5584 23808 5636
rect 24032 5627 24084 5636
rect 24032 5593 24041 5627
rect 24041 5593 24075 5627
rect 24075 5593 24084 5627
rect 24032 5584 24084 5593
rect 24308 5584 24360 5636
rect 10876 5516 10928 5568
rect 11152 5516 11204 5568
rect 11796 5516 11848 5568
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 19340 5516 19392 5568
rect 19892 5516 19944 5568
rect 20260 5516 20312 5568
rect 21180 5516 21232 5568
rect 26424 5516 26476 5568
rect 5648 5414 5700 5466
rect 5712 5414 5764 5466
rect 5776 5414 5828 5466
rect 5840 5414 5892 5466
rect 14982 5414 15034 5466
rect 15046 5414 15098 5466
rect 15110 5414 15162 5466
rect 15174 5414 15226 5466
rect 24315 5414 24367 5466
rect 24379 5414 24431 5466
rect 24443 5414 24495 5466
rect 24507 5414 24559 5466
rect 3332 5312 3384 5364
rect 5080 5312 5132 5364
rect 6828 5312 6880 5364
rect 8300 5312 8352 5364
rect 11060 5312 11112 5364
rect 12348 5312 12400 5364
rect 14188 5312 14240 5364
rect 14556 5312 14608 5364
rect 15660 5312 15712 5364
rect 17040 5312 17092 5364
rect 20720 5312 20772 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 23480 5312 23532 5364
rect 24676 5355 24728 5364
rect 24676 5321 24685 5355
rect 24685 5321 24719 5355
rect 24719 5321 24728 5355
rect 24676 5312 24728 5321
rect 25872 5355 25924 5364
rect 25872 5321 25881 5355
rect 25881 5321 25915 5355
rect 25915 5321 25924 5355
rect 25872 5312 25924 5321
rect 10692 5244 10744 5296
rect 11612 5244 11664 5296
rect 15384 5244 15436 5296
rect 20076 5244 20128 5296
rect 22836 5244 22888 5296
rect 23756 5244 23808 5296
rect 25780 5244 25832 5296
rect 5448 5176 5500 5228
rect 6276 5176 6328 5228
rect 6920 5176 6972 5228
rect 7012 5176 7064 5228
rect 10876 5176 10928 5228
rect 18604 5219 18656 5228
rect 3792 5108 3844 5160
rect 4068 5108 4120 5160
rect 4712 5151 4764 5160
rect 4712 5117 4721 5151
rect 4721 5117 4755 5151
rect 4755 5117 4764 5151
rect 4712 5108 4764 5117
rect 6092 5108 6144 5160
rect 6552 5108 6604 5160
rect 9312 5151 9364 5160
rect 9312 5117 9321 5151
rect 9321 5117 9355 5151
rect 9355 5117 9364 5151
rect 9312 5108 9364 5117
rect 10140 5108 10192 5160
rect 756 5040 808 5092
rect 2688 5040 2740 5092
rect 3240 5040 3292 5092
rect 2412 5015 2464 5024
rect 2412 4981 2421 5015
rect 2421 4981 2455 5015
rect 2455 4981 2464 5015
rect 2412 4972 2464 4981
rect 2964 4972 3016 5024
rect 3792 4972 3844 5024
rect 6552 5015 6604 5024
rect 6552 4981 6561 5015
rect 6561 4981 6595 5015
rect 6595 4981 6604 5015
rect 6552 4972 6604 4981
rect 8116 5083 8168 5092
rect 8116 5049 8125 5083
rect 8125 5049 8159 5083
rect 8159 5049 8168 5083
rect 8116 5040 8168 5049
rect 11612 5108 11664 5160
rect 11888 5108 11940 5160
rect 13176 5108 13228 5160
rect 14188 5108 14240 5160
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 18972 5176 19024 5228
rect 19892 5176 19944 5228
rect 20996 5176 21048 5228
rect 22468 5176 22520 5228
rect 23204 5176 23256 5228
rect 24124 5176 24176 5228
rect 15568 5108 15620 5160
rect 16948 5108 17000 5160
rect 20536 5108 20588 5160
rect 21088 5108 21140 5160
rect 24032 5151 24084 5160
rect 24032 5117 24041 5151
rect 24041 5117 24075 5151
rect 24075 5117 24084 5151
rect 24032 5108 24084 5117
rect 25872 5108 25924 5160
rect 10968 5040 11020 5092
rect 13084 5040 13136 5092
rect 8024 4972 8076 5024
rect 8300 4972 8352 5024
rect 9128 4972 9180 5024
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 12532 4972 12584 5024
rect 13268 4972 13320 5024
rect 15108 5040 15160 5092
rect 16580 5040 16632 5092
rect 17500 5040 17552 5092
rect 20720 5040 20772 5092
rect 21640 5083 21692 5092
rect 21640 5049 21649 5083
rect 21649 5049 21683 5083
rect 21683 5049 21692 5083
rect 21640 5040 21692 5049
rect 22376 5040 22428 5092
rect 26332 5040 26384 5092
rect 14464 4972 14516 5024
rect 16764 4972 16816 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 18420 5015 18472 5024
rect 18420 4981 18429 5015
rect 18429 4981 18463 5015
rect 18463 4981 18472 5015
rect 18420 4972 18472 4981
rect 18512 5015 18564 5024
rect 18512 4981 18521 5015
rect 18521 4981 18555 5015
rect 18555 4981 18564 5015
rect 19064 5015 19116 5024
rect 18512 4972 18564 4981
rect 19064 4981 19073 5015
rect 19073 4981 19107 5015
rect 19107 4981 19116 5015
rect 19064 4972 19116 4981
rect 19524 4972 19576 5024
rect 20996 5015 21048 5024
rect 20996 4981 21005 5015
rect 21005 4981 21039 5015
rect 21039 4981 21048 5015
rect 20996 4972 21048 4981
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 22008 4972 22060 5024
rect 25044 5015 25096 5024
rect 25044 4981 25053 5015
rect 25053 4981 25087 5015
rect 25087 4981 25096 5015
rect 25044 4972 25096 4981
rect 25136 4972 25188 5024
rect 10315 4870 10367 4922
rect 10379 4870 10431 4922
rect 10443 4870 10495 4922
rect 10507 4870 10559 4922
rect 19648 4870 19700 4922
rect 19712 4870 19764 4922
rect 19776 4870 19828 4922
rect 19840 4870 19892 4922
rect 1952 4811 2004 4820
rect 1952 4777 1961 4811
rect 1961 4777 1995 4811
rect 1995 4777 2004 4811
rect 1952 4768 2004 4777
rect 2688 4768 2740 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3240 4811 3292 4820
rect 3240 4777 3249 4811
rect 3249 4777 3283 4811
rect 3283 4777 3292 4811
rect 3240 4768 3292 4777
rect 5172 4768 5224 4820
rect 8576 4811 8628 4820
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 9680 4768 9732 4820
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 12348 4768 12400 4820
rect 12624 4768 12676 4820
rect 14280 4768 14332 4820
rect 14832 4768 14884 4820
rect 15384 4768 15436 4820
rect 16580 4768 16632 4820
rect 18144 4811 18196 4820
rect 18144 4777 18153 4811
rect 18153 4777 18187 4811
rect 18187 4777 18196 4811
rect 18144 4768 18196 4777
rect 18328 4768 18380 4820
rect 3792 4700 3844 4752
rect 9772 4700 9824 4752
rect 9956 4743 10008 4752
rect 9956 4709 9965 4743
rect 9965 4709 9999 4743
rect 9999 4709 10008 4743
rect 9956 4700 10008 4709
rect 11428 4700 11480 4752
rect 3976 4632 4028 4684
rect 6828 4675 6880 4684
rect 6828 4641 6862 4675
rect 6862 4641 6880 4675
rect 3056 4607 3108 4616
rect 3056 4573 3065 4607
rect 3065 4573 3099 4607
rect 3099 4573 3108 4607
rect 3056 4564 3108 4573
rect 3332 4564 3384 4616
rect 1584 4539 1636 4548
rect 1584 4505 1593 4539
rect 1593 4505 1627 4539
rect 1627 4505 1636 4539
rect 1584 4496 1636 4505
rect 3424 4428 3476 4480
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 6828 4632 6880 4641
rect 10600 4675 10652 4684
rect 10600 4641 10609 4675
rect 10609 4641 10643 4675
rect 10643 4641 10652 4675
rect 10600 4632 10652 4641
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 9772 4564 9824 4616
rect 10140 4564 10192 4616
rect 10692 4607 10744 4616
rect 10692 4573 10701 4607
rect 10701 4573 10735 4607
rect 10735 4573 10744 4607
rect 10692 4564 10744 4573
rect 10784 4607 10836 4616
rect 10784 4573 10793 4607
rect 10793 4573 10827 4607
rect 10827 4573 10836 4607
rect 10784 4564 10836 4573
rect 12716 4632 12768 4684
rect 14004 4675 14056 4684
rect 14004 4641 14013 4675
rect 14013 4641 14047 4675
rect 14047 4641 14056 4675
rect 14004 4632 14056 4641
rect 12348 4607 12400 4616
rect 12348 4573 12357 4607
rect 12357 4573 12391 4607
rect 12391 4573 12400 4607
rect 12348 4564 12400 4573
rect 13176 4607 13228 4616
rect 13176 4573 13185 4607
rect 13185 4573 13219 4607
rect 13219 4573 13228 4607
rect 13176 4564 13228 4573
rect 15108 4700 15160 4752
rect 15292 4700 15344 4752
rect 18696 4768 18748 4820
rect 18880 4811 18932 4820
rect 18880 4777 18889 4811
rect 18889 4777 18923 4811
rect 18923 4777 18932 4811
rect 18880 4768 18932 4777
rect 19524 4768 19576 4820
rect 20076 4811 20128 4820
rect 20076 4777 20085 4811
rect 20085 4777 20119 4811
rect 20119 4777 20128 4811
rect 20076 4768 20128 4777
rect 23020 4768 23072 4820
rect 24032 4768 24084 4820
rect 24124 4811 24176 4820
rect 24124 4777 24133 4811
rect 24133 4777 24167 4811
rect 24167 4777 24176 4811
rect 24124 4768 24176 4777
rect 21364 4700 21416 4752
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 17040 4632 17092 4684
rect 22836 4675 22888 4684
rect 22836 4641 22845 4675
rect 22845 4641 22879 4675
rect 22879 4641 22888 4675
rect 22836 4632 22888 4641
rect 22928 4675 22980 4684
rect 22928 4641 22937 4675
rect 22937 4641 22971 4675
rect 22971 4641 22980 4675
rect 24492 4675 24544 4684
rect 22928 4632 22980 4641
rect 11152 4496 11204 4548
rect 11428 4496 11480 4548
rect 13728 4496 13780 4548
rect 16948 4564 17000 4616
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 17500 4607 17552 4616
rect 17500 4573 17509 4607
rect 17509 4573 17543 4607
rect 17543 4573 17552 4607
rect 17500 4564 17552 4573
rect 20904 4564 20956 4616
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 21916 4564 21968 4616
rect 23020 4607 23072 4616
rect 23020 4573 23029 4607
rect 23029 4573 23063 4607
rect 23063 4573 23072 4607
rect 23020 4564 23072 4573
rect 24492 4641 24501 4675
rect 24501 4641 24535 4675
rect 24535 4641 24544 4675
rect 24492 4632 24544 4641
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 19432 4496 19484 4548
rect 20536 4496 20588 4548
rect 23112 4496 23164 4548
rect 4344 4428 4396 4480
rect 6000 4428 6052 4480
rect 6736 4428 6788 4480
rect 7932 4471 7984 4480
rect 7932 4437 7941 4471
rect 7941 4437 7975 4471
rect 7975 4437 7984 4471
rect 7932 4428 7984 4437
rect 8944 4471 8996 4480
rect 8944 4437 8953 4471
rect 8953 4437 8987 4471
rect 8987 4437 8996 4471
rect 8944 4428 8996 4437
rect 9128 4428 9180 4480
rect 11060 4428 11112 4480
rect 11704 4471 11756 4480
rect 11704 4437 11713 4471
rect 11713 4437 11747 4471
rect 11747 4437 11756 4471
rect 11704 4428 11756 4437
rect 13636 4471 13688 4480
rect 13636 4437 13645 4471
rect 13645 4437 13679 4471
rect 13679 4437 13688 4471
rect 13636 4428 13688 4437
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 15568 4428 15620 4480
rect 20996 4428 21048 4480
rect 22100 4428 22152 4480
rect 23572 4428 23624 4480
rect 24676 4471 24728 4480
rect 24676 4437 24685 4471
rect 24685 4437 24719 4471
rect 24719 4437 24728 4471
rect 24676 4428 24728 4437
rect 24768 4428 24820 4480
rect 26240 4471 26292 4480
rect 26240 4437 26249 4471
rect 26249 4437 26283 4471
rect 26283 4437 26292 4471
rect 26240 4428 26292 4437
rect 5648 4326 5700 4378
rect 5712 4326 5764 4378
rect 5776 4326 5828 4378
rect 5840 4326 5892 4378
rect 14982 4326 15034 4378
rect 15046 4326 15098 4378
rect 15110 4326 15162 4378
rect 15174 4326 15226 4378
rect 24315 4326 24367 4378
rect 24379 4326 24431 4378
rect 24443 4326 24495 4378
rect 24507 4326 24559 4378
rect 2872 4224 2924 4276
rect 4068 4224 4120 4276
rect 4344 4267 4396 4276
rect 4344 4233 4353 4267
rect 4353 4233 4387 4267
rect 4387 4233 4396 4267
rect 4344 4224 4396 4233
rect 10692 4267 10744 4276
rect 10692 4233 10701 4267
rect 10701 4233 10735 4267
rect 10735 4233 10744 4267
rect 10692 4224 10744 4233
rect 11428 4224 11480 4276
rect 2320 4088 2372 4140
rect 3792 4156 3844 4208
rect 3424 4088 3476 4140
rect 12348 4224 12400 4276
rect 18512 4224 18564 4276
rect 18696 4224 18748 4276
rect 20996 4224 21048 4276
rect 22928 4224 22980 4276
rect 24124 4224 24176 4276
rect 6000 4156 6052 4208
rect 9128 4156 9180 4208
rect 5172 4088 5224 4140
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 8668 4088 8720 4140
rect 11888 4156 11940 4208
rect 13636 4156 13688 4208
rect 14188 4199 14240 4208
rect 11244 4088 11296 4140
rect 14188 4165 14197 4199
rect 14197 4165 14231 4199
rect 14231 4165 14240 4199
rect 14188 4156 14240 4165
rect 15936 4156 15988 4208
rect 16304 4156 16356 4208
rect 18052 4156 18104 4208
rect 14740 4131 14792 4140
rect 2688 4020 2740 4072
rect 2780 4020 2832 4072
rect 4068 4020 4120 4072
rect 4252 4020 4304 4072
rect 5080 4020 5132 4072
rect 6552 4020 6604 4072
rect 10968 4020 11020 4072
rect 12624 4020 12676 4072
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 14740 4097 14749 4131
rect 14749 4097 14783 4131
rect 14783 4097 14792 4131
rect 14740 4088 14792 4097
rect 14924 4131 14976 4140
rect 14924 4097 14933 4131
rect 14933 4097 14967 4131
rect 14967 4097 14976 4131
rect 14924 4088 14976 4097
rect 16764 4088 16816 4140
rect 18144 4088 18196 4140
rect 18604 4131 18656 4140
rect 13728 4020 13780 4072
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 16396 4020 16448 4072
rect 18604 4097 18613 4131
rect 18613 4097 18647 4131
rect 18647 4097 18656 4131
rect 18604 4088 18656 4097
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 21364 4156 21416 4208
rect 21732 4131 21784 4140
rect 21732 4097 21741 4131
rect 21741 4097 21775 4131
rect 21775 4097 21784 4131
rect 21732 4088 21784 4097
rect 23480 4088 23532 4140
rect 19432 4063 19484 4072
rect 19432 4029 19441 4063
rect 19441 4029 19475 4063
rect 19475 4029 19484 4063
rect 19432 4020 19484 4029
rect 1676 3995 1728 4004
rect 1676 3961 1685 3995
rect 1685 3961 1719 3995
rect 1719 3961 1728 3995
rect 1676 3952 1728 3961
rect 2504 3952 2556 4004
rect 3884 3952 3936 4004
rect 4804 3995 4856 4004
rect 4804 3961 4813 3995
rect 4813 3961 4847 3995
rect 4847 3961 4856 3995
rect 4804 3952 4856 3961
rect 1768 3927 1820 3936
rect 1768 3893 1777 3927
rect 1777 3893 1811 3927
rect 1811 3893 1820 3927
rect 1768 3884 1820 3893
rect 2688 3884 2740 3936
rect 6000 3884 6052 3936
rect 7932 3952 7984 4004
rect 10600 3952 10652 4004
rect 10876 3952 10928 4004
rect 8208 3927 8260 3936
rect 8208 3893 8217 3927
rect 8217 3893 8251 3927
rect 8251 3893 8260 3927
rect 8208 3884 8260 3893
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 8852 3884 8904 3893
rect 9220 3884 9272 3936
rect 9956 3884 10008 3936
rect 12624 3884 12676 3936
rect 13176 3927 13228 3936
rect 13176 3893 13185 3927
rect 13185 3893 13219 3927
rect 13219 3893 13228 3927
rect 13176 3884 13228 3893
rect 14004 3884 14056 3936
rect 14280 3927 14332 3936
rect 14280 3893 14289 3927
rect 14289 3893 14323 3927
rect 14323 3893 14332 3927
rect 14280 3884 14332 3893
rect 17868 3952 17920 4004
rect 16304 3884 16356 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17040 3884 17092 3936
rect 19248 3952 19300 4004
rect 18328 3884 18380 3936
rect 20720 4020 20772 4072
rect 20812 4020 20864 4072
rect 22008 4020 22060 4072
rect 22560 4020 22612 4072
rect 23020 4020 23072 4072
rect 23572 4020 23624 4072
rect 25228 4063 25280 4072
rect 20168 3952 20220 4004
rect 23756 3952 23808 4004
rect 23940 3952 23992 4004
rect 25228 4029 25237 4063
rect 25237 4029 25271 4063
rect 25271 4029 25280 4063
rect 25228 4020 25280 4029
rect 20720 3927 20772 3936
rect 20720 3893 20729 3927
rect 20729 3893 20763 3927
rect 20763 3893 20772 3927
rect 20720 3884 20772 3893
rect 20812 3884 20864 3936
rect 21180 3927 21232 3936
rect 21180 3893 21189 3927
rect 21189 3893 21223 3927
rect 21223 3893 21232 3927
rect 21180 3884 21232 3893
rect 23020 3884 23072 3936
rect 23480 3927 23532 3936
rect 23480 3893 23489 3927
rect 23489 3893 23523 3927
rect 23523 3893 23532 3927
rect 23480 3884 23532 3893
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 24124 3884 24176 3936
rect 24768 3884 24820 3936
rect 25044 3927 25096 3936
rect 25044 3893 25053 3927
rect 25053 3893 25087 3927
rect 25087 3893 25096 3927
rect 25044 3884 25096 3893
rect 25412 3927 25464 3936
rect 25412 3893 25421 3927
rect 25421 3893 25455 3927
rect 25455 3893 25464 3927
rect 25412 3884 25464 3893
rect 10315 3782 10367 3834
rect 10379 3782 10431 3834
rect 10443 3782 10495 3834
rect 10507 3782 10559 3834
rect 19648 3782 19700 3834
rect 19712 3782 19764 3834
rect 19776 3782 19828 3834
rect 19840 3782 19892 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 2504 3680 2556 3732
rect 2596 3680 2648 3732
rect 3976 3680 4028 3732
rect 5080 3723 5132 3732
rect 5080 3689 5089 3723
rect 5089 3689 5123 3723
rect 5123 3689 5132 3723
rect 5080 3680 5132 3689
rect 6920 3680 6972 3732
rect 9680 3723 9732 3732
rect 3884 3612 3936 3664
rect 4988 3612 5040 3664
rect 9680 3689 9689 3723
rect 9689 3689 9723 3723
rect 9723 3689 9732 3723
rect 9680 3680 9732 3689
rect 9864 3680 9916 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 1400 3587 1452 3596
rect 1400 3553 1409 3587
rect 1409 3553 1443 3587
rect 1443 3553 1452 3587
rect 1400 3544 1452 3553
rect 3976 3544 4028 3596
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 5908 3544 5960 3596
rect 10692 3612 10744 3664
rect 8300 3544 8352 3596
rect 8852 3544 8904 3596
rect 3056 3519 3108 3528
rect 3056 3485 3065 3519
rect 3065 3485 3099 3519
rect 3099 3485 3108 3519
rect 3056 3476 3108 3485
rect 3424 3476 3476 3528
rect 4068 3476 4120 3528
rect 5448 3476 5500 3528
rect 7012 3476 7064 3528
rect 7840 3451 7892 3460
rect 7840 3417 7849 3451
rect 7849 3417 7883 3451
rect 7883 3417 7892 3451
rect 7840 3408 7892 3417
rect 9588 3476 9640 3528
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 12164 3680 12216 3732
rect 12716 3680 12768 3732
rect 13176 3680 13228 3732
rect 13728 3680 13780 3732
rect 14280 3680 14332 3732
rect 15844 3680 15896 3732
rect 16488 3680 16540 3732
rect 17408 3680 17460 3732
rect 17868 3680 17920 3732
rect 20168 3680 20220 3732
rect 21916 3680 21968 3732
rect 22100 3680 22152 3732
rect 22836 3680 22888 3732
rect 24492 3723 24544 3732
rect 24492 3689 24501 3723
rect 24501 3689 24535 3723
rect 24535 3689 24544 3723
rect 24492 3680 24544 3689
rect 25228 3680 25280 3732
rect 11520 3612 11572 3664
rect 14096 3655 14148 3664
rect 14096 3621 14105 3655
rect 14105 3621 14139 3655
rect 14139 3621 14148 3655
rect 14096 3612 14148 3621
rect 15108 3612 15160 3664
rect 18880 3612 18932 3664
rect 19248 3655 19300 3664
rect 19248 3621 19257 3655
rect 19257 3621 19291 3655
rect 19291 3621 19300 3655
rect 19248 3612 19300 3621
rect 19432 3612 19484 3664
rect 20536 3612 20588 3664
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 14924 3544 14976 3596
rect 9128 3408 9180 3460
rect 14832 3476 14884 3528
rect 16580 3544 16632 3596
rect 17592 3544 17644 3596
rect 18052 3544 18104 3596
rect 19064 3544 19116 3596
rect 21272 3587 21324 3596
rect 21272 3553 21281 3587
rect 21281 3553 21315 3587
rect 21315 3553 21324 3587
rect 21272 3544 21324 3553
rect 24308 3612 24360 3664
rect 26240 3655 26292 3664
rect 26240 3621 26249 3655
rect 26249 3621 26283 3655
rect 26283 3621 26292 3655
rect 26240 3612 26292 3621
rect 22836 3587 22888 3596
rect 15384 3476 15436 3528
rect 16764 3476 16816 3528
rect 14556 3408 14608 3460
rect 15016 3408 15068 3460
rect 16672 3408 16724 3460
rect 17776 3519 17828 3528
rect 17776 3485 17785 3519
rect 17785 3485 17819 3519
rect 17819 3485 17828 3519
rect 17776 3476 17828 3485
rect 18972 3476 19024 3528
rect 20996 3476 21048 3528
rect 21364 3519 21416 3528
rect 21364 3485 21373 3519
rect 21373 3485 21407 3519
rect 21407 3485 21416 3519
rect 21364 3476 21416 3485
rect 22836 3553 22845 3587
rect 22845 3553 22879 3587
rect 22879 3553 22888 3587
rect 22836 3544 22888 3553
rect 22928 3587 22980 3596
rect 22928 3553 22937 3587
rect 22937 3553 22971 3587
rect 22971 3553 22980 3587
rect 22928 3544 22980 3553
rect 24952 3544 25004 3596
rect 21640 3476 21692 3528
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 23572 3476 23624 3528
rect 23940 3408 23992 3460
rect 8668 3340 8720 3392
rect 11244 3383 11296 3392
rect 11244 3349 11253 3383
rect 11253 3349 11287 3383
rect 11287 3349 11296 3383
rect 11244 3340 11296 3349
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 13728 3340 13780 3392
rect 17132 3340 17184 3392
rect 18328 3340 18380 3392
rect 19432 3340 19484 3392
rect 20260 3340 20312 3392
rect 23480 3383 23532 3392
rect 23480 3349 23489 3383
rect 23489 3349 23523 3383
rect 23523 3349 23532 3383
rect 23480 3340 23532 3349
rect 24032 3383 24084 3392
rect 24032 3349 24041 3383
rect 24041 3349 24075 3383
rect 24075 3349 24084 3383
rect 24032 3340 24084 3349
rect 25044 3383 25096 3392
rect 25044 3349 25053 3383
rect 25053 3349 25087 3383
rect 25087 3349 25096 3383
rect 25044 3340 25096 3349
rect 5648 3238 5700 3290
rect 5712 3238 5764 3290
rect 5776 3238 5828 3290
rect 5840 3238 5892 3290
rect 14982 3238 15034 3290
rect 15046 3238 15098 3290
rect 15110 3238 15162 3290
rect 15174 3238 15226 3290
rect 24315 3238 24367 3290
rect 24379 3238 24431 3290
rect 24443 3238 24495 3290
rect 24507 3238 24559 3290
rect 1676 3136 1728 3188
rect 3056 3136 3108 3188
rect 3516 3179 3568 3188
rect 3516 3145 3525 3179
rect 3525 3145 3559 3179
rect 3559 3145 3568 3179
rect 3516 3136 3568 3145
rect 3792 3136 3844 3188
rect 6644 3136 6696 3188
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10140 3136 10192 3188
rect 13728 3136 13780 3188
rect 13820 3179 13872 3188
rect 13820 3145 13829 3179
rect 13829 3145 13863 3179
rect 13863 3145 13872 3179
rect 13820 3136 13872 3145
rect 15476 3136 15528 3188
rect 16488 3179 16540 3188
rect 16488 3145 16497 3179
rect 16497 3145 16531 3179
rect 16531 3145 16540 3179
rect 16488 3136 16540 3145
rect 17776 3136 17828 3188
rect 18788 3136 18840 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 20904 3136 20956 3188
rect 4528 3111 4580 3120
rect 4528 3077 4537 3111
rect 4537 3077 4571 3111
rect 4571 3077 4580 3111
rect 4528 3068 4580 3077
rect 4988 3111 5040 3120
rect 4988 3077 4997 3111
rect 4997 3077 5031 3111
rect 5031 3077 5040 3111
rect 4988 3068 5040 3077
rect 5172 3068 5224 3120
rect 7288 3068 7340 3120
rect 9864 3068 9916 3120
rect 2320 3000 2372 3052
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 5264 3000 5316 3052
rect 6460 3000 6512 3052
rect 6644 3000 6696 3052
rect 7012 3000 7064 3052
rect 9404 3000 9456 3052
rect 11060 3000 11112 3052
rect 12440 3068 12492 3120
rect 16764 3068 16816 3120
rect 2872 2932 2924 2984
rect 5356 2932 5408 2984
rect 6092 2932 6144 2984
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 2136 2864 2188 2916
rect 7288 2907 7340 2916
rect 1952 2839 2004 2848
rect 1952 2805 1961 2839
rect 1961 2805 1995 2839
rect 1995 2805 2004 2839
rect 1952 2796 2004 2805
rect 2412 2796 2464 2848
rect 2780 2796 2832 2848
rect 3884 2839 3936 2848
rect 3884 2805 3893 2839
rect 3893 2805 3927 2839
rect 3927 2805 3936 2839
rect 3884 2796 3936 2805
rect 7288 2873 7297 2907
rect 7297 2873 7331 2907
rect 7331 2873 7340 2907
rect 7288 2864 7340 2873
rect 4068 2796 4120 2848
rect 4436 2796 4488 2848
rect 6000 2796 6052 2848
rect 6552 2796 6604 2848
rect 8484 2932 8536 2984
rect 8668 2975 8720 2984
rect 8668 2941 8702 2975
rect 8702 2941 8720 2975
rect 8668 2932 8720 2941
rect 9496 2932 9548 2984
rect 10784 2864 10836 2916
rect 17592 3000 17644 3052
rect 14648 2932 14700 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 15384 2975 15436 2984
rect 15384 2941 15418 2975
rect 15418 2941 15436 2975
rect 15384 2932 15436 2941
rect 18420 2975 18472 2984
rect 18420 2941 18429 2975
rect 18429 2941 18463 2975
rect 18463 2941 18472 2975
rect 18420 2932 18472 2941
rect 18512 2975 18564 2984
rect 18512 2941 18521 2975
rect 18521 2941 18555 2975
rect 18555 2941 18564 2975
rect 20628 3068 20680 3120
rect 21272 3136 21324 3188
rect 21824 3136 21876 3188
rect 23480 3179 23532 3188
rect 23480 3145 23489 3179
rect 23489 3145 23523 3179
rect 23523 3145 23532 3179
rect 23480 3136 23532 3145
rect 24676 3136 24728 3188
rect 24952 3136 25004 3188
rect 20536 3000 20588 3052
rect 18512 2932 18564 2941
rect 20352 2932 20404 2984
rect 22100 3068 22152 3120
rect 23020 3068 23072 3120
rect 23112 3068 23164 3120
rect 24584 3068 24636 3120
rect 25228 3068 25280 3120
rect 21640 3000 21692 3052
rect 22376 3000 22428 3052
rect 23848 3000 23900 3052
rect 23940 3000 23992 3052
rect 22928 2932 22980 2984
rect 23572 2932 23624 2984
rect 25228 2975 25280 2984
rect 25228 2941 25237 2975
rect 25237 2941 25271 2975
rect 25271 2941 25280 2975
rect 25228 2932 25280 2941
rect 8392 2796 8444 2848
rect 8668 2796 8720 2848
rect 9496 2796 9548 2848
rect 11336 2796 11388 2848
rect 13728 2864 13780 2916
rect 15660 2864 15712 2916
rect 21364 2864 21416 2916
rect 22744 2864 22796 2916
rect 23480 2864 23532 2916
rect 12532 2796 12584 2848
rect 14648 2839 14700 2848
rect 14648 2805 14657 2839
rect 14657 2805 14691 2839
rect 14691 2805 14700 2839
rect 14648 2796 14700 2805
rect 15844 2796 15896 2848
rect 20996 2796 21048 2848
rect 21824 2796 21876 2848
rect 23664 2839 23716 2848
rect 23664 2805 23673 2839
rect 23673 2805 23707 2839
rect 23707 2805 23716 2839
rect 23664 2796 23716 2805
rect 25136 2796 25188 2848
rect 26240 2839 26292 2848
rect 26240 2805 26249 2839
rect 26249 2805 26283 2839
rect 26283 2805 26292 2839
rect 26240 2796 26292 2805
rect 10315 2694 10367 2746
rect 10379 2694 10431 2746
rect 10443 2694 10495 2746
rect 10507 2694 10559 2746
rect 19648 2694 19700 2746
rect 19712 2694 19764 2746
rect 19776 2694 19828 2746
rect 19840 2694 19892 2746
rect 2136 2592 2188 2644
rect 3792 2592 3844 2644
rect 3884 2592 3936 2644
rect 4804 2592 4856 2644
rect 6184 2592 6236 2644
rect 6552 2592 6604 2644
rect 3148 2524 3200 2576
rect 1952 2456 2004 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 1768 2320 1820 2372
rect 4436 2456 4488 2508
rect 5080 2456 5132 2508
rect 7380 2592 7432 2644
rect 7840 2592 7892 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 10140 2592 10192 2644
rect 12256 2592 12308 2644
rect 12532 2592 12584 2644
rect 7932 2524 7984 2576
rect 8484 2524 8536 2576
rect 11336 2524 11388 2576
rect 13176 2567 13228 2576
rect 13176 2533 13210 2567
rect 13210 2533 13228 2567
rect 13176 2524 13228 2533
rect 10784 2456 10836 2508
rect 13452 2592 13504 2644
rect 13820 2592 13872 2644
rect 14556 2592 14608 2644
rect 16856 2635 16908 2644
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 17592 2592 17644 2644
rect 18052 2635 18104 2644
rect 18052 2601 18061 2635
rect 18061 2601 18095 2635
rect 18095 2601 18104 2635
rect 18052 2592 18104 2601
rect 21180 2635 21232 2644
rect 21180 2601 21189 2635
rect 21189 2601 21223 2635
rect 21223 2601 21232 2635
rect 21180 2592 21232 2601
rect 21640 2592 21692 2644
rect 21824 2592 21876 2644
rect 23204 2592 23256 2644
rect 23572 2592 23624 2644
rect 24124 2592 24176 2644
rect 24952 2592 25004 2644
rect 25872 2592 25924 2644
rect 14832 2524 14884 2576
rect 16488 2524 16540 2576
rect 15200 2456 15252 2508
rect 15568 2456 15620 2508
rect 18696 2499 18748 2508
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 1952 2295 2004 2304
rect 1952 2261 1961 2295
rect 1961 2261 1995 2295
rect 1995 2261 2004 2295
rect 1952 2252 2004 2261
rect 2872 2252 2924 2304
rect 6276 2252 6328 2304
rect 11244 2252 11296 2304
rect 14464 2252 14516 2304
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 20352 2524 20404 2576
rect 18788 2388 18840 2440
rect 19800 2320 19852 2372
rect 21640 2499 21692 2508
rect 21640 2465 21649 2499
rect 21649 2465 21683 2499
rect 21683 2465 21692 2499
rect 21640 2456 21692 2465
rect 22376 2456 22428 2508
rect 24032 2456 24084 2508
rect 24124 2456 24176 2508
rect 24768 2456 24820 2508
rect 26056 2456 26108 2508
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 23664 2388 23716 2440
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 19892 2252 19944 2304
rect 20904 2295 20956 2304
rect 20904 2261 20913 2295
rect 20913 2261 20947 2295
rect 20947 2261 20956 2295
rect 20904 2252 20956 2261
rect 21640 2252 21692 2304
rect 22928 2295 22980 2304
rect 22928 2261 22937 2295
rect 22937 2261 22971 2295
rect 22971 2261 22980 2295
rect 22928 2252 22980 2261
rect 23848 2252 23900 2304
rect 5648 2150 5700 2202
rect 5712 2150 5764 2202
rect 5776 2150 5828 2202
rect 5840 2150 5892 2202
rect 14982 2150 15034 2202
rect 15046 2150 15098 2202
rect 15110 2150 15162 2202
rect 15174 2150 15226 2202
rect 24315 2150 24367 2202
rect 24379 2150 24431 2202
rect 24443 2150 24495 2202
rect 24507 2150 24559 2202
rect 12900 2048 12952 2100
rect 15384 2048 15436 2100
rect 13268 1980 13320 2032
rect 17132 1980 17184 2032
rect 12072 1572 12124 1624
rect 12532 1572 12584 1624
rect 6552 1504 6604 1556
rect 9220 1504 9272 1556
rect 3424 1436 3476 1488
rect 4528 1436 4580 1488
<< metal2 >>
rect 294 27520 350 28000
rect 846 27520 902 28000
rect 1398 27520 1454 28000
rect 2042 27520 2098 28000
rect 2594 27520 2650 28000
rect 3146 27520 3202 28000
rect 3790 27520 3846 28000
rect 4250 27704 4306 27713
rect 4250 27639 4306 27648
rect 20 21412 72 21418
rect 20 21354 72 21360
rect 32 12374 60 21354
rect 308 12986 336 27520
rect 754 27160 810 27169
rect 754 27095 810 27104
rect 768 21486 796 27095
rect 756 21480 808 21486
rect 756 21422 808 21428
rect 860 21418 888 27520
rect 1306 26616 1362 26625
rect 1306 26551 1362 26560
rect 1214 25936 1270 25945
rect 1214 25871 1270 25880
rect 1122 24848 1178 24857
rect 1122 24783 1178 24792
rect 938 24168 994 24177
rect 938 24103 994 24112
rect 848 21412 900 21418
rect 848 21354 900 21360
rect 952 20602 980 24103
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1136 20058 1164 24783
rect 1228 21894 1256 25871
rect 1216 21888 1268 21894
rect 1216 21830 1268 21836
rect 1320 21690 1348 26551
rect 1412 25242 1440 27520
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 1412 25214 1716 25242
rect 1400 25152 1452 25158
rect 1400 25094 1452 25100
rect 1308 21684 1360 21690
rect 1308 21626 1360 21632
rect 1412 20097 1440 25094
rect 1584 24744 1636 24750
rect 1584 24686 1636 24692
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1504 22930 1532 23462
rect 1596 23322 1624 24686
rect 1688 23322 1716 25214
rect 1780 24886 1808 25842
rect 2056 25242 2084 27520
rect 2136 25356 2188 25362
rect 2136 25298 2188 25304
rect 1872 25214 2084 25242
rect 1768 24880 1820 24886
rect 1768 24822 1820 24828
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1676 23316 1728 23322
rect 1676 23258 1728 23264
rect 1504 22902 1624 22930
rect 1492 22772 1544 22778
rect 1492 22714 1544 22720
rect 1398 20088 1454 20097
rect 1124 20052 1176 20058
rect 1398 20023 1454 20032
rect 1124 19994 1176 20000
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1412 16561 1440 16594
rect 1398 16552 1454 16561
rect 1398 16487 1454 16496
rect 1412 13258 1440 16487
rect 1504 13569 1532 22714
rect 1596 19446 1624 22902
rect 1676 22568 1728 22574
rect 1676 22510 1728 22516
rect 1584 19440 1636 19446
rect 1584 19382 1636 19388
rect 1584 19168 1636 19174
rect 1584 19110 1636 19116
rect 1596 15473 1624 19110
rect 1582 15464 1638 15473
rect 1582 15399 1638 15408
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 1596 14929 1624 15030
rect 1582 14920 1638 14929
rect 1582 14855 1638 14864
rect 1688 14770 1716 22510
rect 1596 14742 1716 14770
rect 1596 13841 1624 14742
rect 1674 14648 1730 14657
rect 1674 14583 1730 14592
rect 1582 13832 1638 13841
rect 1582 13767 1638 13776
rect 1582 13696 1638 13705
rect 1582 13631 1638 13640
rect 1490 13560 1546 13569
rect 1490 13495 1546 13504
rect 1400 13252 1452 13258
rect 1400 13194 1452 13200
rect 296 12980 348 12986
rect 296 12922 348 12928
rect 1504 12696 1532 13495
rect 1412 12668 1532 12696
rect 1412 12458 1440 12668
rect 1490 12608 1546 12617
rect 1490 12543 1546 12552
rect 1320 12430 1440 12458
rect 20 12368 72 12374
rect 20 12310 72 12316
rect 1320 12186 1348 12430
rect 1398 12336 1454 12345
rect 1398 12271 1400 12280
rect 1452 12271 1454 12280
rect 1400 12242 1452 12248
rect 1320 12158 1440 12186
rect 1412 11898 1440 12158
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1398 11520 1454 11529
rect 1398 11455 1454 11464
rect 1412 11218 1440 11455
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 572 8560 624 8566
rect 570 8528 572 8537
rect 624 8528 626 8537
rect 570 8463 626 8472
rect 1412 8430 1440 10367
rect 1504 8634 1532 12543
rect 1596 10810 1624 13631
rect 1688 12442 1716 14583
rect 1780 13734 1808 24006
rect 1872 22778 1900 25214
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 1952 24336 2004 24342
rect 1952 24278 2004 24284
rect 1964 23474 1992 24278
rect 2056 23730 2084 25094
rect 2148 24614 2176 25298
rect 2608 24970 2636 27520
rect 2870 25392 2926 25401
rect 2870 25327 2926 25336
rect 2332 24942 2636 24970
rect 2136 24608 2188 24614
rect 2136 24550 2188 24556
rect 2148 24041 2176 24550
rect 2226 24168 2282 24177
rect 2226 24103 2282 24112
rect 2134 24032 2190 24041
rect 2134 23967 2190 23976
rect 2044 23724 2096 23730
rect 2096 23684 2176 23712
rect 2044 23666 2096 23672
rect 1964 23446 2084 23474
rect 1952 23316 2004 23322
rect 1952 23258 2004 23264
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1860 22500 1912 22506
rect 1860 22442 1912 22448
rect 1872 21146 1900 22442
rect 1860 21140 1912 21146
rect 1860 21082 1912 21088
rect 1860 19304 1912 19310
rect 1860 19246 1912 19252
rect 1872 16046 1900 19246
rect 1964 17921 1992 23258
rect 2056 22234 2084 23446
rect 2044 22228 2096 22234
rect 2044 22170 2096 22176
rect 2148 20602 2176 23684
rect 2240 23594 2268 24103
rect 2228 23588 2280 23594
rect 2228 23530 2280 23536
rect 2240 22506 2268 23530
rect 2332 22574 2360 24942
rect 2504 24744 2556 24750
rect 2502 24712 2504 24721
rect 2780 24744 2832 24750
rect 2556 24712 2558 24721
rect 2502 24647 2558 24656
rect 2608 24704 2780 24732
rect 2410 24440 2466 24449
rect 2410 24375 2412 24384
rect 2464 24375 2466 24384
rect 2412 24346 2464 24352
rect 2424 23610 2452 24346
rect 2504 24200 2556 24206
rect 2504 24142 2556 24148
rect 2516 23730 2544 24142
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2424 23582 2544 23610
rect 2410 23352 2466 23361
rect 2410 23287 2412 23296
rect 2464 23287 2466 23296
rect 2412 23258 2464 23264
rect 2410 23216 2466 23225
rect 2410 23151 2466 23160
rect 2424 23118 2452 23151
rect 2412 23112 2464 23118
rect 2412 23054 2464 23060
rect 2412 22976 2464 22982
rect 2412 22918 2464 22924
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 2228 22500 2280 22506
rect 2228 22442 2280 22448
rect 2424 22166 2452 22918
rect 2412 22160 2464 22166
rect 2412 22102 2464 22108
rect 2320 22092 2372 22098
rect 2320 22034 2372 22040
rect 2332 22001 2360 22034
rect 2412 22024 2464 22030
rect 2318 21992 2374 22001
rect 2412 21966 2464 21972
rect 2318 21927 2374 21936
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2332 21146 2360 21830
rect 2424 21729 2452 21966
rect 2410 21720 2466 21729
rect 2516 21690 2544 23582
rect 2608 22778 2636 24704
rect 2780 24686 2832 24692
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2596 22024 2648 22030
rect 2596 21966 2648 21972
rect 2410 21655 2466 21664
rect 2504 21684 2556 21690
rect 2320 21140 2372 21146
rect 2320 21082 2372 21088
rect 2424 21078 2452 21655
rect 2504 21626 2556 21632
rect 2502 21584 2558 21593
rect 2608 21554 2636 21966
rect 2502 21519 2558 21528
rect 2596 21548 2648 21554
rect 2412 21072 2464 21078
rect 2412 21014 2464 21020
rect 2318 20632 2374 20641
rect 2136 20596 2188 20602
rect 2318 20567 2374 20576
rect 2136 20538 2188 20544
rect 2332 20262 2360 20567
rect 2412 20460 2464 20466
rect 2412 20402 2464 20408
rect 2424 20369 2452 20402
rect 2410 20360 2466 20369
rect 2410 20295 2466 20304
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2332 20058 2360 20198
rect 2320 20052 2372 20058
rect 2372 20012 2452 20040
rect 2320 19994 2372 20000
rect 2320 19712 2372 19718
rect 2320 19654 2372 19660
rect 2044 19440 2096 19446
rect 2044 19382 2096 19388
rect 1950 17912 2006 17921
rect 1950 17847 2006 17856
rect 2056 16658 2084 19382
rect 2136 19304 2188 19310
rect 2134 19272 2136 19281
rect 2188 19272 2190 19281
rect 2134 19207 2190 19216
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 2148 18358 2176 18770
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 2240 18290 2268 18702
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2240 17746 2268 18226
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2136 17332 2188 17338
rect 2240 17320 2268 17682
rect 2188 17292 2268 17320
rect 2136 17274 2188 17280
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1860 16040 1912 16046
rect 1860 15982 1912 15988
rect 1858 15464 1914 15473
rect 1858 15399 1860 15408
rect 1912 15399 1914 15408
rect 1860 15370 1912 15376
rect 1860 14272 1912 14278
rect 1860 14214 1912 14220
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1768 11552 1820 11558
rect 1768 11494 1820 11500
rect 1780 11393 1808 11494
rect 1766 11384 1822 11393
rect 1766 11319 1822 11328
rect 1872 11200 1900 14214
rect 1964 13870 1992 16526
rect 2044 15904 2096 15910
rect 2044 15846 2096 15852
rect 2056 15065 2084 15846
rect 2042 15056 2098 15065
rect 2042 14991 2098 15000
rect 2044 14816 2096 14822
rect 2044 14758 2096 14764
rect 2056 13977 2084 14758
rect 2148 14414 2176 16934
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2240 15366 2268 15914
rect 2228 15360 2280 15366
rect 2226 15328 2228 15337
rect 2280 15328 2282 15337
rect 2226 15263 2282 15272
rect 2332 14618 2360 19654
rect 2424 19417 2452 20012
rect 2410 19408 2466 19417
rect 2410 19343 2466 19352
rect 2412 19304 2464 19310
rect 2412 19246 2464 19252
rect 2424 18766 2452 19246
rect 2412 18760 2464 18766
rect 2412 18702 2464 18708
rect 2516 18578 2544 21519
rect 2596 21490 2648 21496
rect 2608 20942 2636 21490
rect 2596 20936 2648 20942
rect 2596 20878 2648 20884
rect 2608 20466 2636 20878
rect 2700 20777 2728 24550
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 2792 22982 2820 23462
rect 2884 23322 2912 25327
rect 3056 25220 3108 25226
rect 3056 25162 3108 25168
rect 3068 24954 3096 25162
rect 3056 24948 3108 24954
rect 3056 24890 3108 24896
rect 2964 24676 3016 24682
rect 2964 24618 3016 24624
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 2884 22778 2912 23258
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 2780 22704 2832 22710
rect 2780 22646 2832 22652
rect 2686 20768 2742 20777
rect 2686 20703 2742 20712
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2608 19938 2636 20402
rect 2608 19910 2728 19938
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2608 18970 2636 19790
rect 2700 19378 2728 19910
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2596 18964 2648 18970
rect 2596 18906 2648 18912
rect 2424 18550 2544 18578
rect 2424 16590 2452 18550
rect 2596 16788 2648 16794
rect 2596 16730 2648 16736
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 2424 16153 2452 16390
rect 2410 16144 2466 16153
rect 2516 16114 2544 16662
rect 2410 16079 2466 16088
rect 2504 16108 2556 16114
rect 2424 15570 2452 16079
rect 2504 16050 2556 16056
rect 2412 15564 2464 15570
rect 2412 15506 2464 15512
rect 2608 15450 2636 16730
rect 2700 16640 2728 19110
rect 2792 17785 2820 22646
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2884 20602 2912 20810
rect 2872 20596 2924 20602
rect 2872 20538 2924 20544
rect 2870 20088 2926 20097
rect 2870 20023 2926 20032
rect 2884 19990 2912 20023
rect 2872 19984 2924 19990
rect 2872 19926 2924 19932
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2884 18222 2912 19450
rect 2976 19009 3004 24618
rect 3068 23610 3096 24890
rect 3160 24857 3188 27520
rect 3240 25492 3292 25498
rect 3240 25434 3292 25440
rect 3146 24848 3202 24857
rect 3146 24783 3202 24792
rect 3148 24064 3200 24070
rect 3148 24006 3200 24012
rect 3160 23730 3188 24006
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3068 23582 3188 23610
rect 3056 22976 3108 22982
rect 3056 22918 3108 22924
rect 3068 21962 3096 22918
rect 3160 22438 3188 23582
rect 3148 22432 3200 22438
rect 3148 22374 3200 22380
rect 3056 21956 3108 21962
rect 3056 21898 3108 21904
rect 3252 21321 3280 25434
rect 3424 25356 3476 25362
rect 3424 25298 3476 25304
rect 3436 24818 3464 25298
rect 3516 25152 3568 25158
rect 3516 25094 3568 25100
rect 3700 25152 3752 25158
rect 3700 25094 3752 25100
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3332 24200 3384 24206
rect 3332 24142 3384 24148
rect 3424 24200 3476 24206
rect 3424 24142 3476 24148
rect 3344 23526 3372 24142
rect 3332 23520 3384 23526
rect 3332 23462 3384 23468
rect 3344 23322 3372 23462
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 3436 23225 3464 24142
rect 3528 23866 3556 25094
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3422 23216 3478 23225
rect 3422 23151 3424 23160
rect 3476 23151 3478 23160
rect 3424 23122 3476 23128
rect 3436 23091 3464 23122
rect 3330 23080 3386 23089
rect 3330 23015 3386 23024
rect 3344 22409 3372 23015
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3330 22400 3386 22409
rect 3330 22335 3386 22344
rect 3238 21312 3294 21321
rect 3238 21247 3294 21256
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3160 20534 3188 21082
rect 3148 20528 3200 20534
rect 3148 20470 3200 20476
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 3056 19304 3108 19310
rect 3054 19272 3056 19281
rect 3108 19272 3110 19281
rect 3054 19207 3110 19216
rect 2962 19000 3018 19009
rect 3160 18970 3188 19751
rect 3332 19168 3384 19174
rect 3332 19110 3384 19116
rect 2962 18935 3018 18944
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2884 17814 2912 18158
rect 2976 17882 3004 18634
rect 3160 18426 3188 18906
rect 3240 18760 3292 18766
rect 3240 18702 3292 18708
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3252 18358 3280 18702
rect 3344 18630 3372 19110
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3146 17912 3202 17921
rect 2964 17876 3016 17882
rect 3146 17847 3202 17856
rect 2964 17818 3016 17824
rect 2872 17808 2924 17814
rect 2778 17776 2834 17785
rect 2872 17750 2924 17756
rect 2778 17711 2834 17720
rect 2884 17626 2912 17750
rect 2792 17598 2912 17626
rect 2792 16794 2820 17598
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2884 17066 2912 17478
rect 3054 17096 3110 17105
rect 2872 17060 2924 17066
rect 3054 17031 3110 17040
rect 2872 17002 2924 17008
rect 2962 16960 3018 16969
rect 2962 16895 3018 16904
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2700 16612 2820 16640
rect 2792 16572 2820 16612
rect 2976 16590 3004 16895
rect 3068 16658 3096 17031
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16584 3016 16590
rect 2792 16544 2912 16572
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 15910 2728 16390
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2516 15422 2636 15450
rect 2410 14648 2466 14657
rect 2320 14612 2372 14618
rect 2410 14583 2412 14592
rect 2320 14554 2372 14560
rect 2464 14583 2466 14592
rect 2412 14554 2464 14560
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2042 13968 2098 13977
rect 2148 13938 2176 14350
rect 2228 14000 2280 14006
rect 2228 13942 2280 13948
rect 2042 13903 2098 13912
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 2042 13832 2098 13841
rect 1964 13258 1992 13806
rect 2042 13767 2098 13776
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 2056 13138 2084 13767
rect 2148 13530 2176 13874
rect 2136 13524 2188 13530
rect 2136 13466 2188 13472
rect 2240 13394 2268 13942
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2056 13110 2176 13138
rect 2042 13016 2098 13025
rect 2042 12951 2044 12960
rect 2096 12951 2098 12960
rect 2044 12922 2096 12928
rect 2148 12714 2176 13110
rect 2136 12708 2188 12714
rect 2136 12650 2188 12656
rect 2148 11694 2176 12650
rect 2136 11688 2188 11694
rect 2240 11665 2268 13330
rect 2332 12170 2360 13670
rect 2424 13530 2452 14554
rect 2412 13524 2464 13530
rect 2412 13466 2464 13472
rect 2412 12640 2464 12646
rect 2410 12608 2412 12617
rect 2464 12608 2466 12617
rect 2410 12543 2466 12552
rect 2424 12374 2452 12543
rect 2516 12374 2544 15422
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2608 13734 2636 15302
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2700 13546 2728 15846
rect 2884 15162 2912 16544
rect 2964 16526 3016 16532
rect 2976 16250 3004 16526
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3056 16108 3108 16114
rect 3056 16050 3108 16056
rect 2964 15564 3016 15570
rect 2964 15506 3016 15512
rect 2976 15348 3004 15506
rect 3068 15502 3096 16050
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2976 15320 3096 15348
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2962 15056 3018 15065
rect 2962 14991 3018 15000
rect 2976 14958 3004 14991
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 3068 14890 3096 15320
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2884 14550 2912 14758
rect 2872 14544 2924 14550
rect 2870 14512 2872 14521
rect 2924 14512 2926 14521
rect 2780 14476 2832 14482
rect 2870 14447 2926 14456
rect 2780 14418 2832 14424
rect 2792 14074 2820 14418
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 3068 13705 3096 14826
rect 3054 13696 3110 13705
rect 3054 13631 3110 13640
rect 2608 13518 2728 13546
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2424 11762 2452 12174
rect 2412 11756 2464 11762
rect 2412 11698 2464 11704
rect 2136 11630 2188 11636
rect 2226 11656 2282 11665
rect 2148 11354 2176 11630
rect 2226 11591 2282 11600
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 1780 11172 1900 11200
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1780 10441 1808 11172
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1766 10432 1822 10441
rect 1766 10367 1822 10376
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 8945 1808 9318
rect 1766 8936 1822 8945
rect 1676 8900 1728 8906
rect 1766 8871 1822 8880
rect 1676 8842 1728 8848
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1582 7848 1638 7857
rect 1412 7041 1440 7822
rect 1582 7783 1638 7792
rect 1492 7744 1544 7750
rect 1492 7686 1544 7692
rect 1398 7032 1454 7041
rect 1398 6967 1454 6976
rect 1504 6916 1532 7686
rect 1596 7546 1624 7783
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1688 7313 1716 8842
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1674 7304 1730 7313
rect 1674 7239 1730 7248
rect 1412 6888 1532 6916
rect 756 5092 808 5098
rect 756 5034 808 5040
rect 768 4457 796 5034
rect 754 4448 810 4457
rect 754 4383 810 4392
rect 1412 3602 1440 6888
rect 1780 5914 1808 8774
rect 1872 8401 1900 11018
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 10033 2084 10406
rect 2042 10024 2098 10033
rect 2042 9959 2098 9968
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1964 9489 1992 9862
rect 2148 9518 2176 11018
rect 2410 10296 2466 10305
rect 2516 10266 2544 11222
rect 2608 10985 2636 13518
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2700 12850 2728 13398
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3068 12986 3096 13262
rect 2780 12980 2832 12986
rect 2780 12922 2832 12928
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2688 12844 2740 12850
rect 2688 12786 2740 12792
rect 2792 12442 2820 12922
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 3160 12306 3188 17847
rect 3344 14618 3372 18566
rect 3436 18426 3464 22918
rect 3528 22574 3556 23802
rect 3712 23526 3740 25094
rect 3804 24857 3832 27520
rect 4160 25356 4212 25362
rect 4160 25298 4212 25304
rect 3976 25152 4028 25158
rect 3976 25094 4028 25100
rect 3790 24848 3846 24857
rect 3790 24783 3846 24792
rect 3790 23760 3846 23769
rect 3790 23695 3846 23704
rect 3700 23520 3752 23526
rect 3700 23462 3752 23468
rect 3608 23248 3660 23254
rect 3712 23225 3740 23462
rect 3608 23190 3660 23196
rect 3698 23216 3754 23225
rect 3620 23089 3648 23190
rect 3698 23151 3754 23160
rect 3606 23080 3662 23089
rect 3606 23015 3608 23024
rect 3660 23015 3662 23024
rect 3608 22986 3660 22992
rect 3700 22772 3752 22778
rect 3700 22714 3752 22720
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 3514 22264 3570 22273
rect 3514 22199 3570 22208
rect 3528 21690 3556 22199
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 3620 21486 3648 21830
rect 3516 21480 3568 21486
rect 3516 21422 3568 21428
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 3528 21321 3556 21422
rect 3608 21344 3660 21350
rect 3514 21312 3570 21321
rect 3608 21286 3660 21292
rect 3514 21247 3570 21256
rect 3620 20806 3648 21286
rect 3608 20800 3660 20806
rect 3608 20742 3660 20748
rect 3516 20528 3568 20534
rect 3620 20505 3648 20742
rect 3712 20602 3740 22714
rect 3700 20596 3752 20602
rect 3700 20538 3752 20544
rect 3516 20470 3568 20476
rect 3606 20496 3662 20505
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3436 17678 3464 18362
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17082 3464 17614
rect 3528 17338 3556 20470
rect 3804 20482 3832 23695
rect 3882 23488 3938 23497
rect 3882 23423 3938 23432
rect 3896 22545 3924 23423
rect 3882 22536 3938 22545
rect 3882 22471 3938 22480
rect 3884 21888 3936 21894
rect 3988 21865 4016 25094
rect 4172 24818 4200 25298
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4264 24206 4292 27639
rect 4342 27520 4398 28000
rect 4894 27520 4950 28000
rect 5538 27520 5594 28000
rect 6090 27520 6146 28000
rect 6642 27520 6698 28000
rect 7286 27520 7342 28000
rect 7838 27520 7894 28000
rect 8390 27520 8446 28000
rect 9034 27520 9090 28000
rect 9586 27520 9642 28000
rect 10138 27520 10194 28000
rect 10782 27520 10838 28000
rect 11334 27520 11390 28000
rect 11886 27520 11942 28000
rect 12530 27520 12586 28000
rect 13082 27520 13138 28000
rect 13634 27520 13690 28000
rect 14278 27520 14334 28000
rect 14830 27520 14886 28000
rect 15382 27520 15438 28000
rect 16026 27520 16082 28000
rect 16578 27520 16634 28000
rect 17130 27520 17186 28000
rect 17774 27520 17830 28000
rect 18326 27520 18382 28000
rect 18878 27520 18934 28000
rect 19522 27520 19578 28000
rect 20074 27520 20130 28000
rect 20626 27520 20682 28000
rect 21270 27520 21326 28000
rect 21822 27520 21878 28000
rect 22374 27520 22430 28000
rect 23018 27520 23074 28000
rect 23570 27520 23626 28000
rect 23846 27704 23902 27713
rect 23846 27639 23902 27648
rect 4252 24200 4304 24206
rect 4252 24142 4304 24148
rect 4068 24132 4120 24138
rect 4068 24074 4120 24080
rect 4080 22166 4108 24074
rect 4160 24064 4212 24070
rect 4160 24006 4212 24012
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 4172 22098 4200 24006
rect 4264 23322 4292 24142
rect 4252 23316 4304 23322
rect 4252 23258 4304 23264
rect 4250 22672 4306 22681
rect 4250 22607 4306 22616
rect 4160 22092 4212 22098
rect 4160 22034 4212 22040
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3884 21830 3936 21836
rect 3974 21856 4030 21865
rect 3896 20874 3924 21830
rect 3974 21791 4030 21800
rect 4080 21146 4108 21966
rect 4068 21140 4120 21146
rect 4068 21082 4120 21088
rect 3976 21004 4028 21010
rect 3976 20946 4028 20952
rect 3884 20868 3936 20874
rect 3884 20810 3936 20816
rect 3606 20431 3662 20440
rect 3712 20454 3832 20482
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3712 17270 3740 20454
rect 3792 20392 3844 20398
rect 3792 20334 3844 20340
rect 3804 19718 3832 20334
rect 3896 19922 3924 20810
rect 3988 19990 4016 20946
rect 4264 20641 4292 22607
rect 4356 22386 4384 27520
rect 4710 26208 4766 26217
rect 4710 26143 4766 26152
rect 4436 24880 4488 24886
rect 4436 24822 4488 24828
rect 4448 24614 4476 24822
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4448 23730 4476 24550
rect 4436 23724 4488 23730
rect 4436 23666 4488 23672
rect 4448 22982 4476 23666
rect 4528 23316 4580 23322
rect 4528 23258 4580 23264
rect 4436 22976 4488 22982
rect 4436 22918 4488 22924
rect 4448 22506 4476 22918
rect 4436 22500 4488 22506
rect 4436 22442 4488 22448
rect 4356 22358 4476 22386
rect 4250 20632 4306 20641
rect 4250 20567 4306 20576
rect 4342 20224 4398 20233
rect 4342 20159 4398 20168
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 4066 19952 4122 19961
rect 3884 19916 3936 19922
rect 4066 19887 4068 19896
rect 3884 19858 3936 19864
rect 4120 19887 4122 19896
rect 4068 19858 4120 19864
rect 3884 19780 3936 19786
rect 3884 19722 3936 19728
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19446 3832 19654
rect 3792 19440 3844 19446
rect 3792 19382 3844 19388
rect 3804 19242 3832 19382
rect 3896 19378 3924 19722
rect 4080 19514 4108 19858
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3884 19372 3936 19378
rect 3884 19314 3936 19320
rect 3792 19236 3844 19242
rect 3792 19178 3844 19184
rect 3896 18970 3924 19314
rect 3884 18964 3936 18970
rect 3884 18906 3936 18912
rect 3882 18864 3938 18873
rect 3882 18799 3884 18808
rect 3936 18799 3938 18808
rect 3884 18770 3936 18776
rect 4160 18760 4212 18766
rect 3988 18720 4160 18748
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 3896 17882 3924 17983
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3436 17054 3556 17082
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16726 3464 16934
rect 3528 16794 3556 17054
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3436 15910 3464 16662
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3240 14068 3292 14074
rect 3240 14010 3292 14016
rect 3252 13530 3280 14010
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3436 13326 3464 15846
rect 3528 15026 3556 16730
rect 3608 16584 3660 16590
rect 3608 16526 3660 16532
rect 3620 15910 3648 16526
rect 3712 16130 3740 17206
rect 3792 17060 3844 17066
rect 3792 17002 3844 17008
rect 3804 16794 3832 17002
rect 3882 16824 3938 16833
rect 3792 16788 3844 16794
rect 3882 16759 3938 16768
rect 3792 16730 3844 16736
rect 3712 16102 3832 16130
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3608 15904 3660 15910
rect 3606 15872 3608 15881
rect 3660 15872 3662 15881
rect 3606 15807 3662 15816
rect 3712 15706 3740 15982
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3804 15638 3832 16102
rect 3896 15910 3924 16759
rect 3988 16046 4016 18720
rect 4160 18702 4212 18708
rect 4068 18624 4120 18630
rect 4068 18566 4120 18572
rect 4080 16697 4108 18566
rect 4264 17241 4292 19654
rect 4250 17232 4306 17241
rect 4250 17167 4306 17176
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3804 15094 3832 15574
rect 4068 15496 4120 15502
rect 4356 15450 4384 20159
rect 4068 15438 4120 15444
rect 4080 15178 4108 15438
rect 4264 15422 4384 15450
rect 4080 15150 4200 15178
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3528 14550 3556 14962
rect 3516 14544 3568 14550
rect 3516 14486 3568 14492
rect 3528 14006 3556 14486
rect 3700 14068 3752 14074
rect 3700 14010 3752 14016
rect 3516 14000 3568 14006
rect 3516 13942 3568 13948
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3620 12986 3648 13330
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 2870 12200 2926 12209
rect 2870 12135 2926 12144
rect 2688 12096 2740 12102
rect 2688 12038 2740 12044
rect 2778 12064 2834 12073
rect 2700 11098 2728 12038
rect 2778 11999 2834 12008
rect 2792 11354 2820 11999
rect 2884 11354 2912 12135
rect 3160 12102 3188 12242
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11898 3188 12038
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2700 11070 2820 11098
rect 2792 10996 2820 11070
rect 2594 10976 2650 10985
rect 2792 10968 3096 10996
rect 2594 10911 2650 10920
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2778 10296 2834 10305
rect 2410 10231 2466 10240
rect 2504 10260 2556 10266
rect 2424 10146 2452 10231
rect 2504 10202 2556 10208
rect 2596 10260 2648 10266
rect 2778 10231 2834 10240
rect 2872 10260 2924 10266
rect 2596 10202 2648 10208
rect 2608 10146 2636 10202
rect 2424 10118 2636 10146
rect 2424 9994 2452 10118
rect 2792 10033 2820 10231
rect 2872 10202 2924 10208
rect 2778 10024 2834 10033
rect 2412 9988 2464 9994
rect 2778 9959 2834 9968
rect 2412 9930 2464 9936
rect 2318 9752 2374 9761
rect 2318 9687 2374 9696
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2136 9512 2188 9518
rect 1950 9480 2006 9489
rect 2136 9454 2188 9460
rect 1950 9415 2006 9424
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 1964 8090 1992 9415
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2056 8430 2084 8910
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 2042 6760 2098 6769
rect 2042 6695 2098 6704
rect 2056 6458 2084 6695
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2056 6254 2084 6394
rect 2148 6338 2176 9454
rect 2240 9178 2268 9522
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2226 7440 2282 7449
rect 2332 7410 2360 9687
rect 2502 9480 2558 9489
rect 2778 9480 2834 9489
rect 2502 9415 2504 9424
rect 2556 9415 2558 9424
rect 2700 9438 2778 9466
rect 2504 9386 2556 9392
rect 2700 9178 2728 9438
rect 2778 9415 2834 9424
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2596 9104 2648 9110
rect 2596 9046 2648 9052
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2410 8120 2466 8129
rect 2410 8055 2412 8064
rect 2464 8055 2466 8064
rect 2412 8026 2464 8032
rect 2424 7478 2452 8026
rect 2412 7472 2464 7478
rect 2412 7414 2464 7420
rect 2226 7375 2282 7384
rect 2320 7404 2372 7410
rect 2240 6458 2268 7375
rect 2320 7346 2372 7352
rect 2332 6934 2360 7346
rect 2410 7304 2466 7313
rect 2410 7239 2412 7248
rect 2464 7239 2466 7248
rect 2412 7210 2464 7216
rect 2424 7002 2452 7210
rect 2412 6996 2464 7002
rect 2412 6938 2464 6944
rect 2320 6928 2372 6934
rect 2516 6882 2544 8978
rect 2608 8566 2636 9046
rect 2686 8936 2742 8945
rect 2686 8871 2742 8880
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2700 8242 2728 8871
rect 2884 8548 2912 10202
rect 2976 10062 3004 10474
rect 3068 10130 3096 10968
rect 3344 10606 3372 11630
rect 3528 11354 3556 12174
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3528 11150 3556 11290
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2964 10056 3016 10062
rect 3068 10033 3096 10066
rect 2964 9998 3016 10004
rect 3054 10024 3110 10033
rect 3054 9959 3110 9968
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9586 3096 9862
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2964 9444 3016 9450
rect 2964 9386 3016 9392
rect 2976 8974 3004 9386
rect 3068 9382 3096 9522
rect 3160 9518 3188 10202
rect 3238 9616 3294 9625
rect 3344 9586 3372 10542
rect 3712 10266 3740 14010
rect 4080 13818 4108 15030
rect 4172 14278 4200 15150
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 13938 4200 14214
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 4080 13790 4200 13818
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13433 3832 13670
rect 3790 13424 3846 13433
rect 3790 13359 3846 13368
rect 4172 13326 4200 13790
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4158 13152 4214 13161
rect 4158 13087 4214 13096
rect 3974 12880 4030 12889
rect 3974 12815 3976 12824
rect 4028 12815 4030 12824
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3882 12744 3884 12753
rect 3936 12744 3938 12753
rect 3882 12679 3938 12688
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3988 12481 4016 12582
rect 3974 12472 4030 12481
rect 4172 12442 4200 13087
rect 4264 12850 4292 15422
rect 4342 15328 4398 15337
rect 4342 15263 4398 15272
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 3974 12407 4030 12416
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4158 12200 4214 12209
rect 4158 12135 4160 12144
rect 4212 12135 4214 12144
rect 4160 12106 4212 12112
rect 3790 11928 3846 11937
rect 3790 11863 3846 11872
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3620 9602 3648 9862
rect 3238 9551 3294 9560
rect 3332 9580 3384 9586
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3146 9072 3202 9081
rect 3146 9007 3202 9016
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2884 8520 3004 8548
rect 2700 8214 2820 8242
rect 2792 8090 2820 8214
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2976 8022 3004 8520
rect 3160 8378 3188 9007
rect 3252 8634 3280 9551
rect 3620 9574 3740 9602
rect 3332 9522 3384 9528
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3330 8528 3386 8537
rect 3330 8463 3332 8472
rect 3384 8463 3386 8472
rect 3332 8434 3384 8440
rect 3344 8378 3372 8434
rect 3160 8362 3372 8378
rect 3148 8356 3372 8362
rect 3200 8350 3372 8356
rect 3148 8298 3200 8304
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3252 8090 3280 8230
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2608 7206 2636 7754
rect 3146 7576 3202 7585
rect 3146 7511 3148 7520
rect 3200 7511 3202 7520
rect 3148 7482 3200 7488
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2320 6870 2372 6876
rect 2424 6854 2544 6882
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2148 6310 2268 6338
rect 2332 6322 2360 6598
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 1768 5908 1820 5914
rect 1768 5850 1820 5856
rect 1490 5808 1546 5817
rect 1490 5743 1546 5752
rect 1504 3777 1532 5743
rect 2136 5568 2188 5574
rect 2136 5510 2188 5516
rect 1950 5128 2006 5137
rect 1950 5063 2006 5072
rect 1964 4826 1992 5063
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1582 4584 1638 4593
rect 1582 4519 1584 4528
rect 1636 4519 1638 4528
rect 1584 4490 1636 4496
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1676 4004 1728 4010
rect 1490 3768 1546 3777
rect 1596 3738 1624 3975
rect 1676 3946 1728 3952
rect 1490 3703 1546 3712
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1400 3596 1452 3602
rect 1400 3538 1452 3544
rect 662 3496 718 3505
rect 662 3431 718 3440
rect 202 1728 258 1737
rect 202 1663 258 1672
rect 216 480 244 1663
rect 676 480 704 3431
rect 1412 3097 1440 3538
rect 1688 3194 1716 3946
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1780 3777 1808 3878
rect 1766 3768 1822 3777
rect 1766 3703 1822 3712
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1398 3088 1454 3097
rect 1398 3023 1454 3032
rect 1950 2952 2006 2961
rect 2148 2922 2176 5510
rect 1950 2887 2006 2896
rect 2136 2916 2188 2922
rect 1964 2854 1992 2887
rect 2136 2858 2188 2864
rect 1952 2848 2004 2854
rect 1214 2816 1270 2825
rect 1952 2790 2004 2796
rect 1214 2751 1270 2760
rect 1228 480 1256 2751
rect 2148 2650 2176 2858
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1768 2372 1820 2378
rect 1768 2314 1820 2320
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1596 2145 1624 2246
rect 1582 2136 1638 2145
rect 1582 2071 1638 2080
rect 1780 480 1808 2314
rect 1964 2310 1992 2450
rect 1952 2304 2004 2310
rect 1952 2246 2004 2252
rect 1964 1737 1992 2246
rect 1950 1728 2006 1737
rect 1950 1663 2006 1672
rect 2240 649 2268 6310
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5953 2360 6258
rect 2318 5944 2374 5953
rect 2318 5879 2374 5888
rect 2318 5808 2374 5817
rect 2318 5743 2320 5752
rect 2372 5743 2374 5752
rect 2320 5714 2372 5720
rect 2424 5030 2452 6854
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2412 5024 2464 5030
rect 2412 4966 2464 4972
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2332 3738 2360 4082
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2332 3058 2360 3674
rect 2424 3233 2452 4966
rect 2516 4010 2544 6598
rect 2608 6390 2636 7142
rect 3160 7002 3188 7482
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 2964 6792 3016 6798
rect 2870 6760 2926 6769
rect 2964 6734 3016 6740
rect 2870 6695 2926 6704
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2608 5681 2636 6190
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5817 2728 6054
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2686 5808 2742 5817
rect 2686 5743 2742 5752
rect 2594 5672 2650 5681
rect 2792 5658 2820 5850
rect 2594 5607 2650 5616
rect 2700 5630 2820 5658
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2516 3738 2544 3946
rect 2608 3738 2636 5510
rect 2700 5098 2728 5630
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2688 5092 2740 5098
rect 2688 5034 2740 5040
rect 2792 4842 2820 5510
rect 2700 4826 2820 4842
rect 2884 4826 2912 6695
rect 2976 6390 3004 6734
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2976 5030 3004 5646
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2688 4820 2820 4826
rect 2740 4814 2820 4820
rect 2872 4820 2924 4826
rect 2688 4762 2740 4768
rect 2872 4762 2924 4768
rect 2700 4078 2728 4762
rect 2884 4282 2912 4762
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2410 3224 2466 3233
rect 2410 3159 2466 3168
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2412 2848 2464 2854
rect 2332 2808 2412 2836
rect 2226 640 2282 649
rect 2226 575 2282 584
rect 2332 480 2360 2808
rect 2412 2790 2464 2796
rect 2700 2666 2728 3878
rect 2792 2854 2820 4014
rect 3068 3534 3096 4558
rect 3056 3528 3108 3534
rect 3056 3470 3108 3476
rect 2870 3224 2926 3233
rect 3068 3194 3096 3470
rect 2870 3159 2926 3168
rect 3056 3188 3108 3194
rect 2884 2990 2912 3159
rect 3056 3130 3108 3136
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2700 2638 2912 2666
rect 2884 2310 2912 2638
rect 3068 2446 3096 3130
rect 3160 2582 3188 6666
rect 3252 6458 3280 7346
rect 3436 7274 3464 8570
rect 3528 8498 3556 8910
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 8022 3556 8434
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 3344 5370 3372 6054
rect 3436 5710 3464 6122
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 4826 3280 5034
rect 3240 4820 3292 4826
rect 3240 4762 3292 4768
rect 3344 4622 3372 5306
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3436 4486 3464 5646
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 4146 3464 4422
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3436 3534 3464 4082
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3528 3194 3556 7686
rect 3620 7342 3648 9415
rect 3712 7562 3740 9574
rect 3804 8090 3832 11863
rect 3976 11620 4028 11626
rect 3976 11562 4028 11568
rect 3882 11384 3938 11393
rect 3882 11319 3938 11328
rect 3896 10713 3924 11319
rect 3988 11014 4016 11562
rect 4068 11144 4120 11150
rect 4120 11092 4200 11098
rect 4068 11086 4200 11092
rect 4080 11070 4200 11086
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 4066 10976 4122 10985
rect 3882 10704 3938 10713
rect 3882 10639 3938 10648
rect 3896 10198 3924 10639
rect 3988 10470 4016 10950
rect 4066 10911 4122 10920
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3712 7534 3832 7562
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3606 6080 3662 6089
rect 3606 6015 3662 6024
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 480 2912 2246
rect 3160 1601 3188 2518
rect 3146 1592 3202 1601
rect 3146 1527 3202 1536
rect 3424 1488 3476 1494
rect 3424 1430 3476 1436
rect 3436 480 3464 1430
rect 3620 513 3648 6015
rect 3698 5672 3754 5681
rect 3698 5607 3754 5616
rect 3712 921 3740 5607
rect 3804 5166 3832 7534
rect 3792 5160 3844 5166
rect 3792 5102 3844 5108
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4758 3832 4966
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3804 4486 3832 4694
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4214 3832 4422
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3896 4010 3924 8774
rect 3988 7886 4016 10406
rect 4080 8650 4108 10911
rect 4172 10062 4200 11070
rect 4250 10840 4306 10849
rect 4250 10775 4306 10784
rect 4264 10470 4292 10775
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4356 10266 4384 15263
rect 4448 12209 4476 22358
rect 4540 21729 4568 23258
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4526 21720 4582 21729
rect 4526 21655 4582 21664
rect 4540 21146 4568 21655
rect 4632 21350 4660 21966
rect 4620 21344 4672 21350
rect 4620 21286 4672 21292
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4632 20398 4660 21286
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4528 20256 4580 20262
rect 4528 20198 4580 20204
rect 4540 19854 4568 20198
rect 4632 20058 4660 20334
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4540 19310 4568 19790
rect 4618 19408 4674 19417
rect 4618 19343 4674 19352
rect 4528 19304 4580 19310
rect 4528 19246 4580 19252
rect 4540 18970 4568 19246
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4540 18426 4568 18770
rect 4528 18420 4580 18426
rect 4528 18362 4580 18368
rect 4632 17082 4660 19343
rect 4724 17241 4752 26143
rect 4908 25702 4936 27520
rect 4896 25696 4948 25702
rect 4896 25638 4948 25644
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 5080 25220 5132 25226
rect 5080 25162 5132 25168
rect 4988 25152 5040 25158
rect 4988 25094 5040 25100
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4908 24290 4936 24754
rect 5000 24750 5028 25094
rect 4988 24744 5040 24750
rect 4988 24686 5040 24692
rect 5000 24410 5028 24686
rect 5092 24614 5120 25162
rect 5080 24608 5132 24614
rect 5080 24550 5132 24556
rect 4988 24404 5040 24410
rect 4988 24346 5040 24352
rect 4908 24262 5028 24290
rect 4894 22808 4950 22817
rect 4894 22743 4950 22752
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4816 19990 4844 21082
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4816 17649 4844 17682
rect 4802 17640 4858 17649
rect 4802 17575 4858 17584
rect 4710 17232 4766 17241
rect 4710 17167 4766 17176
rect 4632 17054 4844 17082
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 4632 15910 4660 16594
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4632 15570 4660 15846
rect 4620 15564 4672 15570
rect 4540 15524 4620 15552
rect 4540 14890 4568 15524
rect 4620 15506 4672 15512
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4724 14958 4752 15438
rect 4712 14952 4764 14958
rect 4710 14920 4712 14929
rect 4764 14920 4766 14929
rect 4528 14884 4580 14890
rect 4710 14855 4766 14864
rect 4528 14826 4580 14832
rect 4540 14618 4568 14826
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4712 14544 4764 14550
rect 4712 14486 4764 14492
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4434 12200 4490 12209
rect 4434 12135 4490 12144
rect 4434 11384 4490 11393
rect 4434 11319 4436 11328
rect 4488 11319 4490 11328
rect 4436 11290 4488 11296
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4448 10742 4476 11154
rect 4540 10810 4568 13262
rect 4632 11830 4660 13738
rect 4724 13530 4752 14486
rect 4712 13524 4764 13530
rect 4712 13466 4764 13472
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4724 12374 4752 13262
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4710 12200 4766 12209
rect 4710 12135 4766 12144
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4632 11218 4660 11494
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9450 4200 9998
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4356 9178 4384 10202
rect 4632 9761 4660 11154
rect 4724 10266 4752 12135
rect 4816 10606 4844 17054
rect 4908 14793 4936 22743
rect 5000 16454 5028 24262
rect 5092 23361 5120 24550
rect 5184 24274 5212 25230
rect 5264 25220 5316 25226
rect 5264 25162 5316 25168
rect 5172 24268 5224 24274
rect 5172 24210 5224 24216
rect 5170 24032 5226 24041
rect 5170 23967 5226 23976
rect 5078 23352 5134 23361
rect 5078 23287 5134 23296
rect 5080 22092 5132 22098
rect 5080 22034 5132 22040
rect 5092 21690 5120 22034
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5184 21593 5212 23967
rect 5276 22273 5304 25162
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5368 24342 5396 25094
rect 5356 24336 5408 24342
rect 5552 24313 5580 27520
rect 6104 25838 6132 27520
rect 6368 26172 6420 26178
rect 6368 26114 6420 26120
rect 6092 25832 6144 25838
rect 6092 25774 6144 25780
rect 6276 25424 6328 25430
rect 6276 25366 6328 25372
rect 5622 25052 5918 25072
rect 5678 25050 5702 25052
rect 5758 25050 5782 25052
rect 5838 25050 5862 25052
rect 5700 24998 5702 25050
rect 5764 24998 5776 25050
rect 5838 24998 5840 25050
rect 5678 24996 5702 24998
rect 5758 24996 5782 24998
rect 5838 24996 5862 24998
rect 5622 24976 5918 24996
rect 6000 24608 6052 24614
rect 6000 24550 6052 24556
rect 6012 24449 6040 24550
rect 5998 24440 6054 24449
rect 5998 24375 6054 24384
rect 5356 24278 5408 24284
rect 5538 24304 5594 24313
rect 5538 24239 5594 24248
rect 6184 24268 6236 24274
rect 5552 23730 5580 24239
rect 6184 24210 6236 24216
rect 5908 24200 5960 24206
rect 5906 24168 5908 24177
rect 5960 24168 5962 24177
rect 5906 24103 5962 24112
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5622 23964 5918 23984
rect 5678 23962 5702 23964
rect 5758 23962 5782 23964
rect 5838 23962 5862 23964
rect 5700 23910 5702 23962
rect 5764 23910 5776 23962
rect 5838 23910 5840 23962
rect 5678 23908 5702 23910
rect 5758 23908 5782 23910
rect 5838 23908 5862 23910
rect 5622 23888 5918 23908
rect 6012 23730 6040 24006
rect 6090 23896 6146 23905
rect 6196 23866 6224 24210
rect 6090 23831 6146 23840
rect 6184 23860 6236 23866
rect 5540 23724 5592 23730
rect 5540 23666 5592 23672
rect 6000 23724 6052 23730
rect 6000 23666 6052 23672
rect 5448 23248 5500 23254
rect 5448 23190 5500 23196
rect 5538 23216 5594 23225
rect 5460 22574 5488 23190
rect 6012 23186 6040 23666
rect 6104 23594 6132 23831
rect 6184 23802 6236 23808
rect 6092 23588 6144 23594
rect 6092 23530 6144 23536
rect 6288 23474 6316 25366
rect 6104 23446 6316 23474
rect 5538 23151 5594 23160
rect 6000 23180 6052 23186
rect 5552 22778 5580 23151
rect 6000 23122 6052 23128
rect 5622 22876 5918 22896
rect 5678 22874 5702 22876
rect 5758 22874 5782 22876
rect 5838 22874 5862 22876
rect 5700 22822 5702 22874
rect 5764 22822 5776 22874
rect 5838 22822 5840 22874
rect 5678 22820 5702 22822
rect 5758 22820 5782 22822
rect 5838 22820 5862 22822
rect 5622 22800 5918 22820
rect 5540 22772 5592 22778
rect 5540 22714 5592 22720
rect 6012 22642 6040 23122
rect 6000 22636 6052 22642
rect 5920 22596 6000 22624
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5262 22264 5318 22273
rect 5262 22199 5318 22208
rect 5460 21962 5488 22510
rect 5920 22234 5948 22596
rect 6000 22578 6052 22584
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 5908 22228 5960 22234
rect 5908 22170 5960 22176
rect 5448 21956 5500 21962
rect 5448 21898 5500 21904
rect 5622 21788 5918 21808
rect 5678 21786 5702 21788
rect 5758 21786 5782 21788
rect 5838 21786 5862 21788
rect 5700 21734 5702 21786
rect 5764 21734 5776 21786
rect 5838 21734 5840 21786
rect 5678 21732 5702 21734
rect 5758 21732 5782 21734
rect 5838 21732 5862 21734
rect 5622 21712 5918 21732
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5170 21584 5226 21593
rect 5170 21519 5226 21528
rect 5368 20942 5396 21626
rect 5540 21344 5592 21350
rect 5540 21286 5592 21292
rect 5356 20936 5408 20942
rect 5408 20896 5488 20924
rect 5356 20878 5408 20884
rect 5262 20768 5318 20777
rect 5262 20703 5318 20712
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5184 18290 5212 18702
rect 5172 18284 5224 18290
rect 5172 18226 5224 18232
rect 5172 18080 5224 18086
rect 5172 18022 5224 18028
rect 5078 17912 5134 17921
rect 5078 17847 5134 17856
rect 5092 17678 5120 17847
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5092 17338 5120 17614
rect 5080 17332 5132 17338
rect 5080 17274 5132 17280
rect 5078 17232 5134 17241
rect 5078 17167 5134 17176
rect 4988 16448 5040 16454
rect 4988 16390 5040 16396
rect 4986 16144 5042 16153
rect 4986 16079 5042 16088
rect 5000 15745 5028 16079
rect 4986 15736 5042 15745
rect 4986 15671 5042 15680
rect 4894 14784 4950 14793
rect 4894 14719 4950 14728
rect 4988 14000 5040 14006
rect 4894 13968 4950 13977
rect 4988 13942 5040 13948
rect 5092 13954 5120 17167
rect 5184 17105 5212 18022
rect 5170 17096 5226 17105
rect 5170 17031 5226 17040
rect 5276 16776 5304 20703
rect 5460 19972 5488 20896
rect 5552 20874 5580 21286
rect 5540 20868 5592 20874
rect 5540 20810 5592 20816
rect 5622 20700 5918 20720
rect 5678 20698 5702 20700
rect 5758 20698 5782 20700
rect 5838 20698 5862 20700
rect 5700 20646 5702 20698
rect 5764 20646 5776 20698
rect 5838 20646 5840 20698
rect 5678 20644 5702 20646
rect 5758 20644 5782 20646
rect 5838 20644 5862 20646
rect 5622 20624 5918 20644
rect 5724 20392 5776 20398
rect 5722 20360 5724 20369
rect 5776 20360 5778 20369
rect 5722 20295 5778 20304
rect 5540 19984 5592 19990
rect 5460 19944 5540 19972
rect 5540 19926 5592 19932
rect 5448 19712 5500 19718
rect 5500 19672 5580 19700
rect 5448 19654 5500 19660
rect 5552 18970 5580 19672
rect 5622 19612 5918 19632
rect 5678 19610 5702 19612
rect 5758 19610 5782 19612
rect 5838 19610 5862 19612
rect 5700 19558 5702 19610
rect 5764 19558 5776 19610
rect 5838 19558 5840 19610
rect 5678 19556 5702 19558
rect 5758 19556 5782 19558
rect 5838 19556 5862 19558
rect 5622 19536 5918 19556
rect 5632 19168 5684 19174
rect 5632 19110 5684 19116
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5644 18902 5672 19110
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 5644 18714 5672 18838
rect 5552 18686 5672 18714
rect 5552 18426 5580 18686
rect 5622 18524 5918 18544
rect 5678 18522 5702 18524
rect 5758 18522 5782 18524
rect 5838 18522 5862 18524
rect 5700 18470 5702 18522
rect 5764 18470 5776 18522
rect 5838 18470 5840 18522
rect 5678 18468 5702 18470
rect 5758 18468 5782 18470
rect 5838 18468 5862 18470
rect 5622 18448 5918 18468
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5538 18184 5594 18193
rect 5538 18119 5540 18128
rect 5592 18119 5594 18128
rect 5540 18090 5592 18096
rect 5552 18034 5580 18090
rect 5460 18006 5580 18034
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5460 17882 5488 18006
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5356 17808 5408 17814
rect 5644 17785 5672 18022
rect 5630 17776 5686 17785
rect 5356 17750 5408 17756
rect 5184 16748 5304 16776
rect 5184 14074 5212 16748
rect 5262 16688 5318 16697
rect 5262 16623 5318 16632
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4894 13903 4950 13912
rect 4908 13530 4936 13903
rect 5000 13841 5028 13942
rect 5092 13926 5212 13954
rect 4986 13832 5042 13841
rect 4986 13767 5042 13776
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4988 13456 5040 13462
rect 4908 13404 4988 13410
rect 5184 13410 5212 13926
rect 5276 13682 5304 16623
rect 5368 13802 5396 17750
rect 5460 17734 5630 17762
rect 5460 17338 5488 17734
rect 5630 17711 5686 17720
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5552 17202 5580 17546
rect 5622 17436 5918 17456
rect 5678 17434 5702 17436
rect 5758 17434 5782 17436
rect 5838 17434 5862 17436
rect 5700 17382 5702 17434
rect 5764 17382 5776 17434
rect 5838 17382 5840 17434
rect 5678 17380 5702 17382
rect 5758 17380 5782 17382
rect 5838 17380 5862 17382
rect 5622 17360 5918 17380
rect 5630 17232 5686 17241
rect 5540 17196 5592 17202
rect 5630 17167 5686 17176
rect 5540 17138 5592 17144
rect 5552 16794 5580 17138
rect 5644 17134 5672 17167
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5460 15638 5488 16390
rect 5552 16250 5580 16730
rect 5622 16348 5918 16368
rect 5678 16346 5702 16348
rect 5758 16346 5782 16348
rect 5838 16346 5862 16348
rect 5700 16294 5702 16346
rect 5764 16294 5776 16346
rect 5838 16294 5840 16346
rect 5678 16292 5702 16294
rect 5758 16292 5782 16294
rect 5838 16292 5862 16294
rect 5622 16272 5918 16292
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5632 16176 5684 16182
rect 5630 16144 5632 16153
rect 5684 16144 5686 16153
rect 5630 16079 5686 16088
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 15632 5500 15638
rect 5552 15609 5580 15846
rect 5448 15574 5500 15580
rect 5538 15600 5594 15609
rect 5460 15473 5488 15574
rect 5538 15535 5594 15544
rect 5446 15464 5502 15473
rect 5446 15399 5502 15408
rect 5446 15328 5502 15337
rect 5502 15286 5580 15314
rect 5446 15263 5502 15272
rect 5552 14906 5580 15286
rect 5622 15260 5918 15280
rect 5678 15258 5702 15260
rect 5758 15258 5782 15260
rect 5838 15258 5862 15260
rect 5700 15206 5702 15258
rect 5764 15206 5776 15258
rect 5838 15206 5840 15258
rect 5678 15204 5702 15206
rect 5758 15204 5782 15206
rect 5838 15204 5862 15206
rect 5622 15184 5918 15204
rect 5552 14878 5672 14906
rect 5540 14816 5592 14822
rect 5446 14784 5502 14793
rect 5540 14758 5592 14764
rect 5446 14719 5502 14728
rect 5460 13870 5488 14719
rect 5552 14550 5580 14758
rect 5540 14544 5592 14550
rect 5540 14486 5592 14492
rect 5644 14482 5672 14878
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5356 13796 5408 13802
rect 5356 13738 5408 13744
rect 5446 13696 5502 13705
rect 5276 13654 5396 13682
rect 4908 13398 5040 13404
rect 4908 13382 5028 13398
rect 5175 13382 5212 13410
rect 5264 13388 5316 13394
rect 4908 13025 4936 13382
rect 5175 13376 5203 13382
rect 5092 13348 5203 13376
rect 4894 13016 4950 13025
rect 4894 12951 4950 12960
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4908 12442 4936 12582
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 10266 4844 10542
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4618 9752 4674 9761
rect 4618 9687 4674 9696
rect 4724 9636 4752 10202
rect 4802 10160 4858 10169
rect 4802 10095 4858 10104
rect 4632 9608 4752 9636
rect 4632 9178 4660 9608
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4724 9058 4752 9318
rect 4816 9110 4844 10095
rect 4252 9036 4304 9042
rect 4252 8978 4304 8984
rect 4632 9030 4752 9058
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4080 8634 4200 8650
rect 4080 8628 4212 8634
rect 4080 8622 4160 8628
rect 4160 8570 4212 8576
rect 4066 8392 4122 8401
rect 4264 8362 4292 8978
rect 4528 8560 4580 8566
rect 4528 8502 4580 8508
rect 4066 8327 4122 8336
rect 4252 8356 4304 8362
rect 4080 7954 4108 8327
rect 4252 8298 4304 8304
rect 4342 7984 4398 7993
rect 4068 7948 4120 7954
rect 4342 7919 4398 7928
rect 4068 7890 4120 7896
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 4356 7041 4384 7919
rect 4540 7041 4568 8502
rect 4632 7410 4660 9030
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 7954 4752 8434
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4724 7410 4752 7890
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4342 7032 4398 7041
rect 4342 6967 4398 6976
rect 4526 7032 4582 7041
rect 4526 6967 4582 6976
rect 3974 6896 4030 6905
rect 4540 6866 4568 6967
rect 3974 6831 4030 6840
rect 4068 6860 4120 6866
rect 3988 4690 4016 6831
rect 4068 6802 4120 6808
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4080 6662 4108 6802
rect 4632 6798 4660 7346
rect 4712 7200 4764 7206
rect 4710 7168 4712 7177
rect 4764 7168 4766 7177
rect 4710 7103 4766 7112
rect 4724 7002 4752 7103
rect 4712 6996 4764 7002
rect 4712 6938 4764 6944
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4080 5681 4108 6598
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4356 5914 4384 6190
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4252 5704 4304 5710
rect 4066 5672 4122 5681
rect 4252 5646 4304 5652
rect 4066 5607 4122 5616
rect 4068 5160 4120 5166
rect 4068 5102 4120 5108
rect 3976 4684 4028 4690
rect 3976 4626 4028 4632
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 3896 3670 3924 3946
rect 3988 3738 4016 4626
rect 4080 4282 4108 5102
rect 4068 4276 4120 4282
rect 4068 4218 4120 4224
rect 4066 4176 4122 4185
rect 4066 4111 4122 4120
rect 4080 4078 4108 4111
rect 4264 4078 4292 5646
rect 4712 5160 4764 5166
rect 4710 5128 4712 5137
rect 4764 5128 4766 5137
rect 4710 5063 4766 5072
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4356 4282 4384 4422
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4816 4010 4844 9046
rect 4908 9024 4936 11766
rect 5000 9489 5028 12786
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 5092 9178 5120 13348
rect 5264 13330 5316 13336
rect 5276 13297 5304 13330
rect 5262 13288 5318 13297
rect 5262 13223 5318 13232
rect 5368 13138 5396 13654
rect 5446 13631 5502 13640
rect 5460 13326 5488 13631
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5276 13110 5396 13138
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5184 12073 5212 12786
rect 5170 12064 5226 12073
rect 5170 11999 5226 12008
rect 5170 11248 5226 11257
rect 5170 11183 5226 11192
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 4908 8996 5028 9024
rect 4894 8936 4950 8945
rect 4894 8871 4950 8880
rect 4908 8430 4936 8871
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 8090 4936 8366
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 5000 7274 5028 8996
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 5092 5370 5120 9114
rect 5184 7546 5212 11183
rect 5276 10810 5304 13110
rect 5460 12918 5488 13262
rect 5448 12912 5500 12918
rect 5552 12900 5580 14214
rect 5622 14172 5918 14192
rect 5678 14170 5702 14172
rect 5758 14170 5782 14172
rect 5838 14170 5862 14172
rect 5700 14118 5702 14170
rect 5764 14118 5776 14170
rect 5838 14118 5840 14170
rect 5678 14116 5702 14118
rect 5758 14116 5782 14118
rect 5838 14116 5862 14118
rect 5622 14096 5918 14116
rect 6012 13394 6040 22374
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 5622 13084 5918 13104
rect 5678 13082 5702 13084
rect 5758 13082 5782 13084
rect 5838 13082 5862 13084
rect 5700 13030 5702 13082
rect 5764 13030 5776 13082
rect 5838 13030 5840 13082
rect 5678 13028 5702 13030
rect 5758 13028 5782 13030
rect 5838 13028 5862 13030
rect 5622 13008 5918 13028
rect 5552 12872 5672 12900
rect 5448 12854 5500 12860
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5368 12102 5396 12582
rect 5460 12374 5488 12650
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5644 12306 5672 12872
rect 6012 12850 6040 13126
rect 6000 12844 6052 12850
rect 6000 12786 6052 12792
rect 5816 12708 5868 12714
rect 5816 12650 5868 12656
rect 5632 12300 5684 12306
rect 5632 12242 5684 12248
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5368 11914 5396 12038
rect 5368 11886 5488 11914
rect 5460 11257 5488 11886
rect 5446 11248 5502 11257
rect 5356 11212 5408 11218
rect 5446 11183 5502 11192
rect 5356 11154 5408 11160
rect 5368 10810 5396 11154
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5262 9208 5318 9217
rect 5262 9143 5318 9152
rect 5276 9110 5304 9143
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 5264 8832 5316 8838
rect 5262 8800 5264 8809
rect 5316 8800 5318 8809
rect 5262 8735 5318 8744
rect 5356 8424 5408 8430
rect 5356 8366 5408 8372
rect 5368 7954 5396 8366
rect 5460 8362 5488 10950
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5356 7948 5408 7954
rect 5408 7908 5488 7936
rect 5356 7890 5408 7896
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5184 7342 5212 7482
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5460 7274 5488 7908
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 6225 5212 6598
rect 5170 6216 5226 6225
rect 5170 6151 5226 6160
rect 5354 6216 5410 6225
rect 5460 6186 5488 7210
rect 5354 6151 5410 6160
rect 5448 6180 5500 6186
rect 5172 6112 5224 6118
rect 5172 6054 5224 6060
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5184 5914 5212 6054
rect 5276 5914 5304 6054
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5184 4826 5212 5850
rect 5172 4820 5224 4826
rect 5224 4780 5304 4808
rect 5172 4762 5224 4768
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 5092 3738 5120 4014
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 3884 3664 3936 3670
rect 4988 3664 5040 3670
rect 3884 3606 3936 3612
rect 4526 3632 4582 3641
rect 3976 3596 4028 3602
rect 4988 3606 5040 3612
rect 4526 3567 4528 3576
rect 3976 3538 4028 3544
rect 4580 3567 4582 3576
rect 4528 3538 4580 3544
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3804 2650 3832 3130
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3896 2650 3924 2790
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3698 912 3754 921
rect 3698 847 3754 856
rect 3606 504 3662 513
rect 202 0 258 480
rect 662 0 718 480
rect 1214 0 1270 480
rect 1766 0 1822 480
rect 2318 0 2374 480
rect 2870 0 2926 480
rect 3422 0 3478 480
rect 3988 480 4016 3538
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4080 3058 4108 3470
rect 4540 3126 4568 3538
rect 5000 3505 5028 3606
rect 4986 3496 5042 3505
rect 4986 3431 5042 3440
rect 5000 3126 5028 3431
rect 5184 3233 5212 4082
rect 5170 3224 5226 3233
rect 5170 3159 5226 3168
rect 5184 3126 5212 3159
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4068 2848 4120 2854
rect 4066 2816 4068 2825
rect 4436 2848 4488 2854
rect 4120 2816 4122 2825
rect 4436 2790 4488 2796
rect 4066 2751 4122 2760
rect 4448 2514 4476 2790
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4448 1306 4476 2450
rect 4540 1494 4568 3062
rect 5276 3058 5304 4780
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5368 2990 5396 6151
rect 5448 6122 5500 6128
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 5234 5488 5646
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5460 3534 5488 4082
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 4802 2680 4858 2689
rect 4802 2615 4804 2624
rect 4856 2615 4858 2624
rect 4804 2586 4856 2592
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4528 1488 4580 1494
rect 4528 1430 4580 1436
rect 4448 1278 4568 1306
rect 4540 480 4568 1278
rect 5092 480 5120 2450
rect 5552 1442 5580 12174
rect 5828 12170 5856 12650
rect 6000 12640 6052 12646
rect 6000 12582 6052 12588
rect 5816 12164 5868 12170
rect 5816 12106 5868 12112
rect 5622 11996 5918 12016
rect 5678 11994 5702 11996
rect 5758 11994 5782 11996
rect 5838 11994 5862 11996
rect 5700 11942 5702 11994
rect 5764 11942 5776 11994
rect 5838 11942 5840 11994
rect 5678 11940 5702 11942
rect 5758 11940 5782 11942
rect 5838 11940 5862 11942
rect 5622 11920 5918 11940
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5644 11286 5672 11630
rect 5632 11280 5684 11286
rect 5632 11222 5684 11228
rect 5622 10908 5918 10928
rect 5678 10906 5702 10908
rect 5758 10906 5782 10908
rect 5838 10906 5862 10908
rect 5700 10854 5702 10906
rect 5764 10854 5776 10906
rect 5838 10854 5840 10906
rect 5678 10852 5702 10854
rect 5758 10852 5782 10854
rect 5838 10852 5862 10854
rect 5622 10832 5918 10852
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 10266 5764 10610
rect 5814 10568 5870 10577
rect 5814 10503 5870 10512
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5828 9994 5856 10503
rect 5906 10432 5962 10441
rect 5906 10367 5962 10376
rect 5920 10266 5948 10367
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5622 9820 5918 9840
rect 5678 9818 5702 9820
rect 5758 9818 5782 9820
rect 5838 9818 5862 9820
rect 5700 9766 5702 9818
rect 5764 9766 5776 9818
rect 5838 9766 5840 9818
rect 5678 9764 5702 9766
rect 5758 9764 5782 9766
rect 5838 9764 5862 9766
rect 5622 9744 5918 9764
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 8906 5948 9318
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5622 8732 5918 8752
rect 5678 8730 5702 8732
rect 5758 8730 5782 8732
rect 5838 8730 5862 8732
rect 5700 8678 5702 8730
rect 5764 8678 5776 8730
rect 5838 8678 5840 8730
rect 5678 8676 5702 8678
rect 5758 8676 5782 8678
rect 5838 8676 5862 8678
rect 5622 8656 5918 8676
rect 5622 7644 5918 7664
rect 5678 7642 5702 7644
rect 5758 7642 5782 7644
rect 5838 7642 5862 7644
rect 5700 7590 5702 7642
rect 5764 7590 5776 7642
rect 5838 7590 5840 7642
rect 5678 7588 5702 7590
rect 5758 7588 5782 7590
rect 5838 7588 5862 7590
rect 5622 7568 5918 7588
rect 5814 6896 5870 6905
rect 5814 6831 5816 6840
rect 5868 6831 5870 6840
rect 5816 6802 5868 6808
rect 6012 6798 6040 12582
rect 6000 6792 6052 6798
rect 5630 6760 5686 6769
rect 6000 6734 6052 6740
rect 5630 6695 5632 6704
rect 5684 6695 5686 6704
rect 5632 6666 5684 6672
rect 5622 6556 5918 6576
rect 5678 6554 5702 6556
rect 5758 6554 5782 6556
rect 5838 6554 5862 6556
rect 5700 6502 5702 6554
rect 5764 6502 5776 6554
rect 5838 6502 5840 6554
rect 5678 6500 5702 6502
rect 5758 6500 5782 6502
rect 5838 6500 5862 6502
rect 5622 6480 5918 6500
rect 6012 6458 6040 6734
rect 6104 6730 6132 23446
rect 6380 23338 6408 26114
rect 6656 25378 6684 27520
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 6656 25350 6776 25378
rect 6458 25120 6514 25129
rect 6458 25055 6514 25064
rect 6196 23310 6408 23338
rect 6196 12918 6224 23310
rect 6366 22536 6422 22545
rect 6366 22471 6422 22480
rect 6380 22250 6408 22471
rect 6288 22222 6408 22250
rect 6288 21434 6316 22222
rect 6366 22128 6422 22137
rect 6366 22063 6368 22072
rect 6420 22063 6422 22072
rect 6368 22034 6420 22040
rect 6472 21536 6500 25055
rect 6644 24948 6696 24954
rect 6644 24890 6696 24896
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6564 23866 6592 24142
rect 6552 23860 6604 23866
rect 6552 23802 6604 23808
rect 6656 22234 6684 24890
rect 6748 24177 6776 25350
rect 6734 24168 6790 24177
rect 6734 24103 6790 24112
rect 6736 22500 6788 22506
rect 6736 22442 6788 22448
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6748 22098 6776 22442
rect 6736 22092 6788 22098
rect 6736 22034 6788 22040
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6564 21690 6592 21966
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6552 21684 6604 21690
rect 6552 21626 6604 21632
rect 6472 21508 6776 21536
rect 6288 21406 6684 21434
rect 6368 21344 6420 21350
rect 6368 21286 6420 21292
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6380 21078 6408 21286
rect 6368 21072 6420 21078
rect 6368 21014 6420 21020
rect 6276 21004 6328 21010
rect 6276 20946 6328 20952
rect 6288 20602 6316 20946
rect 6276 20596 6328 20602
rect 6276 20538 6328 20544
rect 6380 20398 6408 21014
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20602 6500 20878
rect 6564 20777 6592 21286
rect 6550 20768 6606 20777
rect 6550 20703 6606 20712
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6368 20392 6420 20398
rect 6368 20334 6420 20340
rect 6366 20088 6422 20097
rect 6366 20023 6422 20032
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6288 19378 6316 19858
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6288 18902 6316 19110
rect 6276 18896 6328 18902
rect 6276 18838 6328 18844
rect 6288 18426 6316 18838
rect 6276 18420 6328 18426
rect 6276 18362 6328 18368
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6288 17882 6316 18226
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6288 17066 6316 17818
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6380 16658 6408 20023
rect 6460 19984 6512 19990
rect 6460 19926 6512 19932
rect 6472 19514 6500 19926
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6472 18902 6500 19450
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6564 17814 6592 19858
rect 6656 18873 6684 21406
rect 6642 18864 6698 18873
rect 6642 18799 6698 18808
rect 6644 18080 6696 18086
rect 6644 18022 6696 18028
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6460 17536 6512 17542
rect 6458 17504 6460 17513
rect 6512 17504 6514 17513
rect 6458 17439 6514 17448
rect 6472 16833 6500 17439
rect 6564 17377 6592 17614
rect 6656 17542 6684 18022
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6550 17368 6606 17377
rect 6550 17303 6606 17312
rect 6564 16998 6592 17303
rect 6656 17134 6684 17478
rect 6644 17128 6696 17134
rect 6644 17070 6696 17076
rect 6552 16992 6604 16998
rect 6552 16934 6604 16940
rect 6458 16824 6514 16833
rect 6458 16759 6514 16768
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6276 16584 6328 16590
rect 6328 16532 6408 16538
rect 6276 16526 6408 16532
rect 6288 16510 6408 16526
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6288 15706 6316 16186
rect 6380 15910 6408 16510
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 6274 15328 6330 15337
rect 6274 15263 6330 15272
rect 6288 15162 6316 15263
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6274 14648 6330 14657
rect 6274 14583 6276 14592
rect 6328 14583 6330 14592
rect 6276 14554 6328 14560
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6288 13870 6316 14214
rect 6472 13920 6500 16594
rect 6564 16425 6592 16934
rect 6550 16416 6606 16425
rect 6550 16351 6606 16360
rect 6552 15904 6604 15910
rect 6656 15892 6684 17070
rect 6604 15864 6684 15892
rect 6552 15846 6604 15852
rect 6564 15570 6592 15846
rect 6552 15564 6604 15570
rect 6552 15506 6604 15512
rect 6564 14822 6592 15506
rect 6552 14816 6604 14822
rect 6748 14793 6776 21508
rect 6840 20641 6868 21830
rect 6932 20913 6960 25910
rect 7104 25152 7156 25158
rect 7104 25094 7156 25100
rect 7116 24750 7144 25094
rect 7300 24857 7328 27520
rect 7852 25498 7880 27520
rect 7840 25492 7892 25498
rect 7840 25434 7892 25440
rect 7378 25392 7434 25401
rect 7378 25327 7434 25336
rect 7286 24848 7342 24857
rect 7286 24783 7342 24792
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7286 24712 7342 24721
rect 7286 24647 7342 24656
rect 7300 24614 7328 24647
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 7196 24268 7248 24274
rect 7196 24210 7248 24216
rect 7012 23520 7064 23526
rect 7010 23488 7012 23497
rect 7064 23488 7066 23497
rect 7010 23423 7066 23432
rect 7208 23322 7236 24210
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7208 22438 7236 22918
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7104 22160 7156 22166
rect 7208 22137 7236 22374
rect 7104 22102 7156 22108
rect 7194 22128 7250 22137
rect 7012 22092 7064 22098
rect 7012 22034 7064 22040
rect 6918 20904 6974 20913
rect 6918 20839 6974 20848
rect 6826 20632 6882 20641
rect 6826 20567 6882 20576
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6826 20496 6882 20505
rect 6826 20431 6828 20440
rect 6880 20431 6882 20440
rect 6828 20402 6880 20408
rect 6932 20058 6960 20538
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6840 17898 6868 19790
rect 7024 19310 7052 22034
rect 7116 21486 7144 22102
rect 7194 22063 7250 22072
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7300 21146 7328 24006
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7196 20800 7248 20806
rect 7196 20742 7248 20748
rect 7102 20496 7158 20505
rect 7102 20431 7158 20440
rect 7116 19854 7144 20431
rect 7208 20097 7236 20742
rect 7194 20088 7250 20097
rect 7194 20023 7250 20032
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7024 18737 7052 19110
rect 7010 18728 7066 18737
rect 7010 18663 7066 18672
rect 7102 18456 7158 18465
rect 7102 18391 7158 18400
rect 6840 17870 7052 17898
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6932 17241 6960 17614
rect 6918 17232 6974 17241
rect 6918 17167 6974 17176
rect 6932 15162 6960 17167
rect 7024 16726 7052 17870
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7010 16008 7066 16017
rect 7010 15943 7066 15952
rect 7024 15910 7052 15943
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6552 14758 6604 14764
rect 6734 14784 6790 14793
rect 6380 13892 6500 13920
rect 6276 13864 6328 13870
rect 6276 13806 6328 13812
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6182 12744 6238 12753
rect 6288 12730 6316 13806
rect 6380 12889 6408 13892
rect 6564 13818 6592 14758
rect 6918 14784 6974 14793
rect 6734 14719 6790 14728
rect 6840 14742 6918 14770
rect 6840 14482 6868 14742
rect 6918 14719 6974 14728
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 7010 14376 7066 14385
rect 7010 14311 7012 14320
rect 7064 14311 7066 14320
rect 7012 14282 7064 14288
rect 6472 13802 6592 13818
rect 6460 13796 6592 13802
rect 6512 13790 6592 13796
rect 6460 13738 6512 13744
rect 6472 13326 6500 13738
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6564 13462 6592 13670
rect 6552 13456 6604 13462
rect 6604 13416 6684 13444
rect 6552 13398 6604 13404
rect 6460 13320 6512 13326
rect 6512 13280 6592 13308
rect 6460 13262 6512 13268
rect 6460 12912 6512 12918
rect 6366 12880 6422 12889
rect 6460 12854 6512 12860
rect 6366 12815 6422 12824
rect 6238 12702 6316 12730
rect 6182 12679 6238 12688
rect 6196 10198 6224 12679
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11898 6316 12174
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6472 11744 6500 12854
rect 6564 12646 6592 13280
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6288 11716 6500 11744
rect 6288 11014 6316 11716
rect 6564 11694 6592 12582
rect 6656 12374 6684 13416
rect 6828 12640 6880 12646
rect 7116 12628 7144 18391
rect 7392 18170 7420 25327
rect 7852 25242 7880 25434
rect 7760 25214 7880 25242
rect 8116 25288 8168 25294
rect 8116 25230 8168 25236
rect 8024 25220 8076 25226
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7470 23760 7526 23769
rect 7470 23695 7472 23704
rect 7524 23695 7526 23704
rect 7472 23666 7524 23672
rect 7576 22642 7604 24006
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7760 22522 7788 25214
rect 8024 25162 8076 25168
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7484 22494 7788 22522
rect 7484 19825 7512 22494
rect 7564 22092 7616 22098
rect 7564 22034 7616 22040
rect 7576 21894 7604 22034
rect 7564 21888 7616 21894
rect 7564 21830 7616 21836
rect 7576 21486 7604 21830
rect 7654 21720 7710 21729
rect 7654 21655 7656 21664
rect 7708 21655 7710 21664
rect 7656 21626 7708 21632
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7576 20244 7604 21422
rect 7656 20936 7708 20942
rect 7654 20904 7656 20913
rect 7748 20936 7800 20942
rect 7708 20904 7710 20913
rect 7748 20878 7800 20884
rect 7654 20839 7710 20848
rect 7760 20602 7788 20878
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7656 20256 7708 20262
rect 7576 20216 7656 20244
rect 7656 20198 7708 20204
rect 7470 19816 7526 19825
rect 7470 19751 7526 19760
rect 7668 19378 7696 20198
rect 7760 20058 7788 20402
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7472 19168 7524 19174
rect 7472 19110 7524 19116
rect 7484 18737 7512 19110
rect 7746 18864 7802 18873
rect 7656 18828 7708 18834
rect 7746 18799 7802 18808
rect 7656 18770 7708 18776
rect 7470 18728 7526 18737
rect 7470 18663 7526 18672
rect 7668 18222 7696 18770
rect 7656 18216 7708 18222
rect 7392 18142 7604 18170
rect 7656 18158 7708 18164
rect 7472 18080 7524 18086
rect 7470 18048 7472 18057
rect 7524 18048 7526 18057
rect 7470 17983 7526 17992
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7208 15706 7236 16390
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7208 14958 7236 15642
rect 7470 15464 7526 15473
rect 7470 15399 7526 15408
rect 7484 15026 7512 15399
rect 7472 15020 7524 15026
rect 7472 14962 7524 14968
rect 7196 14952 7248 14958
rect 7196 14894 7248 14900
rect 7380 14884 7432 14890
rect 7380 14826 7432 14832
rect 7196 12912 7248 12918
rect 7196 12854 7248 12860
rect 6828 12582 6880 12588
rect 6932 12600 7144 12628
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6656 12238 6684 12310
rect 6840 12306 6868 12582
rect 6828 12300 6880 12306
rect 6828 12242 6880 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6552 11688 6604 11694
rect 6458 11656 6514 11665
rect 6552 11630 6604 11636
rect 6458 11591 6514 11600
rect 6472 11354 6500 11591
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6458 11248 6514 11257
rect 6458 11183 6514 11192
rect 6368 11076 6420 11082
rect 6368 11018 6420 11024
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6274 10840 6330 10849
rect 6274 10775 6330 10784
rect 6288 10674 6316 10775
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6276 10532 6328 10538
rect 6276 10474 6328 10480
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6196 9722 6224 10134
rect 6184 9716 6236 9722
rect 6184 9658 6236 9664
rect 6288 9602 6316 10474
rect 6196 9574 6316 9602
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6000 6452 6052 6458
rect 6000 6394 6052 6400
rect 5908 6384 5960 6390
rect 5908 6326 5960 6332
rect 5920 5710 5948 6326
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5622 5468 5918 5488
rect 5678 5466 5702 5468
rect 5758 5466 5782 5468
rect 5838 5466 5862 5468
rect 5700 5414 5702 5466
rect 5764 5414 5776 5466
rect 5838 5414 5840 5466
rect 5678 5412 5702 5414
rect 5758 5412 5782 5414
rect 5838 5412 5862 5414
rect 5622 5392 5918 5412
rect 6104 5166 6132 6666
rect 6092 5160 6144 5166
rect 6092 5102 6144 5108
rect 6090 4856 6146 4865
rect 6090 4791 6146 4800
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5622 4380 5918 4400
rect 5678 4378 5702 4380
rect 5758 4378 5782 4380
rect 5838 4378 5862 4380
rect 5700 4326 5702 4378
rect 5764 4326 5776 4378
rect 5838 4326 5840 4378
rect 5678 4324 5702 4326
rect 5758 4324 5782 4326
rect 5838 4324 5862 4326
rect 5622 4304 5918 4324
rect 6012 4214 6040 4422
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5908 3596 5960 3602
rect 6012 3584 6040 3878
rect 5960 3556 6040 3584
rect 5908 3538 5960 3544
rect 5622 3292 5918 3312
rect 5678 3290 5702 3292
rect 5758 3290 5782 3292
rect 5838 3290 5862 3292
rect 5700 3238 5702 3290
rect 5764 3238 5776 3290
rect 5838 3238 5840 3290
rect 5678 3236 5702 3238
rect 5758 3236 5782 3238
rect 5838 3236 5862 3238
rect 5622 3216 5918 3236
rect 6012 2854 6040 3556
rect 6104 2990 6132 4791
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6196 2650 6224 9574
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6288 8401 6316 8774
rect 6274 8392 6330 8401
rect 6274 8327 6330 8336
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6288 7750 6316 8230
rect 6380 8022 6408 11018
rect 6472 9897 6500 11183
rect 6564 10810 6592 11290
rect 6552 10804 6604 10810
rect 6552 10746 6604 10752
rect 6550 10160 6606 10169
rect 6550 10095 6552 10104
rect 6604 10095 6606 10104
rect 6552 10066 6604 10072
rect 6656 10062 6684 12038
rect 6748 11665 6776 12106
rect 6734 11656 6790 11665
rect 6734 11591 6790 11600
rect 6840 11529 6868 12242
rect 6826 11520 6882 11529
rect 6826 11455 6882 11464
rect 6932 11370 6960 12600
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6748 11342 6960 11370
rect 6644 10056 6696 10062
rect 6642 10024 6644 10033
rect 6696 10024 6698 10033
rect 6642 9959 6698 9968
rect 6458 9888 6514 9897
rect 6458 9823 6514 9832
rect 6642 9752 6698 9761
rect 6460 9716 6512 9722
rect 6642 9687 6698 9696
rect 6460 9658 6512 9664
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6276 7744 6328 7750
rect 6276 7686 6328 7692
rect 6288 5953 6316 7686
rect 6380 7546 6408 7958
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6380 6730 6408 7482
rect 6368 6724 6420 6730
rect 6368 6666 6420 6672
rect 6380 6390 6408 6666
rect 6368 6384 6420 6390
rect 6368 6326 6420 6332
rect 6274 5944 6330 5953
rect 6274 5879 6276 5888
rect 6328 5879 6330 5888
rect 6276 5850 6328 5856
rect 6288 5234 6316 5850
rect 6368 5772 6420 5778
rect 6368 5714 6420 5720
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6380 5137 6408 5714
rect 6366 5128 6422 5137
rect 6366 5063 6422 5072
rect 6380 4185 6408 5063
rect 6366 4176 6422 4185
rect 6366 4111 6422 4120
rect 6472 3058 6500 9658
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8498 6592 8978
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6550 8392 6606 8401
rect 6550 8327 6606 8336
rect 6564 5846 6592 8327
rect 6552 5840 6604 5846
rect 6552 5782 6604 5788
rect 6656 5778 6684 9687
rect 6748 9625 6776 11342
rect 7024 11064 7052 12378
rect 7104 12232 7156 12238
rect 7102 12200 7104 12209
rect 7156 12200 7158 12209
rect 7102 12135 7158 12144
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 6932 11036 7052 11064
rect 6932 10690 6960 11036
rect 7010 10976 7066 10985
rect 7010 10911 7066 10920
rect 6840 10662 6960 10690
rect 6734 9616 6790 9625
rect 6734 9551 6790 9560
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6748 8362 6776 8978
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6840 7002 6868 10662
rect 7024 10146 7052 10911
rect 7116 10169 7144 12038
rect 7208 11626 7236 12854
rect 7288 12640 7340 12646
rect 7288 12582 7340 12588
rect 7300 12442 7328 12582
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7288 12300 7340 12306
rect 7288 12242 7340 12248
rect 7300 11937 7328 12242
rect 7286 11928 7342 11937
rect 7286 11863 7342 11872
rect 7196 11620 7248 11626
rect 7248 11580 7328 11608
rect 7196 11562 7248 11568
rect 7300 11354 7328 11580
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7196 11280 7248 11286
rect 7196 11222 7248 11228
rect 6932 10118 7052 10146
rect 7102 10160 7158 10169
rect 6932 9722 6960 10118
rect 7102 10095 7158 10104
rect 7208 10010 7236 11222
rect 7300 11150 7328 11290
rect 7288 11144 7340 11150
rect 7288 11086 7340 11092
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7024 9982 7236 10010
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 7024 9353 7052 9982
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7010 9344 7066 9353
rect 7010 9279 7066 9288
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6840 6458 6868 6938
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6734 6352 6790 6361
rect 6734 6287 6790 6296
rect 6748 5914 6776 6287
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 7024 5846 7052 9279
rect 7208 8634 7236 9522
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 8344 7328 10134
rect 7116 8316 7328 8344
rect 7116 8242 7144 8316
rect 7116 8214 7236 8242
rect 7208 8090 7236 8214
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7194 7984 7250 7993
rect 7194 7919 7250 7928
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6564 5166 6592 5646
rect 6932 5386 6960 5714
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6840 5370 6960 5386
rect 6828 5364 6960 5370
rect 6880 5358 6960 5364
rect 6828 5306 6880 5312
rect 7024 5234 7052 5510
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6564 5030 6592 5102
rect 6552 5024 6604 5030
rect 6552 4966 6604 4972
rect 6564 4622 6592 4966
rect 6642 4720 6698 4729
rect 6642 4655 6698 4664
rect 6828 4684 6880 4690
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6564 4078 6592 4558
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6656 3194 6684 4655
rect 6828 4626 6880 4632
rect 6736 4480 6788 4486
rect 6840 4457 6868 4626
rect 6736 4422 6788 4428
rect 6826 4448 6882 4457
rect 6748 4298 6776 4422
rect 6826 4383 6882 4392
rect 6932 4298 6960 5170
rect 6748 4270 6868 4298
rect 6932 4270 7052 4298
rect 6840 4128 6868 4270
rect 6840 4100 6960 4128
rect 6932 3738 6960 4100
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 7024 3534 7052 4270
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 6734 3360 6790 3369
rect 6734 3295 6790 3304
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2650 6592 2790
rect 6184 2644 6236 2650
rect 6184 2586 6236 2592
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6276 2304 6328 2310
rect 6274 2272 6276 2281
rect 6328 2272 6330 2281
rect 5622 2204 5918 2224
rect 6274 2207 6330 2216
rect 5678 2202 5702 2204
rect 5758 2202 5782 2204
rect 5838 2202 5862 2204
rect 5700 2150 5702 2202
rect 5764 2150 5776 2202
rect 5838 2150 5840 2202
rect 5678 2148 5702 2150
rect 5758 2148 5782 2150
rect 5838 2148 5862 2150
rect 5622 2128 5918 2148
rect 6550 1592 6606 1601
rect 6550 1527 6552 1536
rect 6604 1527 6606 1536
rect 6552 1498 6604 1504
rect 5552 1414 5672 1442
rect 5644 480 5672 1414
rect 6656 762 6684 2994
rect 6196 734 6684 762
rect 6196 480 6224 734
rect 6748 480 6776 3295
rect 7024 3058 7052 3470
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7208 2990 7236 7919
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7300 6458 7328 6802
rect 7288 6452 7340 6458
rect 7288 6394 7340 6400
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7300 3126 7328 5782
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7300 2922 7328 3062
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7392 2650 7420 14826
rect 7484 14618 7512 14962
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 7484 10742 7512 12242
rect 7576 11218 7604 18142
rect 7668 12374 7696 18158
rect 7760 14890 7788 18799
rect 7852 18290 7880 24618
rect 7944 18902 7972 25094
rect 8036 24954 8064 25162
rect 8024 24948 8076 24954
rect 8024 24890 8076 24896
rect 8128 24886 8156 25230
rect 8300 25220 8352 25226
rect 8300 25162 8352 25168
rect 8116 24880 8168 24886
rect 8116 24822 8168 24828
rect 8128 24614 8156 24822
rect 8312 24614 8340 25162
rect 8404 24834 8432 27520
rect 8944 25152 8996 25158
rect 8944 25094 8996 25100
rect 8404 24806 8708 24834
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8116 24608 8168 24614
rect 8300 24608 8352 24614
rect 8116 24550 8168 24556
rect 8220 24568 8300 24596
rect 8022 23080 8078 23089
rect 8022 23015 8024 23024
rect 8076 23015 8078 23024
rect 8024 22986 8076 22992
rect 8128 22506 8156 24550
rect 8116 22500 8168 22506
rect 8116 22442 8168 22448
rect 8220 21962 8248 24568
rect 8300 24550 8352 24556
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8312 22778 8340 23598
rect 8300 22772 8352 22778
rect 8300 22714 8352 22720
rect 8312 22166 8340 22714
rect 8300 22160 8352 22166
rect 8300 22102 8352 22108
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 8312 21418 8340 21898
rect 8300 21412 8352 21418
rect 8300 21354 8352 21360
rect 8024 21140 8076 21146
rect 8024 21082 8076 21088
rect 8036 20058 8064 21082
rect 8312 21010 8340 21354
rect 8404 21185 8432 24686
rect 8576 23520 8628 23526
rect 8576 23462 8628 23468
rect 8482 23352 8538 23361
rect 8482 23287 8538 23296
rect 8496 23118 8524 23287
rect 8588 23254 8616 23462
rect 8576 23248 8628 23254
rect 8576 23190 8628 23196
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8496 22273 8524 23054
rect 8482 22264 8538 22273
rect 8482 22199 8538 22208
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8390 21176 8446 21185
rect 8390 21111 8446 21120
rect 8300 21004 8352 21010
rect 8300 20946 8352 20952
rect 8496 20874 8524 21966
rect 8588 21729 8616 22102
rect 8574 21720 8630 21729
rect 8574 21655 8630 21664
rect 8574 21584 8630 21593
rect 8574 21519 8630 21528
rect 8484 20868 8536 20874
rect 8484 20810 8536 20816
rect 8588 20482 8616 21519
rect 8496 20454 8616 20482
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 8036 18970 8064 19790
rect 8312 19786 8340 20198
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 7944 18222 7972 18838
rect 8128 18630 8156 19178
rect 8312 18766 8340 19722
rect 8496 18970 8524 20454
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8300 18760 8352 18766
rect 8352 18720 8432 18748
rect 8300 18702 8352 18708
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 8128 18170 8156 18566
rect 8404 18358 8432 18720
rect 8392 18352 8444 18358
rect 8206 18320 8262 18329
rect 8392 18294 8444 18300
rect 8206 18255 8208 18264
rect 8260 18255 8262 18264
rect 8208 18226 8260 18232
rect 8128 18142 8248 18170
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7944 16794 7972 17002
rect 8036 16794 8064 17478
rect 8220 16998 8248 18142
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8208 16992 8260 16998
rect 8206 16960 8208 16969
rect 8260 16960 8262 16969
rect 8206 16895 8262 16904
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 8312 15994 8340 17682
rect 8404 17610 8432 18294
rect 8496 18290 8524 18906
rect 8588 18766 8616 20334
rect 8680 19689 8708 24806
rect 8956 24750 8984 25094
rect 8944 24744 8996 24750
rect 8944 24686 8996 24692
rect 9048 24041 9076 27520
rect 9128 26104 9180 26110
rect 9128 26046 9180 26052
rect 9034 24032 9090 24041
rect 9034 23967 9090 23976
rect 9036 23044 9088 23050
rect 9036 22986 9088 22992
rect 8758 22672 8814 22681
rect 8758 22607 8814 22616
rect 8772 19922 8800 22607
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8864 21690 8892 22442
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 9048 21146 9076 22986
rect 9140 22080 9168 26046
rect 9496 25968 9548 25974
rect 9494 25936 9496 25945
rect 9548 25936 9550 25945
rect 9494 25871 9550 25880
rect 9496 25832 9548 25838
rect 9494 25800 9496 25809
rect 9548 25800 9550 25809
rect 9494 25735 9550 25744
rect 9312 24064 9364 24070
rect 9312 24006 9364 24012
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9324 23594 9352 24006
rect 9508 23633 9536 24006
rect 9494 23624 9550 23633
rect 9312 23588 9364 23594
rect 9494 23559 9550 23568
rect 9312 23530 9364 23536
rect 9324 23118 9352 23530
rect 9494 23216 9550 23225
rect 9494 23151 9496 23160
rect 9548 23151 9550 23160
rect 9496 23122 9548 23128
rect 9312 23112 9364 23118
rect 9312 23054 9364 23060
rect 9324 22234 9352 23054
rect 9312 22228 9364 22234
rect 9312 22170 9364 22176
rect 9600 22114 9628 27520
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9876 24886 9904 25298
rect 10060 25226 10088 26182
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 9864 24880 9916 24886
rect 9678 24848 9734 24857
rect 10152 24857 10180 27520
rect 10796 25770 10824 27520
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 10968 25832 11020 25838
rect 10968 25774 11020 25780
rect 10784 25764 10836 25770
rect 10784 25706 10836 25712
rect 10289 25596 10585 25616
rect 10345 25594 10369 25596
rect 10425 25594 10449 25596
rect 10505 25594 10529 25596
rect 10367 25542 10369 25594
rect 10431 25542 10443 25594
rect 10505 25542 10507 25594
rect 10345 25540 10369 25542
rect 10425 25540 10449 25542
rect 10505 25540 10529 25542
rect 10289 25520 10585 25540
rect 10796 25344 10824 25706
rect 10874 25528 10930 25537
rect 10980 25498 11008 25774
rect 10874 25463 10930 25472
rect 10968 25492 11020 25498
rect 10704 25316 10824 25344
rect 9864 24822 9916 24828
rect 10138 24848 10194 24857
rect 9678 24783 9734 24792
rect 9956 24812 10008 24818
rect 9692 24410 9720 24783
rect 10138 24783 10194 24792
rect 9956 24754 10008 24760
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 9772 24608 9824 24614
rect 9772 24550 9824 24556
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23361 9720 23462
rect 9678 23352 9734 23361
rect 9784 23322 9812 24550
rect 9678 23287 9734 23296
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9678 22400 9734 22409
rect 9678 22335 9734 22344
rect 9508 22086 9628 22114
rect 9140 22052 9352 22080
rect 9126 21448 9182 21457
rect 9126 21383 9182 21392
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 8760 19916 8812 19922
rect 8760 19858 8812 19864
rect 9140 19802 9168 21383
rect 9218 20904 9274 20913
rect 9218 20839 9274 20848
rect 9048 19774 9168 19802
rect 8666 19680 8722 19689
rect 8666 19615 8722 19624
rect 8850 19680 8906 19689
rect 8850 19615 8906 19624
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18426 8616 18702
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8484 18284 8536 18290
rect 8484 18226 8536 18232
rect 8760 17808 8812 17814
rect 8760 17750 8812 17756
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8392 17604 8444 17610
rect 8392 17546 8444 17552
rect 8680 17338 8708 17614
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8680 16794 8708 17274
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8482 16688 8538 16697
rect 8482 16623 8484 16632
rect 8536 16623 8538 16632
rect 8484 16594 8536 16600
rect 8588 16046 8616 16730
rect 8666 16416 8722 16425
rect 8666 16351 8722 16360
rect 8680 16114 8708 16351
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8128 15966 8340 15994
rect 8392 16040 8444 16046
rect 8576 16040 8628 16046
rect 8392 15982 8444 15988
rect 8482 16008 8538 16017
rect 7838 15600 7894 15609
rect 7838 15535 7894 15544
rect 7748 14884 7800 14890
rect 7748 14826 7800 14832
rect 7852 14346 7880 15535
rect 8036 15473 8064 15914
rect 8128 15745 8156 15966
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 8114 15736 8170 15745
rect 8114 15671 8116 15680
rect 8168 15671 8170 15680
rect 8116 15642 8168 15648
rect 8128 15611 8156 15642
rect 8022 15464 8078 15473
rect 8022 15399 8024 15408
rect 8076 15399 8078 15408
rect 8024 15370 8076 15376
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 7930 14648 7986 14657
rect 7930 14583 7986 14592
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7746 13560 7802 13569
rect 7852 13530 7880 13806
rect 7746 13495 7802 13504
rect 7840 13524 7892 13530
rect 7760 12753 7788 13495
rect 7840 13466 7892 13472
rect 7746 12744 7802 12753
rect 7746 12679 7802 12688
rect 7656 12368 7708 12374
rect 7656 12310 7708 12316
rect 7838 12336 7894 12345
rect 7748 12300 7800 12306
rect 7838 12271 7894 12280
rect 7748 12242 7800 12248
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 11558 7696 12174
rect 7656 11552 7708 11558
rect 7656 11494 7708 11500
rect 7564 11212 7616 11218
rect 7564 11154 7616 11160
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7472 10736 7524 10742
rect 7472 10678 7524 10684
rect 7576 10554 7604 10950
rect 7484 10526 7604 10554
rect 7484 8809 7512 10526
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 9761 7604 10406
rect 7562 9752 7618 9761
rect 7562 9687 7618 9696
rect 7668 9586 7696 11494
rect 7760 11257 7788 12242
rect 7746 11248 7802 11257
rect 7746 11183 7802 11192
rect 7760 10266 7788 11183
rect 7852 11082 7880 12271
rect 7944 11286 7972 14583
rect 8036 14498 8064 14894
rect 8036 14470 8156 14498
rect 8022 13560 8078 13569
rect 8022 13495 8078 13504
rect 8036 12481 8064 13495
rect 8022 12472 8078 12481
rect 8128 12442 8156 14470
rect 8022 12407 8078 12416
rect 8116 12436 8168 12442
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7930 10976 7986 10985
rect 7930 10911 7986 10920
rect 7838 10704 7894 10713
rect 7838 10639 7894 10648
rect 7852 10538 7880 10639
rect 7944 10606 7972 10911
rect 7932 10600 7984 10606
rect 7932 10542 7984 10548
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7852 10198 7880 10474
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7840 10192 7892 10198
rect 7840 10134 7892 10140
rect 7944 9586 7972 10202
rect 8036 9654 8064 12407
rect 8116 12378 8168 12384
rect 8220 12288 8248 15846
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8312 15026 8340 15370
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8404 14482 8432 15982
rect 8576 15982 8628 15988
rect 8482 15943 8538 15952
rect 8496 15570 8524 15943
rect 8680 15638 8708 16050
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8496 15162 8524 15506
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8588 14890 8616 15302
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8392 14476 8444 14482
rect 8392 14418 8444 14424
rect 8298 13832 8354 13841
rect 8298 13767 8354 13776
rect 8312 13138 8340 13767
rect 8404 13258 8432 14418
rect 8588 14006 8616 14826
rect 8772 14498 8800 17750
rect 8864 15706 8892 19615
rect 8942 19544 8998 19553
rect 8942 19479 8998 19488
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8864 15201 8892 15642
rect 8850 15192 8906 15201
rect 8850 15127 8852 15136
rect 8904 15127 8906 15136
rect 8852 15098 8904 15104
rect 8864 15067 8892 15098
rect 8772 14470 8892 14498
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8666 13968 8722 13977
rect 8588 13705 8616 13942
rect 8666 13903 8722 13912
rect 8574 13696 8630 13705
rect 8574 13631 8630 13640
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8312 13110 8616 13138
rect 8390 13016 8446 13025
rect 8390 12951 8392 12960
rect 8444 12951 8446 12960
rect 8484 12980 8536 12986
rect 8392 12922 8444 12928
rect 8484 12922 8536 12928
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8128 12260 8248 12288
rect 8128 11393 8156 12260
rect 8206 12200 8262 12209
rect 8206 12135 8262 12144
rect 8114 11384 8170 11393
rect 8220 11354 8248 12135
rect 8114 11319 8170 11328
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11234 8340 12310
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8220 11206 8340 11234
rect 8128 10538 8156 11154
rect 8220 11014 8248 11206
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8208 11008 8260 11014
rect 8208 10950 8260 10956
rect 8208 10736 8260 10742
rect 8260 10684 8340 10690
rect 8208 10678 8340 10684
rect 8220 10662 8340 10678
rect 8116 10532 8168 10538
rect 8116 10474 8168 10480
rect 8114 10296 8170 10305
rect 8114 10231 8116 10240
rect 8168 10231 8170 10240
rect 8116 10202 8168 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 8024 9648 8076 9654
rect 8024 9590 8076 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7470 8800 7526 8809
rect 7470 8735 7526 8744
rect 7484 8401 7512 8735
rect 7668 8498 7696 9318
rect 8128 9178 8156 9930
rect 8220 9722 8248 9998
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9172 8168 9178
rect 8116 9114 8168 9120
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7656 8492 7708 8498
rect 7656 8434 7708 8440
rect 7470 8392 7526 8401
rect 7760 8362 7788 8774
rect 8220 8401 8248 9658
rect 8312 9110 8340 10662
rect 8404 10062 8432 11086
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8206 8392 8262 8401
rect 7470 8327 7526 8336
rect 7748 8356 7800 8362
rect 8206 8327 8262 8336
rect 7748 8298 7800 8304
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 7206 7512 7822
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 5001 7512 7142
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7576 2530 7604 8026
rect 7760 8022 7788 8298
rect 7748 8016 7800 8022
rect 7746 7984 7748 7993
rect 7800 7984 7802 7993
rect 7746 7919 7802 7928
rect 8404 7818 8432 9862
rect 8496 8820 8524 12922
rect 8588 12442 8616 13110
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8588 9382 8616 11494
rect 8680 9518 8708 13903
rect 8772 13530 8800 14350
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 8758 13424 8814 13433
rect 8758 13359 8814 13368
rect 8772 11898 8800 13359
rect 8864 12986 8892 14470
rect 8956 13818 8984 19479
rect 9048 17814 9076 19774
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9140 18222 9168 19654
rect 9232 18426 9260 20839
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9036 17672 9088 17678
rect 9036 17614 9088 17620
rect 9048 16658 9076 17614
rect 9218 16688 9274 16697
rect 9036 16652 9088 16658
rect 9218 16623 9274 16632
rect 9036 16594 9088 16600
rect 9232 16114 9260 16623
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 9048 14278 9076 14826
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9036 14272 9088 14278
rect 9232 14249 9260 14282
rect 9036 14214 9088 14220
rect 9218 14240 9274 14249
rect 9048 13938 9076 14214
rect 9218 14175 9274 14184
rect 9232 14074 9260 14175
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9036 13932 9088 13938
rect 9036 13874 9088 13880
rect 8956 13790 9168 13818
rect 9036 13252 9088 13258
rect 9036 13194 9088 13200
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8864 12345 8892 12582
rect 8850 12336 8906 12345
rect 8850 12271 8906 12280
rect 8956 12238 8984 12786
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8850 12064 8906 12073
rect 8850 11999 8906 12008
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8758 11656 8814 11665
rect 8758 11591 8814 11600
rect 8772 10266 8800 11591
rect 8864 10577 8892 11999
rect 9048 10690 9076 13194
rect 9140 10826 9168 13790
rect 9220 12640 9272 12646
rect 9218 12608 9220 12617
rect 9272 12608 9274 12617
rect 9218 12543 9274 12552
rect 9140 10798 9260 10826
rect 9048 10662 9168 10690
rect 8944 10600 8996 10606
rect 8850 10568 8906 10577
rect 8944 10542 8996 10548
rect 8850 10503 8906 10512
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8864 9926 8892 10406
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8668 9512 8720 9518
rect 8668 9454 8720 9460
rect 8576 9376 8628 9382
rect 8576 9318 8628 9324
rect 8496 8792 8800 8820
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8392 7812 8444 7818
rect 8392 7754 8444 7760
rect 7654 7576 7710 7585
rect 7654 7511 7656 7520
rect 7708 7511 7710 7520
rect 7656 7482 7708 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 6866 8064 7346
rect 8128 7206 8156 7754
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8024 6860 8076 6866
rect 8024 6802 8076 6808
rect 8128 6769 8156 7142
rect 8220 6882 8248 7686
rect 8392 6928 8444 6934
rect 8220 6854 8340 6882
rect 8392 6870 8444 6876
rect 8312 6798 8340 6854
rect 8300 6792 8352 6798
rect 8114 6760 8170 6769
rect 8300 6734 8352 6740
rect 8114 6695 8170 6704
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 8036 6497 8064 6598
rect 8022 6488 8078 6497
rect 8022 6423 8078 6432
rect 8220 6186 8248 6666
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8220 5914 8248 6122
rect 8312 5914 8340 6734
rect 8404 6361 8432 6870
rect 8390 6352 8446 6361
rect 8390 6287 8446 6296
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8220 5817 8248 5850
rect 8206 5808 8262 5817
rect 8206 5743 8262 5752
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8220 5545 8248 5646
rect 8206 5536 8262 5545
rect 8206 5471 8262 5480
rect 8114 5128 8170 5137
rect 8114 5063 8116 5072
rect 8168 5063 8170 5072
rect 8116 5034 8168 5040
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 4010 7972 4422
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7838 3496 7894 3505
rect 7838 3431 7840 3440
rect 7892 3431 7894 3440
rect 7840 3402 7892 3408
rect 7852 3108 7880 3402
rect 7852 3080 7972 3108
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7300 2502 7604 2530
rect 6918 1592 6974 1601
rect 6918 1527 6974 1536
rect 3606 439 3662 448
rect 3974 0 4030 480
rect 4526 0 4582 480
rect 5078 0 5134 480
rect 5630 0 5686 480
rect 6182 0 6238 480
rect 6734 0 6790 480
rect 6932 377 6960 1527
rect 7300 480 7328 2502
rect 7852 480 7880 2586
rect 7944 2582 7972 3080
rect 7932 2576 7984 2582
rect 7932 2518 7984 2524
rect 8036 513 8064 4966
rect 8220 3942 8248 5471
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 8312 5030 8340 5306
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8496 4468 8524 8599
rect 8666 8528 8722 8537
rect 8666 8463 8722 8472
rect 8680 7954 8708 8463
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 7478 8616 7822
rect 8680 7546 8708 7890
rect 8668 7540 8720 7546
rect 8668 7482 8720 7488
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8588 7002 8616 7414
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8680 6798 8708 6831
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8772 6118 8800 8792
rect 8864 8537 8892 9522
rect 8850 8528 8906 8537
rect 8850 8463 8906 8472
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8574 4856 8630 4865
rect 8574 4791 8576 4800
rect 8628 4791 8630 4800
rect 8576 4762 8628 4768
rect 8772 4536 8800 6054
rect 8312 4440 8524 4468
rect 8680 4508 8800 4536
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8312 3602 8340 4440
rect 8574 4176 8630 4185
rect 8680 4146 8708 4508
rect 8864 4434 8892 7278
rect 8956 6254 8984 10542
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8772 4406 8892 4434
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8574 4111 8630 4120
rect 8668 4140 8720 4146
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8312 2650 8340 3538
rect 8390 3224 8446 3233
rect 8390 3159 8446 3168
rect 8404 2961 8432 3159
rect 8484 2984 8536 2990
rect 8390 2952 8446 2961
rect 8484 2926 8536 2932
rect 8390 2887 8446 2896
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8022 504 8078 513
rect 6918 368 6974 377
rect 6918 303 6974 312
rect 7286 0 7342 480
rect 7838 0 7894 480
rect 8404 480 8432 2790
rect 8496 2582 8524 2926
rect 8588 2836 8616 4111
rect 8668 4082 8720 4088
rect 8772 3482 8800 4406
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 3602 8892 3878
rect 8956 3777 8984 4422
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8772 3454 8892 3482
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 2990 8708 3334
rect 8668 2984 8720 2990
rect 8666 2952 8668 2961
rect 8720 2952 8722 2961
rect 8666 2887 8722 2896
rect 8668 2848 8720 2854
rect 8588 2808 8668 2836
rect 8668 2790 8720 2796
rect 8864 2666 8892 3454
rect 8864 2638 8984 2666
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8956 480 8984 2638
rect 9048 1601 9076 10474
rect 9140 5409 9168 10662
rect 9232 9217 9260 10798
rect 9324 10538 9352 22052
rect 9508 21894 9536 22086
rect 9588 22024 9640 22030
rect 9588 21966 9640 21972
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9600 21842 9628 21966
rect 9692 21962 9720 22335
rect 9876 22098 9904 24686
rect 9968 24342 9996 24754
rect 10289 24508 10585 24528
rect 10345 24506 10369 24508
rect 10425 24506 10449 24508
rect 10505 24506 10529 24508
rect 10367 24454 10369 24506
rect 10431 24454 10443 24506
rect 10505 24454 10507 24506
rect 10345 24452 10369 24454
rect 10425 24452 10449 24454
rect 10505 24452 10529 24454
rect 10289 24432 10585 24452
rect 9956 24336 10008 24342
rect 9956 24278 10008 24284
rect 9968 24070 9996 24278
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 9956 24064 10008 24070
rect 9956 24006 10008 24012
rect 9968 23866 9996 24006
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 9968 22778 9996 23802
rect 10520 23662 10548 24142
rect 10598 24032 10654 24041
rect 10598 23967 10654 23976
rect 10612 23780 10640 23967
rect 10704 23905 10732 25316
rect 10888 25129 10916 25463
rect 10968 25434 11020 25440
rect 11060 25492 11112 25498
rect 11060 25434 11112 25440
rect 11072 25378 11100 25434
rect 10980 25350 11100 25378
rect 11256 25362 11284 25978
rect 11244 25356 11296 25362
rect 10980 25294 11008 25350
rect 11244 25298 11296 25304
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10874 25120 10930 25129
rect 10874 25055 10930 25064
rect 11072 24614 11100 25230
rect 11348 24834 11376 27520
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11348 24806 11744 24834
rect 11610 24712 11666 24721
rect 11610 24647 11666 24656
rect 11060 24608 11112 24614
rect 11060 24550 11112 24556
rect 11072 24313 11100 24550
rect 11336 24336 11388 24342
rect 11058 24304 11114 24313
rect 11336 24278 11388 24284
rect 11058 24239 11114 24248
rect 11244 24064 11296 24070
rect 11244 24006 11296 24012
rect 10690 23896 10746 23905
rect 10690 23831 10746 23840
rect 10968 23792 11020 23798
rect 10612 23752 10732 23780
rect 10508 23656 10560 23662
rect 10508 23598 10560 23604
rect 10289 23420 10585 23440
rect 10345 23418 10369 23420
rect 10425 23418 10449 23420
rect 10505 23418 10529 23420
rect 10367 23366 10369 23418
rect 10431 23366 10443 23418
rect 10505 23366 10507 23418
rect 10345 23364 10369 23366
rect 10425 23364 10449 23366
rect 10505 23364 10529 23366
rect 10289 23344 10585 23364
rect 10140 23316 10192 23322
rect 10140 23258 10192 23264
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9968 22166 9996 22374
rect 10152 22234 10180 23258
rect 10289 22332 10585 22352
rect 10345 22330 10369 22332
rect 10425 22330 10449 22332
rect 10505 22330 10529 22332
rect 10367 22278 10369 22330
rect 10431 22278 10443 22330
rect 10505 22278 10507 22330
rect 10345 22276 10369 22278
rect 10425 22276 10449 22278
rect 10505 22276 10529 22278
rect 10289 22256 10585 22276
rect 10704 22234 10732 23752
rect 10874 23760 10930 23769
rect 10968 23734 11020 23740
rect 10874 23695 10930 23704
rect 10784 23656 10836 23662
rect 10784 23598 10836 23604
rect 10796 22982 10824 23598
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10140 22228 10192 22234
rect 10140 22170 10192 22176
rect 10692 22228 10744 22234
rect 10692 22170 10744 22176
rect 9956 22160 10008 22166
rect 9956 22102 10008 22108
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9680 21956 9732 21962
rect 9680 21898 9732 21904
rect 9600 21814 9720 21842
rect 9692 21321 9720 21814
rect 9784 21418 9812 22034
rect 9862 21992 9918 22001
rect 9862 21927 9918 21936
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 9678 21312 9734 21321
rect 9734 21270 9812 21298
rect 9678 21247 9734 21256
rect 9692 21187 9720 21247
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9588 20868 9640 20874
rect 9588 20810 9640 20816
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9416 19990 9444 20742
rect 9600 20602 9628 20810
rect 9588 20596 9640 20602
rect 9588 20538 9640 20544
rect 9692 20482 9720 21014
rect 9508 20466 9720 20482
rect 9508 20460 9732 20466
rect 9508 20454 9680 20460
rect 9404 19984 9456 19990
rect 9404 19926 9456 19932
rect 9416 19378 9444 19926
rect 9508 19718 9536 20454
rect 9680 20402 9732 20408
rect 9692 20371 9720 20402
rect 9678 20224 9734 20233
rect 9678 20159 9734 20168
rect 9692 19922 9720 20159
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9784 19802 9812 21270
rect 9876 20058 9904 21927
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9600 19774 9812 19802
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 19514 9536 19654
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9404 19372 9456 19378
rect 9404 19314 9456 19320
rect 9600 19258 9628 19774
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9508 19230 9628 19258
rect 9404 18964 9456 18970
rect 9404 18906 9456 18912
rect 9416 18290 9444 18906
rect 9508 18850 9536 19230
rect 9588 18964 9640 18970
rect 9692 18952 9720 19654
rect 9640 18924 9720 18952
rect 9588 18906 9640 18912
rect 9508 18822 9720 18850
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9600 18222 9628 18362
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9692 18034 9720 18822
rect 9600 18006 9720 18034
rect 9494 17640 9550 17649
rect 9494 17575 9550 17584
rect 9404 17060 9456 17066
rect 9404 17002 9456 17008
rect 9416 16794 9444 17002
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9402 16552 9458 16561
rect 9402 16487 9458 16496
rect 9416 15706 9444 16487
rect 9508 15706 9536 17575
rect 9600 17082 9628 18006
rect 9678 17912 9734 17921
rect 9678 17847 9734 17856
rect 9784 17864 9812 19654
rect 9862 19408 9918 19417
rect 9862 19343 9918 19352
rect 9876 18970 9904 19343
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9876 18222 9904 18770
rect 9968 18329 9996 22102
rect 10704 21554 10732 22170
rect 10796 22030 10824 22918
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10692 21548 10744 21554
rect 10692 21490 10744 21496
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10060 20806 10088 21422
rect 10796 21350 10824 21830
rect 10784 21344 10836 21350
rect 10784 21286 10836 21292
rect 10289 21244 10585 21264
rect 10345 21242 10369 21244
rect 10425 21242 10449 21244
rect 10505 21242 10529 21244
rect 10367 21190 10369 21242
rect 10431 21190 10443 21242
rect 10505 21190 10507 21242
rect 10345 21188 10369 21190
rect 10425 21188 10449 21190
rect 10505 21188 10529 21190
rect 10138 21176 10194 21185
rect 10289 21168 10585 21188
rect 10138 21111 10194 21120
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10060 20262 10088 20742
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10060 18834 10088 20198
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 10152 18714 10180 21111
rect 10888 20602 10916 23695
rect 10980 23254 11008 23734
rect 11256 23730 11284 24006
rect 11244 23724 11296 23730
rect 11244 23666 11296 23672
rect 11242 23624 11298 23633
rect 11242 23559 11298 23568
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 10968 23248 11020 23254
rect 11164 23225 11192 23462
rect 10968 23190 11020 23196
rect 11150 23216 11206 23225
rect 11060 23180 11112 23186
rect 11150 23151 11206 23160
rect 11060 23122 11112 23128
rect 11072 22817 11100 23122
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11058 22808 11114 22817
rect 11164 22778 11192 23054
rect 11058 22743 11114 22752
rect 11152 22772 11204 22778
rect 11072 22710 11100 22743
rect 11152 22714 11204 22720
rect 11256 22710 11284 23559
rect 11060 22704 11112 22710
rect 11060 22646 11112 22652
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11256 22574 11284 22646
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 11150 22128 11206 22137
rect 11150 22063 11206 22072
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 10980 21486 11008 21966
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10784 20392 10836 20398
rect 10888 20380 10916 20538
rect 10980 20534 11008 21286
rect 11072 21049 11100 21558
rect 11058 21040 11114 21049
rect 11058 20975 11114 20984
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10836 20352 10916 20380
rect 10784 20334 10836 20340
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10289 20156 10585 20176
rect 10345 20154 10369 20156
rect 10425 20154 10449 20156
rect 10505 20154 10529 20156
rect 10367 20102 10369 20154
rect 10431 20102 10443 20154
rect 10505 20102 10507 20154
rect 10345 20100 10369 20102
rect 10425 20100 10449 20102
rect 10505 20100 10529 20102
rect 10289 20080 10585 20100
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10244 19417 10272 19858
rect 10322 19816 10378 19825
rect 10322 19751 10378 19760
rect 10230 19408 10286 19417
rect 10230 19343 10286 19352
rect 10336 19281 10364 19751
rect 10600 19712 10652 19718
rect 10704 19700 10732 20198
rect 10652 19672 10732 19700
rect 10600 19654 10652 19660
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10322 19272 10378 19281
rect 10322 19207 10378 19216
rect 10289 19068 10585 19088
rect 10345 19066 10369 19068
rect 10425 19066 10449 19068
rect 10505 19066 10529 19068
rect 10367 19014 10369 19066
rect 10431 19014 10443 19066
rect 10505 19014 10507 19066
rect 10345 19012 10369 19014
rect 10425 19012 10449 19014
rect 10505 19012 10529 19014
rect 10289 18992 10585 19012
rect 10060 18686 10180 18714
rect 9954 18320 10010 18329
rect 9954 18255 10010 18264
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9692 17746 9720 17847
rect 9784 17836 9904 17864
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9692 17270 9720 17682
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9600 17054 9720 17082
rect 9586 16552 9642 16561
rect 9586 16487 9642 16496
rect 9600 15881 9628 16487
rect 9692 16046 9720 17054
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9680 15904 9732 15910
rect 9586 15872 9642 15881
rect 9680 15846 9732 15852
rect 9586 15807 9642 15816
rect 9692 15745 9720 15846
rect 9678 15736 9734 15745
rect 9404 15700 9456 15706
rect 9404 15642 9456 15648
rect 9496 15700 9548 15706
rect 9678 15671 9734 15680
rect 9496 15642 9548 15648
rect 9496 14816 9548 14822
rect 9496 14758 9548 14764
rect 9678 14784 9734 14793
rect 9508 14278 9536 14758
rect 9678 14719 9734 14728
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9508 13802 9536 14214
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 13530 9536 13738
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9588 13320 9640 13326
rect 9588 13262 9640 13268
rect 9600 12918 9628 13262
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 9508 12458 9536 12650
rect 9416 12430 9536 12458
rect 9312 10532 9364 10538
rect 9312 10474 9364 10480
rect 9310 10432 9366 10441
rect 9310 10367 9366 10376
rect 9324 10062 9352 10367
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9416 9625 9444 12430
rect 9600 12306 9628 12854
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11218 9628 11562
rect 9692 11354 9720 14719
rect 9770 14104 9826 14113
rect 9770 14039 9826 14048
rect 9784 13705 9812 14039
rect 9770 13696 9826 13705
rect 9770 13631 9826 13640
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9784 12889 9812 13330
rect 9770 12880 9826 12889
rect 9876 12866 9904 17836
rect 9956 17128 10008 17134
rect 9956 17070 10008 17076
rect 9968 16794 9996 17070
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 10060 15586 10088 18686
rect 10289 17980 10585 18000
rect 10345 17978 10369 17980
rect 10425 17978 10449 17980
rect 10505 17978 10529 17980
rect 10367 17926 10369 17978
rect 10431 17926 10443 17978
rect 10505 17926 10507 17978
rect 10345 17924 10369 17926
rect 10425 17924 10449 17926
rect 10505 17924 10529 17926
rect 10289 17904 10585 17924
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10244 17338 10272 17614
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10244 17048 10272 17274
rect 10152 17020 10272 17048
rect 10152 16726 10180 17020
rect 10289 16892 10585 16912
rect 10345 16890 10369 16892
rect 10425 16890 10449 16892
rect 10505 16890 10529 16892
rect 10367 16838 10369 16890
rect 10431 16838 10443 16890
rect 10505 16838 10507 16890
rect 10345 16836 10369 16838
rect 10425 16836 10449 16838
rect 10505 16836 10529 16838
rect 10289 16816 10585 16836
rect 10704 16776 10732 19450
rect 10612 16748 10732 16776
rect 10140 16720 10192 16726
rect 10140 16662 10192 16668
rect 10152 16114 10180 16662
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 16250 10364 16594
rect 10612 16266 10640 16748
rect 10796 16504 10824 20334
rect 10874 20224 10930 20233
rect 10874 20159 10930 20168
rect 10888 18154 10916 20159
rect 10980 19514 11008 20470
rect 11072 20058 11100 20975
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11164 19514 11192 22063
rect 11348 20058 11376 24278
rect 11520 24200 11572 24206
rect 11518 24168 11520 24177
rect 11572 24168 11574 24177
rect 11518 24103 11574 24112
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23730 11468 24006
rect 11518 23760 11574 23769
rect 11428 23724 11480 23730
rect 11518 23695 11574 23704
rect 11428 23666 11480 23672
rect 11426 23080 11482 23089
rect 11426 23015 11482 23024
rect 11440 22778 11468 23015
rect 11428 22772 11480 22778
rect 11428 22714 11480 22720
rect 11532 22658 11560 23695
rect 11440 22630 11560 22658
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11336 19848 11388 19854
rect 11336 19790 11388 19796
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 11152 19508 11204 19514
rect 11152 19450 11204 19456
rect 11348 19378 11376 19790
rect 11440 19666 11468 22630
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11532 21690 11560 22034
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11624 21026 11652 24647
rect 11532 20998 11652 21026
rect 11532 20330 11560 20998
rect 11612 20936 11664 20942
rect 11610 20904 11612 20913
rect 11664 20904 11666 20913
rect 11610 20839 11666 20848
rect 11520 20324 11572 20330
rect 11520 20266 11572 20272
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11440 19638 11560 19666
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11164 18358 11192 18838
rect 11152 18352 11204 18358
rect 11152 18294 11204 18300
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10874 18048 10930 18057
rect 10874 17983 10930 17992
rect 10888 17882 10916 17983
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10796 16476 10916 16504
rect 10324 16244 10376 16250
rect 10612 16238 10732 16266
rect 10324 16186 10376 16192
rect 10140 16108 10192 16114
rect 10140 16050 10192 16056
rect 10152 15706 10180 16050
rect 10289 15804 10585 15824
rect 10345 15802 10369 15804
rect 10425 15802 10449 15804
rect 10505 15802 10529 15804
rect 10367 15750 10369 15802
rect 10431 15750 10443 15802
rect 10505 15750 10507 15802
rect 10345 15748 10369 15750
rect 10425 15748 10449 15750
rect 10505 15748 10529 15750
rect 10289 15728 10585 15748
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10060 15558 10180 15586
rect 10048 14408 10100 14414
rect 10048 14350 10100 14356
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 13841 9996 14214
rect 9954 13832 10010 13841
rect 9954 13767 10010 13776
rect 9954 13560 10010 13569
rect 9954 13495 9956 13504
rect 10008 13495 10010 13504
rect 9956 13466 10008 13472
rect 9954 13152 10010 13161
rect 10060 13138 10088 14350
rect 10152 13512 10180 15558
rect 10508 15360 10560 15366
rect 10506 15328 10508 15337
rect 10560 15328 10562 15337
rect 10506 15263 10562 15272
rect 10289 14716 10585 14736
rect 10345 14714 10369 14716
rect 10425 14714 10449 14716
rect 10505 14714 10529 14716
rect 10367 14662 10369 14714
rect 10431 14662 10443 14714
rect 10505 14662 10507 14714
rect 10345 14660 10369 14662
rect 10425 14660 10449 14662
rect 10505 14660 10529 14662
rect 10289 14640 10585 14660
rect 10704 14600 10732 16238
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10796 15570 10824 16186
rect 10784 15564 10836 15570
rect 10784 15506 10836 15512
rect 10796 15162 10824 15506
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10796 14890 10824 15098
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10612 14572 10732 14600
rect 10612 13802 10640 14572
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10600 13796 10652 13802
rect 10600 13738 10652 13744
rect 10289 13628 10585 13648
rect 10345 13626 10369 13628
rect 10425 13626 10449 13628
rect 10505 13626 10529 13628
rect 10367 13574 10369 13626
rect 10431 13574 10443 13626
rect 10505 13574 10507 13626
rect 10345 13572 10369 13574
rect 10425 13572 10449 13574
rect 10505 13572 10529 13574
rect 10289 13552 10585 13572
rect 10152 13484 10272 13512
rect 10138 13288 10194 13297
rect 10138 13223 10194 13232
rect 10010 13110 10088 13138
rect 9954 13087 10010 13096
rect 9968 12986 9996 13087
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 9876 12838 10088 12866
rect 9770 12815 9826 12824
rect 9784 12442 9812 12815
rect 9956 12776 10008 12782
rect 9862 12744 9918 12753
rect 9956 12718 10008 12724
rect 9862 12679 9918 12688
rect 9876 12646 9904 12679
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9876 12442 9904 12582
rect 9772 12436 9824 12442
rect 9772 12378 9824 12384
rect 9864 12436 9916 12442
rect 9864 12378 9916 12384
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 11098 9720 11154
rect 9508 11070 9720 11098
rect 9402 9616 9458 9625
rect 9402 9551 9458 9560
rect 9402 9480 9458 9489
rect 9402 9415 9404 9424
rect 9456 9415 9458 9424
rect 9404 9386 9456 9392
rect 9218 9208 9274 9217
rect 9218 9143 9274 9152
rect 9312 9172 9364 9178
rect 9126 5400 9182 5409
rect 9126 5335 9182 5344
rect 9140 5030 9168 5335
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9140 3466 9168 4150
rect 9232 3942 9260 9143
rect 9416 9160 9444 9386
rect 9364 9132 9444 9160
rect 9312 9114 9364 9120
rect 9324 8634 9352 9114
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9312 5160 9364 5166
rect 9310 5128 9312 5137
rect 9364 5128 9366 5137
rect 9310 5063 9366 5072
rect 9416 5012 9444 7210
rect 9324 4984 9444 5012
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 9324 2281 9352 4984
rect 9402 4720 9458 4729
rect 9402 4655 9458 4664
rect 9416 3058 9444 4655
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9310 2272 9366 2281
rect 9310 2207 9366 2216
rect 9034 1592 9090 1601
rect 9034 1527 9090 1536
rect 9218 1592 9274 1601
rect 9218 1527 9220 1536
rect 9272 1527 9274 1536
rect 9220 1498 9272 1504
rect 9416 1465 9444 2994
rect 9508 2990 9536 11070
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10690 9720 10950
rect 9600 10674 9720 10690
rect 9600 10668 9732 10674
rect 9600 10662 9680 10668
rect 9600 10198 9628 10662
rect 9680 10610 9732 10616
rect 9678 10568 9734 10577
rect 9678 10503 9734 10512
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9692 10130 9720 10503
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 9586 9616 9642 9625
rect 9586 9551 9642 9560
rect 9600 9518 9628 9551
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 8090 9628 9318
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9692 8022 9720 8910
rect 9784 8498 9812 12242
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9772 8356 9824 8362
rect 9772 8298 9824 8304
rect 9784 8090 9812 8298
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7342 9628 7754
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 9600 6882 9628 7278
rect 9600 6854 9720 6882
rect 9692 4826 9720 6854
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9784 5778 9812 6054
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4758 9812 5714
rect 9772 4752 9824 4758
rect 9772 4694 9824 4700
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9692 3738 9720 3975
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9784 3618 9812 4558
rect 9876 3738 9904 12242
rect 9968 10266 9996 12718
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9954 10024 10010 10033
rect 9954 9959 10010 9968
rect 9968 8634 9996 9959
rect 9956 8628 10008 8634
rect 9956 8570 10008 8576
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9968 8090 9996 8434
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9968 7002 9996 8026
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9968 5574 9996 6734
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9956 4752 10008 4758
rect 9954 4720 9956 4729
rect 10008 4720 10010 4729
rect 9954 4655 10010 4664
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9692 3590 9812 3618
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9402 1456 9458 1465
rect 9402 1391 9458 1400
rect 9508 480 9536 2790
rect 9600 1329 9628 3470
rect 9586 1320 9642 1329
rect 9586 1255 9642 1264
rect 8022 439 8078 448
rect 8390 0 8446 480
rect 8942 0 8998 480
rect 9494 0 9550 480
rect 9692 105 9720 3590
rect 9770 3496 9826 3505
rect 9770 3431 9826 3440
rect 9784 3194 9812 3431
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9876 3126 9904 3674
rect 9968 3369 9996 3878
rect 9954 3360 10010 3369
rect 9954 3295 10010 3304
rect 9864 3120 9916 3126
rect 9864 3062 9916 3068
rect 10060 480 10088 12838
rect 10152 10266 10180 13223
rect 10244 12782 10272 13484
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10322 13288 10378 13297
rect 10322 13223 10378 13232
rect 10232 12776 10284 12782
rect 10336 12753 10364 13223
rect 10612 12850 10640 13330
rect 10796 13190 10824 14418
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10508 12776 10560 12782
rect 10232 12718 10284 12724
rect 10322 12744 10378 12753
rect 10322 12679 10378 12688
rect 10506 12744 10508 12753
rect 10560 12744 10562 12753
rect 10506 12679 10562 12688
rect 10692 12708 10744 12714
rect 10692 12650 10744 12656
rect 10289 12540 10585 12560
rect 10345 12538 10369 12540
rect 10425 12538 10449 12540
rect 10505 12538 10529 12540
rect 10367 12486 10369 12538
rect 10431 12486 10443 12538
rect 10505 12486 10507 12538
rect 10345 12484 10369 12486
rect 10425 12484 10449 12486
rect 10505 12484 10529 12486
rect 10289 12464 10585 12484
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10428 11898 10456 12174
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10289 11452 10585 11472
rect 10345 11450 10369 11452
rect 10425 11450 10449 11452
rect 10505 11450 10529 11452
rect 10367 11398 10369 11450
rect 10431 11398 10443 11450
rect 10505 11398 10507 11450
rect 10345 11396 10369 11398
rect 10425 11396 10449 11398
rect 10505 11396 10529 11398
rect 10289 11376 10585 11396
rect 10506 11112 10562 11121
rect 10506 11047 10508 11056
rect 10560 11047 10562 11056
rect 10508 11018 10560 11024
rect 10289 10364 10585 10384
rect 10345 10362 10369 10364
rect 10425 10362 10449 10364
rect 10505 10362 10529 10364
rect 10367 10310 10369 10362
rect 10431 10310 10443 10362
rect 10505 10310 10507 10362
rect 10345 10308 10369 10310
rect 10425 10308 10449 10310
rect 10505 10308 10529 10310
rect 10289 10288 10585 10308
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 10289 9276 10585 9296
rect 10345 9274 10369 9276
rect 10425 9274 10449 9276
rect 10505 9274 10529 9276
rect 10367 9222 10369 9274
rect 10431 9222 10443 9274
rect 10505 9222 10507 9274
rect 10345 9220 10369 9222
rect 10425 9220 10449 9222
rect 10505 9220 10529 9222
rect 10289 9200 10585 9220
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 10152 8294 10180 8978
rect 10244 8634 10272 9046
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10152 7410 10180 8230
rect 10289 8188 10585 8208
rect 10345 8186 10369 8188
rect 10425 8186 10449 8188
rect 10505 8186 10529 8188
rect 10367 8134 10369 8186
rect 10431 8134 10443 8186
rect 10505 8134 10507 8186
rect 10345 8132 10369 8134
rect 10425 8132 10449 8134
rect 10505 8132 10529 8134
rect 10289 8112 10585 8132
rect 10704 8090 10732 12650
rect 10796 12481 10824 13126
rect 10888 12782 10916 16476
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10980 12714 11008 18158
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 16674 11100 18022
rect 11164 16998 11192 18294
rect 11256 18170 11284 19246
rect 11348 18970 11376 19314
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11348 18290 11376 18906
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11256 18142 11376 18170
rect 11244 18080 11296 18086
rect 11242 18048 11244 18057
rect 11296 18048 11298 18057
rect 11242 17983 11298 17992
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16697 11192 16934
rect 11063 16646 11100 16674
rect 11150 16688 11206 16697
rect 11063 16572 11091 16646
rect 11150 16623 11206 16632
rect 11063 16544 11100 16572
rect 11072 16504 11100 16544
rect 11072 16476 11192 16504
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 11072 15026 11100 15574
rect 11164 15162 11192 16476
rect 11256 16425 11284 17478
rect 11242 16416 11298 16425
rect 11242 16351 11298 16360
rect 11242 15736 11298 15745
rect 11348 15722 11376 18142
rect 11440 17882 11468 19450
rect 11532 19174 11560 19638
rect 11624 19446 11652 19994
rect 11612 19440 11664 19446
rect 11612 19382 11664 19388
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11532 18952 11560 19110
rect 11716 19009 11744 24806
rect 11808 23798 11836 25162
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11900 23361 11928 27520
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11992 24818 12020 25842
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 11980 24812 12032 24818
rect 11980 24754 12032 24760
rect 11992 24682 12020 24754
rect 11980 24676 12032 24682
rect 11980 24618 12032 24624
rect 11886 23352 11942 23361
rect 11886 23287 11942 23296
rect 11796 23248 11848 23254
rect 11796 23190 11848 23196
rect 11808 22438 11836 23190
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11980 22432 12032 22438
rect 11980 22374 12032 22380
rect 11808 19718 11836 22374
rect 11888 21548 11940 21554
rect 11888 21490 11940 21496
rect 11900 21350 11928 21490
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20466 11928 21286
rect 11888 20460 11940 20466
rect 11888 20402 11940 20408
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11702 19000 11758 19009
rect 11532 18924 11652 18952
rect 11758 18958 11836 18986
rect 11702 18935 11758 18944
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11532 18426 11560 18770
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11440 16522 11468 17818
rect 11428 16516 11480 16522
rect 11428 16458 11480 16464
rect 11426 16416 11482 16425
rect 11426 16351 11482 16360
rect 11298 15694 11376 15722
rect 11242 15671 11298 15680
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 14618 11100 14962
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14612 11112 14618
rect 11060 14554 11112 14560
rect 11072 14414 11100 14554
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11072 14074 11100 14350
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13977 11192 14758
rect 11150 13968 11206 13977
rect 11150 13903 11206 13912
rect 11256 13818 11284 15671
rect 11440 15609 11468 16351
rect 11426 15600 11482 15609
rect 11426 15535 11482 15544
rect 11428 15156 11480 15162
rect 11428 15098 11480 15104
rect 11334 15056 11390 15065
rect 11334 14991 11390 15000
rect 11348 14618 11376 14991
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11060 13796 11112 13802
rect 11060 13738 11112 13744
rect 11164 13790 11284 13818
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10876 12640 10928 12646
rect 11072 12594 11100 13738
rect 11164 12646 11192 13790
rect 11336 13524 11388 13530
rect 11440 13512 11468 15098
rect 11388 13484 11468 13512
rect 11336 13466 11388 13472
rect 11242 13288 11298 13297
rect 11242 13223 11244 13232
rect 11296 13223 11298 13232
rect 11244 13194 11296 13200
rect 11348 12850 11376 13466
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 10876 12582 10928 12588
rect 10782 12472 10838 12481
rect 10782 12407 10838 12416
rect 10888 12356 10916 12582
rect 10796 12328 10916 12356
rect 10980 12566 11100 12594
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 10796 11286 10824 12328
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 9897 10824 11086
rect 10888 10198 10916 11494
rect 10876 10192 10928 10198
rect 10876 10134 10928 10140
rect 10782 9888 10838 9897
rect 10782 9823 10838 9832
rect 10796 9178 10824 9823
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10888 8838 10916 10134
rect 10876 8832 10928 8838
rect 10796 8780 10876 8786
rect 10796 8774 10928 8780
rect 10796 8758 10916 8774
rect 10796 8498 10824 8758
rect 10980 8514 11008 12566
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 11072 11558 11100 12242
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11150 11248 11206 11257
rect 11150 11183 11206 11192
rect 11164 10810 11192 11183
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11164 10606 11192 10746
rect 11256 10674 11284 11086
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 9994 11100 10406
rect 11348 10266 11376 12582
rect 11336 10260 11388 10266
rect 11164 10220 11336 10248
rect 11164 10062 11192 10220
rect 11336 10202 11388 10208
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11164 9722 11192 9998
rect 11256 9722 11284 10066
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10888 8486 11008 8514
rect 10784 8288 10836 8294
rect 10784 8230 10836 8236
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10704 7546 10732 8026
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10796 7478 10824 8230
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10796 7342 10824 7414
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10784 7200 10836 7206
rect 10690 7168 10746 7177
rect 10289 7100 10585 7120
rect 10784 7142 10836 7148
rect 10690 7103 10746 7112
rect 10345 7098 10369 7100
rect 10425 7098 10449 7100
rect 10505 7098 10529 7100
rect 10367 7046 10369 7098
rect 10431 7046 10443 7098
rect 10505 7046 10507 7098
rect 10345 7044 10369 7046
rect 10425 7044 10449 7046
rect 10505 7044 10529 7046
rect 10138 7032 10194 7041
rect 10289 7024 10585 7044
rect 10704 6984 10732 7103
rect 10194 6976 10732 6984
rect 10138 6967 10732 6976
rect 10152 6956 10732 6967
rect 10796 6934 10824 7142
rect 10784 6928 10836 6934
rect 10784 6870 10836 6876
rect 10414 6624 10470 6633
rect 10414 6559 10470 6568
rect 10428 6458 10456 6559
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10428 6254 10456 6394
rect 10888 6390 10916 8486
rect 10968 8424 11020 8430
rect 11020 8372 11100 8378
rect 10968 8366 11100 8372
rect 10980 8350 11100 8366
rect 10966 8256 11022 8265
rect 10966 8191 11022 8200
rect 10876 6384 10928 6390
rect 10876 6326 10928 6332
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10784 6112 10836 6118
rect 10690 6080 10746 6089
rect 10289 6012 10585 6032
rect 10784 6054 10836 6060
rect 10690 6015 10746 6024
rect 10345 6010 10369 6012
rect 10425 6010 10449 6012
rect 10505 6010 10529 6012
rect 10367 5958 10369 6010
rect 10431 5958 10443 6010
rect 10505 5958 10507 6010
rect 10345 5956 10369 5958
rect 10425 5956 10449 5958
rect 10505 5956 10529 5958
rect 10289 5936 10585 5956
rect 10704 5817 10732 6015
rect 10796 5953 10824 6054
rect 10782 5944 10838 5953
rect 10782 5879 10838 5888
rect 10876 5840 10928 5846
rect 10690 5808 10746 5817
rect 10876 5782 10928 5788
rect 10690 5743 10746 5752
rect 10888 5574 10916 5782
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10152 4622 10180 5102
rect 10289 4924 10585 4944
rect 10345 4922 10369 4924
rect 10425 4922 10449 4924
rect 10505 4922 10529 4924
rect 10367 4870 10369 4922
rect 10431 4870 10443 4922
rect 10505 4870 10507 4922
rect 10345 4868 10369 4870
rect 10425 4868 10449 4870
rect 10505 4868 10529 4870
rect 10289 4848 10585 4868
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10612 4010 10640 4626
rect 10704 4622 10732 5238
rect 10888 5234 10916 5510
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10796 4865 10824 4966
rect 10782 4856 10838 4865
rect 10782 4791 10838 4800
rect 10888 4706 10916 5170
rect 10980 5098 11008 8191
rect 11072 8090 11100 8350
rect 11164 8294 11192 9658
rect 11334 9072 11390 9081
rect 11244 9036 11296 9042
rect 11334 9007 11390 9016
rect 11244 8978 11296 8984
rect 11256 8634 11284 8978
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11164 7342 11192 7958
rect 11256 7954 11284 8570
rect 11244 7948 11296 7954
rect 11244 7890 11296 7896
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11164 6322 11192 6802
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 11164 5574 11192 6258
rect 11152 5568 11204 5574
rect 11152 5510 11204 5516
rect 11150 5400 11206 5409
rect 11060 5364 11112 5370
rect 11150 5335 11206 5344
rect 11060 5306 11112 5312
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10796 4678 10916 4706
rect 10796 4622 10824 4678
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 10704 4282 10732 4558
rect 10692 4276 10744 4282
rect 10692 4218 10744 4224
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10690 3904 10746 3913
rect 10289 3836 10585 3856
rect 10690 3839 10746 3848
rect 10345 3834 10369 3836
rect 10425 3834 10449 3836
rect 10505 3834 10529 3836
rect 10367 3782 10369 3834
rect 10431 3782 10443 3834
rect 10505 3782 10507 3834
rect 10345 3780 10369 3782
rect 10425 3780 10449 3782
rect 10505 3780 10529 3782
rect 10289 3760 10585 3780
rect 10704 3670 10732 3839
rect 10796 3738 10824 4558
rect 11164 4554 11192 5335
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11150 4448 11206 4457
rect 11072 4185 11100 4422
rect 11150 4383 11206 4392
rect 11058 4176 11114 4185
rect 11058 4111 11114 4120
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10152 3194 10180 3470
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10289 2748 10585 2768
rect 10345 2746 10369 2748
rect 10425 2746 10449 2748
rect 10505 2746 10529 2748
rect 10367 2694 10369 2746
rect 10431 2694 10443 2746
rect 10505 2694 10507 2746
rect 10345 2692 10369 2694
rect 10425 2692 10449 2694
rect 10505 2692 10529 2694
rect 10138 2680 10194 2689
rect 10289 2672 10585 2692
rect 10138 2615 10140 2624
rect 10192 2615 10194 2624
rect 10140 2586 10192 2592
rect 10704 1442 10732 3295
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10796 2514 10824 2858
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10888 2009 10916 3946
rect 10980 3777 11008 4014
rect 10966 3768 11022 3777
rect 10966 3703 11022 3712
rect 11072 3058 11100 4111
rect 11164 3602 11192 4383
rect 11242 4312 11298 4321
rect 11242 4247 11298 4256
rect 11256 4146 11284 4247
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11348 3482 11376 9007
rect 11440 4758 11468 12922
rect 11532 12646 11560 18158
rect 11624 12646 11652 18924
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 17066 11744 17546
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11716 16794 11744 17002
rect 11704 16788 11756 16794
rect 11704 16730 11756 16736
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11716 15892 11744 16458
rect 11808 16017 11836 18958
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 17338 11928 18362
rect 11888 17332 11940 17338
rect 11888 17274 11940 17280
rect 11794 16008 11850 16017
rect 11794 15943 11850 15952
rect 11716 15864 11836 15892
rect 11702 14512 11758 14521
rect 11702 14447 11704 14456
rect 11756 14447 11758 14456
rect 11704 14418 11756 14424
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 12986 11744 13262
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11518 11656 11574 11665
rect 11518 11591 11574 11600
rect 11532 11354 11560 11591
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 11520 11008 11572 11014
rect 11716 10985 11744 12650
rect 11520 10950 11572 10956
rect 11702 10976 11758 10985
rect 11532 9382 11560 10950
rect 11702 10911 11758 10920
rect 11716 10742 11744 10911
rect 11704 10736 11756 10742
rect 11704 10678 11756 10684
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11532 8634 11560 9318
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11624 5302 11652 9318
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11716 7410 11744 7686
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 6662 11744 7346
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11808 5658 11836 15864
rect 11886 14240 11942 14249
rect 11886 14175 11942 14184
rect 11900 12374 11928 14175
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11886 11384 11942 11393
rect 11886 11319 11888 11328
rect 11940 11319 11942 11328
rect 11888 11290 11940 11296
rect 11886 10160 11942 10169
rect 11886 10095 11888 10104
rect 11940 10095 11942 10104
rect 11888 10066 11940 10072
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11900 7546 11928 7890
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11900 6458 11928 7482
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 6118 11928 6394
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11808 5630 11928 5658
rect 11796 5568 11848 5574
rect 11716 5528 11796 5556
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11440 4282 11468 4490
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11624 4060 11652 5102
rect 11716 4570 11744 5528
rect 11796 5510 11848 5516
rect 11900 5166 11928 5630
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11888 5024 11940 5030
rect 11794 4992 11850 5001
rect 11888 4966 11940 4972
rect 11794 4927 11850 4936
rect 11808 4826 11836 4927
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11716 4542 11836 4570
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11716 4185 11744 4422
rect 11702 4176 11758 4185
rect 11702 4111 11758 4120
rect 11624 4032 11744 4060
rect 11520 3664 11572 3670
rect 11518 3632 11520 3641
rect 11572 3632 11574 3641
rect 11716 3618 11744 4032
rect 11518 3567 11574 3576
rect 11624 3590 11744 3618
rect 11164 3454 11376 3482
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10874 2000 10930 2009
rect 10874 1935 10930 1944
rect 10612 1414 10732 1442
rect 10612 480 10640 1414
rect 11164 480 11192 3454
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 3097 11284 3334
rect 11624 3108 11652 3590
rect 11704 3528 11756 3534
rect 11808 3516 11836 4542
rect 11900 4321 11928 4966
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11756 3488 11836 3516
rect 11704 3470 11756 3476
rect 11716 3233 11744 3470
rect 11702 3224 11758 3233
rect 11702 3159 11758 3168
rect 11242 3088 11298 3097
rect 11624 3080 11744 3108
rect 11242 3023 11298 3032
rect 11334 2952 11390 2961
rect 11334 2887 11390 2896
rect 11348 2854 11376 2887
rect 11336 2848 11388 2854
rect 11242 2816 11298 2825
rect 11336 2790 11388 2796
rect 11242 2751 11298 2760
rect 11256 2310 11284 2751
rect 11348 2582 11376 2790
rect 11336 2576 11388 2582
rect 11336 2518 11388 2524
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11256 1193 11284 2246
rect 11242 1184 11298 1193
rect 11242 1119 11298 1128
rect 11716 480 11744 3080
rect 11900 1057 11928 4150
rect 11992 1170 12020 22374
rect 12084 21146 12112 24890
rect 12176 23202 12204 25910
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12268 24818 12296 25094
rect 12256 24812 12308 24818
rect 12256 24754 12308 24760
rect 12360 24750 12388 24781
rect 12348 24744 12400 24750
rect 12452 24698 12480 25366
rect 12544 24750 12572 27520
rect 13096 25378 13124 27520
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13096 25350 13308 25378
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 12624 24812 12676 24818
rect 12624 24754 12676 24760
rect 12400 24692 12480 24698
rect 12348 24686 12480 24692
rect 12532 24744 12584 24750
rect 12532 24686 12584 24692
rect 12360 24670 12480 24686
rect 12256 24200 12308 24206
rect 12256 24142 12308 24148
rect 12268 23866 12296 24142
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12360 23769 12388 24670
rect 12346 23760 12402 23769
rect 12346 23695 12402 23704
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12360 23474 12388 23598
rect 12360 23446 12480 23474
rect 12176 23174 12388 23202
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12176 22778 12204 23054
rect 12254 22808 12310 22817
rect 12164 22772 12216 22778
rect 12254 22743 12310 22752
rect 12164 22714 12216 22720
rect 12176 22642 12204 22714
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12268 22234 12296 22743
rect 12256 22228 12308 22234
rect 12256 22170 12308 22176
rect 12360 21593 12388 23174
rect 12452 22778 12480 23446
rect 12544 22982 12572 23598
rect 12636 23594 12664 24754
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12532 22976 12584 22982
rect 12532 22918 12584 22924
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12636 22234 12664 23530
rect 12728 22574 12756 24550
rect 13096 24410 13124 25230
rect 13176 24676 13228 24682
rect 13176 24618 13228 24624
rect 13084 24404 13136 24410
rect 13084 24346 13136 24352
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12820 23225 12848 23258
rect 12806 23216 12862 23225
rect 12806 23151 12862 23160
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12728 22234 12756 22510
rect 12912 22234 12940 22578
rect 13004 22506 13032 24006
rect 13096 23322 13124 24346
rect 13188 23497 13216 24618
rect 13280 24138 13308 25350
rect 13358 24848 13414 24857
rect 13358 24783 13414 24792
rect 13372 24274 13400 24783
rect 13464 24410 13492 25842
rect 13542 24984 13598 24993
rect 13648 24970 13676 27520
rect 14186 25800 14242 25809
rect 14186 25735 14242 25744
rect 14004 25696 14056 25702
rect 14004 25638 14056 25644
rect 13648 24942 13768 24970
rect 13542 24919 13598 24928
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13360 24268 13412 24274
rect 13360 24210 13412 24216
rect 13464 24206 13492 24346
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13174 23488 13230 23497
rect 13174 23423 13230 23432
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13096 22778 13124 23258
rect 13084 22772 13136 22778
rect 13084 22714 13136 22720
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 13096 22438 13124 22714
rect 13280 22545 13308 24074
rect 13556 23338 13584 24919
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13648 24206 13676 24754
rect 13740 24698 13768 24942
rect 13740 24670 13860 24698
rect 14016 24682 14044 25638
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13740 24449 13768 24550
rect 13726 24440 13782 24449
rect 13726 24375 13782 24384
rect 13832 24290 13860 24670
rect 14004 24676 14056 24682
rect 14004 24618 14056 24624
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13740 24262 13860 24290
rect 13912 24268 13964 24274
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13648 23866 13676 24142
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13740 23338 13768 24262
rect 13912 24210 13964 24216
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13464 23310 13584 23338
rect 13648 23310 13768 23338
rect 13360 22568 13412 22574
rect 13266 22536 13322 22545
rect 13360 22510 13412 22516
rect 13266 22471 13322 22480
rect 13084 22432 13136 22438
rect 13084 22374 13136 22380
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13082 22264 13138 22273
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12624 22228 12676 22234
rect 12624 22170 12676 22176
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12900 22228 12952 22234
rect 13082 22199 13138 22208
rect 12900 22170 12952 22176
rect 12452 21690 12480 22170
rect 12990 22128 13046 22137
rect 12990 22063 13046 22072
rect 12530 21720 12586 21729
rect 12440 21684 12492 21690
rect 12530 21655 12586 21664
rect 12900 21684 12952 21690
rect 12440 21626 12492 21632
rect 12346 21584 12402 21593
rect 12544 21570 12572 21655
rect 12900 21626 12952 21632
rect 12346 21519 12402 21528
rect 12452 21542 12572 21570
rect 12254 21176 12310 21185
rect 12072 21140 12124 21146
rect 12254 21111 12310 21120
rect 12072 21082 12124 21088
rect 12070 20768 12126 20777
rect 12070 20703 12126 20712
rect 12084 20233 12112 20703
rect 12164 20256 12216 20262
rect 12070 20224 12126 20233
rect 12164 20198 12216 20204
rect 12070 20159 12126 20168
rect 12176 19961 12204 20198
rect 12162 19952 12218 19961
rect 12268 19922 12296 21111
rect 12162 19887 12218 19896
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12268 19514 12296 19858
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12070 17776 12126 17785
rect 12070 17711 12126 17720
rect 12084 17610 12112 17711
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12360 16538 12388 21519
rect 12452 19446 12480 21542
rect 12716 21072 12768 21078
rect 12622 21040 12678 21049
rect 12532 21004 12584 21010
rect 12716 21014 12768 21020
rect 12622 20975 12624 20984
rect 12532 20946 12584 20952
rect 12676 20975 12678 20984
rect 12624 20946 12676 20952
rect 12544 20602 12572 20946
rect 12728 20942 12756 21014
rect 12716 20936 12768 20942
rect 12622 20904 12678 20913
rect 12768 20896 12848 20924
rect 12716 20878 12768 20884
rect 12622 20839 12678 20848
rect 12532 20596 12584 20602
rect 12532 20538 12584 20544
rect 12636 20534 12664 20839
rect 12820 20602 12848 20896
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12912 20398 12940 21626
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12900 20392 12952 20398
rect 12900 20334 12952 20340
rect 12636 20262 12664 20334
rect 12624 20256 12676 20262
rect 12530 20224 12586 20233
rect 12624 20198 12676 20204
rect 12530 20159 12586 20168
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12544 19394 12572 20159
rect 12912 20058 12940 20334
rect 12900 20052 12952 20058
rect 12900 19994 12952 20000
rect 12624 19984 12676 19990
rect 12624 19926 12676 19932
rect 12636 19514 12664 19926
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12624 19508 12676 19514
rect 12624 19450 12676 19456
rect 12544 19366 12756 19394
rect 12820 19378 12848 19858
rect 12912 19689 12940 19994
rect 12898 19680 12954 19689
rect 12898 19615 12954 19624
rect 13004 19496 13032 22063
rect 13096 19825 13124 22199
rect 13280 20618 13308 22374
rect 13372 21894 13400 22510
rect 13464 22438 13492 23310
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13556 22234 13584 23122
rect 13648 22964 13676 23310
rect 13832 23202 13860 23462
rect 13924 23254 13952 24210
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13740 23174 13860 23202
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13740 23118 13768 23174
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13648 22936 13768 22964
rect 13740 22273 13768 22936
rect 13912 22704 13964 22710
rect 13912 22646 13964 22652
rect 13726 22264 13782 22273
rect 13544 22228 13596 22234
rect 13726 22199 13782 22208
rect 13544 22170 13596 22176
rect 13820 22160 13872 22166
rect 13820 22102 13872 22108
rect 13360 21888 13412 21894
rect 13360 21830 13412 21836
rect 13372 21486 13400 21830
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13636 21412 13688 21418
rect 13636 21354 13688 21360
rect 13648 21078 13676 21354
rect 13728 21140 13780 21146
rect 13832 21128 13860 22102
rect 13780 21100 13860 21128
rect 13728 21082 13780 21088
rect 13636 21072 13688 21078
rect 13636 21014 13688 21020
rect 13280 20590 13584 20618
rect 13358 20496 13414 20505
rect 13358 20431 13414 20440
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13082 19816 13138 19825
rect 13082 19751 13138 19760
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 12995 19468 13032 19496
rect 12900 19440 12952 19446
rect 12995 19428 13023 19468
rect 13096 19446 13124 19654
rect 13084 19440 13136 19446
rect 12995 19400 13032 19428
rect 12900 19382 12952 19388
rect 12532 19304 12584 19310
rect 12530 19272 12532 19281
rect 12584 19272 12586 19281
rect 12530 19207 12586 19216
rect 12544 18970 12572 19207
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12438 18728 12494 18737
rect 12494 18686 12572 18714
rect 12438 18663 12494 18672
rect 12544 18465 12572 18686
rect 12530 18456 12586 18465
rect 12530 18391 12586 18400
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12544 17542 12572 17750
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12360 16510 12480 16538
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 12084 12628 12112 15982
rect 12452 15706 12480 16510
rect 12544 16250 12572 17478
rect 12624 17060 12676 17066
rect 12624 17002 12676 17008
rect 12636 16454 12664 17002
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 14550 12296 15302
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12256 14544 12308 14550
rect 12256 14486 12308 14492
rect 12440 14544 12492 14550
rect 12440 14486 12492 14492
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12176 14074 12204 14350
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12452 13938 12480 14486
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12544 13802 12572 14758
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13252 12400 13258
rect 12348 13194 12400 13200
rect 12360 13025 12388 13194
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12256 12776 12308 12782
rect 12308 12736 12388 12764
rect 12256 12718 12308 12724
rect 12084 12600 12296 12628
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11558 12112 11766
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 11286 12112 11494
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12070 10976 12126 10985
rect 12070 10911 12126 10920
rect 12084 10033 12112 10911
rect 12070 10024 12126 10033
rect 12070 9959 12126 9968
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 8022 12112 8774
rect 12072 8016 12124 8022
rect 12072 7958 12124 7964
rect 12084 7002 12112 7958
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12084 6905 12112 6938
rect 12070 6896 12126 6905
rect 12070 6831 12126 6840
rect 12176 4672 12204 12174
rect 12268 10713 12296 12600
rect 12254 10704 12310 10713
rect 12254 10639 12310 10648
rect 12360 9722 12388 12736
rect 12452 12209 12480 13330
rect 12636 13326 12664 16390
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12728 12628 12756 19366
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12820 18834 12848 19314
rect 12912 18902 12940 19382
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12820 18154 12848 18770
rect 12912 18290 12940 18838
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12808 18148 12860 18154
rect 12808 18090 12860 18096
rect 12808 17740 12860 17746
rect 12808 17682 12860 17688
rect 12820 16794 12848 17682
rect 12898 17232 12954 17241
rect 12898 17167 12954 17176
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12912 14074 12940 17167
rect 13004 16114 13032 19400
rect 13084 19382 13136 19388
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 13096 18426 13124 18770
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13096 15994 13124 18226
rect 13004 15966 13124 15994
rect 13004 14618 13032 15966
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12806 13968 12862 13977
rect 12806 13903 12862 13912
rect 12992 13932 13044 13938
rect 12820 13394 12848 13903
rect 12992 13874 13044 13880
rect 12900 13864 12952 13870
rect 12898 13832 12900 13841
rect 12952 13832 12954 13841
rect 12898 13767 12954 13776
rect 13004 13462 13032 13874
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12992 13320 13044 13326
rect 13096 13297 13124 14758
rect 12992 13262 13044 13268
rect 13082 13288 13138 13297
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12728 12600 12848 12628
rect 12438 12200 12494 12209
rect 12494 12158 12756 12186
rect 12438 12135 12494 12144
rect 12440 12096 12492 12102
rect 12440 12038 12492 12044
rect 12452 11642 12480 12038
rect 12622 11928 12678 11937
rect 12622 11863 12678 11872
rect 12452 11626 12572 11642
rect 12452 11620 12584 11626
rect 12452 11614 12532 11620
rect 12452 11150 12480 11614
rect 12532 11562 12584 11568
rect 12636 11393 12664 11863
rect 12622 11384 12678 11393
rect 12622 11319 12678 11328
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12544 10266 12572 11154
rect 12636 10810 12664 11319
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9722 12480 9998
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12544 9586 12572 10066
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8090 12388 8842
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12268 5710 12296 6802
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12360 5370 12388 5714
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12084 4644 12204 4672
rect 12084 2417 12112 4644
rect 12360 4622 12388 4762
rect 12348 4616 12400 4622
rect 12176 4564 12348 4570
rect 12176 4558 12400 4564
rect 12176 4542 12388 4558
rect 12176 3738 12204 4542
rect 12348 4276 12400 4282
rect 12348 4218 12400 4224
rect 12360 4049 12388 4218
rect 12346 4040 12402 4049
rect 12346 3975 12402 3984
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12452 3369 12480 8910
rect 12544 6458 12572 9522
rect 12636 8634 12664 9522
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12544 5642 12572 6054
rect 12622 5944 12678 5953
rect 12622 5879 12624 5888
rect 12676 5879 12678 5888
rect 12624 5850 12676 5856
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 12544 5030 12572 5578
rect 12622 5400 12678 5409
rect 12622 5335 12678 5344
rect 12636 5148 12664 5335
rect 12728 5250 12756 12158
rect 12820 11642 12848 12600
rect 12912 12209 12940 12922
rect 12898 12200 12954 12209
rect 12898 12135 12954 12144
rect 12912 11801 12940 12135
rect 12898 11792 12954 11801
rect 12898 11727 12954 11736
rect 12820 11614 12940 11642
rect 12808 10124 12860 10130
rect 12912 10112 12940 11614
rect 13004 10849 13032 13262
rect 13082 13223 13138 13232
rect 13096 11370 13124 13223
rect 13188 12866 13216 20198
rect 13266 20088 13322 20097
rect 13266 20023 13322 20032
rect 13280 19378 13308 20023
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13280 18970 13308 19314
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13372 18222 13400 20431
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 18426 13492 20334
rect 13556 19258 13584 20590
rect 13648 20058 13676 21014
rect 13636 20052 13688 20058
rect 13636 19994 13688 20000
rect 13820 19780 13872 19786
rect 13820 19722 13872 19728
rect 13832 19666 13860 19722
rect 13740 19638 13860 19666
rect 13556 19230 13676 19258
rect 13740 19242 13768 19638
rect 13544 19168 13596 19174
rect 13544 19110 13596 19116
rect 13556 18630 13584 19110
rect 13648 18766 13676 19230
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13360 18216 13412 18222
rect 13360 18158 13412 18164
rect 13648 18086 13676 18702
rect 13728 18624 13780 18630
rect 13780 18584 13860 18612
rect 13728 18566 13780 18572
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13280 17241 13308 17614
rect 13266 17232 13322 17241
rect 13266 17167 13322 17176
rect 13268 16584 13320 16590
rect 13268 16526 13320 16532
rect 13280 16017 13308 16526
rect 13266 16008 13322 16017
rect 13266 15943 13322 15952
rect 13280 15638 13308 15943
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 13372 15450 13400 18022
rect 13832 17882 13860 18584
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13648 17066 13676 17614
rect 13636 17060 13688 17066
rect 13636 17002 13688 17008
rect 13452 16720 13504 16726
rect 13452 16662 13504 16668
rect 13280 15422 13400 15450
rect 13464 15434 13492 16662
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13452 15428 13504 15434
rect 13280 13734 13308 15422
rect 13452 15370 13504 15376
rect 13360 15360 13412 15366
rect 13464 15337 13492 15370
rect 13360 15302 13412 15308
rect 13450 15328 13506 15337
rect 13372 14890 13400 15302
rect 13450 15263 13506 15272
rect 13556 15162 13584 15642
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13280 12986 13308 13262
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13188 12838 13308 12866
rect 13176 12640 13228 12646
rect 13174 12608 13176 12617
rect 13228 12608 13230 12617
rect 13174 12543 13230 12552
rect 13188 12238 13216 12543
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11529 13216 12038
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13096 11342 13216 11370
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12990 10840 13046 10849
rect 12990 10775 13046 10784
rect 13096 10674 13124 11222
rect 13188 10713 13216 11342
rect 13174 10704 13230 10713
rect 13084 10668 13136 10674
rect 13174 10639 13230 10648
rect 13084 10610 13136 10616
rect 13280 10248 13308 12838
rect 12860 10084 12940 10112
rect 13188 10220 13308 10248
rect 12808 10066 12860 10072
rect 13084 10056 13136 10062
rect 13084 9998 13136 10004
rect 13096 9722 13124 9998
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12820 8974 12848 9318
rect 13188 9178 13216 10220
rect 13372 10112 13400 14554
rect 13464 14074 13492 14962
rect 13542 14920 13598 14929
rect 13648 14906 13676 17002
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13832 16810 13860 16934
rect 13740 16782 13860 16810
rect 13740 16590 13768 16782
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13740 16250 13768 16526
rect 13832 16425 13860 16594
rect 13818 16416 13874 16425
rect 13818 16351 13874 16360
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13726 15736 13782 15745
rect 13726 15671 13782 15680
rect 13740 15638 13768 15671
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13740 15348 13768 15574
rect 13832 15473 13860 15846
rect 13818 15464 13874 15473
rect 13818 15399 13874 15408
rect 13740 15320 13860 15348
rect 13832 15026 13860 15320
rect 13924 15162 13952 22646
rect 14016 22030 14044 23802
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14004 20256 14056 20262
rect 14004 20198 14056 20204
rect 14016 19825 14044 20198
rect 14002 19816 14058 19825
rect 14002 19751 14058 19760
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 14016 17814 14044 18226
rect 14108 18154 14136 24550
rect 14200 21418 14228 25735
rect 14292 24857 14320 27520
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14278 24848 14334 24857
rect 14384 24818 14412 25094
rect 14278 24783 14334 24792
rect 14372 24812 14424 24818
rect 14372 24754 14424 24760
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14476 24342 14504 24550
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14278 23080 14334 23089
rect 14278 23015 14334 23024
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 14292 21146 14320 23015
rect 14384 21690 14412 24210
rect 14476 24070 14504 24278
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14476 23866 14504 24006
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14660 23633 14688 24550
rect 14646 23624 14702 23633
rect 14646 23559 14702 23568
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22574 14504 22918
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14556 22160 14608 22166
rect 14476 22120 14556 22148
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14384 21593 14412 21626
rect 14370 21584 14426 21593
rect 14370 21519 14426 21528
rect 14476 21350 14504 22120
rect 14556 22102 14608 22108
rect 14660 22001 14688 22510
rect 14646 21992 14702 22001
rect 14568 21950 14646 21978
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14278 20904 14334 20913
rect 14278 20839 14334 20848
rect 14186 20632 14242 20641
rect 14186 20567 14242 20576
rect 14096 18148 14148 18154
rect 14096 18090 14148 18096
rect 14108 17814 14136 18090
rect 14004 17808 14056 17814
rect 14004 17750 14056 17756
rect 14096 17808 14148 17814
rect 14096 17750 14148 17756
rect 14200 17762 14228 20567
rect 14292 19310 14320 20839
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14384 20369 14412 20538
rect 14370 20360 14426 20369
rect 14476 20346 14504 21082
rect 14568 20466 14596 21950
rect 14646 21927 14702 21936
rect 14752 21010 14780 25094
rect 14844 24274 14872 27520
rect 15396 25786 15424 27520
rect 15396 25758 15976 25786
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 14956 25052 15252 25072
rect 15012 25050 15036 25052
rect 15092 25050 15116 25052
rect 15172 25050 15196 25052
rect 15034 24998 15036 25050
rect 15098 24998 15110 25050
rect 15172 24998 15174 25050
rect 15012 24996 15036 24998
rect 15092 24996 15116 24998
rect 15172 24996 15196 24998
rect 14956 24976 15252 24996
rect 15304 24886 15332 25298
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15016 24880 15068 24886
rect 15292 24880 15344 24886
rect 15068 24840 15240 24868
rect 15016 24822 15068 24828
rect 15212 24342 15240 24840
rect 15292 24822 15344 24828
rect 15108 24336 15160 24342
rect 15106 24304 15108 24313
rect 15200 24336 15252 24342
rect 15160 24304 15162 24313
rect 14832 24268 14884 24274
rect 15200 24278 15252 24284
rect 15106 24239 15162 24248
rect 15292 24268 15344 24274
rect 14832 24210 14884 24216
rect 15292 24210 15344 24216
rect 14830 24168 14886 24177
rect 14830 24103 14832 24112
rect 14884 24103 14886 24112
rect 14832 24074 14884 24080
rect 14956 23964 15252 23984
rect 15012 23962 15036 23964
rect 15092 23962 15116 23964
rect 15172 23962 15196 23964
rect 15034 23910 15036 23962
rect 15098 23910 15110 23962
rect 15172 23910 15174 23962
rect 15012 23908 15036 23910
rect 15092 23908 15116 23910
rect 15172 23908 15196 23910
rect 14956 23888 15252 23908
rect 15200 23792 15252 23798
rect 15198 23760 15200 23769
rect 15252 23760 15254 23769
rect 15304 23746 15332 24210
rect 15254 23718 15332 23746
rect 15198 23695 15254 23704
rect 15396 23186 15424 25230
rect 15488 24410 15516 25638
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 15752 24812 15804 24818
rect 15752 24754 15804 24760
rect 15660 24608 15712 24614
rect 15660 24550 15712 24556
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15474 23352 15530 23361
rect 15580 23322 15608 23598
rect 15474 23287 15530 23296
rect 15568 23316 15620 23322
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 14956 22876 15252 22896
rect 15012 22874 15036 22876
rect 15092 22874 15116 22876
rect 15172 22874 15196 22876
rect 15034 22822 15036 22874
rect 15098 22822 15110 22874
rect 15172 22822 15174 22874
rect 15012 22820 15036 22822
rect 15092 22820 15116 22822
rect 15172 22820 15196 22822
rect 14956 22800 15252 22820
rect 15396 22817 15424 23122
rect 15488 22953 15516 23287
rect 15568 23258 15620 23264
rect 15474 22944 15530 22953
rect 15474 22879 15530 22888
rect 15382 22808 15438 22817
rect 15580 22778 15608 23258
rect 15382 22743 15438 22752
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15568 22636 15620 22642
rect 15568 22578 15620 22584
rect 15292 22432 15344 22438
rect 15292 22374 15344 22380
rect 15304 22030 15332 22374
rect 15292 22024 15344 22030
rect 15292 21966 15344 21972
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 21146 14872 21830
rect 14956 21788 15252 21808
rect 15012 21786 15036 21788
rect 15092 21786 15116 21788
rect 15172 21786 15196 21788
rect 15034 21734 15036 21786
rect 15098 21734 15110 21786
rect 15172 21734 15174 21786
rect 15012 21732 15036 21734
rect 15092 21732 15116 21734
rect 15172 21732 15196 21734
rect 14956 21712 15252 21732
rect 15304 21486 15332 21966
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 15212 21026 15240 21286
rect 14740 21004 14792 21010
rect 15212 20998 15332 21026
rect 14740 20946 14792 20952
rect 14648 20800 14700 20806
rect 14648 20742 14700 20748
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14476 20330 14596 20346
rect 14476 20324 14608 20330
rect 14476 20318 14556 20324
rect 14370 20295 14426 20304
rect 14556 20266 14608 20272
rect 14372 20256 14424 20262
rect 14660 20210 14688 20742
rect 14372 20198 14424 20204
rect 14384 19786 14412 20198
rect 14476 20182 14688 20210
rect 14372 19780 14424 19786
rect 14372 19722 14424 19728
rect 14476 19718 14504 20182
rect 14752 20074 14780 20946
rect 14832 20800 14884 20806
rect 14832 20742 14884 20748
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14660 20046 14780 20074
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14476 19378 14504 19654
rect 14568 19514 14596 19994
rect 14556 19508 14608 19514
rect 14556 19450 14608 19456
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14292 18222 14320 19246
rect 14568 18766 14596 19450
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14280 18216 14332 18222
rect 14384 18193 14412 18566
rect 14568 18426 14596 18702
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14280 18158 14332 18164
rect 14370 18184 14426 18193
rect 14370 18119 14426 18128
rect 14200 17734 14320 17762
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14016 16114 14044 17614
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 14004 16108 14056 16114
rect 14004 16050 14056 16056
rect 14002 16008 14058 16017
rect 14002 15943 14004 15952
rect 14056 15943 14058 15952
rect 14004 15914 14056 15920
rect 14004 15496 14056 15502
rect 14004 15438 14056 15444
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 14016 15094 14044 15438
rect 14108 15314 14136 17478
rect 14186 17096 14242 17105
rect 14186 17031 14242 17040
rect 14200 16794 14228 17031
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14108 15286 14228 15314
rect 14094 15192 14150 15201
rect 14094 15127 14150 15136
rect 14004 15088 14056 15094
rect 14004 15030 14056 15036
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13598 14878 13676 14906
rect 13728 14884 13780 14890
rect 13542 14855 13598 14864
rect 13556 14618 13584 14855
rect 13728 14826 13780 14832
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13740 14362 13768 14826
rect 14016 14464 14044 15030
rect 14108 14618 14136 15127
rect 14200 14958 14228 15286
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14016 14436 14136 14464
rect 13740 14334 14044 14362
rect 13452 14068 13504 14074
rect 13452 14010 13504 14016
rect 13464 13938 13492 14010
rect 13452 13932 13504 13938
rect 13452 13874 13504 13880
rect 13464 13326 13492 13874
rect 13820 13864 13872 13870
rect 13820 13806 13872 13812
rect 13728 13796 13780 13802
rect 13728 13738 13780 13744
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13452 13320 13504 13326
rect 13452 13262 13504 13268
rect 13464 12918 13492 13262
rect 13452 12912 13504 12918
rect 13452 12854 13504 12860
rect 13648 12850 13676 13466
rect 13740 12866 13768 13738
rect 13832 12986 13860 13806
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13297 13952 13670
rect 13910 13288 13966 13297
rect 13910 13223 13966 13232
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13636 12844 13688 12850
rect 13740 12838 13860 12866
rect 13636 12786 13688 12792
rect 13542 12744 13598 12753
rect 13542 12679 13598 12688
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13280 10084 13400 10112
rect 13280 9382 13308 10084
rect 13464 10044 13492 12582
rect 13556 12306 13584 12679
rect 13728 12368 13780 12374
rect 13726 12336 13728 12345
rect 13832 12356 13860 12838
rect 13780 12336 13782 12345
rect 13832 12328 13952 12356
rect 13544 12300 13596 12306
rect 13726 12271 13782 12280
rect 13544 12242 13596 12248
rect 13556 11898 13584 12242
rect 13636 12232 13688 12238
rect 13636 12174 13688 12180
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13648 11626 13676 12174
rect 13636 11620 13688 11626
rect 13636 11562 13688 11568
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10674 13584 11154
rect 13648 10985 13676 11562
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13832 11286 13860 11494
rect 13820 11280 13872 11286
rect 13820 11222 13872 11228
rect 13726 11112 13782 11121
rect 13726 11047 13728 11056
rect 13780 11047 13782 11056
rect 13728 11018 13780 11024
rect 13634 10976 13690 10985
rect 13634 10911 13690 10920
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13372 10016 13492 10044
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13176 9172 13228 9178
rect 13176 9114 13228 9120
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 13188 8634 13216 9114
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13082 8256 13138 8265
rect 13082 8191 13138 8200
rect 12806 6760 12862 6769
rect 12806 6695 12808 6704
rect 12860 6695 12862 6704
rect 12808 6666 12860 6672
rect 12728 5222 13032 5250
rect 12636 5120 12940 5148
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12256 2644 12308 2650
rect 12256 2586 12308 2592
rect 12268 2417 12296 2586
rect 12070 2408 12126 2417
rect 12070 2343 12126 2352
rect 12254 2408 12310 2417
rect 12254 2343 12310 2352
rect 12070 1864 12126 1873
rect 12070 1799 12126 1808
rect 12084 1630 12112 1799
rect 12072 1624 12124 1630
rect 12072 1566 12124 1572
rect 12452 1465 12480 3062
rect 12544 2854 12572 4966
rect 12622 4856 12678 4865
rect 12622 4791 12624 4800
rect 12676 4791 12678 4800
rect 12624 4762 12676 4768
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12624 4072 12676 4078
rect 12622 4040 12624 4049
rect 12676 4040 12678 4049
rect 12622 3975 12678 3984
rect 12624 3936 12676 3942
rect 12728 3924 12756 4626
rect 12676 3896 12756 3924
rect 12806 3904 12862 3913
rect 12624 3878 12676 3884
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 2650 12572 2790
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12636 2009 12664 3878
rect 12806 3839 12862 3848
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 2553 12756 3674
rect 12820 3369 12848 3839
rect 12806 3360 12862 3369
rect 12806 3295 12862 3304
rect 12714 2544 12770 2553
rect 12714 2479 12770 2488
rect 12912 2106 12940 5120
rect 12900 2100 12952 2106
rect 12900 2042 12952 2048
rect 12622 2000 12678 2009
rect 12622 1935 12678 1944
rect 12530 1864 12586 1873
rect 12530 1799 12586 1808
rect 12544 1630 12572 1799
rect 12532 1624 12584 1630
rect 12532 1566 12584 1572
rect 12438 1456 12494 1465
rect 12438 1391 12494 1400
rect 11992 1142 12296 1170
rect 11886 1048 11942 1057
rect 11886 983 11942 992
rect 12268 480 12296 1142
rect 13004 898 13032 5222
rect 13096 5098 13124 8191
rect 13188 5409 13216 8570
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13280 5914 13308 6734
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13174 5400 13230 5409
rect 13174 5335 13230 5344
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 13188 4622 13216 5102
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13176 4616 13228 4622
rect 13174 4584 13176 4593
rect 13228 4584 13230 4593
rect 13174 4519 13230 4528
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3777 13124 4014
rect 13176 3936 13228 3942
rect 13174 3904 13176 3913
rect 13228 3904 13230 3913
rect 13174 3839 13230 3848
rect 13082 3768 13138 3777
rect 13188 3738 13216 3839
rect 13082 3703 13138 3712
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 13174 2680 13230 2689
rect 13174 2615 13230 2624
rect 13188 2582 13216 2615
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 2038 13308 4966
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 12820 870 13032 898
rect 12820 480 12848 870
rect 13372 480 13400 10016
rect 13452 9920 13504 9926
rect 13450 9888 13452 9897
rect 13504 9888 13506 9897
rect 13450 9823 13506 9832
rect 13556 9330 13584 10610
rect 13740 10606 13768 11018
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13832 10742 13860 10950
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13728 10464 13780 10470
rect 13780 10412 13860 10418
rect 13728 10406 13860 10412
rect 13740 10390 13860 10406
rect 13634 10296 13690 10305
rect 13634 10231 13690 10240
rect 13648 9926 13676 10231
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13464 9302 13584 9330
rect 13464 8294 13492 9302
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13556 9110 13584 9143
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13556 8634 13584 9046
rect 13740 8974 13768 9522
rect 13832 9110 13860 10390
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13728 8832 13780 8838
rect 13728 8774 13780 8780
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13740 8362 13768 8774
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13636 8288 13688 8294
rect 13636 8230 13688 8236
rect 13464 8090 13492 8230
rect 13452 8084 13504 8090
rect 13504 8044 13584 8072
rect 13452 8026 13504 8032
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7342 13492 7686
rect 13556 7546 13584 8044
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13450 5808 13506 5817
rect 13450 5743 13506 5752
rect 13464 4049 13492 5743
rect 13648 5273 13676 8230
rect 13740 6118 13768 8298
rect 13924 8090 13952 12328
rect 14016 9178 14044 14334
rect 14108 13530 14136 14436
rect 14292 14346 14320 17734
rect 14554 17504 14610 17513
rect 14554 17439 14610 17448
rect 14568 16794 14596 17439
rect 14556 16788 14608 16794
rect 14556 16730 14608 16736
rect 14370 16144 14426 16153
rect 14370 16079 14426 16088
rect 14384 15706 14412 16079
rect 14464 16040 14516 16046
rect 14464 15982 14516 15988
rect 14372 15700 14424 15706
rect 14372 15642 14424 15648
rect 14476 15042 14504 15982
rect 14660 15586 14688 20046
rect 14844 19242 14872 20742
rect 14956 20700 15252 20720
rect 15012 20698 15036 20700
rect 15092 20698 15116 20700
rect 15172 20698 15196 20700
rect 15034 20646 15036 20698
rect 15098 20646 15110 20698
rect 15172 20646 15174 20698
rect 15012 20644 15036 20646
rect 15092 20644 15116 20646
rect 15172 20644 15196 20646
rect 14956 20624 15252 20644
rect 14924 20528 14976 20534
rect 14922 20496 14924 20505
rect 14976 20496 14978 20505
rect 14922 20431 14978 20440
rect 15106 20496 15162 20505
rect 15304 20482 15332 20998
rect 15106 20431 15162 20440
rect 15212 20454 15332 20482
rect 15120 20058 15148 20431
rect 15212 20262 15240 20454
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 15212 20097 15240 20198
rect 15198 20088 15254 20097
rect 15108 20052 15160 20058
rect 15198 20023 15254 20032
rect 15108 19994 15160 20000
rect 15120 19802 15148 19994
rect 15120 19774 15332 19802
rect 14956 19612 15252 19632
rect 15012 19610 15036 19612
rect 15092 19610 15116 19612
rect 15172 19610 15196 19612
rect 15034 19558 15036 19610
rect 15098 19558 15110 19610
rect 15172 19558 15174 19610
rect 15012 19556 15036 19558
rect 15092 19556 15116 19558
rect 15172 19556 15196 19558
rect 14956 19536 15252 19556
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14936 18612 14964 19314
rect 15304 19242 15332 19774
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 14844 18584 14964 18612
rect 14738 18456 14794 18465
rect 14738 18391 14794 18400
rect 14752 18193 14780 18391
rect 14738 18184 14794 18193
rect 14738 18119 14794 18128
rect 14844 16794 14872 18584
rect 14956 18524 15252 18544
rect 15012 18522 15036 18524
rect 15092 18522 15116 18524
rect 15172 18522 15196 18524
rect 15034 18470 15036 18522
rect 15098 18470 15110 18522
rect 15172 18470 15174 18522
rect 15012 18468 15036 18470
rect 15092 18468 15116 18470
rect 15172 18468 15196 18470
rect 14956 18448 15252 18468
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15120 17678 15148 18158
rect 15108 17672 15160 17678
rect 15108 17614 15160 17620
rect 14956 17436 15252 17456
rect 15012 17434 15036 17436
rect 15092 17434 15116 17436
rect 15172 17434 15196 17436
rect 15034 17382 15036 17434
rect 15098 17382 15110 17434
rect 15172 17382 15174 17434
rect 15012 17380 15036 17382
rect 15092 17380 15116 17382
rect 15172 17380 15196 17382
rect 14956 17360 15252 17380
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14924 16720 14976 16726
rect 14922 16688 14924 16697
rect 14976 16688 14978 16697
rect 14922 16623 14978 16632
rect 14738 16552 14794 16561
rect 15120 16538 15148 16934
rect 15304 16674 15332 18770
rect 15396 18057 15424 21490
rect 15580 20788 15608 22578
rect 15672 20913 15700 24550
rect 15764 24070 15792 24754
rect 15856 24750 15884 25094
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15948 24449 15976 25758
rect 15934 24440 15990 24449
rect 15934 24375 15990 24384
rect 15752 24064 15804 24070
rect 15752 24006 15804 24012
rect 15764 22642 15792 24006
rect 16040 23712 16068 27520
rect 16592 26246 16620 27520
rect 16580 26240 16632 26246
rect 16580 26182 16632 26188
rect 17144 25480 17172 27520
rect 17408 26172 17460 26178
rect 17408 26114 17460 26120
rect 17052 25452 17172 25480
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 15856 23684 16068 23712
rect 15752 22636 15804 22642
rect 15752 22578 15804 22584
rect 15752 22160 15804 22166
rect 15752 22102 15804 22108
rect 15764 21434 15792 22102
rect 15856 21554 15884 23684
rect 15934 23624 15990 23633
rect 16132 23576 16160 25094
rect 16486 24984 16542 24993
rect 16486 24919 16542 24928
rect 16396 24880 16448 24886
rect 16396 24822 16448 24828
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 15934 23559 15990 23568
rect 15948 23050 15976 23559
rect 16040 23548 16160 23576
rect 15936 23044 15988 23050
rect 15936 22986 15988 22992
rect 15934 22944 15990 22953
rect 15934 22879 15990 22888
rect 15948 22273 15976 22879
rect 15934 22264 15990 22273
rect 15934 22199 15990 22208
rect 15936 22092 15988 22098
rect 15936 22034 15988 22040
rect 15844 21548 15896 21554
rect 15844 21490 15896 21496
rect 15764 21406 15884 21434
rect 15752 20936 15804 20942
rect 15658 20904 15714 20913
rect 15752 20878 15804 20884
rect 15658 20839 15714 20848
rect 15580 20760 15700 20788
rect 15474 20632 15530 20641
rect 15474 20567 15530 20576
rect 15488 20534 15516 20567
rect 15476 20528 15528 20534
rect 15476 20470 15528 20476
rect 15566 19680 15622 19689
rect 15566 19615 15622 19624
rect 15580 19310 15608 19615
rect 15568 19304 15620 19310
rect 15672 19281 15700 20760
rect 15764 20398 15792 20878
rect 15752 20392 15804 20398
rect 15752 20334 15804 20340
rect 15856 20244 15884 21406
rect 15948 21350 15976 22034
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 20942 15976 21286
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15764 20216 15884 20244
rect 15568 19246 15620 19252
rect 15658 19272 15714 19281
rect 15580 18970 15608 19246
rect 15658 19207 15714 19216
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15476 18828 15528 18834
rect 15476 18770 15528 18776
rect 15488 18086 15516 18770
rect 15658 18456 15714 18465
rect 15658 18391 15714 18400
rect 15476 18080 15528 18086
rect 15382 18048 15438 18057
rect 15476 18022 15528 18028
rect 15382 17983 15438 17992
rect 15382 17640 15438 17649
rect 15382 17575 15438 17584
rect 15396 17202 15424 17575
rect 15488 17542 15516 18022
rect 15568 17808 15620 17814
rect 15568 17750 15620 17756
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15488 16998 15516 17478
rect 15580 17270 15608 17750
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15304 16646 15424 16674
rect 15120 16510 15332 16538
rect 14738 16487 14794 16496
rect 14752 15706 14780 16487
rect 14956 16348 15252 16368
rect 15012 16346 15036 16348
rect 15092 16346 15116 16348
rect 15172 16346 15196 16348
rect 15034 16294 15036 16346
rect 15098 16294 15110 16346
rect 15172 16294 15174 16346
rect 15012 16292 15036 16294
rect 15092 16292 15116 16294
rect 15172 16292 15196 16294
rect 14956 16272 15252 16292
rect 15304 15978 15332 16510
rect 15292 15972 15344 15978
rect 15292 15914 15344 15920
rect 15016 15904 15068 15910
rect 14830 15872 14886 15881
rect 15200 15904 15252 15910
rect 15016 15846 15068 15852
rect 15198 15872 15200 15881
rect 15252 15872 15254 15881
rect 14830 15807 14886 15816
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14660 15558 14780 15586
rect 14384 15014 14504 15042
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14188 13728 14240 13734
rect 14384 13705 14412 15014
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14188 13670 14240 13676
rect 14370 13696 14426 13705
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14108 12986 14136 13330
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12714 14228 13670
rect 14370 13631 14426 13640
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14384 12646 14412 13631
rect 14476 12866 14504 14894
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14568 14385 14596 14486
rect 14554 14376 14610 14385
rect 14554 14311 14610 14320
rect 14554 13560 14610 13569
rect 14554 13495 14556 13504
rect 14608 13495 14610 13504
rect 14556 13466 14608 13472
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14568 13002 14596 13330
rect 14648 13184 14700 13190
rect 14646 13152 14648 13161
rect 14700 13152 14702 13161
rect 14646 13087 14702 13096
rect 14568 12974 14688 13002
rect 14476 12838 14596 12866
rect 14660 12850 14688 12974
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14568 12345 14596 12838
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14660 12442 14688 12786
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14554 12336 14610 12345
rect 14554 12271 14610 12280
rect 14096 12164 14148 12170
rect 14096 12106 14148 12112
rect 14108 11354 14136 12106
rect 14280 12096 14332 12102
rect 14278 12064 14280 12073
rect 14332 12064 14334 12073
rect 14278 11999 14334 12008
rect 14200 11830 14228 11861
rect 14188 11824 14240 11830
rect 14186 11792 14188 11801
rect 14240 11792 14242 11801
rect 14186 11727 14242 11736
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14108 10674 14136 11290
rect 14096 10668 14148 10674
rect 14096 10610 14148 10616
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 14200 7936 14228 11727
rect 14752 11354 14780 15558
rect 14844 14618 14872 15807
rect 15028 15609 15056 15846
rect 15198 15807 15254 15816
rect 15014 15600 15070 15609
rect 15014 15535 15070 15544
rect 14956 15260 15252 15280
rect 15012 15258 15036 15260
rect 15092 15258 15116 15260
rect 15172 15258 15196 15260
rect 15034 15206 15036 15258
rect 15098 15206 15110 15258
rect 15172 15206 15174 15258
rect 15012 15204 15036 15206
rect 15092 15204 15116 15206
rect 15172 15204 15196 15206
rect 14956 15184 15252 15204
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 15108 14544 15160 14550
rect 15396 14532 15424 16646
rect 15488 16402 15516 16934
rect 15488 16374 15608 16402
rect 15474 16280 15530 16289
rect 15474 16215 15530 16224
rect 15160 14504 15424 14532
rect 15108 14486 15160 14492
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 14956 14172 15252 14192
rect 15012 14170 15036 14172
rect 15092 14170 15116 14172
rect 15172 14170 15196 14172
rect 15034 14118 15036 14170
rect 15098 14118 15110 14170
rect 15172 14118 15174 14170
rect 15012 14116 15036 14118
rect 15092 14116 15116 14118
rect 15172 14116 15196 14118
rect 14956 14096 15252 14116
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 13569 14964 13806
rect 14922 13560 14978 13569
rect 14922 13495 14978 13504
rect 14830 13288 14886 13297
rect 14830 13223 14832 13232
rect 14884 13223 14886 13232
rect 14832 13194 14884 13200
rect 14844 12782 14872 13194
rect 14956 13084 15252 13104
rect 15012 13082 15036 13084
rect 15092 13082 15116 13084
rect 15172 13082 15196 13084
rect 15034 13030 15036 13082
rect 15098 13030 15110 13082
rect 15172 13030 15174 13082
rect 15012 13028 15036 13030
rect 15092 13028 15116 13030
rect 15172 13028 15196 13030
rect 14956 13008 15252 13028
rect 15304 12986 15332 14350
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15016 12640 15068 12646
rect 15014 12608 15016 12617
rect 15068 12608 15070 12617
rect 15014 12543 15070 12552
rect 14832 12436 14884 12442
rect 14832 12378 14884 12384
rect 14740 11348 14792 11354
rect 14740 11290 14792 11296
rect 14648 11280 14700 11286
rect 14646 11248 14648 11257
rect 14700 11248 14702 11257
rect 14646 11183 14702 11192
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14278 9208 14334 9217
rect 14278 9143 14334 9152
rect 13924 7908 14228 7936
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13832 7002 13860 7686
rect 13820 6996 13872 7002
rect 13820 6938 13872 6944
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13726 5944 13782 5953
rect 13726 5879 13782 5888
rect 13740 5778 13768 5879
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13832 5658 13860 6938
rect 13740 5630 13860 5658
rect 13634 5264 13690 5273
rect 13634 5199 13690 5208
rect 13740 5148 13768 5630
rect 13556 5120 13768 5148
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 13450 2816 13506 2825
rect 13450 2751 13506 2760
rect 13464 2650 13492 2751
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13556 2145 13584 5120
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13648 4214 13676 4422
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13740 4078 13768 4490
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13740 3738 13768 4014
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13648 3097 13676 3334
rect 13740 3194 13768 3334
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13634 3088 13690 3097
rect 13634 3023 13690 3032
rect 13832 2961 13860 3130
rect 13818 2952 13874 2961
rect 13728 2916 13780 2922
rect 13818 2887 13874 2896
rect 13728 2858 13780 2864
rect 13740 2666 13768 2858
rect 13740 2650 13860 2666
rect 13740 2644 13872 2650
rect 13740 2638 13820 2644
rect 13820 2586 13872 2592
rect 13542 2136 13598 2145
rect 13542 2071 13598 2080
rect 13924 480 13952 7908
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6254 14136 6734
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14108 5914 14136 6190
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 14200 5370 14228 7754
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14200 5166 14228 5306
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 14292 4826 14320 9143
rect 14384 7818 14412 10950
rect 14462 10840 14518 10849
rect 14462 10775 14518 10784
rect 14476 10062 14504 10775
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 10305 14596 10542
rect 14554 10296 14610 10305
rect 14554 10231 14556 10240
rect 14608 10231 14610 10240
rect 14556 10202 14608 10208
rect 14568 10171 14596 10202
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14476 8634 14504 9998
rect 14648 9036 14700 9042
rect 14648 8978 14700 8984
rect 14660 8809 14688 8978
rect 14646 8800 14702 8809
rect 14646 8735 14702 8744
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14752 7857 14780 11154
rect 14738 7848 14794 7857
rect 14372 7812 14424 7818
rect 14738 7783 14794 7792
rect 14372 7754 14424 7760
rect 14738 7576 14794 7585
rect 14738 7511 14794 7520
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14280 4820 14332 4826
rect 14200 4780 14280 4808
rect 14004 4684 14056 4690
rect 14004 4626 14056 4632
rect 14016 3942 14044 4626
rect 14200 4214 14228 4780
rect 14280 4762 14332 4768
rect 14278 4312 14334 4321
rect 14278 4247 14334 4256
rect 14188 4208 14240 4214
rect 14094 4176 14150 4185
rect 14188 4150 14240 4156
rect 14094 4111 14150 4120
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 2961 14044 3878
rect 14108 3670 14136 4111
rect 14292 3942 14320 4247
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3738 14320 3878
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14002 2952 14058 2961
rect 14002 2887 14058 2896
rect 14016 1737 14044 2887
rect 14002 1728 14058 1737
rect 14002 1663 14058 1672
rect 14384 480 14412 7346
rect 14752 6866 14780 7511
rect 14844 7410 14872 12378
rect 14956 11996 15252 12016
rect 15012 11994 15036 11996
rect 15092 11994 15116 11996
rect 15172 11994 15196 11996
rect 15034 11942 15036 11994
rect 15098 11942 15110 11994
rect 15172 11942 15174 11994
rect 15012 11940 15036 11942
rect 15092 11940 15116 11942
rect 15172 11940 15196 11942
rect 14956 11920 15252 11940
rect 15290 11248 15346 11257
rect 15290 11183 15292 11192
rect 15344 11183 15346 11192
rect 15292 11154 15344 11160
rect 14956 10908 15252 10928
rect 15012 10906 15036 10908
rect 15092 10906 15116 10908
rect 15172 10906 15196 10908
rect 15034 10854 15036 10906
rect 15098 10854 15110 10906
rect 15172 10854 15174 10906
rect 15012 10852 15036 10854
rect 15092 10852 15116 10854
rect 15172 10852 15196 10854
rect 14956 10832 15252 10852
rect 15198 10704 15254 10713
rect 15198 10639 15254 10648
rect 15212 10266 15240 10639
rect 15382 10568 15438 10577
rect 15382 10503 15438 10512
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 14956 9820 15252 9840
rect 15012 9818 15036 9820
rect 15092 9818 15116 9820
rect 15172 9818 15196 9820
rect 15034 9766 15036 9818
rect 15098 9766 15110 9818
rect 15172 9766 15174 9818
rect 15012 9764 15036 9766
rect 15092 9764 15116 9766
rect 15172 9764 15196 9766
rect 14956 9744 15252 9764
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 9178 15332 9658
rect 15396 9518 15424 10503
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15382 9344 15438 9353
rect 15382 9279 15438 9288
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 14956 8732 15252 8752
rect 15012 8730 15036 8732
rect 15092 8730 15116 8732
rect 15172 8730 15196 8732
rect 15034 8678 15036 8730
rect 15098 8678 15110 8730
rect 15172 8678 15174 8730
rect 15012 8676 15036 8678
rect 15092 8676 15116 8678
rect 15172 8676 15196 8678
rect 14956 8656 15252 8676
rect 15304 8634 15332 9114
rect 15396 9081 15424 9279
rect 15488 9110 15516 16215
rect 15580 15706 15608 16374
rect 15672 15745 15700 18391
rect 15764 17218 15792 20216
rect 15948 19922 15976 20742
rect 16040 20058 16068 23548
rect 16224 23474 16252 24278
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16132 23446 16252 23474
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 15936 19916 15988 19922
rect 15936 19858 15988 19864
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15856 19378 15884 19790
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15948 19174 15976 19858
rect 15936 19168 15988 19174
rect 15934 19136 15936 19145
rect 15988 19136 15990 19145
rect 15934 19071 15990 19080
rect 15948 19045 15976 19071
rect 16040 18970 16068 19994
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 16132 18698 16160 23446
rect 16316 23338 16344 23734
rect 16224 23310 16344 23338
rect 16224 20942 16252 23310
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16316 21690 16344 22918
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16304 21412 16356 21418
rect 16304 21354 16356 21360
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 15844 18624 15896 18630
rect 15842 18592 15844 18601
rect 15896 18592 15898 18601
rect 15842 18527 15898 18536
rect 15856 18222 15884 18527
rect 16120 18352 16172 18358
rect 16120 18294 16172 18300
rect 15844 18216 15896 18222
rect 16132 18170 16160 18294
rect 15844 18158 15896 18164
rect 16040 18142 16160 18170
rect 16040 17814 16068 18142
rect 16118 18048 16174 18057
rect 16118 17983 16174 17992
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16132 17338 16160 17983
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 15764 17190 16160 17218
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15752 16652 15804 16658
rect 15752 16594 15804 16600
rect 15658 15736 15714 15745
rect 15568 15700 15620 15706
rect 15658 15671 15714 15680
rect 15568 15642 15620 15648
rect 15580 15570 15608 15642
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 14958 15608 15506
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15580 14482 15608 14894
rect 15764 14657 15792 16594
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15948 16250 15976 16526
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15750 14648 15806 14657
rect 15750 14583 15806 14592
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15844 14340 15896 14346
rect 15844 14282 15896 14288
rect 15856 13870 15884 14282
rect 15934 14104 15990 14113
rect 15934 14039 15990 14048
rect 15844 13864 15896 13870
rect 15764 13824 15844 13852
rect 15566 13424 15622 13433
rect 15566 13359 15622 13368
rect 15580 12986 15608 13359
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15764 12442 15792 13824
rect 15844 13806 15896 13812
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13530 15884 13670
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15948 13410 15976 14039
rect 16040 13802 16068 16730
rect 16028 13796 16080 13802
rect 16028 13738 16080 13744
rect 15856 13382 15976 13410
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15580 11286 15608 11630
rect 15672 11626 15700 12038
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15568 11280 15620 11286
rect 15568 11222 15620 11228
rect 15580 10538 15608 11222
rect 15672 10742 15700 11562
rect 15750 11384 15806 11393
rect 15750 11319 15752 11328
rect 15804 11319 15806 11328
rect 15752 11290 15804 11296
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15476 9104 15528 9110
rect 15382 9072 15438 9081
rect 15476 9046 15528 9052
rect 15382 9007 15438 9016
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15488 8514 15516 9046
rect 15580 8838 15608 10474
rect 15672 9722 15700 10678
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9897 15792 9998
rect 15750 9888 15806 9897
rect 15750 9823 15806 9832
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15750 9616 15806 9625
rect 15750 9551 15806 9560
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 15672 8945 15700 9318
rect 15658 8936 15714 8945
rect 15658 8871 15714 8880
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8566 15608 8774
rect 15764 8634 15792 9551
rect 15856 9489 15884 13382
rect 15934 13288 15990 13297
rect 15934 13223 15936 13232
rect 15988 13223 15990 13232
rect 15936 13194 15988 13200
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 16040 10849 16068 12922
rect 16132 10985 16160 17190
rect 16224 15910 16252 20742
rect 16316 16522 16344 21354
rect 16408 17490 16436 24822
rect 16500 23798 16528 24919
rect 16776 24177 16804 25094
rect 16856 24608 16908 24614
rect 16960 24596 16988 25230
rect 16908 24568 16988 24596
rect 16856 24550 16908 24556
rect 16762 24168 16818 24177
rect 16762 24103 16818 24112
rect 16580 24064 16632 24070
rect 16580 24006 16632 24012
rect 16488 23792 16540 23798
rect 16488 23734 16540 23740
rect 16488 23656 16540 23662
rect 16488 23598 16540 23604
rect 16500 23118 16528 23598
rect 16592 23225 16620 24006
rect 16672 23316 16724 23322
rect 16672 23258 16724 23264
rect 16578 23216 16634 23225
rect 16578 23151 16634 23160
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16500 22438 16528 23054
rect 16684 22953 16712 23258
rect 16670 22944 16726 22953
rect 16670 22879 16726 22888
rect 16488 22432 16540 22438
rect 16488 22374 16540 22380
rect 16486 22264 16542 22273
rect 16486 22199 16542 22208
rect 16500 20806 16528 22199
rect 16670 21992 16726 22001
rect 16670 21927 16672 21936
rect 16724 21927 16726 21936
rect 16672 21898 16724 21904
rect 16776 21486 16804 24103
rect 16868 22574 16896 24550
rect 16948 24336 17000 24342
rect 16946 24304 16948 24313
rect 17000 24304 17002 24313
rect 16946 24239 17002 24248
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 16960 23526 16988 24074
rect 16948 23520 17000 23526
rect 16948 23462 17000 23468
rect 16960 23254 16988 23462
rect 17052 23361 17080 25452
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 17144 24750 17172 25298
rect 17224 25288 17276 25294
rect 17224 25230 17276 25236
rect 17236 24750 17264 25230
rect 17132 24744 17184 24750
rect 17130 24712 17132 24721
rect 17224 24744 17276 24750
rect 17184 24712 17186 24721
rect 17224 24686 17276 24692
rect 17130 24647 17186 24656
rect 17130 24440 17186 24449
rect 17130 24375 17186 24384
rect 17038 23352 17094 23361
rect 17038 23287 17094 23296
rect 16948 23248 17000 23254
rect 16948 23190 17000 23196
rect 16856 22568 16908 22574
rect 16854 22536 16856 22545
rect 16908 22536 16910 22545
rect 16854 22471 16910 22480
rect 16960 22098 16988 23190
rect 17038 22808 17094 22817
rect 17038 22743 17040 22752
rect 17092 22743 17094 22752
rect 17040 22714 17092 22720
rect 16948 22092 17000 22098
rect 16948 22034 17000 22040
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16856 21412 16908 21418
rect 16856 21354 16908 21360
rect 16868 21146 16896 21354
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16580 21072 16632 21078
rect 16580 21014 16632 21020
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16592 20618 16620 21014
rect 16960 21010 16988 22034
rect 16948 21004 17000 21010
rect 16948 20946 17000 20952
rect 16500 20602 16620 20618
rect 16488 20596 16620 20602
rect 16540 20590 16620 20596
rect 16488 20538 16540 20544
rect 16762 20496 16818 20505
rect 16960 20466 16988 20946
rect 16762 20431 16818 20440
rect 16948 20460 17000 20466
rect 16776 20398 16804 20431
rect 16948 20402 17000 20408
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16776 20058 16804 20334
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16868 19961 16896 20266
rect 16854 19952 16910 19961
rect 16854 19887 16910 19896
rect 16486 19816 16542 19825
rect 16960 19802 16988 20402
rect 16868 19786 16988 19802
rect 16486 19751 16542 19760
rect 16856 19780 16988 19786
rect 16500 18465 16528 19751
rect 16908 19774 16988 19780
rect 16856 19722 16908 19728
rect 16868 19514 16896 19722
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16960 19310 16988 19654
rect 16948 19304 17000 19310
rect 16946 19272 16948 19281
rect 17000 19272 17002 19281
rect 16946 19207 17002 19216
rect 17040 19236 17092 19242
rect 17040 19178 17092 19184
rect 16486 18456 16542 18465
rect 16486 18391 16542 18400
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16500 18193 16528 18294
rect 16486 18184 16542 18193
rect 16486 18119 16542 18128
rect 16672 17536 16724 17542
rect 16408 17462 16620 17490
rect 16672 17478 16724 17484
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16833 16436 16934
rect 16394 16824 16450 16833
rect 16592 16794 16620 17462
rect 16394 16759 16450 16768
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16684 16561 16712 17478
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16670 16552 16726 16561
rect 16304 16516 16356 16522
rect 16670 16487 16726 16496
rect 16856 16516 16908 16522
rect 16304 16458 16356 16464
rect 16394 16416 16450 16425
rect 16394 16351 16450 16360
rect 16408 16250 16436 16351
rect 16684 16289 16712 16487
rect 16856 16458 16908 16464
rect 16764 16448 16816 16454
rect 16764 16390 16816 16396
rect 16670 16280 16726 16289
rect 16396 16244 16448 16250
rect 16670 16215 16726 16224
rect 16396 16186 16448 16192
rect 16304 16108 16356 16114
rect 16304 16050 16356 16056
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16316 15570 16344 16050
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16304 15564 16356 15570
rect 16304 15506 16356 15512
rect 16210 14920 16266 14929
rect 16210 14855 16266 14864
rect 16224 14074 16252 14855
rect 16316 14618 16344 15506
rect 16578 15056 16634 15065
rect 16578 14991 16634 15000
rect 16488 14884 16540 14890
rect 16488 14826 16540 14832
rect 16304 14612 16356 14618
rect 16304 14554 16356 14560
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16408 14074 16436 14418
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16224 13977 16252 14010
rect 16210 13968 16266 13977
rect 16210 13903 16266 13912
rect 16224 13852 16252 13903
rect 16500 13870 16528 14826
rect 16304 13864 16356 13870
rect 16224 13824 16304 13852
rect 16304 13806 16356 13812
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16316 12986 16344 13330
rect 16500 13326 16528 13806
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16394 12744 16450 12753
rect 16394 12679 16450 12688
rect 16408 12646 16436 12679
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16394 12472 16450 12481
rect 16500 12442 16528 13262
rect 16394 12407 16450 12416
rect 16488 12436 16540 12442
rect 16408 12374 16436 12407
rect 16488 12378 16540 12384
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16592 12102 16620 14991
rect 16684 12714 16712 15846
rect 16776 15162 16804 16390
rect 16868 15910 16896 16458
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16868 14618 16896 14758
rect 16856 14612 16908 14618
rect 16856 14554 16908 14560
rect 16868 14521 16896 14554
rect 16854 14512 16910 14521
rect 16854 14447 16910 14456
rect 16960 14396 16988 16934
rect 16868 14368 16988 14396
rect 16762 12880 16818 12889
rect 16762 12815 16818 12824
rect 16776 12782 16804 12815
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16672 12436 16724 12442
rect 16672 12378 16724 12384
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16224 11801 16252 12038
rect 16210 11792 16266 11801
rect 16210 11727 16266 11736
rect 16684 11234 16712 12378
rect 16868 11898 16896 14368
rect 17052 13977 17080 19178
rect 17038 13968 17094 13977
rect 17038 13903 17094 13912
rect 16946 13832 17002 13841
rect 16946 13767 17002 13776
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16776 11286 16804 11630
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16500 11206 16712 11234
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16118 10976 16174 10985
rect 16118 10911 16174 10920
rect 16026 10840 16082 10849
rect 15948 10798 16026 10826
rect 15948 9654 15976 10798
rect 16026 10775 16082 10784
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15936 9648 15988 9654
rect 15936 9590 15988 9596
rect 15842 9480 15898 9489
rect 15898 9438 15976 9466
rect 15842 9415 15898 9424
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 9081 15884 9318
rect 15842 9072 15898 9081
rect 15842 9007 15898 9016
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15120 8486 15516 8514
rect 15568 8560 15620 8566
rect 15620 8508 15700 8514
rect 15568 8502 15700 8508
rect 15580 8486 15700 8502
rect 15120 8090 15148 8486
rect 15566 8392 15622 8401
rect 15566 8327 15568 8336
rect 15620 8327 15622 8336
rect 15568 8298 15620 8304
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 14956 7644 15252 7664
rect 15012 7642 15036 7644
rect 15092 7642 15116 7644
rect 15172 7642 15196 7644
rect 15034 7590 15036 7642
rect 15098 7590 15110 7642
rect 15172 7590 15174 7642
rect 15012 7588 15036 7590
rect 15092 7588 15116 7590
rect 15172 7588 15196 7590
rect 14956 7568 15252 7588
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14556 6384 14608 6390
rect 14554 6352 14556 6361
rect 14752 6361 14780 6598
rect 14608 6352 14610 6361
rect 14554 6287 14610 6296
rect 14738 6352 14794 6361
rect 14738 6287 14794 6296
rect 14462 6216 14518 6225
rect 14462 6151 14518 6160
rect 14476 6118 14504 6151
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14568 5370 14596 5782
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 4593 14504 4966
rect 14462 4584 14518 4593
rect 14462 4519 14518 4528
rect 14660 4078 14688 6054
rect 14844 5642 14872 7142
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 14922 6896 14978 6905
rect 14922 6831 14978 6840
rect 15120 6848 15148 6938
rect 15200 6860 15252 6866
rect 14936 6798 14964 6831
rect 15120 6820 15200 6848
rect 15200 6802 15252 6808
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15014 6760 15070 6769
rect 15014 6695 15016 6704
rect 15068 6695 15070 6704
rect 15016 6666 15068 6672
rect 14956 6556 15252 6576
rect 15012 6554 15036 6556
rect 15092 6554 15116 6556
rect 15172 6554 15196 6556
rect 15034 6502 15036 6554
rect 15098 6502 15110 6554
rect 15172 6502 15174 6554
rect 15012 6500 15036 6502
rect 15092 6500 15116 6502
rect 15172 6500 15196 6502
rect 14956 6480 15252 6500
rect 15382 6488 15438 6497
rect 15028 6432 15382 6440
rect 15028 6423 15438 6432
rect 15476 6452 15528 6458
rect 15028 6412 15424 6423
rect 15028 5817 15056 6412
rect 15476 6394 15528 6400
rect 15384 6112 15436 6118
rect 15106 6080 15162 6089
rect 15290 6080 15346 6089
rect 15162 6038 15240 6066
rect 15106 6015 15162 6024
rect 15212 5817 15240 6038
rect 15384 6054 15436 6060
rect 15290 6015 15346 6024
rect 15304 5914 15332 6015
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15014 5808 15070 5817
rect 15014 5743 15070 5752
rect 15198 5808 15254 5817
rect 15198 5743 15254 5752
rect 15108 5704 15160 5710
rect 15160 5664 15332 5692
rect 15108 5646 15160 5652
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14752 4146 14780 5510
rect 14844 4826 14872 5578
rect 14956 5468 15252 5488
rect 15012 5466 15036 5468
rect 15092 5466 15116 5468
rect 15172 5466 15196 5468
rect 15034 5414 15036 5466
rect 15098 5414 15110 5466
rect 15172 5414 15174 5466
rect 15012 5412 15036 5414
rect 15092 5412 15116 5414
rect 15172 5412 15196 5414
rect 14956 5392 15252 5412
rect 15108 5092 15160 5098
rect 15108 5034 15160 5040
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 15120 4758 15148 5034
rect 15304 4758 15332 5664
rect 15396 5302 15424 6054
rect 15384 5296 15436 5302
rect 15384 5238 15436 5244
rect 15396 4826 15424 5238
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 14956 4380 15252 4400
rect 15012 4378 15036 4380
rect 15092 4378 15116 4380
rect 15172 4378 15196 4380
rect 15034 4326 15036 4378
rect 15098 4326 15110 4378
rect 15172 4326 15174 4378
rect 15012 4324 15036 4326
rect 15092 4324 15116 4326
rect 15172 4324 15196 4326
rect 14956 4304 15252 4324
rect 15304 4162 15332 4422
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 15120 4134 15332 4162
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14738 3632 14794 3641
rect 14936 3602 14964 4082
rect 15120 3670 15148 4134
rect 15488 4060 15516 6394
rect 15580 5914 15608 8026
rect 15672 8022 15700 8486
rect 15660 8016 15712 8022
rect 15660 7958 15712 7964
rect 15672 7546 15700 7958
rect 15856 7698 15884 8570
rect 15764 7670 15884 7698
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15672 7002 15700 7482
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15764 6746 15792 7670
rect 15842 7576 15898 7585
rect 15842 7511 15844 7520
rect 15896 7511 15898 7520
rect 15844 7482 15896 7488
rect 15764 6718 15884 6746
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15672 5370 15700 5714
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15580 4486 15608 5102
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15304 4032 15516 4060
rect 15108 3664 15160 3670
rect 15014 3632 15070 3641
rect 14738 3567 14794 3576
rect 14924 3596 14976 3602
rect 14556 3460 14608 3466
rect 14556 3402 14608 3408
rect 14568 2650 14596 3402
rect 14646 3360 14702 3369
rect 14646 3295 14702 3304
rect 14660 2990 14688 3295
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14648 2848 14700 2854
rect 14646 2816 14648 2825
rect 14700 2816 14702 2825
rect 14646 2751 14702 2760
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14462 2544 14518 2553
rect 14462 2479 14518 2488
rect 14476 2310 14504 2479
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14752 1442 14780 3567
rect 15108 3606 15160 3612
rect 15014 3567 15070 3576
rect 14924 3538 14976 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14844 2582 14872 3470
rect 15028 3466 15056 3567
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14956 3292 15252 3312
rect 15012 3290 15036 3292
rect 15092 3290 15116 3292
rect 15172 3290 15196 3292
rect 15034 3238 15036 3290
rect 15098 3238 15110 3290
rect 15172 3238 15174 3290
rect 15012 3236 15036 3238
rect 15092 3236 15116 3238
rect 15172 3236 15196 3238
rect 14956 3216 15252 3236
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15120 2802 15148 2926
rect 15304 2836 15332 4032
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15396 2990 15424 3470
rect 15474 3224 15530 3233
rect 15474 3159 15476 3168
rect 15528 3159 15530 3168
rect 15476 3130 15528 3136
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15198 2816 15254 2825
rect 15120 2774 15198 2802
rect 15304 2808 15424 2836
rect 15198 2751 15254 2760
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 15212 2514 15240 2751
rect 15396 2666 15424 2808
rect 15396 2638 15516 2666
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14956 2204 15252 2224
rect 15012 2202 15036 2204
rect 15092 2202 15116 2204
rect 15172 2202 15196 2204
rect 15034 2150 15036 2202
rect 15098 2150 15110 2202
rect 15172 2150 15174 2202
rect 15012 2148 15036 2150
rect 15092 2148 15116 2150
rect 15172 2148 15196 2150
rect 14956 2128 15252 2148
rect 15382 2136 15438 2145
rect 15382 2071 15384 2080
rect 15436 2071 15438 2080
rect 15384 2042 15436 2048
rect 14752 1414 14964 1442
rect 14936 480 14964 1414
rect 15488 480 15516 2638
rect 15580 2514 15608 4422
rect 15672 3913 15700 5306
rect 15764 4049 15792 6598
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15658 3904 15714 3913
rect 15658 3839 15714 3848
rect 15856 3738 15884 6718
rect 15948 4214 15976 9438
rect 15936 4208 15988 4214
rect 15936 4150 15988 4156
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15660 2916 15712 2922
rect 15660 2858 15712 2864
rect 15672 2825 15700 2858
rect 15856 2854 15884 3674
rect 15844 2848 15896 2854
rect 15658 2816 15714 2825
rect 15844 2790 15896 2796
rect 15658 2751 15714 2760
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 16040 480 16068 10474
rect 16132 8786 16160 10911
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 10198 16252 10406
rect 16212 10192 16264 10198
rect 16212 10134 16264 10140
rect 16224 9586 16252 10134
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16316 9722 16344 10066
rect 16396 10056 16448 10062
rect 16394 10024 16396 10033
rect 16448 10024 16450 10033
rect 16394 9959 16450 9968
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16408 9586 16436 9959
rect 16212 9580 16264 9586
rect 16212 9522 16264 9528
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16316 8922 16344 9522
rect 16500 9450 16528 11206
rect 16776 10810 16804 11222
rect 16868 11218 16896 11494
rect 16856 11212 16908 11218
rect 16856 11154 16908 11160
rect 16764 10804 16816 10810
rect 16764 10746 16816 10752
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16488 9444 16540 9450
rect 16488 9386 16540 9392
rect 16316 8894 16436 8922
rect 16302 8800 16358 8809
rect 16132 8758 16252 8786
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 16132 8430 16160 8599
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16224 8090 16252 8758
rect 16302 8735 16358 8744
rect 16212 8084 16264 8090
rect 16212 8026 16264 8032
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16132 6662 16160 7890
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7206 16252 7686
rect 16316 7478 16344 8735
rect 16408 8634 16436 8894
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16592 8378 16620 10542
rect 16868 10198 16896 11154
rect 16960 10266 16988 13767
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 12850 17080 13126
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 17144 11762 17172 24375
rect 17236 24070 17264 24686
rect 17316 24676 17368 24682
rect 17316 24618 17368 24624
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17236 20233 17264 22646
rect 17328 21185 17356 24618
rect 17314 21176 17370 21185
rect 17314 21111 17370 21120
rect 17222 20224 17278 20233
rect 17222 20159 17278 20168
rect 17420 19922 17448 26114
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17682 24168 17738 24177
rect 17512 23526 17540 24142
rect 17682 24103 17684 24112
rect 17736 24103 17738 24112
rect 17684 24074 17736 24080
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17512 22982 17540 23462
rect 17788 23089 17816 27520
rect 18236 26716 18288 26722
rect 18236 26658 18288 26664
rect 17868 25424 17920 25430
rect 17868 25366 17920 25372
rect 17880 24818 17908 25366
rect 18248 25158 18276 26658
rect 18340 25498 18368 27520
rect 18328 25492 18380 25498
rect 18328 25434 18380 25440
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17774 23080 17830 23089
rect 17774 23015 17830 23024
rect 17500 22976 17552 22982
rect 17500 22918 17552 22924
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17788 22234 17816 22374
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17512 21690 17540 21966
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17512 20942 17540 21490
rect 17788 21486 17816 22170
rect 17776 21480 17828 21486
rect 17776 21422 17828 21428
rect 17880 21418 17908 24550
rect 18064 24138 18092 24686
rect 18248 24614 18276 25094
rect 18512 24744 18564 24750
rect 18512 24686 18564 24692
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 18064 24041 18092 24074
rect 18144 24064 18196 24070
rect 18050 24032 18106 24041
rect 18144 24006 18196 24012
rect 18050 23967 18106 23976
rect 18156 23322 18184 24006
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18144 22092 18196 22098
rect 18144 22034 18196 22040
rect 18050 21448 18106 21457
rect 17868 21412 17920 21418
rect 18050 21383 18106 21392
rect 17868 21354 17920 21360
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17592 21004 17644 21010
rect 17592 20946 17644 20952
rect 17500 20936 17552 20942
rect 17500 20878 17552 20884
rect 17512 20602 17540 20878
rect 17500 20596 17552 20602
rect 17500 20538 17552 20544
rect 17498 20224 17554 20233
rect 17498 20159 17554 20168
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17420 19242 17448 19858
rect 17408 19236 17460 19242
rect 17408 19178 17460 19184
rect 17316 19168 17368 19174
rect 17512 19145 17540 20159
rect 17604 19718 17632 20946
rect 17880 20618 17908 21014
rect 17880 20590 18000 20618
rect 17774 20360 17830 20369
rect 17774 20295 17776 20304
rect 17828 20295 17830 20304
rect 17776 20266 17828 20272
rect 17682 20088 17738 20097
rect 17682 20023 17738 20032
rect 17696 19922 17724 20023
rect 17684 19916 17736 19922
rect 17684 19858 17736 19864
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17316 19110 17368 19116
rect 17498 19136 17554 19145
rect 17328 18465 17356 19110
rect 17498 19071 17554 19080
rect 17512 18970 17540 19071
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17314 18456 17370 18465
rect 17420 18426 17448 18770
rect 17314 18391 17370 18400
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17222 17232 17278 17241
rect 17222 17167 17278 17176
rect 17236 12918 17264 17167
rect 17420 16946 17448 18362
rect 17604 17882 17632 19654
rect 17696 19174 17724 19858
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17592 17876 17644 17882
rect 17592 17818 17644 17824
rect 17498 17776 17554 17785
rect 17498 17711 17554 17720
rect 17512 17338 17540 17711
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17512 17134 17540 17274
rect 17604 17202 17632 17478
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17328 16918 17448 16946
rect 17328 15706 17356 16918
rect 17604 16810 17632 17138
rect 17696 16998 17724 19110
rect 17868 18760 17920 18766
rect 17774 18728 17830 18737
rect 17868 18702 17920 18708
rect 17774 18663 17830 18672
rect 17788 18193 17816 18663
rect 17880 18426 17908 18702
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17774 18184 17830 18193
rect 17774 18119 17830 18128
rect 17972 17882 18000 20590
rect 18064 20398 18092 21383
rect 18156 21146 18184 22034
rect 18144 21140 18196 21146
rect 18144 21082 18196 21088
rect 18144 21004 18196 21010
rect 18144 20946 18196 20952
rect 18052 20392 18104 20398
rect 18052 20334 18104 20340
rect 18064 19825 18092 20334
rect 18050 19816 18106 19825
rect 18050 19751 18106 19760
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17338 17908 17682
rect 18064 17678 18092 18022
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 18064 17270 18092 17614
rect 18052 17264 18104 17270
rect 18052 17206 18104 17212
rect 17684 16992 17736 16998
rect 18052 16992 18104 16998
rect 17684 16934 17736 16940
rect 17958 16960 18014 16969
rect 18052 16934 18104 16940
rect 17958 16895 18014 16904
rect 17408 16788 17460 16794
rect 17604 16782 17724 16810
rect 17408 16730 17460 16736
rect 17420 16182 17448 16730
rect 17696 16590 17724 16782
rect 17868 16788 17920 16794
rect 17868 16730 17920 16736
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17316 15700 17368 15706
rect 17316 15642 17368 15648
rect 17328 15201 17356 15642
rect 17314 15192 17370 15201
rect 17314 15127 17370 15136
rect 17314 13696 17370 13705
rect 17314 13631 17370 13640
rect 17328 13530 17356 13631
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17420 13025 17448 16118
rect 17696 16114 17724 16526
rect 17880 16250 17908 16730
rect 17972 16522 18000 16895
rect 18064 16697 18092 16934
rect 18156 16726 18184 20946
rect 18248 18290 18276 24550
rect 18328 22636 18380 22642
rect 18328 22578 18380 22584
rect 18340 22030 18368 22578
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18418 21992 18474 22001
rect 18340 21690 18368 21966
rect 18418 21927 18474 21936
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18432 21350 18460 21927
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18524 21010 18552 24686
rect 18616 24410 18644 25094
rect 18892 24585 18920 27520
rect 19432 25968 19484 25974
rect 19432 25910 19484 25916
rect 18972 25900 19024 25906
rect 18972 25842 19024 25848
rect 18878 24576 18934 24585
rect 18878 24511 18934 24520
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18512 21004 18564 21010
rect 18512 20946 18564 20952
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18236 18080 18288 18086
rect 18236 18022 18288 18028
rect 18144 16720 18196 16726
rect 18050 16688 18106 16697
rect 18144 16662 18196 16668
rect 18050 16623 18106 16632
rect 17960 16516 18012 16522
rect 17960 16458 18012 16464
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17684 16108 17736 16114
rect 17684 16050 17736 16056
rect 17592 15904 17644 15910
rect 17592 15846 17644 15852
rect 17604 14414 17632 15846
rect 17696 15706 17724 16050
rect 17972 15994 18000 16458
rect 18052 16448 18104 16454
rect 18050 16416 18052 16425
rect 18104 16416 18106 16425
rect 18050 16351 18106 16360
rect 18064 16114 18092 16351
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17972 15966 18092 15994
rect 18064 15745 18092 15966
rect 18142 15872 18198 15881
rect 18142 15807 18198 15816
rect 18050 15736 18106 15745
rect 17684 15700 17736 15706
rect 17960 15700 18012 15706
rect 17736 15660 17816 15688
rect 17684 15642 17736 15648
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17696 15162 17724 15506
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17788 14550 17816 15660
rect 18050 15671 18106 15680
rect 17960 15642 18012 15648
rect 17972 15178 18000 15642
rect 18156 15434 18184 15807
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17880 15162 18000 15178
rect 17868 15156 18000 15162
rect 17920 15150 18000 15156
rect 17868 15098 17920 15104
rect 18064 14890 18092 15302
rect 18248 14958 18276 18022
rect 18340 16794 18368 19994
rect 18420 19916 18472 19922
rect 18420 19858 18472 19864
rect 18432 19174 18460 19858
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18432 18873 18460 19110
rect 18524 18970 18552 20742
rect 18616 20058 18644 23530
rect 18708 22778 18736 23598
rect 18786 23488 18842 23497
rect 18786 23423 18842 23432
rect 18696 22772 18748 22778
rect 18696 22714 18748 22720
rect 18708 22574 18736 22714
rect 18696 22568 18748 22574
rect 18696 22510 18748 22516
rect 18800 22420 18828 23423
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18708 22392 18828 22420
rect 18604 20052 18656 20058
rect 18604 19994 18656 20000
rect 18604 19168 18656 19174
rect 18604 19110 18656 19116
rect 18512 18964 18564 18970
rect 18512 18906 18564 18912
rect 18418 18864 18474 18873
rect 18418 18799 18474 18808
rect 18512 18624 18564 18630
rect 18512 18566 18564 18572
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18432 16969 18460 18226
rect 18524 17921 18552 18566
rect 18616 18193 18644 19110
rect 18602 18184 18658 18193
rect 18602 18119 18658 18128
rect 18602 18048 18658 18057
rect 18602 17983 18658 17992
rect 18510 17912 18566 17921
rect 18510 17847 18566 17856
rect 18418 16960 18474 16969
rect 18418 16895 18474 16904
rect 18418 16824 18474 16833
rect 18328 16788 18380 16794
rect 18418 16759 18474 16768
rect 18328 16730 18380 16736
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 18340 15706 18368 16390
rect 18432 16046 18460 16759
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18432 15638 18460 15982
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18510 15464 18566 15473
rect 18510 15399 18566 15408
rect 18524 15042 18552 15399
rect 18616 15348 18644 17983
rect 18708 17218 18736 22392
rect 18892 21962 18920 22918
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18892 21554 18920 21898
rect 18880 21548 18932 21554
rect 18880 21490 18932 21496
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18800 20210 18828 21286
rect 18984 21146 19012 25842
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19352 25294 19380 25706
rect 19064 25288 19116 25294
rect 19064 25230 19116 25236
rect 19156 25288 19208 25294
rect 19156 25230 19208 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19076 24954 19104 25230
rect 19064 24948 19116 24954
rect 19064 24890 19116 24896
rect 19168 24818 19196 25230
rect 19444 25140 19472 25910
rect 19352 25112 19472 25140
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19168 24274 19196 24754
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 19352 24138 19380 25112
rect 19536 24834 19564 27520
rect 20088 26194 20116 27520
rect 20088 26166 20208 26194
rect 20074 26072 20130 26081
rect 20074 26007 20130 26016
rect 20088 25673 20116 26007
rect 20074 25664 20130 25673
rect 19622 25596 19918 25616
rect 20074 25599 20130 25608
rect 19678 25594 19702 25596
rect 19758 25594 19782 25596
rect 19838 25594 19862 25596
rect 19700 25542 19702 25594
rect 19764 25542 19776 25594
rect 19838 25542 19840 25594
rect 19678 25540 19702 25542
rect 19758 25540 19782 25542
rect 19838 25540 19862 25542
rect 19622 25520 19918 25540
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19720 24886 19748 25094
rect 19444 24806 19564 24834
rect 19708 24880 19760 24886
rect 20180 24834 20208 26166
rect 20352 26036 20404 26042
rect 20352 25978 20404 25984
rect 19708 24822 19760 24828
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19338 23216 19394 23225
rect 19338 23151 19340 23160
rect 19392 23151 19394 23160
rect 19340 23122 19392 23128
rect 19248 23044 19300 23050
rect 19248 22986 19300 22992
rect 19156 22568 19208 22574
rect 19156 22510 19208 22516
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 19076 21146 19104 22442
rect 19168 22234 19196 22510
rect 19260 22409 19288 22986
rect 19340 22432 19392 22438
rect 19246 22400 19302 22409
rect 19340 22374 19392 22380
rect 19246 22335 19302 22344
rect 19156 22228 19208 22234
rect 19156 22170 19208 22176
rect 19248 21548 19300 21554
rect 19352 21536 19380 22374
rect 19300 21508 19380 21536
rect 19248 21490 19300 21496
rect 18972 21140 19024 21146
rect 18972 21082 19024 21088
rect 19064 21140 19116 21146
rect 19116 21100 19196 21128
rect 19064 21082 19116 21088
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18892 20369 18920 20946
rect 18984 20602 19012 21082
rect 19064 20936 19116 20942
rect 19064 20878 19116 20884
rect 19168 20890 19196 21100
rect 19260 21078 19288 21490
rect 19338 21176 19394 21185
rect 19338 21111 19394 21120
rect 19248 21072 19300 21078
rect 19248 21014 19300 21020
rect 18972 20596 19024 20602
rect 18972 20538 19024 20544
rect 18878 20360 18934 20369
rect 18878 20295 18934 20304
rect 18800 20182 18920 20210
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18800 18426 18828 19722
rect 18892 19156 18920 20182
rect 19076 19938 19104 20878
rect 19168 20862 19288 20890
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 19168 20534 19196 20742
rect 19156 20528 19208 20534
rect 19156 20470 19208 20476
rect 19260 20398 19288 20862
rect 19352 20618 19380 21111
rect 19444 20806 19472 24806
rect 19720 24682 19748 24822
rect 20088 24806 20208 24834
rect 19982 24712 20038 24721
rect 19708 24676 19760 24682
rect 19982 24647 20038 24656
rect 19708 24618 19760 24624
rect 19524 24608 19576 24614
rect 19524 24550 19576 24556
rect 19536 24313 19564 24550
rect 19622 24508 19918 24528
rect 19678 24506 19702 24508
rect 19758 24506 19782 24508
rect 19838 24506 19862 24508
rect 19700 24454 19702 24506
rect 19764 24454 19776 24506
rect 19838 24454 19840 24506
rect 19678 24452 19702 24454
rect 19758 24452 19782 24454
rect 19838 24452 19862 24454
rect 19622 24432 19918 24452
rect 19996 24410 20024 24647
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19522 24304 19578 24313
rect 19522 24239 19578 24248
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19720 23594 19748 24210
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19708 23588 19760 23594
rect 19708 23530 19760 23536
rect 19524 23520 19576 23526
rect 19524 23462 19576 23468
rect 19536 23118 19564 23462
rect 19622 23420 19918 23440
rect 19678 23418 19702 23420
rect 19758 23418 19782 23420
rect 19838 23418 19862 23420
rect 19700 23366 19702 23418
rect 19764 23366 19776 23418
rect 19838 23366 19840 23418
rect 19678 23364 19702 23366
rect 19758 23364 19782 23366
rect 19838 23364 19862 23366
rect 19622 23344 19918 23364
rect 19524 23112 19576 23118
rect 19524 23054 19576 23060
rect 19536 22574 19564 23054
rect 19996 22574 20024 24074
rect 20088 22817 20116 24806
rect 20168 24676 20220 24682
rect 20168 24618 20220 24624
rect 20180 24313 20208 24618
rect 20260 24608 20312 24614
rect 20260 24550 20312 24556
rect 20272 24449 20300 24550
rect 20258 24440 20314 24449
rect 20258 24375 20314 24384
rect 20166 24304 20222 24313
rect 20166 24239 20222 24248
rect 20364 24206 20392 25978
rect 20640 24834 20668 27520
rect 20810 25800 20866 25809
rect 20810 25735 20866 25744
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20548 24806 20668 24834
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20352 24200 20404 24206
rect 20352 24142 20404 24148
rect 20180 23186 20208 24142
rect 20456 24138 20484 24754
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20350 24032 20406 24041
rect 20350 23967 20406 23976
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20168 23180 20220 23186
rect 20168 23122 20220 23128
rect 20166 22944 20222 22953
rect 20166 22879 20222 22888
rect 20074 22808 20130 22817
rect 20074 22743 20130 22752
rect 19524 22568 19576 22574
rect 19524 22510 19576 22516
rect 19984 22568 20036 22574
rect 19984 22510 20036 22516
rect 20074 22400 20130 22409
rect 19622 22332 19918 22352
rect 20074 22335 20130 22344
rect 19678 22330 19702 22332
rect 19758 22330 19782 22332
rect 19838 22330 19862 22332
rect 19700 22278 19702 22330
rect 19764 22278 19776 22330
rect 19838 22278 19840 22330
rect 19678 22276 19702 22278
rect 19758 22276 19782 22278
rect 19838 22276 19862 22278
rect 19622 22256 19918 22276
rect 20088 22166 20116 22335
rect 19616 22160 19668 22166
rect 19616 22102 19668 22108
rect 20076 22160 20128 22166
rect 20076 22102 20128 22108
rect 19524 22092 19576 22098
rect 19524 22034 19576 22040
rect 19536 21350 19564 22034
rect 19628 21486 19656 22102
rect 19616 21480 19668 21486
rect 20076 21480 20128 21486
rect 19616 21422 19668 21428
rect 19706 21448 19762 21457
rect 20076 21422 20128 21428
rect 19706 21383 19708 21392
rect 19760 21383 19762 21392
rect 19708 21354 19760 21360
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19984 21344 20036 21350
rect 19984 21286 20036 21292
rect 19622 21244 19918 21264
rect 19678 21242 19702 21244
rect 19758 21242 19782 21244
rect 19838 21242 19862 21244
rect 19700 21190 19702 21242
rect 19764 21190 19776 21242
rect 19838 21190 19840 21242
rect 19678 21188 19702 21190
rect 19758 21188 19782 21190
rect 19838 21188 19862 21190
rect 19622 21168 19918 21188
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19352 20590 19472 20618
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19340 20052 19392 20058
rect 19340 19994 19392 20000
rect 19076 19910 19196 19938
rect 19168 19854 19196 19910
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19248 19712 19300 19718
rect 19248 19654 19300 19660
rect 19260 19174 19288 19654
rect 19352 19310 19380 19994
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18972 19168 19024 19174
rect 18892 19128 18972 19156
rect 18972 19110 19024 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19340 19168 19392 19174
rect 19444 19145 19472 20590
rect 19536 20330 19564 21014
rect 19996 20777 20024 21286
rect 19982 20768 20038 20777
rect 19982 20703 20038 20712
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19536 20058 19564 20266
rect 19622 20156 19918 20176
rect 19678 20154 19702 20156
rect 19758 20154 19782 20156
rect 19838 20154 19862 20156
rect 19700 20102 19702 20154
rect 19764 20102 19776 20154
rect 19838 20102 19840 20154
rect 19678 20100 19702 20102
rect 19758 20100 19782 20102
rect 19838 20100 19862 20102
rect 19622 20080 19918 20100
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19982 19816 20038 19825
rect 19982 19751 20038 19760
rect 19996 19310 20024 19751
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19340 19110 19392 19116
rect 19430 19136 19486 19145
rect 18984 18698 19012 19110
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 18788 18420 18840 18426
rect 18788 18362 18840 18368
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18984 17513 19012 18090
rect 18970 17504 19026 17513
rect 18970 17439 19026 17448
rect 18708 17190 19104 17218
rect 18972 16720 19024 16726
rect 18972 16662 19024 16668
rect 18984 16425 19012 16662
rect 18970 16416 19026 16425
rect 18970 16351 19026 16360
rect 18984 16250 19012 16351
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18708 15502 18736 16050
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18616 15320 19012 15348
rect 18524 15014 18644 15042
rect 18236 14952 18288 14958
rect 18236 14894 18288 14900
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 17776 14544 17828 14550
rect 18064 14498 18092 14826
rect 17776 14486 17828 14492
rect 17592 14408 17644 14414
rect 17592 14350 17644 14356
rect 17788 14074 17816 14486
rect 17880 14470 18092 14498
rect 17880 14278 17908 14470
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17776 14068 17828 14074
rect 17776 14010 17828 14016
rect 17880 13870 17908 14214
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17866 13696 17922 13705
rect 17866 13631 17922 13640
rect 17880 13530 17908 13631
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17406 13016 17462 13025
rect 17406 12951 17462 12960
rect 17224 12912 17276 12918
rect 17224 12854 17276 12860
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17222 12336 17278 12345
rect 17222 12271 17224 12280
rect 17276 12271 17278 12280
rect 17224 12242 17276 12248
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 17052 10062 17080 10542
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16408 8350 16620 8378
rect 16672 8356 16724 8362
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16224 7041 16252 7142
rect 16210 7032 16266 7041
rect 16210 6967 16266 6976
rect 16316 6934 16344 7142
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 5710 16160 6598
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16304 4208 16356 4214
rect 16304 4150 16356 4156
rect 16316 3942 16344 4150
rect 16408 4078 16436 8350
rect 16672 8298 16724 8304
rect 16684 8090 16712 8298
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16776 7018 16804 8774
rect 16592 6990 16804 7018
rect 16486 6624 16542 6633
rect 16486 6559 16542 6568
rect 16500 6458 16528 6559
rect 16488 6452 16540 6458
rect 16488 6394 16540 6400
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 16500 4808 16528 6122
rect 16592 5914 16620 6990
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16592 5098 16620 5850
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16580 4820 16632 4826
rect 16500 4780 16580 4808
rect 16396 4072 16448 4078
rect 16396 4014 16448 4020
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16500 3738 16528 4780
rect 16580 4762 16632 4768
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16500 2582 16528 3130
rect 16488 2576 16540 2582
rect 16488 2518 16540 2524
rect 16210 912 16266 921
rect 16210 847 16266 856
rect 9678 96 9734 105
rect 9678 31 9734 40
rect 10046 0 10102 480
rect 10598 0 10654 480
rect 11150 0 11206 480
rect 11702 0 11758 480
rect 12254 0 12310 480
rect 12806 0 12862 480
rect 13358 0 13414 480
rect 13910 0 13966 480
rect 14370 0 14426 480
rect 14922 0 14978 480
rect 15474 0 15530 480
rect 16026 0 16082 480
rect 16224 377 16252 847
rect 16592 480 16620 3538
rect 16684 3466 16712 6598
rect 16776 5914 16804 6802
rect 17130 6760 17186 6769
rect 17130 6695 17186 6704
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16854 6352 16910 6361
rect 17052 6322 17080 6598
rect 17144 6497 17172 6695
rect 17130 6488 17186 6497
rect 17130 6423 17186 6432
rect 16854 6287 16910 6296
rect 17040 6316 17092 6322
rect 16868 6254 16896 6287
rect 17040 6258 17092 6264
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16764 5908 16816 5914
rect 16764 5850 16816 5856
rect 16960 5710 16988 6054
rect 17052 5846 17080 6258
rect 17144 6186 17172 6423
rect 17132 6180 17184 6186
rect 17132 6122 17184 6128
rect 17040 5840 17092 5846
rect 17040 5782 17092 5788
rect 16948 5704 17000 5710
rect 16948 5646 17000 5652
rect 16960 5166 16988 5646
rect 17052 5370 17080 5782
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16948 5160 17000 5166
rect 16948 5102 17000 5108
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16776 4690 16804 4966
rect 17236 4808 17264 12038
rect 17420 11558 17448 12174
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17314 11384 17370 11393
rect 17420 11354 17448 11494
rect 17314 11319 17370 11328
rect 17408 11348 17460 11354
rect 17328 9058 17356 11319
rect 17408 11290 17460 11296
rect 17512 11257 17540 12106
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17512 10266 17540 11183
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17408 9376 17460 9382
rect 17406 9344 17408 9353
rect 17460 9344 17462 9353
rect 17406 9279 17462 9288
rect 17604 9217 17632 12854
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17696 12345 17724 12378
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17868 12232 17920 12238
rect 17774 12200 17830 12209
rect 17868 12174 17920 12180
rect 17774 12135 17830 12144
rect 17684 11756 17736 11762
rect 17684 11698 17736 11704
rect 17590 9208 17646 9217
rect 17590 9143 17646 9152
rect 17328 9030 17632 9058
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17144 4780 17264 4808
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 16776 4146 16804 4626
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16776 3534 16804 4082
rect 16960 3942 16988 4558
rect 17052 4457 17080 4626
rect 17038 4448 17094 4457
rect 17038 4383 17094 4392
rect 17052 3942 17080 4383
rect 16948 3936 17000 3942
rect 16946 3904 16948 3913
rect 17040 3936 17092 3942
rect 17000 3904 17002 3913
rect 17040 3878 17092 3884
rect 16946 3839 17002 3848
rect 16764 3528 16816 3534
rect 16764 3470 16816 3476
rect 16672 3460 16724 3466
rect 16672 3402 16724 3408
rect 16776 3126 16804 3470
rect 16764 3120 16816 3126
rect 16764 3062 16816 3068
rect 16854 2680 16910 2689
rect 16854 2615 16856 2624
rect 16908 2615 16910 2624
rect 16856 2586 16908 2592
rect 16670 2544 16726 2553
rect 16670 2479 16726 2488
rect 16684 2281 16712 2479
rect 16670 2272 16726 2281
rect 16670 2207 16726 2216
rect 17052 785 17080 3878
rect 17144 3482 17172 4780
rect 17328 4622 17356 6122
rect 17500 5092 17552 5098
rect 17500 5034 17552 5040
rect 17512 4622 17540 5034
rect 17316 4616 17368 4622
rect 17500 4616 17552 4622
rect 17316 4558 17368 4564
rect 17420 4576 17500 4604
rect 17420 3738 17448 4576
rect 17500 4558 17552 4564
rect 17498 4040 17554 4049
rect 17498 3975 17554 3984
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17144 3454 17448 3482
rect 17144 3398 17172 3454
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 17132 2032 17184 2038
rect 17132 1974 17184 1980
rect 17038 776 17094 785
rect 17038 711 17094 720
rect 17144 480 17172 1974
rect 17420 1737 17448 3454
rect 17406 1728 17462 1737
rect 17406 1663 17462 1672
rect 17512 1442 17540 3975
rect 17604 3602 17632 9030
rect 17696 7954 17724 11698
rect 17788 11393 17816 12135
rect 17774 11384 17830 11393
rect 17774 11319 17830 11328
rect 17880 10713 17908 12174
rect 17866 10704 17922 10713
rect 17866 10639 17922 10648
rect 17972 10538 18000 13738
rect 18248 13530 18276 14894
rect 18512 14816 18564 14822
rect 18512 14758 18564 14764
rect 18524 14385 18552 14758
rect 18510 14376 18566 14385
rect 18510 14311 18566 14320
rect 18328 13728 18380 13734
rect 18328 13670 18380 13676
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18340 13433 18368 13670
rect 18510 13560 18566 13569
rect 18510 13495 18566 13504
rect 18326 13424 18382 13433
rect 18326 13359 18382 13368
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12782 18092 13262
rect 18052 12776 18104 12782
rect 18052 12718 18104 12724
rect 18064 12646 18092 12718
rect 18432 12646 18460 13330
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18420 12640 18472 12646
rect 18420 12582 18472 12588
rect 18064 12102 18092 12582
rect 18432 12442 18460 12582
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 18064 11694 18092 12038
rect 18052 11688 18104 11694
rect 18052 11630 18104 11636
rect 18524 11354 18552 13495
rect 18616 12986 18644 15014
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18786 14648 18842 14657
rect 18786 14583 18788 14592
rect 18840 14583 18842 14592
rect 18788 14554 18840 14560
rect 18892 14550 18920 14826
rect 18880 14544 18932 14550
rect 18880 14486 18932 14492
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 18420 11008 18472 11014
rect 18420 10950 18472 10956
rect 18326 10840 18382 10849
rect 18326 10775 18328 10784
rect 18380 10775 18382 10784
rect 18328 10746 18380 10752
rect 17960 10532 18012 10538
rect 17960 10474 18012 10480
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17788 9625 17816 10202
rect 17866 10160 17922 10169
rect 17866 10095 17868 10104
rect 17920 10095 17922 10104
rect 17868 10066 17920 10072
rect 17774 9616 17830 9625
rect 17774 9551 17830 9560
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17788 8090 17816 8910
rect 17868 8832 17920 8838
rect 17868 8774 17920 8780
rect 17880 8129 17908 8774
rect 17866 8120 17922 8129
rect 17776 8084 17828 8090
rect 17866 8055 17922 8064
rect 17776 8026 17828 8032
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17696 7546 17724 7890
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17972 6882 18000 9046
rect 18064 8945 18092 10406
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18050 8936 18106 8945
rect 18050 8871 18106 8880
rect 18156 8090 18184 8978
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18156 7546 18184 8026
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18248 7342 18276 10406
rect 18432 10305 18460 10950
rect 18510 10840 18566 10849
rect 18510 10775 18566 10784
rect 18524 10674 18552 10775
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18418 10296 18474 10305
rect 18418 10231 18420 10240
rect 18472 10231 18474 10240
rect 18420 10202 18472 10208
rect 18432 9586 18460 10202
rect 18524 9722 18552 10610
rect 18512 9716 18564 9722
rect 18512 9658 18564 9664
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18420 9376 18472 9382
rect 18418 9344 18420 9353
rect 18512 9376 18564 9382
rect 18472 9344 18474 9353
rect 18512 9318 18564 9324
rect 18418 9279 18474 9288
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8362 18368 8910
rect 18524 8401 18552 9318
rect 18510 8392 18566 8401
rect 18328 8356 18380 8362
rect 18510 8327 18566 8336
rect 18328 8298 18380 8304
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 17972 6854 18184 6882
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17880 3738 17908 3946
rect 17868 3732 17920 3738
rect 17972 3720 18000 6734
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4214 18092 4966
rect 18156 4826 18184 6854
rect 18144 4820 18196 4826
rect 18144 4762 18196 4768
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 17920 3692 18000 3720
rect 18050 3768 18106 3777
rect 18050 3703 18106 3712
rect 17868 3674 17920 3680
rect 18064 3602 18092 3703
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17776 3528 17828 3534
rect 18156 3482 18184 4082
rect 17776 3470 17828 3476
rect 17788 3194 17816 3470
rect 18064 3454 18184 3482
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17604 2650 17632 2994
rect 18064 2961 18092 3454
rect 18050 2952 18106 2961
rect 18050 2887 18106 2896
rect 18064 2650 18092 2887
rect 18248 2836 18276 7142
rect 18340 6322 18368 8298
rect 18616 8294 18644 12650
rect 18696 11144 18748 11150
rect 18696 11086 18748 11092
rect 18708 10674 18736 11086
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 10266 18736 10610
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18800 10146 18828 14350
rect 18984 12306 19012 15320
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18972 12164 19024 12170
rect 18972 12106 19024 12112
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18892 11937 18920 12038
rect 18878 11928 18934 11937
rect 18878 11863 18934 11872
rect 18880 11076 18932 11082
rect 18984 11064 19012 12106
rect 18932 11036 19012 11064
rect 18880 11018 18932 11024
rect 18708 10118 18828 10146
rect 18604 8288 18656 8294
rect 18604 8230 18656 8236
rect 18708 8022 18736 10118
rect 18788 9920 18840 9926
rect 18788 9862 18840 9868
rect 18696 8016 18748 8022
rect 18696 7958 18748 7964
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18616 7002 18644 7890
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18708 7410 18736 7754
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18604 6996 18656 7002
rect 18604 6938 18656 6944
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18512 6112 18564 6118
rect 18510 6080 18512 6089
rect 18564 6080 18566 6089
rect 18510 6015 18566 6024
rect 18326 5944 18382 5953
rect 18326 5879 18382 5888
rect 18340 5642 18368 5879
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18418 5536 18474 5545
rect 18418 5471 18474 5480
rect 18432 5030 18460 5471
rect 18602 5264 18658 5273
rect 18602 5199 18604 5208
rect 18656 5199 18658 5208
rect 18604 5170 18656 5176
rect 18420 5024 18472 5030
rect 18418 4992 18420 5001
rect 18512 5024 18564 5030
rect 18472 4992 18474 5001
rect 18512 4966 18564 4972
rect 18418 4927 18474 4936
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18340 3942 18368 4762
rect 18524 4593 18552 4966
rect 18602 4856 18658 4865
rect 18708 4826 18736 7142
rect 18602 4791 18658 4800
rect 18696 4820 18748 4826
rect 18510 4584 18566 4593
rect 18510 4519 18566 4528
rect 18524 4282 18552 4519
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 18616 4146 18644 4791
rect 18696 4762 18748 4768
rect 18708 4282 18736 4762
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18328 3392 18380 3398
rect 18418 3360 18474 3369
rect 18380 3340 18418 3346
rect 18328 3334 18418 3340
rect 18340 3318 18418 3334
rect 18418 3295 18474 3304
rect 18432 2990 18460 3295
rect 18800 3194 18828 9862
rect 18892 7274 18920 11018
rect 19076 10470 19104 17190
rect 19168 16674 19196 18566
rect 19260 16794 19288 19110
rect 19352 18766 19380 19110
rect 19430 19071 19486 19080
rect 19622 19068 19918 19088
rect 19678 19066 19702 19068
rect 19758 19066 19782 19068
rect 19838 19066 19862 19068
rect 19700 19014 19702 19066
rect 19764 19014 19776 19066
rect 19838 19014 19840 19066
rect 19678 19012 19702 19014
rect 19758 19012 19782 19014
rect 19838 19012 19862 19014
rect 19622 18992 19918 19012
rect 19996 18970 20024 19246
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18426 19380 18702
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19536 18465 19564 18566
rect 19522 18456 19578 18465
rect 19340 18420 19392 18426
rect 19522 18391 19578 18400
rect 19708 18420 19760 18426
rect 19340 18362 19392 18368
rect 19708 18362 19760 18368
rect 19338 18320 19394 18329
rect 19338 18255 19394 18264
rect 19343 18244 19380 18255
rect 19343 18204 19371 18244
rect 19720 18222 19748 18362
rect 19708 18216 19760 18222
rect 19343 18176 19564 18204
rect 19536 18086 19564 18176
rect 19614 18184 19670 18193
rect 19708 18158 19760 18164
rect 19614 18119 19616 18128
rect 19668 18119 19670 18128
rect 19616 18090 19668 18096
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19352 17134 19380 18022
rect 19622 17980 19918 18000
rect 19678 17978 19702 17980
rect 19758 17978 19782 17980
rect 19838 17978 19862 17980
rect 19700 17926 19702 17978
rect 19764 17926 19776 17978
rect 19838 17926 19840 17978
rect 19678 17924 19702 17926
rect 19758 17924 19782 17926
rect 19838 17924 19862 17926
rect 19622 17904 19918 17924
rect 19996 17785 20024 18906
rect 19982 17776 20038 17785
rect 19982 17711 20038 17720
rect 19430 17504 19486 17513
rect 19430 17439 19486 17448
rect 19340 17128 19392 17134
rect 19340 17070 19392 17076
rect 19248 16788 19300 16794
rect 19248 16730 19300 16736
rect 19168 16658 19360 16674
rect 19168 16652 19392 16658
rect 19168 16646 19340 16652
rect 19332 16612 19340 16646
rect 19340 16594 19392 16600
rect 19156 16584 19208 16590
rect 19156 16526 19208 16532
rect 19168 15910 19196 16526
rect 19444 16114 19472 17439
rect 19522 17368 19578 17377
rect 19522 17303 19578 17312
rect 19536 16250 19564 17303
rect 19984 17060 20036 17066
rect 19984 17002 20036 17008
rect 19622 16892 19918 16912
rect 19678 16890 19702 16892
rect 19758 16890 19782 16892
rect 19838 16890 19862 16892
rect 19700 16838 19702 16890
rect 19764 16838 19776 16890
rect 19838 16838 19840 16890
rect 19678 16836 19702 16838
rect 19758 16836 19782 16838
rect 19838 16836 19862 16838
rect 19622 16816 19918 16836
rect 19996 16726 20024 17002
rect 19984 16720 20036 16726
rect 19984 16662 20036 16668
rect 19996 16522 20024 16662
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 19890 16280 19946 16289
rect 19524 16244 19576 16250
rect 19890 16215 19946 16224
rect 19524 16186 19576 16192
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19156 15904 19208 15910
rect 19156 15846 19208 15852
rect 19154 15736 19210 15745
rect 19154 15671 19210 15680
rect 19168 13734 19196 15671
rect 19340 14952 19392 14958
rect 19246 14920 19302 14929
rect 19340 14894 19392 14900
rect 19246 14855 19302 14864
rect 19260 14414 19288 14855
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19260 14113 19288 14350
rect 19246 14104 19302 14113
rect 19246 14039 19248 14048
rect 19300 14039 19302 14048
rect 19248 14010 19300 14016
rect 19260 13979 19288 14010
rect 19352 13938 19380 14894
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19156 13728 19208 13734
rect 19444 13705 19472 16050
rect 19524 15904 19576 15910
rect 19904 15892 19932 16215
rect 19982 16144 20038 16153
rect 19982 16079 20038 16088
rect 19996 16046 20024 16079
rect 19984 16040 20036 16046
rect 19984 15982 20036 15988
rect 19904 15864 20024 15892
rect 19524 15846 19576 15852
rect 19536 15434 19564 15846
rect 19622 15804 19918 15824
rect 19678 15802 19702 15804
rect 19758 15802 19782 15804
rect 19838 15802 19862 15804
rect 19700 15750 19702 15802
rect 19764 15750 19776 15802
rect 19838 15750 19840 15802
rect 19678 15748 19702 15750
rect 19758 15748 19782 15750
rect 19838 15748 19862 15750
rect 19622 15728 19918 15748
rect 19996 15570 20024 15864
rect 19984 15564 20036 15570
rect 19984 15506 20036 15512
rect 19524 15428 19576 15434
rect 19524 15370 19576 15376
rect 19982 15056 20038 15065
rect 19982 14991 20038 15000
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19536 14464 19564 14894
rect 19622 14716 19918 14736
rect 19678 14714 19702 14716
rect 19758 14714 19782 14716
rect 19838 14714 19862 14716
rect 19700 14662 19702 14714
rect 19764 14662 19776 14714
rect 19838 14662 19840 14714
rect 19678 14660 19702 14662
rect 19758 14660 19782 14662
rect 19838 14660 19862 14662
rect 19622 14640 19918 14660
rect 19616 14476 19668 14482
rect 19536 14436 19616 14464
rect 19616 14418 19668 14424
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 13802 19564 14214
rect 19524 13796 19576 13802
rect 19524 13738 19576 13744
rect 19156 13670 19208 13676
rect 19430 13696 19486 13705
rect 19430 13631 19486 13640
rect 19536 13190 19564 13738
rect 19622 13628 19918 13648
rect 19678 13626 19702 13628
rect 19758 13626 19782 13628
rect 19838 13626 19862 13628
rect 19700 13574 19702 13626
rect 19764 13574 19776 13626
rect 19838 13574 19840 13626
rect 19678 13572 19702 13574
rect 19758 13572 19782 13574
rect 19838 13572 19862 13574
rect 19622 13552 19918 13572
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19996 13138 20024 14991
rect 20088 14278 20116 21422
rect 20180 15706 20208 22879
rect 20272 19258 20300 23802
rect 20364 22817 20392 23967
rect 20456 23730 20484 24074
rect 20444 23724 20496 23730
rect 20444 23666 20496 23672
rect 20456 23322 20484 23666
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20444 23180 20496 23186
rect 20444 23122 20496 23128
rect 20350 22808 20406 22817
rect 20350 22743 20406 22752
rect 20352 22092 20404 22098
rect 20352 22034 20404 22040
rect 20364 21146 20392 22034
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 20272 19230 20392 19258
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18834 20300 19110
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 17882 20300 18770
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 16794 20300 17614
rect 20260 16788 20312 16794
rect 20260 16730 20312 16736
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20364 15586 20392 19230
rect 20180 15558 20392 15586
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19720 13025 19748 13126
rect 19996 13110 20116 13138
rect 19522 13016 19578 13025
rect 19522 12951 19578 12960
rect 19706 13016 19762 13025
rect 19706 12951 19762 12960
rect 19984 12980 20036 12986
rect 19432 12776 19484 12782
rect 19432 12718 19484 12724
rect 19340 12708 19392 12714
rect 19340 12650 19392 12656
rect 19352 12220 19380 12650
rect 19444 12617 19472 12718
rect 19430 12608 19486 12617
rect 19430 12543 19486 12552
rect 19432 12232 19484 12238
rect 19352 12192 19432 12220
rect 19432 12174 19484 12180
rect 19444 11830 19472 12174
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19340 11552 19392 11558
rect 19340 11494 19392 11500
rect 19430 11520 19486 11529
rect 19246 11112 19302 11121
rect 19156 11076 19208 11082
rect 19246 11047 19302 11056
rect 19156 11018 19208 11024
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18970 10024 19026 10033
rect 18970 9959 19026 9968
rect 18984 9654 19012 9959
rect 19064 9920 19116 9926
rect 19064 9862 19116 9868
rect 18972 9648 19024 9654
rect 18972 9590 19024 9596
rect 19076 9489 19104 9862
rect 19062 9480 19118 9489
rect 19062 9415 19118 9424
rect 19064 9376 19116 9382
rect 19064 9318 19116 9324
rect 19076 8838 19104 9318
rect 19168 9081 19196 11018
rect 19154 9072 19210 9081
rect 19154 9007 19210 9016
rect 19260 8906 19288 11047
rect 19352 9353 19380 11494
rect 19430 11455 19486 11464
rect 19444 11354 19472 11455
rect 19432 11348 19484 11354
rect 19536 11336 19564 12951
rect 19984 12922 20036 12928
rect 19622 12540 19918 12560
rect 19678 12538 19702 12540
rect 19758 12538 19782 12540
rect 19838 12538 19862 12540
rect 19700 12486 19702 12538
rect 19764 12486 19776 12538
rect 19838 12486 19840 12538
rect 19678 12484 19702 12486
rect 19758 12484 19782 12486
rect 19838 12484 19862 12486
rect 19622 12464 19918 12484
rect 19708 12164 19760 12170
rect 19708 12106 19760 12112
rect 19720 11694 19748 12106
rect 19996 11830 20024 12922
rect 20088 12850 20116 13110
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20088 12102 20116 12242
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 20088 11898 20116 12038
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 19984 11824 20036 11830
rect 19984 11766 20036 11772
rect 19708 11688 19760 11694
rect 19708 11630 19760 11636
rect 19622 11452 19918 11472
rect 19678 11450 19702 11452
rect 19758 11450 19782 11452
rect 19838 11450 19862 11452
rect 19700 11398 19702 11450
rect 19764 11398 19776 11450
rect 19838 11398 19840 11450
rect 19678 11396 19702 11398
rect 19758 11396 19782 11398
rect 19838 11396 19862 11398
rect 19622 11376 19918 11396
rect 20076 11348 20128 11354
rect 19536 11308 19656 11336
rect 19432 11290 19484 11296
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19444 10742 19472 11154
rect 19522 10976 19578 10985
rect 19522 10911 19578 10920
rect 19432 10736 19484 10742
rect 19432 10678 19484 10684
rect 19536 10674 19564 10911
rect 19524 10668 19576 10674
rect 19524 10610 19576 10616
rect 19628 10554 19656 11308
rect 20076 11290 20128 11296
rect 20088 11121 20116 11290
rect 20074 11112 20130 11121
rect 19984 11076 20036 11082
rect 20074 11047 20130 11056
rect 19984 11018 20036 11024
rect 19536 10526 19656 10554
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19444 10033 19472 10202
rect 19430 10024 19486 10033
rect 19430 9959 19486 9968
rect 19536 9654 19564 10526
rect 19622 10364 19918 10384
rect 19678 10362 19702 10364
rect 19758 10362 19782 10364
rect 19838 10362 19862 10364
rect 19700 10310 19702 10362
rect 19764 10310 19776 10362
rect 19838 10310 19840 10362
rect 19678 10308 19702 10310
rect 19758 10308 19782 10310
rect 19838 10308 19862 10310
rect 19622 10288 19918 10308
rect 19996 10248 20024 11018
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 20088 10305 20116 10678
rect 19904 10220 20024 10248
rect 20074 10296 20130 10305
rect 20074 10231 20130 10240
rect 19616 10056 19668 10062
rect 19616 9998 19668 10004
rect 19628 9722 19656 9998
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 19432 9648 19484 9654
rect 19430 9616 19432 9625
rect 19524 9648 19576 9654
rect 19484 9616 19486 9625
rect 19524 9590 19576 9596
rect 19904 9586 19932 10220
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19430 9551 19486 9560
rect 19616 9580 19668 9586
rect 19444 9450 19472 9551
rect 19616 9522 19668 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19628 9364 19656 9522
rect 20088 9518 20116 9862
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19338 9344 19394 9353
rect 19338 9279 19394 9288
rect 19536 9336 19656 9364
rect 19984 9376 20036 9382
rect 19248 8900 19300 8906
rect 19248 8842 19300 8848
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 19076 8673 19104 8774
rect 19062 8664 19118 8673
rect 19062 8599 19118 8608
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19156 8288 19208 8294
rect 19156 8230 19208 8236
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18880 7268 18932 7274
rect 18880 7210 18932 7216
rect 18984 6934 19012 7958
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 18972 6928 19024 6934
rect 18972 6870 19024 6876
rect 18880 6316 18932 6322
rect 18880 6258 18932 6264
rect 18892 5846 18920 6258
rect 18880 5840 18932 5846
rect 18880 5782 18932 5788
rect 18984 5692 19012 6870
rect 19076 5846 19104 7278
rect 19168 7206 19196 8230
rect 19246 7848 19302 7857
rect 19246 7783 19302 7792
rect 19260 7274 19288 7783
rect 19248 7268 19300 7274
rect 19248 7210 19300 7216
rect 19156 7200 19208 7206
rect 19156 7142 19208 7148
rect 19352 6780 19380 8502
rect 19430 8120 19486 8129
rect 19430 8055 19432 8064
rect 19484 8055 19486 8064
rect 19536 8072 19564 9336
rect 19984 9318 20036 9324
rect 19622 9276 19918 9296
rect 19678 9274 19702 9276
rect 19758 9274 19782 9276
rect 19838 9274 19862 9276
rect 19700 9222 19702 9274
rect 19764 9222 19776 9274
rect 19838 9222 19840 9274
rect 19678 9220 19702 9222
rect 19758 9220 19782 9222
rect 19838 9220 19862 9222
rect 19622 9200 19918 9220
rect 19892 8832 19944 8838
rect 19890 8800 19892 8809
rect 19944 8800 19946 8809
rect 19890 8735 19946 8744
rect 19890 8664 19946 8673
rect 19890 8599 19946 8608
rect 19904 8276 19932 8599
rect 19996 8430 20024 9318
rect 20076 9036 20128 9042
rect 20076 8978 20128 8984
rect 20088 8673 20116 8978
rect 20074 8664 20130 8673
rect 20074 8599 20076 8608
rect 20128 8599 20130 8608
rect 20076 8570 20128 8576
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19904 8248 20116 8276
rect 19622 8188 19918 8208
rect 19678 8186 19702 8188
rect 19758 8186 19782 8188
rect 19838 8186 19862 8188
rect 19700 8134 19702 8186
rect 19764 8134 19776 8186
rect 19838 8134 19840 8186
rect 19678 8132 19702 8134
rect 19758 8132 19782 8134
rect 19838 8132 19862 8134
rect 19622 8112 19918 8132
rect 20088 8129 20116 8248
rect 20074 8120 20130 8129
rect 19536 8044 19656 8072
rect 20074 8055 20130 8064
rect 19432 8026 19484 8032
rect 19444 7002 19472 8026
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19536 7546 19564 7890
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19628 7188 19656 8044
rect 19890 7984 19946 7993
rect 19890 7919 19892 7928
rect 19944 7919 19946 7928
rect 19984 7948 20036 7954
rect 19892 7890 19944 7896
rect 19984 7890 20036 7896
rect 19904 7410 19932 7890
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19996 7274 20024 7890
rect 20074 7848 20130 7857
rect 20074 7783 20076 7792
rect 20128 7783 20130 7792
rect 20076 7754 20128 7760
rect 20088 7342 20116 7754
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 19536 7160 19656 7188
rect 19432 6996 19484 7002
rect 19432 6938 19484 6944
rect 19536 6882 19564 7160
rect 19622 7100 19918 7120
rect 19678 7098 19702 7100
rect 19758 7098 19782 7100
rect 19838 7098 19862 7100
rect 19700 7046 19702 7098
rect 19764 7046 19776 7098
rect 19838 7046 19840 7098
rect 19678 7044 19702 7046
rect 19758 7044 19782 7046
rect 19838 7044 19862 7046
rect 19622 7024 19918 7044
rect 19536 6854 19748 6882
rect 19616 6792 19668 6798
rect 19352 6752 19616 6780
rect 19616 6734 19668 6740
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19524 6656 19576 6662
rect 19524 6598 19576 6604
rect 19168 6254 19196 6598
rect 19248 6452 19300 6458
rect 19300 6412 19472 6440
rect 19248 6394 19300 6400
rect 19338 6352 19394 6361
rect 19444 6338 19472 6412
rect 19536 6361 19564 6598
rect 19522 6352 19578 6361
rect 19444 6310 19522 6338
rect 19338 6287 19394 6296
rect 19522 6287 19578 6296
rect 19352 6254 19380 6287
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19340 6248 19392 6254
rect 19628 6202 19656 6734
rect 19720 6390 19748 6854
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 19996 6322 20024 6598
rect 19984 6316 20036 6322
rect 19984 6258 20036 6264
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 19340 6190 19392 6196
rect 19444 6174 19656 6202
rect 19444 5914 19472 6174
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19536 5914 19564 6054
rect 19622 6012 19918 6032
rect 19678 6010 19702 6012
rect 19758 6010 19782 6012
rect 19838 6010 19862 6012
rect 19700 5958 19702 6010
rect 19764 5958 19776 6010
rect 19838 5958 19840 6010
rect 19678 5956 19702 5958
rect 19758 5956 19782 5958
rect 19838 5956 19862 5958
rect 19622 5936 19918 5956
rect 19432 5908 19484 5914
rect 19432 5850 19484 5856
rect 19524 5908 19576 5914
rect 19524 5850 19576 5856
rect 19064 5840 19116 5846
rect 19064 5782 19116 5788
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 18892 5664 19012 5692
rect 18892 4826 18920 5664
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18892 3670 18920 4762
rect 18880 3664 18932 3670
rect 18880 3606 18932 3612
rect 18984 3534 19012 5170
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 4865 19104 4966
rect 19062 4856 19118 4865
rect 19062 4791 19118 4800
rect 19248 4004 19300 4010
rect 19248 3946 19300 3952
rect 19260 3670 19288 3946
rect 19248 3664 19300 3670
rect 19246 3632 19248 3641
rect 19300 3632 19302 3641
rect 19064 3596 19116 3602
rect 19246 3567 19302 3576
rect 19064 3538 19116 3544
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 19076 3194 19104 3538
rect 18788 3188 18840 3194
rect 18788 3130 18840 3136
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 18510 3088 18566 3097
rect 18510 3023 18566 3032
rect 18524 2990 18552 3023
rect 18420 2984 18472 2990
rect 18420 2926 18472 2932
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18248 2808 18460 2836
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 1601 18368 2246
rect 18326 1592 18382 1601
rect 18326 1527 18382 1536
rect 18234 1456 18290 1465
rect 17512 1414 17724 1442
rect 17222 912 17278 921
rect 17222 847 17278 856
rect 16210 368 16266 377
rect 16210 303 16266 312
rect 16578 0 16634 480
rect 17130 0 17186 480
rect 17236 105 17264 847
rect 17696 480 17724 1414
rect 18234 1391 18290 1400
rect 18248 480 18276 1391
rect 17222 96 17278 105
rect 17222 31 17278 40
rect 17682 0 17738 480
rect 18234 0 18290 480
rect 18432 241 18460 2808
rect 18786 2816 18842 2825
rect 18786 2751 18842 2760
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18708 2145 18736 2450
rect 18800 2446 18828 2751
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 18510 2136 18566 2145
rect 18510 2071 18566 2080
rect 18694 2136 18750 2145
rect 18694 2071 18750 2080
rect 18524 1714 18552 2071
rect 18602 1728 18658 1737
rect 18524 1686 18602 1714
rect 18602 1663 18658 1672
rect 18786 1456 18842 1465
rect 18786 1391 18842 1400
rect 18800 480 18828 1391
rect 19352 480 19380 5510
rect 19444 5273 19472 5714
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19430 5264 19486 5273
rect 19904 5234 19932 5510
rect 19430 5199 19486 5208
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19522 5128 19578 5137
rect 19522 5063 19578 5072
rect 19536 5030 19564 5063
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4826 19564 4966
rect 19622 4924 19918 4944
rect 19678 4922 19702 4924
rect 19758 4922 19782 4924
rect 19838 4922 19862 4924
rect 19700 4870 19702 4922
rect 19764 4870 19776 4922
rect 19838 4870 19840 4922
rect 19678 4868 19702 4870
rect 19758 4868 19782 4870
rect 19838 4868 19862 4870
rect 19622 4848 19918 4868
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19444 4078 19472 4490
rect 19432 4072 19484 4078
rect 19432 4014 19484 4020
rect 19622 3836 19918 3856
rect 19678 3834 19702 3836
rect 19758 3834 19782 3836
rect 19838 3834 19862 3836
rect 19700 3782 19702 3834
rect 19764 3782 19776 3834
rect 19838 3782 19840 3834
rect 19678 3780 19702 3782
rect 19758 3780 19782 3782
rect 19838 3780 19862 3782
rect 19430 3768 19486 3777
rect 19622 3760 19918 3780
rect 19430 3703 19486 3712
rect 19444 3670 19472 3703
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19432 3392 19484 3398
rect 19432 3334 19484 3340
rect 19444 2825 19472 3334
rect 19430 2816 19486 2825
rect 19430 2751 19486 2760
rect 19622 2748 19918 2768
rect 19678 2746 19702 2748
rect 19758 2746 19782 2748
rect 19838 2746 19862 2748
rect 19700 2694 19702 2746
rect 19764 2694 19776 2746
rect 19838 2694 19840 2746
rect 19678 2692 19702 2694
rect 19758 2692 19782 2694
rect 19838 2692 19862 2694
rect 19622 2672 19918 2692
rect 19798 2408 19854 2417
rect 19798 2343 19800 2352
rect 19852 2343 19854 2352
rect 19800 2314 19852 2320
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 19904 480 19932 2246
rect 18418 232 18474 241
rect 18418 167 18474 176
rect 18786 0 18842 480
rect 19338 0 19394 480
rect 19890 0 19946 480
rect 19996 377 20024 6054
rect 20088 5302 20116 6258
rect 20180 6066 20208 15558
rect 20352 15360 20404 15366
rect 20350 15328 20352 15337
rect 20404 15328 20406 15337
rect 20350 15263 20406 15272
rect 20364 14890 20392 15263
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 20456 14414 20484 23122
rect 20548 22030 20576 24806
rect 20628 24608 20680 24614
rect 20628 24550 20680 24556
rect 20640 24342 20668 24550
rect 20628 24336 20680 24342
rect 20628 24278 20680 24284
rect 20640 23866 20668 24278
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20720 23588 20772 23594
rect 20720 23530 20772 23536
rect 20640 23066 20668 23530
rect 20732 23322 20760 23530
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20824 23202 20852 25735
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 20902 24168 20958 24177
rect 20902 24103 20904 24112
rect 20956 24103 20958 24112
rect 20904 24074 20956 24080
rect 21008 23526 21036 24822
rect 21100 24614 21128 25298
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 21088 24608 21140 24614
rect 21088 24550 21140 24556
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 20824 23174 21036 23202
rect 20904 23112 20956 23118
rect 20640 23038 20852 23066
rect 20904 23054 20956 23060
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 20626 22808 20682 22817
rect 20626 22743 20682 22752
rect 20640 22137 20668 22743
rect 20626 22128 20682 22137
rect 20626 22063 20682 22072
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 20548 21554 20576 21830
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20548 20466 20576 21490
rect 20640 21486 20668 22063
rect 20732 22030 20760 22918
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20628 21480 20680 21486
rect 20628 21422 20680 21428
rect 20640 21078 20668 21422
rect 20732 21146 20760 21966
rect 20720 21140 20772 21146
rect 20720 21082 20772 21088
rect 20628 21072 20680 21078
rect 20628 21014 20680 21020
rect 20824 20992 20852 23038
rect 20916 22710 20944 23054
rect 21008 22710 21036 23174
rect 20904 22704 20956 22710
rect 20902 22672 20904 22681
rect 20996 22704 21048 22710
rect 20956 22672 20958 22681
rect 20996 22646 21048 22652
rect 20902 22607 20958 22616
rect 20904 22568 20956 22574
rect 20904 22510 20956 22516
rect 20916 22012 20944 22510
rect 21100 22409 21128 24550
rect 21086 22400 21142 22409
rect 21086 22335 21142 22344
rect 21192 22148 21220 24686
rect 21284 23633 21312 27520
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21376 24410 21404 25774
rect 21836 25378 21864 27520
rect 22008 26444 22060 26450
rect 22008 26386 22060 26392
rect 21836 25350 21956 25378
rect 21822 24848 21878 24857
rect 21822 24783 21878 24792
rect 21836 24614 21864 24783
rect 21824 24608 21876 24614
rect 21824 24550 21876 24556
rect 21364 24404 21416 24410
rect 21364 24346 21416 24352
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21560 23866 21588 24210
rect 21928 23866 21956 25350
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21270 23624 21326 23633
rect 21270 23559 21326 23568
rect 21560 23338 21588 23802
rect 22020 23594 22048 26386
rect 22388 25498 22416 27520
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22836 25288 22888 25294
rect 22836 25230 22888 25236
rect 22466 25120 22522 25129
rect 22466 25055 22522 25064
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21560 23310 21772 23338
rect 21640 23180 21692 23186
rect 21640 23122 21692 23128
rect 21456 23112 21508 23118
rect 21456 23054 21508 23060
rect 21546 23080 21602 23089
rect 21468 22642 21496 23054
rect 21546 23015 21602 23024
rect 21456 22636 21508 22642
rect 21456 22578 21508 22584
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21183 22120 21220 22148
rect 21183 22012 21211 22120
rect 20916 21984 21036 22012
rect 21183 21984 21220 22012
rect 20732 20964 20852 20992
rect 20732 20890 20760 20964
rect 20640 20862 20760 20890
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20812 20868 20864 20874
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 20369 20576 20402
rect 20534 20360 20590 20369
rect 20534 20295 20590 20304
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20548 20058 20576 20198
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20548 19378 20576 19994
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20640 19258 20668 20862
rect 20812 20810 20864 20816
rect 20824 20534 20852 20810
rect 20812 20528 20864 20534
rect 20916 20505 20944 20878
rect 20812 20470 20864 20476
rect 20902 20496 20958 20505
rect 20824 19922 20852 20470
rect 20902 20431 20958 20440
rect 20902 20224 20958 20233
rect 20902 20159 20958 20168
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20548 19230 20668 19258
rect 20548 17921 20576 19230
rect 20628 19168 20680 19174
rect 20626 19136 20628 19145
rect 20680 19136 20682 19145
rect 20626 19071 20682 19080
rect 20732 18034 20760 19450
rect 20824 19446 20852 19858
rect 20812 19440 20864 19446
rect 20812 19382 20864 19388
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20824 18426 20852 18838
rect 20916 18737 20944 20159
rect 20902 18728 20958 18737
rect 20902 18663 20958 18672
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20640 18006 20760 18034
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20534 17912 20590 17921
rect 20534 17847 20590 17856
rect 20640 17814 20668 18006
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20628 17808 20680 17814
rect 20548 17768 20628 17796
rect 20548 16114 20576 17768
rect 20628 17750 20680 17756
rect 20732 17746 20760 17847
rect 20720 17740 20772 17746
rect 20720 17682 20772 17688
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20732 17490 20760 17546
rect 20640 17462 20760 17490
rect 20640 17338 20668 17462
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20640 16794 20668 17274
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20824 16726 20852 18022
rect 20916 17746 20944 18663
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 20904 17536 20956 17542
rect 20902 17504 20904 17513
rect 20956 17504 20958 17513
rect 20902 17439 20958 17448
rect 20904 16992 20956 16998
rect 20902 16960 20904 16969
rect 20956 16960 20958 16969
rect 20902 16895 20958 16904
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20812 16720 20864 16726
rect 20718 16688 20774 16697
rect 20812 16662 20864 16668
rect 20718 16623 20774 16632
rect 20732 16250 20760 16623
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15638 20576 16050
rect 20732 16046 20760 16186
rect 20720 16040 20772 16046
rect 20720 15982 20772 15988
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20536 15632 20588 15638
rect 20536 15574 20588 15580
rect 20640 15450 20668 15914
rect 20720 15632 20772 15638
rect 20718 15600 20720 15609
rect 20772 15600 20774 15609
rect 20718 15535 20774 15544
rect 20824 15502 20852 16526
rect 20916 16153 20944 16730
rect 20902 16144 20958 16153
rect 20902 16079 20958 16088
rect 20904 15904 20956 15910
rect 20902 15872 20904 15881
rect 20956 15872 20958 15881
rect 20902 15807 20958 15816
rect 21008 15688 21036 21984
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 21100 21049 21128 21830
rect 21086 21040 21142 21049
rect 21086 20975 21142 20984
rect 21100 20505 21128 20975
rect 21086 20496 21142 20505
rect 21086 20431 21142 20440
rect 21088 18760 21140 18766
rect 21088 18702 21140 18708
rect 21100 17882 21128 18702
rect 21088 17876 21140 17882
rect 21088 17818 21140 17824
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 15978 21128 17682
rect 21088 15972 21140 15978
rect 21088 15914 21140 15920
rect 21192 15858 21220 21984
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 21284 21554 21312 21898
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21270 21448 21326 21457
rect 21270 21383 21326 21392
rect 21284 18902 21312 21383
rect 21376 18970 21404 22374
rect 21468 22234 21496 22578
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21468 21690 21496 22170
rect 21456 21684 21508 21690
rect 21456 21626 21508 21632
rect 21468 20602 21496 21626
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21456 19916 21508 19922
rect 21456 19858 21508 19864
rect 21468 19514 21496 19858
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21364 18964 21416 18970
rect 21364 18906 21416 18912
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21362 18864 21418 18873
rect 21362 18799 21418 18808
rect 21376 18426 21404 18799
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21376 18222 21404 18362
rect 21364 18216 21416 18222
rect 21364 18158 21416 18164
rect 21560 18170 21588 23015
rect 21652 21894 21680 23122
rect 21744 22817 21772 23310
rect 21822 23080 21878 23089
rect 21822 23015 21824 23024
rect 21876 23015 21878 23024
rect 21824 22986 21876 22992
rect 21730 22808 21786 22817
rect 21730 22743 21786 22752
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21640 21344 21692 21350
rect 21640 21286 21692 21292
rect 21652 20777 21680 21286
rect 21744 21146 21772 22510
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21836 21418 21864 21966
rect 21928 21593 21956 23462
rect 22020 23322 22048 23530
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 22020 22574 22048 23258
rect 22100 22976 22152 22982
rect 22100 22918 22152 22924
rect 22008 22568 22060 22574
rect 22008 22510 22060 22516
rect 21914 21584 21970 21593
rect 21914 21519 21970 21528
rect 22112 21434 22140 22918
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21928 21406 22140 21434
rect 21732 21140 21784 21146
rect 21732 21082 21784 21088
rect 21638 20768 21694 20777
rect 21638 20703 21694 20712
rect 21744 20398 21772 21082
rect 21836 20806 21864 21354
rect 21928 21350 21956 21406
rect 21916 21344 21968 21350
rect 21916 21286 21968 21292
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21640 20392 21692 20398
rect 21638 20360 21640 20369
rect 21732 20392 21784 20398
rect 21692 20360 21694 20369
rect 21732 20334 21784 20340
rect 21638 20295 21694 20304
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21652 19689 21680 20198
rect 21638 19680 21694 19689
rect 21638 19615 21694 19624
rect 21836 18766 21864 20742
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21928 18698 21956 21286
rect 22204 21078 22232 22034
rect 22480 21962 22508 25055
rect 22652 24268 22704 24274
rect 22652 24210 22704 24216
rect 22664 23526 22692 24210
rect 22652 23520 22704 23526
rect 22652 23462 22704 23468
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22296 21554 22324 21830
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22192 21072 22244 21078
rect 22192 21014 22244 21020
rect 22204 20602 22232 21014
rect 22296 20618 22324 21490
rect 22468 21072 22520 21078
rect 22468 21014 22520 21020
rect 22192 20596 22244 20602
rect 22296 20590 22416 20618
rect 22192 20538 22244 20544
rect 22204 19786 22232 20538
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22296 20058 22324 20402
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22388 19786 22416 20590
rect 22480 20398 22508 21014
rect 22468 20392 22520 20398
rect 22466 20360 22468 20369
rect 22520 20360 22522 20369
rect 22466 20295 22522 20304
rect 22192 19780 22244 19786
rect 22192 19722 22244 19728
rect 22376 19780 22428 19786
rect 22376 19722 22428 19728
rect 22008 19712 22060 19718
rect 22060 19660 22140 19666
rect 22008 19654 22140 19660
rect 22020 19638 22140 19654
rect 22112 19174 22140 19638
rect 22282 19544 22338 19553
rect 22282 19479 22338 19488
rect 22100 19168 22152 19174
rect 22100 19110 22152 19116
rect 21916 18692 21968 18698
rect 21916 18634 21968 18640
rect 21732 18624 21784 18630
rect 21732 18566 21784 18572
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21272 18148 21324 18154
rect 21560 18142 21680 18170
rect 21272 18090 21324 18096
rect 21284 17814 21312 18090
rect 21652 18086 21680 18142
rect 21548 18080 21600 18086
rect 21546 18048 21548 18057
rect 21640 18080 21692 18086
rect 21600 18048 21602 18057
rect 21640 18022 21692 18028
rect 21546 17983 21602 17992
rect 21272 17808 21324 17814
rect 21272 17750 21324 17756
rect 21548 17536 21600 17542
rect 21600 17484 21680 17490
rect 21548 17478 21680 17484
rect 21560 17462 21680 17478
rect 21456 16992 21508 16998
rect 21376 16940 21456 16946
rect 21376 16934 21508 16940
rect 21546 16960 21602 16969
rect 21376 16918 21496 16934
rect 21376 16726 21404 16918
rect 21546 16895 21602 16904
rect 21454 16824 21510 16833
rect 21454 16759 21510 16768
rect 21364 16720 21416 16726
rect 21362 16688 21364 16697
rect 21416 16688 21418 16697
rect 21272 16652 21324 16658
rect 21362 16623 21418 16632
rect 21272 16594 21324 16600
rect 21284 16182 21312 16594
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 21192 15830 21404 15858
rect 21270 15736 21326 15745
rect 21008 15660 21220 15688
rect 21270 15671 21326 15680
rect 20902 15600 20958 15609
rect 20902 15535 20958 15544
rect 20996 15564 21048 15570
rect 20812 15496 20864 15502
rect 20640 15422 20760 15450
rect 20812 15438 20864 15444
rect 20628 15360 20680 15366
rect 20628 15302 20680 15308
rect 20732 15314 20760 15422
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20272 11098 20300 14350
rect 20444 14272 20496 14278
rect 20444 14214 20496 14220
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20350 13152 20406 13161
rect 20350 13087 20406 13096
rect 20364 12442 20392 13087
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20456 11558 20484 14214
rect 20548 14074 20576 14214
rect 20640 14074 20668 15302
rect 20732 15286 20852 15314
rect 20718 15192 20774 15201
rect 20718 15127 20774 15136
rect 20732 15026 20760 15127
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20718 14512 20774 14521
rect 20718 14447 20774 14456
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20628 14068 20680 14074
rect 20628 14010 20680 14016
rect 20732 13938 20760 14447
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20534 13832 20590 13841
rect 20534 13767 20590 13776
rect 20444 11552 20496 11558
rect 20444 11494 20496 11500
rect 20272 11070 20392 11098
rect 20260 11008 20312 11014
rect 20260 10950 20312 10956
rect 20272 10674 20300 10950
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20272 9586 20300 9998
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 8974 20300 9522
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20272 6497 20300 8570
rect 20364 8022 20392 11070
rect 20444 9988 20496 9994
rect 20444 9930 20496 9936
rect 20352 8016 20404 8022
rect 20350 7984 20352 7993
rect 20404 7984 20406 7993
rect 20456 7954 20484 9930
rect 20350 7919 20406 7928
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20444 7744 20496 7750
rect 20350 7712 20406 7721
rect 20444 7686 20496 7692
rect 20350 7647 20406 7656
rect 20364 7041 20392 7647
rect 20350 7032 20406 7041
rect 20350 6967 20406 6976
rect 20350 6760 20406 6769
rect 20350 6695 20352 6704
rect 20404 6695 20406 6704
rect 20352 6666 20404 6672
rect 20258 6488 20314 6497
rect 20258 6423 20314 6432
rect 20260 6384 20312 6390
rect 20260 6326 20312 6332
rect 20272 6186 20300 6326
rect 20260 6180 20312 6186
rect 20260 6122 20312 6128
rect 20180 6038 20392 6066
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 20088 4826 20116 5238
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20074 4176 20130 4185
rect 20074 4111 20076 4120
rect 20128 4111 20130 4120
rect 20076 4082 20128 4088
rect 20168 4004 20220 4010
rect 20168 3946 20220 3952
rect 20180 3738 20208 3946
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20180 2417 20208 3674
rect 20272 3398 20300 5510
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20364 2990 20392 6038
rect 20352 2984 20404 2990
rect 20352 2926 20404 2932
rect 20364 2582 20392 2926
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 20166 2408 20222 2417
rect 20166 2343 20222 2352
rect 20456 480 20484 7686
rect 20548 5166 20576 13767
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20640 12374 20668 13330
rect 20824 13326 20852 15286
rect 20916 13530 20944 15535
rect 20996 15506 21048 15512
rect 21008 14550 21036 15506
rect 21086 15464 21142 15473
rect 21086 15399 21142 15408
rect 21100 14618 21128 15399
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20996 14544 21048 14550
rect 20996 14486 21048 14492
rect 21088 14476 21140 14482
rect 21088 14418 21140 14424
rect 20994 14104 21050 14113
rect 21100 14074 21128 14418
rect 20994 14039 21050 14048
rect 21088 14068 21140 14074
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20720 13184 20772 13190
rect 20720 13126 20772 13132
rect 20732 12442 20760 13126
rect 20824 12986 20852 13262
rect 21008 13172 21036 14039
rect 21088 14010 21140 14016
rect 21100 13977 21128 14010
rect 21086 13968 21142 13977
rect 21086 13903 21142 13912
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 20916 13144 21036 13172
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 20812 12776 20864 12782
rect 20810 12744 20812 12753
rect 20864 12744 20866 12753
rect 20810 12679 20866 12688
rect 20812 12640 20864 12646
rect 20812 12582 20864 12588
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20628 12368 20680 12374
rect 20628 12310 20680 12316
rect 20718 12200 20774 12209
rect 20718 12135 20774 12144
rect 20626 11792 20682 11801
rect 20626 11727 20682 11736
rect 20640 11694 20668 11727
rect 20732 11694 20760 12135
rect 20824 12073 20852 12582
rect 20810 12064 20866 12073
rect 20810 11999 20866 12008
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20626 11520 20682 11529
rect 20626 11455 20682 11464
rect 20640 9722 20668 11455
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 9926 20760 11086
rect 20824 11014 20852 11562
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20916 10538 20944 13144
rect 20996 12844 21048 12850
rect 20996 12786 21048 12792
rect 21008 11286 21036 12786
rect 21100 11354 21128 13767
rect 21088 11348 21140 11354
rect 21088 11290 21140 11296
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21008 10810 21036 11222
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21192 10690 21220 15660
rect 21284 13530 21312 15671
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21284 13394 21312 13466
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21270 12200 21326 12209
rect 21270 12135 21326 12144
rect 21008 10662 21220 10690
rect 20904 10532 20956 10538
rect 20904 10474 20956 10480
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20720 9920 20772 9926
rect 20718 9888 20720 9897
rect 20772 9888 20774 9897
rect 20718 9823 20774 9832
rect 20916 9722 20944 10066
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20640 8537 20668 9522
rect 20718 9480 20774 9489
rect 20718 9415 20774 9424
rect 20732 9178 20760 9415
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20626 8528 20682 8537
rect 20732 8498 20760 9114
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20626 8463 20682 8472
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20824 8378 20852 9046
rect 20640 8350 20852 8378
rect 20640 7546 20668 8350
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 7886 20760 8230
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20626 6760 20682 6769
rect 20732 6746 20760 7686
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 20824 6866 20852 7414
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20732 6718 20852 6746
rect 20626 6695 20682 6704
rect 20640 6390 20668 6695
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20628 6384 20680 6390
rect 20628 6326 20680 6332
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 20548 4321 20576 4490
rect 20534 4312 20590 4321
rect 20534 4247 20590 4256
rect 20536 3664 20588 3670
rect 20536 3606 20588 3612
rect 20548 3058 20576 3606
rect 20640 3126 20668 6326
rect 20732 6254 20760 6598
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20720 5772 20772 5778
rect 20720 5714 20772 5720
rect 20732 5370 20760 5714
rect 20824 5642 20852 6718
rect 20812 5636 20864 5642
rect 20812 5578 20864 5584
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20732 4078 20760 5034
rect 20916 4706 20944 9658
rect 21008 7857 21036 10662
rect 21088 10532 21140 10538
rect 21088 10474 21140 10480
rect 21100 7886 21128 10474
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21192 9518 21220 10406
rect 21284 9654 21312 12135
rect 21376 11898 21404 15830
rect 21468 14464 21496 16759
rect 21560 15706 21588 16895
rect 21548 15700 21600 15706
rect 21548 15642 21600 15648
rect 21468 14436 21588 14464
rect 21454 13560 21510 13569
rect 21560 13530 21588 14436
rect 21454 13495 21510 13504
rect 21548 13524 21600 13530
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 21468 11744 21496 13495
rect 21548 13466 21600 13472
rect 21548 13388 21600 13394
rect 21548 13330 21600 13336
rect 21376 11716 21496 11744
rect 21376 10266 21404 11716
rect 21560 11694 21588 13330
rect 21652 12866 21680 17462
rect 21744 15570 21772 18566
rect 22204 18290 22232 18566
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21836 15881 21864 18090
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 22020 17542 22048 18022
rect 22204 17542 22232 18226
rect 22296 17762 22324 19479
rect 22388 19378 22416 19722
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22388 18970 22416 19314
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22388 17882 22416 18906
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22296 17734 22416 17762
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22192 17536 22244 17542
rect 22192 17478 22244 17484
rect 22100 17196 22152 17202
rect 22204 17184 22232 17478
rect 22204 17156 22324 17184
rect 22100 17138 22152 17144
rect 22112 16522 22140 17138
rect 22192 17060 22244 17066
rect 22192 17002 22244 17008
rect 22100 16516 22152 16522
rect 22100 16458 22152 16464
rect 22112 16114 22140 16458
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 21822 15872 21878 15881
rect 21822 15807 21878 15816
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21928 15434 21956 16050
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 22020 15094 22048 15506
rect 22008 15088 22060 15094
rect 22008 15030 22060 15036
rect 21916 14816 21968 14822
rect 21730 14784 21786 14793
rect 21916 14758 21968 14764
rect 21730 14719 21786 14728
rect 21744 12986 21772 14719
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21836 14074 21864 14554
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21928 13977 21956 14758
rect 22020 14482 22048 15030
rect 22112 14958 22140 15642
rect 22100 14952 22152 14958
rect 22100 14894 22152 14900
rect 22008 14476 22060 14482
rect 22060 14436 22140 14464
rect 22008 14418 22060 14424
rect 22008 14340 22060 14346
rect 22008 14282 22060 14288
rect 21914 13968 21970 13977
rect 21914 13903 21970 13912
rect 22020 13852 22048 14282
rect 22112 14074 22140 14436
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22100 13864 22152 13870
rect 22020 13824 22100 13852
rect 22100 13806 22152 13812
rect 21916 13728 21968 13734
rect 21916 13670 21968 13676
rect 22100 13728 22152 13734
rect 22100 13670 22152 13676
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21652 12838 21772 12866
rect 21744 12730 21772 12838
rect 21744 12702 21864 12730
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21652 11898 21680 12174
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21548 11688 21600 11694
rect 21454 11656 21510 11665
rect 21548 11630 21600 11636
rect 21454 11591 21456 11600
rect 21508 11591 21510 11600
rect 21456 11562 21508 11568
rect 21560 11354 21588 11630
rect 21744 11558 21772 12242
rect 21732 11552 21784 11558
rect 21732 11494 21784 11500
rect 21548 11348 21600 11354
rect 21548 11290 21600 11296
rect 21640 11008 21692 11014
rect 21640 10950 21692 10956
rect 21546 10704 21602 10713
rect 21652 10674 21680 10950
rect 21546 10639 21602 10648
rect 21640 10668 21692 10674
rect 21560 10606 21588 10639
rect 21640 10610 21692 10616
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 10266 21588 10542
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21652 10062 21680 10610
rect 21732 10532 21784 10538
rect 21732 10474 21784 10480
rect 21640 10056 21692 10062
rect 21362 10024 21418 10033
rect 21640 9998 21692 10004
rect 21744 9994 21772 10474
rect 21362 9959 21418 9968
rect 21732 9988 21784 9994
rect 21272 9648 21324 9654
rect 21272 9590 21324 9596
rect 21180 9512 21232 9518
rect 21178 9480 21180 9489
rect 21232 9480 21234 9489
rect 21178 9415 21234 9424
rect 21178 9344 21234 9353
rect 21178 9279 21234 9288
rect 21192 9178 21220 9279
rect 21376 9217 21404 9959
rect 21732 9930 21784 9936
rect 21640 9920 21692 9926
rect 21836 9874 21864 12702
rect 21928 11558 21956 13670
rect 22112 13190 22140 13670
rect 22204 13394 22232 17002
rect 22296 16726 22324 17156
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22296 16250 22324 16662
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22296 15094 22324 16186
rect 22284 15088 22336 15094
rect 22284 15030 22336 15036
rect 22284 14816 22336 14822
rect 22284 14758 22336 14764
rect 22296 14618 22324 14758
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22388 14498 22416 17734
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 15162 22508 17070
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22296 14470 22416 14498
rect 22468 14544 22520 14550
rect 22468 14486 22520 14492
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 22296 13274 22324 14470
rect 22376 13796 22428 13802
rect 22376 13738 22428 13744
rect 22388 13394 22416 13738
rect 22480 13734 22508 14486
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22376 13388 22428 13394
rect 22376 13330 22428 13336
rect 22388 13297 22416 13330
rect 22204 13246 22324 13274
rect 22374 13288 22430 13297
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22008 12640 22060 12646
rect 22008 12582 22060 12588
rect 22020 12442 22048 12582
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 22112 12374 22140 13126
rect 22100 12368 22152 12374
rect 22100 12310 22152 12316
rect 22006 12064 22062 12073
rect 22006 11999 22062 12008
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21928 11354 21956 11494
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 21916 10736 21968 10742
rect 21914 10704 21916 10713
rect 21968 10704 21970 10713
rect 21914 10639 21970 10648
rect 22020 10538 22048 11999
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 22112 10810 22140 11222
rect 22100 10804 22152 10810
rect 22100 10746 22152 10752
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 22020 10248 22048 10474
rect 21640 9862 21692 9868
rect 21652 9586 21680 9862
rect 21744 9846 21864 9874
rect 21928 10220 22048 10248
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21652 9353 21680 9522
rect 21638 9344 21694 9353
rect 21638 9279 21694 9288
rect 21362 9208 21418 9217
rect 21180 9172 21232 9178
rect 21362 9143 21364 9152
rect 21180 9114 21232 9120
rect 21416 9143 21418 9152
rect 21546 9208 21602 9217
rect 21546 9143 21602 9152
rect 21364 9114 21416 9120
rect 21560 9110 21588 9143
rect 21548 9104 21600 9110
rect 21548 9046 21600 9052
rect 21548 8900 21600 8906
rect 21548 8842 21600 8848
rect 21454 8800 21510 8809
rect 21454 8735 21510 8744
rect 21270 8528 21326 8537
rect 21270 8463 21326 8472
rect 21180 7948 21232 7954
rect 21180 7890 21232 7896
rect 21088 7880 21140 7886
rect 20994 7848 21050 7857
rect 21088 7822 21140 7828
rect 20994 7783 21050 7792
rect 20996 6996 21048 7002
rect 20996 6938 21048 6944
rect 21008 6458 21036 6938
rect 21086 6760 21142 6769
rect 21086 6695 21142 6704
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21100 5642 21128 6695
rect 21192 6662 21220 7890
rect 21284 7546 21312 8463
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 21272 7200 21324 7206
rect 21376 7188 21404 7822
rect 21324 7160 21404 7188
rect 21272 7142 21324 7148
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21178 6488 21234 6497
rect 21178 6423 21180 6432
rect 21232 6423 21234 6432
rect 21180 6394 21232 6400
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21088 5636 21140 5642
rect 21088 5578 21140 5584
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21008 5030 21036 5170
rect 21100 5166 21128 5578
rect 21192 5574 21220 6258
rect 21180 5568 21232 5574
rect 21180 5510 21232 5516
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 20996 5024 21048 5030
rect 21180 5024 21232 5030
rect 20996 4966 21048 4972
rect 21178 4992 21180 5001
rect 21232 4992 21234 5001
rect 21008 4729 21036 4966
rect 21178 4927 21234 4936
rect 21284 4842 21312 7142
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21376 6322 21404 6666
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21362 5944 21418 5953
rect 21362 5879 21364 5888
rect 21416 5879 21418 5888
rect 21364 5850 21416 5856
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 5409 21404 5646
rect 21362 5400 21418 5409
rect 21362 5335 21418 5344
rect 21100 4814 21312 4842
rect 20824 4678 20944 4706
rect 20994 4720 21050 4729
rect 20824 4457 20852 4678
rect 20994 4655 21050 4664
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20810 4448 20866 4457
rect 20810 4383 20866 4392
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 20812 4072 20864 4078
rect 20812 4014 20864 4020
rect 20824 3942 20852 4014
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20812 3936 20864 3942
rect 20916 3913 20944 4558
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21008 4282 21036 4422
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 20812 3878 20864 3884
rect 20902 3904 20958 3913
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20732 1873 20760 3878
rect 20824 2553 20852 3878
rect 20902 3839 20958 3848
rect 20916 3194 20944 3839
rect 20994 3768 21050 3777
rect 20994 3703 21050 3712
rect 21008 3534 21036 3703
rect 20996 3528 21048 3534
rect 20996 3470 21048 3476
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21100 3074 21128 4814
rect 21376 4758 21404 5335
rect 21364 4752 21416 4758
rect 21364 4694 21416 4700
rect 21270 4312 21326 4321
rect 21270 4247 21326 4256
rect 21180 3936 21232 3942
rect 21180 3878 21232 3884
rect 21192 3777 21220 3878
rect 21178 3768 21234 3777
rect 21178 3703 21234 3712
rect 21284 3602 21312 4247
rect 21376 4214 21404 4694
rect 21364 4208 21416 4214
rect 21364 4150 21416 4156
rect 21272 3596 21324 3602
rect 21272 3538 21324 3544
rect 21284 3194 21312 3538
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 20916 3046 21128 3074
rect 20810 2544 20866 2553
rect 20810 2479 20866 2488
rect 20916 2394 20944 3046
rect 21376 2922 21404 3470
rect 21364 2916 21416 2922
rect 21364 2858 21416 2864
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21086 2816 21142 2825
rect 20824 2366 20944 2394
rect 20718 1864 20774 1873
rect 20718 1799 20774 1808
rect 19982 368 20038 377
rect 19982 303 20038 312
rect 20442 0 20498 480
rect 20824 105 20852 2366
rect 20904 2304 20956 2310
rect 20902 2272 20904 2281
rect 20956 2272 20958 2281
rect 20902 2207 20958 2216
rect 21008 2145 21036 2790
rect 21086 2751 21142 2760
rect 20994 2136 21050 2145
rect 20994 2071 21050 2080
rect 21100 1170 21128 2751
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21192 2553 21220 2586
rect 21178 2544 21234 2553
rect 21178 2479 21234 2488
rect 21008 1142 21128 1170
rect 21468 1170 21496 8735
rect 21560 8634 21588 8842
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21744 8362 21772 9846
rect 21928 9518 21956 10220
rect 22204 10130 22232 13246
rect 22374 13223 22430 13232
rect 22282 12608 22338 12617
rect 22282 12543 22338 12552
rect 22296 10520 22324 12543
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22374 12064 22430 12073
rect 22374 11999 22430 12008
rect 22388 11354 22416 11999
rect 22480 11762 22508 12310
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22480 11218 22508 11698
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22296 10492 22416 10520
rect 22282 10432 22338 10441
rect 22282 10367 22338 10376
rect 22296 10266 22324 10367
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22008 10124 22060 10130
rect 22008 10066 22060 10072
rect 22192 10124 22244 10130
rect 22192 10066 22244 10072
rect 22020 10010 22048 10066
rect 22388 10010 22416 10492
rect 22466 10432 22522 10441
rect 22466 10367 22522 10376
rect 22020 9982 22416 10010
rect 22204 9586 22232 9982
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 21916 9512 21968 9518
rect 21916 9454 21968 9460
rect 21928 9178 21956 9454
rect 21916 9172 21968 9178
rect 21916 9114 21968 9120
rect 22008 9036 22060 9042
rect 22008 8978 22060 8984
rect 22020 8809 22048 8978
rect 22192 8832 22244 8838
rect 21822 8800 21878 8809
rect 21822 8735 21878 8744
rect 22006 8800 22062 8809
rect 22192 8774 22244 8780
rect 22006 8735 22062 8744
rect 21732 8356 21784 8362
rect 21732 8298 21784 8304
rect 21836 8294 21864 8735
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 21638 7848 21694 7857
rect 21560 7750 21588 7822
rect 21638 7783 21694 7792
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21546 6488 21602 6497
rect 21546 6423 21602 6432
rect 21560 6390 21588 6423
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21560 6254 21588 6326
rect 21652 6254 21680 7783
rect 21732 7744 21784 7750
rect 21732 7686 21784 7692
rect 21744 7206 21772 7686
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21548 6248 21600 6254
rect 21548 6190 21600 6196
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21548 5840 21600 5846
rect 21548 5782 21600 5788
rect 21560 5409 21588 5782
rect 21652 5642 21680 6054
rect 21744 5681 21772 7142
rect 21836 7002 21864 8230
rect 21916 7336 21968 7342
rect 21916 7278 21968 7284
rect 21824 6996 21876 7002
rect 21928 6984 21956 7278
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 21928 6956 22048 6984
rect 21824 6938 21876 6944
rect 21914 6896 21970 6905
rect 21824 6860 21876 6866
rect 21914 6831 21970 6840
rect 21824 6802 21876 6808
rect 21836 6338 21864 6802
rect 21928 6798 21956 6831
rect 21916 6792 21968 6798
rect 21916 6734 21968 6740
rect 22020 6662 22048 6956
rect 22112 6730 22140 7142
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 21836 6310 21956 6338
rect 21928 6254 21956 6310
rect 21824 6248 21876 6254
rect 21824 6190 21876 6196
rect 21916 6248 21968 6254
rect 22020 6225 22048 6598
rect 21916 6190 21968 6196
rect 22006 6216 22062 6225
rect 21730 5672 21786 5681
rect 21640 5636 21692 5642
rect 21730 5607 21786 5616
rect 21640 5578 21692 5584
rect 21546 5400 21602 5409
rect 21546 5335 21602 5344
rect 21638 5128 21694 5137
rect 21638 5063 21640 5072
rect 21692 5063 21694 5072
rect 21640 5034 21692 5040
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 21560 3233 21588 4558
rect 21732 4140 21784 4146
rect 21652 4100 21732 4128
rect 21652 3534 21680 4100
rect 21732 4082 21784 4088
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21546 3224 21602 3233
rect 21546 3159 21602 3168
rect 21652 3058 21680 3470
rect 21836 3194 21864 6190
rect 22006 6151 22062 6160
rect 22204 5778 22232 8774
rect 22296 6934 22324 9862
rect 22480 8022 22508 10367
rect 22572 8090 22600 22578
rect 22664 21865 22692 23462
rect 22848 23322 22876 25230
rect 23032 24721 23060 27520
rect 23480 26104 23532 26110
rect 23480 26046 23532 26052
rect 23018 24712 23074 24721
rect 23492 24698 23520 26046
rect 23584 24857 23612 27520
rect 23570 24848 23626 24857
rect 23570 24783 23626 24792
rect 23492 24670 23612 24698
rect 23018 24647 23074 24656
rect 23202 24304 23258 24313
rect 23202 24239 23258 24248
rect 22926 23760 22982 23769
rect 22926 23695 22982 23704
rect 22836 23316 22888 23322
rect 22756 23276 22836 23304
rect 22756 22642 22784 23276
rect 22836 23258 22888 23264
rect 22836 23180 22888 23186
rect 22836 23122 22888 23128
rect 22848 23089 22876 23122
rect 22834 23080 22890 23089
rect 22834 23015 22890 23024
rect 22848 22778 22876 23015
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22744 22636 22796 22642
rect 22744 22578 22796 22584
rect 22650 21856 22706 21865
rect 22650 21791 22706 21800
rect 22652 20528 22704 20534
rect 22652 20470 22704 20476
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22664 20262 22692 20470
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22664 19378 22692 20198
rect 22652 19372 22704 19378
rect 22652 19314 22704 19320
rect 22664 18834 22692 19314
rect 22848 19174 22876 20470
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22664 18068 22692 18770
rect 22744 18080 22796 18086
rect 22664 18040 22744 18068
rect 22744 18022 22796 18028
rect 22652 17740 22704 17746
rect 22652 17682 22704 17688
rect 22664 16794 22692 17682
rect 22756 17678 22784 18022
rect 22836 17808 22888 17814
rect 22836 17750 22888 17756
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22756 16998 22784 17614
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22756 16674 22784 16934
rect 22848 16794 22876 17750
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 22664 16646 22784 16674
rect 22664 16590 22692 16646
rect 22652 16584 22704 16590
rect 22652 16526 22704 16532
rect 22664 16250 22692 16526
rect 22742 16416 22798 16425
rect 22742 16351 22798 16360
rect 22652 16244 22704 16250
rect 22652 16186 22704 16192
rect 22664 15638 22692 16186
rect 22652 15632 22704 15638
rect 22652 15574 22704 15580
rect 22652 15088 22704 15094
rect 22652 15030 22704 15036
rect 22664 13326 22692 15030
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22652 13184 22704 13190
rect 22652 13126 22704 13132
rect 22664 12714 22692 13126
rect 22756 12782 22784 16351
rect 22836 15564 22888 15570
rect 22836 15506 22888 15512
rect 22848 15162 22876 15506
rect 22836 15156 22888 15162
rect 22836 15098 22888 15104
rect 22848 14618 22876 15098
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22848 13569 22876 13806
rect 22834 13560 22890 13569
rect 22834 13495 22890 13504
rect 22836 13388 22888 13394
rect 22836 13330 22888 13336
rect 22848 13161 22876 13330
rect 22834 13152 22890 13161
rect 22834 13087 22890 13096
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22652 12708 22704 12714
rect 22652 12650 22704 12656
rect 22664 12442 22692 12650
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22664 9722 22692 9998
rect 22652 9716 22704 9722
rect 22652 9658 22704 9664
rect 22650 9616 22706 9625
rect 22650 9551 22706 9560
rect 22664 9178 22692 9551
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22652 8560 22704 8566
rect 22652 8502 22704 8508
rect 22560 8084 22612 8090
rect 22560 8026 22612 8032
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22388 7002 22416 7890
rect 22572 7546 22600 8026
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22376 6996 22428 7002
rect 22376 6938 22428 6944
rect 22572 6934 22600 7482
rect 22284 6928 22336 6934
rect 22284 6870 22336 6876
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 22560 6928 22612 6934
rect 22560 6870 22612 6876
rect 22376 6384 22428 6390
rect 22282 6352 22338 6361
rect 22376 6326 22428 6332
rect 22282 6287 22338 6296
rect 22296 5914 22324 6287
rect 22388 6186 22416 6326
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22284 5908 22336 5914
rect 22284 5850 22336 5856
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22388 5098 22416 6122
rect 22480 5234 22508 6870
rect 22558 6624 22614 6633
rect 22558 6559 22614 6568
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 22376 5092 22428 5098
rect 22376 5034 22428 5040
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 21928 4049 21956 4558
rect 22020 4078 22048 4966
rect 22100 4480 22152 4486
rect 22100 4422 22152 4428
rect 22008 4072 22060 4078
rect 21914 4040 21970 4049
rect 22008 4014 22060 4020
rect 21914 3975 21970 3984
rect 21928 3738 21956 3975
rect 22112 3738 22140 4422
rect 22572 4321 22600 6559
rect 22558 4312 22614 4321
rect 22558 4247 22614 4256
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 22100 3732 22152 3738
rect 22100 3674 22152 3680
rect 22006 3224 22062 3233
rect 21824 3188 21876 3194
rect 22006 3159 22062 3168
rect 21824 3130 21876 3136
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 21652 2650 21680 2994
rect 21836 2854 21864 3130
rect 22020 3074 22048 3159
rect 22100 3120 22152 3126
rect 22020 3068 22100 3074
rect 22020 3062 22152 3068
rect 22020 3046 22140 3062
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 22098 2952 22154 2961
rect 22098 2887 22154 2896
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21824 2644 21876 2650
rect 21824 2586 21876 2592
rect 21640 2508 21692 2514
rect 21640 2450 21692 2456
rect 21652 2310 21680 2450
rect 21836 2446 21864 2586
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21468 1142 21588 1170
rect 21008 480 21036 1142
rect 21560 480 21588 1142
rect 22112 480 22140 2887
rect 22388 2514 22416 2994
rect 22376 2508 22428 2514
rect 22376 2450 22428 2456
rect 22374 2408 22430 2417
rect 22374 2343 22430 2352
rect 22388 1873 22416 2343
rect 22572 2281 22600 4014
rect 22558 2272 22614 2281
rect 22558 2207 22614 2216
rect 22374 1864 22430 1873
rect 22374 1799 22430 1808
rect 22572 1193 22600 2207
rect 22558 1184 22614 1193
rect 22558 1119 22614 1128
rect 22664 480 22692 8502
rect 22756 7954 22784 12038
rect 22940 11354 22968 23695
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 23032 22438 23060 23054
rect 23110 22808 23166 22817
rect 23110 22743 23166 22752
rect 23020 22432 23072 22438
rect 23020 22374 23072 22380
rect 23032 21418 23060 22374
rect 23020 21412 23072 21418
rect 23020 21354 23072 21360
rect 23020 19168 23072 19174
rect 23020 19110 23072 19116
rect 23032 18970 23060 19110
rect 23020 18964 23072 18970
rect 23020 18906 23072 18912
rect 23032 17746 23060 18906
rect 23020 17740 23072 17746
rect 23020 17682 23072 17688
rect 23020 17264 23072 17270
rect 23124 17252 23152 22743
rect 23216 22234 23244 24239
rect 23480 23248 23532 23254
rect 23478 23216 23480 23225
rect 23532 23216 23534 23225
rect 23478 23151 23534 23160
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23204 22228 23256 22234
rect 23204 22170 23256 22176
rect 23216 21690 23244 22170
rect 23296 22024 23348 22030
rect 23348 21984 23428 22012
rect 23296 21966 23348 21972
rect 23400 21729 23428 21984
rect 23386 21720 23442 21729
rect 23204 21684 23256 21690
rect 23386 21655 23442 21664
rect 23204 21626 23256 21632
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23216 18601 23244 21354
rect 23400 21350 23428 21655
rect 23388 21344 23440 21350
rect 23388 21286 23440 21292
rect 23400 20482 23428 21286
rect 23492 20942 23520 22918
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23584 20890 23612 24670
rect 23860 22794 23888 27639
rect 24122 27520 24178 28000
rect 24766 27520 24822 28000
rect 25318 27520 25374 28000
rect 25870 27520 25926 28000
rect 26514 27520 26570 28000
rect 27066 27520 27122 28000
rect 27618 27520 27674 28000
rect 24030 25936 24086 25945
rect 24030 25871 24086 25880
rect 24044 25537 24072 25871
rect 24030 25528 24086 25537
rect 24030 25463 24086 25472
rect 23940 24744 23992 24750
rect 23940 24686 23992 24692
rect 23952 22953 23980 24686
rect 24136 24410 24164 27520
rect 24780 27282 24808 27520
rect 24688 27254 24808 27282
rect 24214 25936 24270 25945
rect 24214 25871 24270 25880
rect 24228 24886 24256 25871
rect 24688 25702 24716 27254
rect 24766 27160 24822 27169
rect 24766 27095 24822 27104
rect 24780 26722 24808 27095
rect 24768 26716 24820 26722
rect 24768 26658 24820 26664
rect 24766 26616 24822 26625
rect 24766 26551 24822 26560
rect 24780 26450 24808 26551
rect 24768 26444 24820 26450
rect 24768 26386 24820 26392
rect 24676 25696 24728 25702
rect 24676 25638 24728 25644
rect 24872 25430 24900 25461
rect 24860 25424 24912 25430
rect 24858 25392 24860 25401
rect 24912 25392 24914 25401
rect 24858 25327 24914 25336
rect 24289 25052 24585 25072
rect 24345 25050 24369 25052
rect 24425 25050 24449 25052
rect 24505 25050 24529 25052
rect 24367 24998 24369 25050
rect 24431 24998 24443 25050
rect 24505 24998 24507 25050
rect 24345 24996 24369 24998
rect 24425 24996 24449 24998
rect 24505 24996 24529 24998
rect 24289 24976 24585 24996
rect 24768 24948 24820 24954
rect 24768 24890 24820 24896
rect 24216 24880 24268 24886
rect 24780 24857 24808 24890
rect 24216 24822 24268 24828
rect 24766 24848 24822 24857
rect 24766 24783 24822 24792
rect 24214 24712 24270 24721
rect 24214 24647 24270 24656
rect 24228 24614 24256 24647
rect 24216 24608 24268 24614
rect 24216 24550 24268 24556
rect 24674 24440 24730 24449
rect 24124 24404 24176 24410
rect 24674 24375 24676 24384
rect 24124 24346 24176 24352
rect 24728 24375 24730 24384
rect 24676 24346 24728 24352
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24122 24168 24178 24177
rect 24122 24103 24178 24112
rect 23938 22944 23994 22953
rect 23938 22879 23994 22888
rect 23860 22766 23980 22794
rect 24136 22778 24164 24103
rect 24289 23964 24585 23984
rect 24345 23962 24369 23964
rect 24425 23962 24449 23964
rect 24505 23962 24529 23964
rect 24367 23910 24369 23962
rect 24431 23910 24443 23962
rect 24505 23910 24507 23962
rect 24345 23908 24369 23910
rect 24425 23908 24449 23910
rect 24505 23908 24529 23910
rect 24289 23888 24585 23908
rect 24688 23730 24716 24210
rect 24766 23896 24822 23905
rect 24766 23831 24768 23840
rect 24820 23831 24822 23840
rect 24768 23802 24820 23808
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 24676 23724 24728 23730
rect 24676 23666 24728 23672
rect 24320 23497 24348 23666
rect 24766 23624 24822 23633
rect 24766 23559 24822 23568
rect 24492 23520 24544 23526
rect 24306 23488 24362 23497
rect 24306 23423 24362 23432
rect 24490 23488 24492 23497
rect 24544 23488 24546 23497
rect 24490 23423 24546 23432
rect 24780 23322 24808 23559
rect 24768 23316 24820 23322
rect 24768 23258 24820 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24289 22876 24585 22896
rect 24345 22874 24369 22876
rect 24425 22874 24449 22876
rect 24505 22874 24529 22876
rect 24367 22822 24369 22874
rect 24431 22822 24443 22874
rect 24505 22822 24507 22874
rect 24345 22820 24369 22822
rect 24425 22820 24449 22822
rect 24505 22820 24529 22822
rect 24289 22800 24585 22820
rect 23662 22672 23718 22681
rect 23662 22607 23718 22616
rect 23848 22636 23900 22642
rect 23676 22574 23704 22607
rect 23848 22578 23900 22584
rect 23664 22568 23716 22574
rect 23664 22510 23716 22516
rect 23756 22500 23808 22506
rect 23756 22442 23808 22448
rect 23664 21344 23716 21350
rect 23664 21286 23716 21292
rect 23676 21146 23704 21286
rect 23664 21140 23716 21146
rect 23664 21082 23716 21088
rect 23584 20862 23704 20890
rect 23572 20800 23624 20806
rect 23572 20742 23624 20748
rect 23478 20632 23534 20641
rect 23478 20567 23480 20576
rect 23532 20567 23534 20576
rect 23480 20538 23532 20544
rect 23400 20454 23520 20482
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23296 19712 23348 19718
rect 23296 19654 23348 19660
rect 23308 19310 23336 19654
rect 23400 19378 23428 19790
rect 23388 19372 23440 19378
rect 23388 19314 23440 19320
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 23202 18592 23258 18601
rect 23202 18527 23258 18536
rect 23216 17814 23244 18527
rect 23308 18426 23336 19246
rect 23296 18420 23348 18426
rect 23296 18362 23348 18368
rect 23492 18306 23520 20454
rect 23584 19990 23612 20742
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 23676 19394 23704 20862
rect 23584 19366 23704 19394
rect 23584 18358 23612 19366
rect 23662 19272 23718 19281
rect 23662 19207 23718 19216
rect 23676 19174 23704 19207
rect 23664 19168 23716 19174
rect 23664 19110 23716 19116
rect 23308 18278 23520 18306
rect 23572 18352 23624 18358
rect 23572 18294 23624 18300
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23124 17224 23244 17252
rect 23020 17206 23072 17212
rect 23032 13802 23060 17206
rect 23112 14612 23164 14618
rect 23112 14554 23164 14560
rect 23020 13796 23072 13802
rect 23020 13738 23072 13744
rect 23018 13696 23074 13705
rect 23018 13631 23074 13640
rect 23032 13462 23060 13631
rect 23020 13456 23072 13462
rect 23020 13398 23072 13404
rect 23124 13326 23152 14554
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23032 12442 23060 13194
rect 23124 12986 23152 13262
rect 23112 12980 23164 12986
rect 23112 12922 23164 12928
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23020 12436 23072 12442
rect 23020 12378 23072 12384
rect 23124 12306 23152 12718
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 23020 12164 23072 12170
rect 23020 12106 23072 12112
rect 23032 11762 23060 12106
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23032 11354 23060 11698
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22836 11212 22888 11218
rect 22836 11154 22888 11160
rect 22848 10470 22876 11154
rect 22940 10810 22968 11290
rect 23124 11150 23152 11698
rect 23112 11144 23164 11150
rect 23018 11112 23074 11121
rect 23112 11086 23164 11092
rect 23018 11047 23074 11056
rect 22928 10804 22980 10810
rect 22928 10746 22980 10752
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 9926 22876 10406
rect 23032 10266 23060 11047
rect 23124 10810 23152 11086
rect 23112 10804 23164 10810
rect 23112 10746 23164 10752
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22940 9722 22968 10066
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22928 8968 22980 8974
rect 22926 8936 22928 8945
rect 22980 8936 22982 8945
rect 22926 8871 22982 8880
rect 23032 8430 23060 8978
rect 23020 8424 23072 8430
rect 23018 8392 23020 8401
rect 23072 8392 23074 8401
rect 23018 8327 23074 8336
rect 23124 8129 23152 10610
rect 23216 8514 23244 17224
rect 23308 16130 23336 18278
rect 23584 18222 23612 18294
rect 23572 18216 23624 18222
rect 23572 18158 23624 18164
rect 23584 18034 23612 18158
rect 23584 18006 23704 18034
rect 23570 17912 23626 17921
rect 23570 17847 23626 17856
rect 23388 17808 23440 17814
rect 23388 17750 23440 17756
rect 23400 17134 23428 17750
rect 23584 17338 23612 17847
rect 23572 17332 23624 17338
rect 23572 17274 23624 17280
rect 23388 17128 23440 17134
rect 23676 17082 23704 18006
rect 23768 17762 23796 22442
rect 23860 18290 23888 22578
rect 23952 22137 23980 22766
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 24688 22642 24716 23122
rect 24676 22636 24728 22642
rect 24676 22578 24728 22584
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24030 22264 24086 22273
rect 24030 22199 24086 22208
rect 23938 22128 23994 22137
rect 23938 22063 23940 22072
rect 23992 22063 23994 22072
rect 23940 22034 23992 22040
rect 23952 21486 23980 22034
rect 23940 21480 23992 21486
rect 23940 21422 23992 21428
rect 23938 20768 23994 20777
rect 23938 20703 23994 20712
rect 23952 19310 23980 20703
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 23952 18834 23980 19246
rect 23940 18828 23992 18834
rect 23940 18770 23992 18776
rect 23848 18284 23900 18290
rect 23848 18226 23900 18232
rect 23938 18048 23994 18057
rect 23938 17983 23994 17992
rect 23768 17734 23888 17762
rect 23756 17604 23808 17610
rect 23756 17546 23808 17552
rect 23768 17377 23796 17546
rect 23754 17368 23810 17377
rect 23754 17303 23810 17312
rect 23388 17070 23440 17076
rect 23584 17054 23704 17082
rect 23386 16552 23442 16561
rect 23386 16487 23442 16496
rect 23400 16250 23428 16487
rect 23584 16402 23612 17054
rect 23664 16992 23716 16998
rect 23664 16934 23716 16940
rect 23676 16833 23704 16934
rect 23662 16824 23718 16833
rect 23662 16759 23718 16768
rect 23756 16448 23808 16454
rect 23584 16374 23704 16402
rect 23756 16390 23808 16396
rect 23570 16280 23626 16289
rect 23388 16244 23440 16250
rect 23570 16215 23626 16224
rect 23388 16186 23440 16192
rect 23308 16102 23520 16130
rect 23492 16017 23520 16102
rect 23478 16008 23534 16017
rect 23296 15972 23348 15978
rect 23478 15943 23534 15952
rect 23296 15914 23348 15920
rect 23308 14074 23336 15914
rect 23388 15360 23440 15366
rect 23386 15328 23388 15337
rect 23440 15328 23442 15337
rect 23442 15286 23520 15314
rect 23386 15263 23442 15272
rect 23492 15162 23520 15286
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23480 14340 23532 14346
rect 23480 14282 23532 14288
rect 23492 14226 23520 14282
rect 23400 14198 23520 14226
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23294 13968 23350 13977
rect 23294 13903 23350 13912
rect 23308 12170 23336 13903
rect 23400 13530 23428 14198
rect 23480 14000 23532 14006
rect 23584 13977 23612 16215
rect 23676 14929 23704 16374
rect 23662 14920 23718 14929
rect 23662 14855 23718 14864
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23480 13942 23532 13948
rect 23570 13968 23626 13977
rect 23388 13524 23440 13530
rect 23388 13466 23440 13472
rect 23492 13394 23520 13942
rect 23570 13903 23626 13912
rect 23572 13728 23624 13734
rect 23572 13670 23624 13676
rect 23584 13462 23612 13670
rect 23572 13456 23624 13462
rect 23570 13424 23572 13433
rect 23624 13424 23626 13433
rect 23480 13388 23532 13394
rect 23570 13359 23626 13368
rect 23480 13330 23532 13336
rect 23570 13288 23626 13297
rect 23570 13223 23626 13232
rect 23478 13016 23534 13025
rect 23478 12951 23480 12960
rect 23532 12951 23534 12960
rect 23480 12922 23532 12928
rect 23480 12776 23532 12782
rect 23400 12724 23480 12730
rect 23400 12718 23532 12724
rect 23400 12702 23520 12718
rect 23400 12442 23428 12702
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23492 11898 23520 12242
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23296 11348 23348 11354
rect 23296 11290 23348 11296
rect 23308 10674 23336 11290
rect 23492 10962 23520 11494
rect 23400 10934 23520 10962
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 23400 10146 23428 10934
rect 23478 10840 23534 10849
rect 23478 10775 23480 10784
rect 23532 10775 23534 10784
rect 23480 10746 23532 10752
rect 23478 10296 23534 10305
rect 23584 10266 23612 13223
rect 23478 10231 23480 10240
rect 23532 10231 23534 10240
rect 23572 10260 23624 10266
rect 23480 10202 23532 10208
rect 23572 10202 23624 10208
rect 23400 10118 23612 10146
rect 23676 10130 23704 14758
rect 23768 13530 23796 16390
rect 23860 16250 23888 17734
rect 23952 16454 23980 17983
rect 23940 16448 23992 16454
rect 23940 16390 23992 16396
rect 23848 16244 23900 16250
rect 23848 16186 23900 16192
rect 24044 16130 24072 22199
rect 24676 22160 24728 22166
rect 24676 22102 24728 22108
rect 24289 21788 24585 21808
rect 24345 21786 24369 21788
rect 24425 21786 24449 21788
rect 24505 21786 24529 21788
rect 24367 21734 24369 21786
rect 24431 21734 24443 21786
rect 24505 21734 24507 21786
rect 24345 21732 24369 21734
rect 24425 21732 24449 21734
rect 24505 21732 24529 21734
rect 24289 21712 24585 21732
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24136 21078 24164 21490
rect 24688 21400 24716 22102
rect 24228 21372 24716 21400
rect 24124 21072 24176 21078
rect 24124 21014 24176 21020
rect 24124 20800 24176 20806
rect 24124 20742 24176 20748
rect 24136 16250 24164 20742
rect 24228 20330 24256 21372
rect 24674 21312 24730 21321
rect 24674 21247 24730 21256
rect 24289 20700 24585 20720
rect 24345 20698 24369 20700
rect 24425 20698 24449 20700
rect 24505 20698 24529 20700
rect 24367 20646 24369 20698
rect 24431 20646 24443 20698
rect 24505 20646 24507 20698
rect 24345 20644 24369 20646
rect 24425 20644 24449 20646
rect 24505 20644 24529 20646
rect 24289 20624 24585 20644
rect 24308 20460 24360 20466
rect 24308 20402 24360 20408
rect 24216 20324 24268 20330
rect 24216 20266 24268 20272
rect 24320 19990 24348 20402
rect 24688 20210 24716 21247
rect 24780 20618 24808 22471
rect 24872 21622 24900 25327
rect 25332 24177 25360 27520
rect 25780 25220 25832 25226
rect 25780 25162 25832 25168
rect 25792 24562 25820 25162
rect 25884 24721 25912 27520
rect 26054 26208 26110 26217
rect 26054 26143 26110 26152
rect 25962 25528 26018 25537
rect 25962 25463 26018 25472
rect 25870 24712 25926 24721
rect 25870 24647 25926 24656
rect 25792 24534 25912 24562
rect 25318 24168 25374 24177
rect 25318 24103 25374 24112
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 24860 21616 24912 21622
rect 24860 21558 24912 21564
rect 24780 20602 24900 20618
rect 24780 20596 24912 20602
rect 24780 20590 24860 20596
rect 24860 20538 24912 20544
rect 24688 20182 24900 20210
rect 24766 20088 24822 20097
rect 24766 20023 24822 20032
rect 24308 19984 24360 19990
rect 24308 19926 24360 19932
rect 24320 19700 24348 19926
rect 24228 19672 24348 19700
rect 24228 19514 24256 19672
rect 24289 19612 24585 19632
rect 24345 19610 24369 19612
rect 24425 19610 24449 19612
rect 24505 19610 24529 19612
rect 24367 19558 24369 19610
rect 24431 19558 24443 19610
rect 24505 19558 24507 19610
rect 24345 19556 24369 19558
rect 24425 19556 24449 19558
rect 24505 19556 24529 19558
rect 24289 19536 24585 19556
rect 24674 19544 24730 19553
rect 24216 19508 24268 19514
rect 24674 19479 24730 19488
rect 24216 19450 24268 19456
rect 24308 19440 24360 19446
rect 24308 19382 24360 19388
rect 24216 19372 24268 19378
rect 24216 19314 24268 19320
rect 24228 18970 24256 19314
rect 24216 18964 24268 18970
rect 24216 18906 24268 18912
rect 24320 18680 24348 19382
rect 24228 18652 24348 18680
rect 24228 18426 24256 18652
rect 24289 18524 24585 18544
rect 24345 18522 24369 18524
rect 24425 18522 24449 18524
rect 24505 18522 24529 18524
rect 24367 18470 24369 18522
rect 24431 18470 24443 18522
rect 24505 18470 24507 18522
rect 24345 18468 24369 18470
rect 24425 18468 24449 18470
rect 24505 18468 24529 18470
rect 24289 18448 24585 18468
rect 24216 18420 24268 18426
rect 24216 18362 24268 18368
rect 24214 18320 24270 18329
rect 24214 18255 24270 18264
rect 24124 16244 24176 16250
rect 24124 16186 24176 16192
rect 23860 16102 24072 16130
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23768 12918 23796 13466
rect 23756 12912 23808 12918
rect 23756 12854 23808 12860
rect 23754 12608 23810 12617
rect 23754 12543 23810 12552
rect 23768 10130 23796 12543
rect 23860 12374 23888 16102
rect 24136 16046 24164 16186
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 15638 24072 15846
rect 24032 15632 24084 15638
rect 24030 15600 24032 15609
rect 24084 15600 24086 15609
rect 24030 15535 24086 15544
rect 24044 15509 24072 15535
rect 24124 15360 24176 15366
rect 24124 15302 24176 15308
rect 23940 14952 23992 14958
rect 23940 14894 23992 14900
rect 23952 14113 23980 14894
rect 24032 14884 24084 14890
rect 24032 14826 24084 14832
rect 24044 14346 24072 14826
rect 24136 14822 24164 15302
rect 24228 15162 24256 18255
rect 24289 17436 24585 17456
rect 24345 17434 24369 17436
rect 24425 17434 24449 17436
rect 24505 17434 24529 17436
rect 24367 17382 24369 17434
rect 24431 17382 24443 17434
rect 24505 17382 24507 17434
rect 24345 17380 24369 17382
rect 24425 17380 24449 17382
rect 24505 17380 24529 17382
rect 24289 17360 24585 17380
rect 24688 17338 24716 19479
rect 24780 17898 24808 20023
rect 24872 18970 24900 20182
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 24964 18834 24992 22374
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25332 22001 25360 22034
rect 25318 21992 25374 22001
rect 25318 21927 25374 21936
rect 25332 21622 25360 21927
rect 25424 21690 25452 23015
rect 25780 21956 25832 21962
rect 25780 21898 25832 21904
rect 25502 21856 25558 21865
rect 25502 21791 25558 21800
rect 25412 21684 25464 21690
rect 25412 21626 25464 21632
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25136 21480 25188 21486
rect 25136 21422 25188 21428
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25056 20262 25084 20878
rect 25044 20256 25096 20262
rect 25042 20224 25044 20233
rect 25096 20224 25098 20233
rect 25042 20159 25098 20168
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 24952 18828 25004 18834
rect 24952 18770 25004 18776
rect 24964 18426 24992 18770
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 25056 17921 25084 19343
rect 25148 18034 25176 21422
rect 25410 20768 25466 20777
rect 25410 20703 25466 20712
rect 25226 19952 25282 19961
rect 25226 19887 25282 19896
rect 25240 18222 25268 19887
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25332 18154 25360 19246
rect 25424 18426 25452 20703
rect 25516 19174 25544 21791
rect 25594 20496 25650 20505
rect 25594 20431 25650 20440
rect 25608 19174 25636 20431
rect 25504 19168 25556 19174
rect 25504 19110 25556 19116
rect 25596 19168 25648 19174
rect 25596 19110 25648 19116
rect 25594 19000 25650 19009
rect 25594 18935 25650 18944
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25320 18148 25372 18154
rect 25320 18090 25372 18096
rect 25148 18006 25360 18034
rect 25042 17912 25098 17921
rect 24780 17882 24900 17898
rect 24780 17876 24912 17882
rect 24780 17870 24860 17876
rect 25042 17847 25098 17856
rect 24860 17818 24912 17824
rect 25044 17808 25096 17814
rect 25042 17776 25044 17785
rect 25096 17776 25098 17785
rect 25042 17711 25098 17720
rect 25136 17740 25188 17746
rect 25136 17682 25188 17688
rect 24950 17640 25006 17649
rect 24950 17575 25006 17584
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24768 17128 24820 17134
rect 24768 17070 24820 17076
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24289 16348 24585 16368
rect 24345 16346 24369 16348
rect 24425 16346 24449 16348
rect 24505 16346 24529 16348
rect 24367 16294 24369 16346
rect 24431 16294 24443 16346
rect 24505 16294 24507 16346
rect 24345 16292 24369 16294
rect 24425 16292 24449 16294
rect 24505 16292 24529 16294
rect 24289 16272 24585 16292
rect 24306 16008 24362 16017
rect 24306 15943 24362 15952
rect 24320 15609 24348 15943
rect 24490 15736 24546 15745
rect 24490 15671 24492 15680
rect 24544 15671 24546 15680
rect 24492 15642 24544 15648
rect 24306 15600 24362 15609
rect 24306 15535 24362 15544
rect 24289 15260 24585 15280
rect 24345 15258 24369 15260
rect 24425 15258 24449 15260
rect 24505 15258 24529 15260
rect 24367 15206 24369 15258
rect 24431 15206 24443 15258
rect 24505 15206 24507 15258
rect 24345 15204 24369 15206
rect 24425 15204 24449 15206
rect 24505 15204 24529 15206
rect 24289 15184 24585 15204
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24124 14816 24176 14822
rect 24122 14784 24124 14793
rect 24176 14784 24178 14793
rect 24122 14719 24178 14728
rect 24122 14648 24178 14657
rect 24122 14583 24178 14592
rect 24032 14340 24084 14346
rect 24032 14282 24084 14288
rect 24030 14240 24086 14249
rect 24030 14175 24086 14184
rect 23938 14104 23994 14113
rect 24044 14074 24072 14175
rect 23938 14039 23994 14048
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23938 13968 23994 13977
rect 23938 13903 23994 13912
rect 23952 12986 23980 13903
rect 24030 13560 24086 13569
rect 24030 13495 24086 13504
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23940 12640 23992 12646
rect 23940 12582 23992 12588
rect 23848 12368 23900 12374
rect 23848 12310 23900 12316
rect 23848 12164 23900 12170
rect 23848 12106 23900 12112
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23400 9518 23428 9930
rect 23584 9602 23612 10118
rect 23664 10124 23716 10130
rect 23664 10066 23716 10072
rect 23756 10124 23808 10130
rect 23756 10066 23808 10072
rect 23676 9722 23704 10066
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23584 9574 23796 9602
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23296 9376 23348 9382
rect 23296 9318 23348 9324
rect 23308 9081 23336 9318
rect 23386 9208 23442 9217
rect 23386 9143 23442 9152
rect 23294 9072 23350 9081
rect 23294 9007 23350 9016
rect 23400 8906 23428 9143
rect 23388 8900 23440 8906
rect 23388 8842 23440 8848
rect 23662 8528 23718 8537
rect 23216 8486 23336 8514
rect 23202 8392 23258 8401
rect 23202 8327 23204 8336
rect 23256 8327 23258 8336
rect 23204 8298 23256 8304
rect 23110 8120 23166 8129
rect 23110 8055 23166 8064
rect 22926 7984 22982 7993
rect 22744 7948 22796 7954
rect 23308 7954 23336 8486
rect 23572 8492 23624 8498
rect 23662 8463 23718 8472
rect 23572 8434 23624 8440
rect 23480 8356 23532 8362
rect 23400 8316 23480 8344
rect 22926 7919 22982 7928
rect 23296 7948 23348 7954
rect 22744 7890 22796 7896
rect 22756 7206 22784 7890
rect 22836 7812 22888 7818
rect 22836 7754 22888 7760
rect 22744 7200 22796 7206
rect 22742 7168 22744 7177
rect 22796 7168 22798 7177
rect 22742 7103 22798 7112
rect 22742 6216 22798 6225
rect 22742 6151 22744 6160
rect 22796 6151 22798 6160
rect 22744 6122 22796 6128
rect 22848 5846 22876 7754
rect 22940 5914 22968 7919
rect 23296 7890 23348 7896
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 23032 7546 23060 7822
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23296 7744 23348 7750
rect 23296 7686 23348 7692
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23032 6934 23060 7482
rect 23020 6928 23072 6934
rect 23020 6870 23072 6876
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23124 6254 23152 6734
rect 23112 6248 23164 6254
rect 23112 6190 23164 6196
rect 23018 6080 23074 6089
rect 23018 6015 23074 6024
rect 22928 5908 22980 5914
rect 22928 5850 22980 5856
rect 22836 5840 22888 5846
rect 22836 5782 22888 5788
rect 22848 5302 22876 5782
rect 22940 5370 22968 5850
rect 23032 5710 23060 6015
rect 23216 5846 23244 7686
rect 23308 6730 23336 7686
rect 23400 7585 23428 8316
rect 23480 8298 23532 8304
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23386 7576 23442 7585
rect 23386 7511 23442 7520
rect 23492 7041 23520 7822
rect 23478 7032 23534 7041
rect 23478 6967 23534 6976
rect 23388 6860 23440 6866
rect 23440 6820 23520 6848
rect 23388 6802 23440 6808
rect 23296 6724 23348 6730
rect 23296 6666 23348 6672
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23400 6458 23428 6666
rect 23388 6452 23440 6458
rect 23388 6394 23440 6400
rect 23296 6384 23348 6390
rect 23296 6326 23348 6332
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 23020 5704 23072 5710
rect 23020 5646 23072 5652
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 22836 5296 22888 5302
rect 22836 5238 22888 5244
rect 22834 4856 22890 4865
rect 23032 4826 23060 5646
rect 23308 5386 23336 6326
rect 23124 5358 23336 5386
rect 23492 5370 23520 6820
rect 23584 6769 23612 8434
rect 23676 8430 23704 8463
rect 23664 8424 23716 8430
rect 23664 8366 23716 8372
rect 23768 7154 23796 9574
rect 23860 9110 23888 12106
rect 23952 11354 23980 12582
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 24044 10742 24072 13495
rect 24136 12617 24164 14583
rect 24216 14476 24268 14482
rect 24216 14418 24268 14424
rect 24228 13938 24256 14418
rect 24688 14414 24716 16390
rect 24780 15434 24808 17070
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24872 16561 24900 16662
rect 24858 16552 24914 16561
rect 24858 16487 24914 16496
rect 24858 16144 24914 16153
rect 24858 16079 24914 16088
rect 24872 15706 24900 16079
rect 24860 15700 24912 15706
rect 24860 15642 24912 15648
rect 24964 15638 24992 17575
rect 25148 16998 25176 17682
rect 25228 17128 25280 17134
rect 25226 17096 25228 17105
rect 25280 17096 25282 17105
rect 25226 17031 25282 17040
rect 25136 16992 25188 16998
rect 25136 16934 25188 16940
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 15910 25084 16526
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24952 15632 25004 15638
rect 24872 15580 24952 15586
rect 24872 15574 25004 15580
rect 24872 15558 24992 15574
rect 24768 15428 24820 15434
rect 24768 15370 24820 15376
rect 24872 15094 24900 15558
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24860 15088 24912 15094
rect 24860 15030 24912 15036
rect 24964 14958 24992 15438
rect 24952 14952 25004 14958
rect 24766 14920 24822 14929
rect 24952 14894 25004 14900
rect 24766 14855 24822 14864
rect 24676 14408 24728 14414
rect 24676 14350 24728 14356
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24289 14172 24585 14192
rect 24345 14170 24369 14172
rect 24425 14170 24449 14172
rect 24505 14170 24529 14172
rect 24367 14118 24369 14170
rect 24431 14118 24443 14170
rect 24505 14118 24507 14170
rect 24345 14116 24369 14118
rect 24425 14116 24449 14118
rect 24505 14116 24529 14118
rect 24289 14096 24585 14116
rect 24216 13932 24268 13938
rect 24216 13874 24268 13880
rect 24228 13326 24256 13874
rect 24688 13705 24716 14214
rect 24780 13954 24808 14855
rect 24950 14784 25006 14793
rect 24950 14719 25006 14728
rect 24964 14618 24992 14719
rect 24952 14612 25004 14618
rect 24952 14554 25004 14560
rect 24860 14476 24912 14482
rect 24860 14418 24912 14424
rect 24872 14074 24900 14418
rect 24964 14346 24992 14554
rect 24952 14340 25004 14346
rect 24952 14282 25004 14288
rect 24964 14074 24992 14282
rect 24860 14068 24912 14074
rect 24860 14010 24912 14016
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 24780 13926 24900 13954
rect 24872 13870 24900 13926
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24674 13696 24730 13705
rect 24674 13631 24730 13640
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24216 13320 24268 13326
rect 24216 13262 24268 13268
rect 24228 12986 24256 13262
rect 24289 13084 24585 13104
rect 24345 13082 24369 13084
rect 24425 13082 24449 13084
rect 24505 13082 24529 13084
rect 24367 13030 24369 13082
rect 24431 13030 24443 13082
rect 24505 13030 24507 13082
rect 24345 13028 24369 13030
rect 24425 13028 24449 13030
rect 24505 13028 24529 13030
rect 24289 13008 24585 13028
rect 24216 12980 24268 12986
rect 24216 12922 24268 12928
rect 24308 12912 24360 12918
rect 24228 12860 24308 12866
rect 24228 12854 24360 12860
rect 24228 12838 24348 12854
rect 24122 12608 24178 12617
rect 24122 12543 24178 12552
rect 24228 12442 24256 12838
rect 24780 12782 24808 13330
rect 25056 13297 25084 15846
rect 25148 13433 25176 16934
rect 25228 16040 25280 16046
rect 25228 15982 25280 15988
rect 25240 14482 25268 15982
rect 25332 15978 25360 18006
rect 25410 17776 25466 17785
rect 25410 17711 25466 17720
rect 25424 16250 25452 17711
rect 25502 17232 25558 17241
rect 25502 17167 25558 17176
rect 25412 16244 25464 16250
rect 25412 16186 25464 16192
rect 25410 16008 25466 16017
rect 25320 15972 25372 15978
rect 25410 15943 25466 15952
rect 25320 15914 25372 15920
rect 25318 15600 25374 15609
rect 25318 15535 25374 15544
rect 25332 15337 25360 15535
rect 25318 15328 25374 15337
rect 25318 15263 25374 15272
rect 25318 14920 25374 14929
rect 25318 14855 25374 14864
rect 25228 14476 25280 14482
rect 25228 14418 25280 14424
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 13977 25268 14214
rect 25226 13968 25282 13977
rect 25226 13903 25282 13912
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25134 13424 25190 13433
rect 25134 13359 25190 13368
rect 25042 13288 25098 13297
rect 25042 13223 25098 13232
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 24768 12776 24820 12782
rect 24768 12718 24820 12724
rect 24308 12708 24360 12714
rect 24308 12650 24360 12656
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24320 12306 24348 12650
rect 24674 12608 24730 12617
rect 24674 12543 24730 12552
rect 24582 12472 24638 12481
rect 24582 12407 24638 12416
rect 24308 12300 24360 12306
rect 24136 12260 24308 12288
rect 24136 12073 24164 12260
rect 24308 12242 24360 12248
rect 24596 12170 24624 12407
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24122 12064 24178 12073
rect 24122 11999 24178 12008
rect 24289 11996 24585 12016
rect 24345 11994 24369 11996
rect 24425 11994 24449 11996
rect 24505 11994 24529 11996
rect 24367 11942 24369 11994
rect 24431 11942 24443 11994
rect 24505 11942 24507 11994
rect 24345 11940 24369 11942
rect 24425 11940 24449 11942
rect 24505 11940 24529 11942
rect 24122 11928 24178 11937
rect 24289 11920 24585 11940
rect 24122 11863 24178 11872
rect 24136 11354 24164 11863
rect 24584 11824 24636 11830
rect 24584 11766 24636 11772
rect 24216 11552 24268 11558
rect 24596 11529 24624 11766
rect 24216 11494 24268 11500
rect 24582 11520 24638 11529
rect 24124 11348 24176 11354
rect 24124 11290 24176 11296
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24032 10736 24084 10742
rect 23938 10704 23994 10713
rect 24032 10678 24084 10684
rect 23938 10639 23994 10648
rect 23952 10606 23980 10639
rect 23940 10600 23992 10606
rect 23940 10542 23992 10548
rect 24136 10538 24164 11086
rect 24228 11014 24256 11494
rect 24582 11455 24638 11464
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24124 10532 24176 10538
rect 24124 10474 24176 10480
rect 23940 10464 23992 10470
rect 23940 10406 23992 10412
rect 23848 9104 23900 9110
rect 23848 9046 23900 9052
rect 23848 8288 23900 8294
rect 23952 8265 23980 10406
rect 24032 10192 24084 10198
rect 24030 10160 24032 10169
rect 24084 10160 24086 10169
rect 24030 10095 24086 10104
rect 24124 10124 24176 10130
rect 24124 10066 24176 10072
rect 24136 9722 24164 10066
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 24136 8634 24164 8978
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 23848 8230 23900 8236
rect 23938 8256 23994 8265
rect 23860 7342 23888 8230
rect 23938 8191 23994 8200
rect 23848 7336 23900 7342
rect 23848 7278 23900 7284
rect 23768 7126 23888 7154
rect 23756 6996 23808 7002
rect 23756 6938 23808 6944
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23570 6760 23626 6769
rect 23570 6695 23626 6704
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23480 5364 23532 5370
rect 22834 4791 22890 4800
rect 23020 4820 23072 4826
rect 22848 4690 22876 4791
rect 23020 4762 23072 4768
rect 22836 4684 22888 4690
rect 22836 4626 22888 4632
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 22848 3738 22876 4626
rect 22940 4282 22968 4626
rect 23020 4616 23072 4622
rect 23020 4558 23072 4564
rect 22928 4276 22980 4282
rect 22928 4218 22980 4224
rect 23032 4078 23060 4558
rect 23124 4554 23152 5358
rect 23480 5306 23532 5312
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23020 3936 23072 3942
rect 23020 3878 23072 3884
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22836 3596 22888 3602
rect 22836 3538 22888 3544
rect 22928 3596 22980 3602
rect 22928 3538 22980 3544
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22756 2553 22784 2858
rect 22742 2544 22798 2553
rect 22742 2479 22798 2488
rect 22848 2417 22876 3538
rect 22940 2990 22968 3538
rect 23032 3534 23060 3878
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23032 3126 23060 3470
rect 23124 3126 23152 4490
rect 23020 3120 23072 3126
rect 23020 3062 23072 3068
rect 23112 3120 23164 3126
rect 23112 3062 23164 3068
rect 22928 2984 22980 2990
rect 22928 2926 22980 2932
rect 22940 2689 22968 2926
rect 22926 2680 22982 2689
rect 23216 2650 23244 5170
rect 23584 4842 23612 6598
rect 23676 6322 23704 6802
rect 23664 6316 23716 6322
rect 23664 6258 23716 6264
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5914 23704 6054
rect 23664 5908 23716 5914
rect 23664 5850 23716 5856
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 23676 5001 23704 5714
rect 23768 5642 23796 6938
rect 23860 6390 23888 7126
rect 23952 6390 23980 8191
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7002 24072 7686
rect 24228 7478 24256 10950
rect 24289 10908 24585 10928
rect 24345 10906 24369 10908
rect 24425 10906 24449 10908
rect 24505 10906 24529 10908
rect 24367 10854 24369 10906
rect 24431 10854 24443 10906
rect 24505 10854 24507 10906
rect 24345 10852 24369 10854
rect 24425 10852 24449 10854
rect 24505 10852 24529 10854
rect 24289 10832 24585 10852
rect 24289 9820 24585 9840
rect 24345 9818 24369 9820
rect 24425 9818 24449 9820
rect 24505 9818 24529 9820
rect 24367 9766 24369 9818
rect 24431 9766 24443 9818
rect 24505 9766 24507 9818
rect 24345 9764 24369 9766
rect 24425 9764 24449 9766
rect 24505 9764 24529 9766
rect 24289 9744 24585 9764
rect 24688 9654 24716 12543
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 24768 12164 24820 12170
rect 24768 12106 24820 12112
rect 24780 11354 24808 12106
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24872 11801 24900 12038
rect 24858 11792 24914 11801
rect 24858 11727 24914 11736
rect 24964 11694 24992 12242
rect 24952 11688 25004 11694
rect 24950 11656 24952 11665
rect 25004 11656 25006 11665
rect 24950 11591 25006 11600
rect 24858 11520 24914 11529
rect 24858 11455 24914 11464
rect 24768 11348 24820 11354
rect 24768 11290 24820 11296
rect 24780 10266 24808 11290
rect 24768 10260 24820 10266
rect 24768 10202 24820 10208
rect 24872 10146 24900 11455
rect 24950 11384 25006 11393
rect 24950 11319 25006 11328
rect 24780 10118 24900 10146
rect 24964 10130 24992 11319
rect 24952 10124 25004 10130
rect 24676 9648 24728 9654
rect 24582 9616 24638 9625
rect 24676 9590 24728 9596
rect 24582 9551 24638 9560
rect 24596 9466 24624 9551
rect 24596 9438 24716 9466
rect 24398 9344 24454 9353
rect 24398 9279 24454 9288
rect 24412 9178 24440 9279
rect 24400 9172 24452 9178
rect 24400 9114 24452 9120
rect 24688 8809 24716 9438
rect 24780 9178 24808 10118
rect 24952 10066 25004 10072
rect 24860 9512 24912 9518
rect 24858 9480 24860 9489
rect 24912 9480 24914 9489
rect 24858 9415 24914 9424
rect 24768 9172 24820 9178
rect 24768 9114 24820 9120
rect 24858 9072 24914 9081
rect 24858 9007 24860 9016
rect 24912 9007 24914 9016
rect 24860 8978 24912 8984
rect 24674 8800 24730 8809
rect 24289 8732 24585 8752
rect 24674 8735 24730 8744
rect 24345 8730 24369 8732
rect 24425 8730 24449 8732
rect 24505 8730 24529 8732
rect 24367 8678 24369 8730
rect 24431 8678 24443 8730
rect 24505 8678 24507 8730
rect 24345 8676 24369 8678
rect 24425 8676 24449 8678
rect 24505 8676 24529 8678
rect 24289 8656 24585 8676
rect 24860 8560 24912 8566
rect 24858 8528 24860 8537
rect 24912 8528 24914 8537
rect 24858 8463 24914 8472
rect 25056 7954 25084 13126
rect 25240 12782 25268 13670
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25228 12232 25280 12238
rect 25148 12192 25228 12220
rect 25148 11762 25176 12192
rect 25228 12174 25280 12180
rect 25332 11898 25360 14855
rect 25424 12986 25452 15943
rect 25516 14074 25544 17167
rect 25608 16794 25636 18935
rect 25792 17746 25820 21898
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 25780 17536 25832 17542
rect 25780 17478 25832 17484
rect 25688 17332 25740 17338
rect 25688 17274 25740 17280
rect 25596 16788 25648 16794
rect 25596 16730 25648 16736
rect 25594 15328 25650 15337
rect 25594 15263 25650 15272
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25608 13326 25636 15263
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25504 13184 25556 13190
rect 25504 13126 25556 13132
rect 25596 13184 25648 13190
rect 25596 13126 25648 13132
rect 25412 12980 25464 12986
rect 25412 12922 25464 12928
rect 25516 12889 25544 13126
rect 25502 12880 25558 12889
rect 25502 12815 25558 12824
rect 25412 12776 25464 12782
rect 25412 12718 25464 12724
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25424 11778 25452 12718
rect 25608 12714 25636 13126
rect 25596 12708 25648 12714
rect 25596 12650 25648 12656
rect 25502 12472 25558 12481
rect 25502 12407 25558 12416
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25332 11750 25452 11778
rect 25148 11354 25176 11698
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25228 11280 25280 11286
rect 25228 11222 25280 11228
rect 25134 10976 25190 10985
rect 25134 10911 25190 10920
rect 25148 10266 25176 10911
rect 25240 10810 25268 11222
rect 25332 11150 25360 11750
rect 25412 11280 25464 11286
rect 25410 11248 25412 11257
rect 25464 11248 25466 11257
rect 25410 11183 25466 11192
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25410 10976 25466 10985
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25332 10033 25360 10950
rect 25410 10911 25466 10920
rect 25424 10470 25452 10911
rect 25412 10464 25464 10470
rect 25412 10406 25464 10412
rect 25318 10024 25374 10033
rect 25318 9959 25374 9968
rect 25134 9208 25190 9217
rect 25134 9143 25190 9152
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 25044 7948 25096 7954
rect 25044 7890 25096 7896
rect 24289 7644 24585 7664
rect 24345 7642 24369 7644
rect 24425 7642 24449 7644
rect 24505 7642 24529 7644
rect 24367 7590 24369 7642
rect 24431 7590 24443 7642
rect 24505 7590 24507 7642
rect 24345 7588 24369 7590
rect 24425 7588 24449 7590
rect 24505 7588 24529 7590
rect 24289 7568 24585 7588
rect 24780 7546 24808 7890
rect 24952 7744 25004 7750
rect 24952 7686 25004 7692
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24216 7472 24268 7478
rect 24216 7414 24268 7420
rect 24768 7336 24820 7342
rect 24768 7278 24820 7284
rect 24124 7200 24176 7206
rect 24176 7160 24256 7188
rect 24124 7142 24176 7148
rect 24032 6996 24084 7002
rect 24032 6938 24084 6944
rect 24032 6860 24084 6866
rect 24032 6802 24084 6808
rect 24044 6458 24072 6802
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 23848 6384 23900 6390
rect 23848 6326 23900 6332
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 24124 6316 24176 6322
rect 24124 6258 24176 6264
rect 23848 6180 23900 6186
rect 23848 6122 23900 6128
rect 23756 5636 23808 5642
rect 23756 5578 23808 5584
rect 23756 5296 23808 5302
rect 23754 5264 23756 5273
rect 23808 5264 23810 5273
rect 23754 5199 23810 5208
rect 23662 4992 23718 5001
rect 23662 4927 23718 4936
rect 23308 4814 23612 4842
rect 22926 2615 22982 2624
rect 23204 2644 23256 2650
rect 23204 2586 23256 2592
rect 22834 2408 22890 2417
rect 22834 2343 22890 2352
rect 22928 2304 22980 2310
rect 22928 2246 22980 2252
rect 22940 1465 22968 2246
rect 22926 1456 22982 1465
rect 22926 1391 22982 1400
rect 23308 1170 23336 4814
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23480 4140 23532 4146
rect 23480 4082 23532 4088
rect 23492 3942 23520 4082
rect 23584 4078 23612 4422
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 23756 4004 23808 4010
rect 23756 3946 23808 3952
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23492 3505 23520 3878
rect 23572 3528 23624 3534
rect 23478 3496 23534 3505
rect 23572 3470 23624 3476
rect 23478 3431 23534 3440
rect 23480 3392 23532 3398
rect 23478 3360 23480 3369
rect 23532 3360 23534 3369
rect 23478 3295 23534 3304
rect 23478 3224 23534 3233
rect 23478 3159 23480 3168
rect 23532 3159 23534 3168
rect 23480 3130 23532 3136
rect 23492 2922 23520 3130
rect 23584 2990 23612 3470
rect 23676 3369 23704 3878
rect 23662 3360 23718 3369
rect 23662 3295 23718 3304
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23584 2650 23612 2926
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23572 2644 23624 2650
rect 23572 2586 23624 2592
rect 23676 2446 23704 2790
rect 23664 2440 23716 2446
rect 23664 2382 23716 2388
rect 23216 1142 23336 1170
rect 23216 480 23244 1142
rect 23768 480 23796 3946
rect 23860 3058 23888 6122
rect 23938 6080 23994 6089
rect 23938 6015 23994 6024
rect 23952 4010 23980 6015
rect 24030 5672 24086 5681
rect 24030 5607 24032 5616
rect 24084 5607 24086 5616
rect 24032 5578 24084 5584
rect 24030 5536 24086 5545
rect 24030 5471 24086 5480
rect 24044 5166 24072 5471
rect 24136 5234 24164 6258
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24032 5160 24084 5166
rect 24032 5102 24084 5108
rect 24044 4826 24072 5102
rect 24136 4826 24164 5170
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 24122 4720 24178 4729
rect 24122 4655 24178 4664
rect 24136 4282 24164 4655
rect 24124 4276 24176 4282
rect 24124 4218 24176 4224
rect 23940 4004 23992 4010
rect 23940 3946 23992 3952
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 23938 3768 23994 3777
rect 23938 3703 23994 3712
rect 23952 3466 23980 3703
rect 23940 3460 23992 3466
rect 23940 3402 23992 3408
rect 23952 3058 23980 3402
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23940 3052 23992 3058
rect 23940 2994 23992 3000
rect 24044 2514 24072 3334
rect 24136 2650 24164 3878
rect 24124 2644 24176 2650
rect 24124 2586 24176 2592
rect 24032 2508 24084 2514
rect 24032 2450 24084 2456
rect 24124 2508 24176 2514
rect 24124 2450 24176 2456
rect 23848 2304 23900 2310
rect 23846 2272 23848 2281
rect 23900 2272 23902 2281
rect 23846 2207 23902 2216
rect 24136 1057 24164 2450
rect 24228 1442 24256 7160
rect 24780 7002 24808 7278
rect 24964 7041 24992 7686
rect 25056 7546 25084 7890
rect 25044 7540 25096 7546
rect 25044 7482 25096 7488
rect 24950 7032 25006 7041
rect 24768 6996 24820 7002
rect 24950 6967 25006 6976
rect 24768 6938 24820 6944
rect 24766 6896 24822 6905
rect 24766 6831 24822 6840
rect 24289 6556 24585 6576
rect 24345 6554 24369 6556
rect 24425 6554 24449 6556
rect 24505 6554 24529 6556
rect 24367 6502 24369 6554
rect 24431 6502 24443 6554
rect 24505 6502 24507 6554
rect 24345 6500 24369 6502
rect 24425 6500 24449 6502
rect 24505 6500 24529 6502
rect 24289 6480 24585 6500
rect 24780 6497 24808 6831
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24766 6488 24822 6497
rect 24766 6423 24822 6432
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24320 6186 24348 6326
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24766 6216 24822 6225
rect 24308 6180 24360 6186
rect 24308 6122 24360 6128
rect 24320 5642 24348 6122
rect 24688 5710 24716 6190
rect 24766 6151 24822 6160
rect 24676 5704 24728 5710
rect 24676 5646 24728 5652
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24289 5468 24585 5488
rect 24345 5466 24369 5468
rect 24425 5466 24449 5468
rect 24505 5466 24529 5468
rect 24367 5414 24369 5466
rect 24431 5414 24443 5466
rect 24505 5414 24507 5466
rect 24345 5412 24369 5414
rect 24425 5412 24449 5414
rect 24505 5412 24529 5414
rect 24289 5392 24585 5412
rect 24688 5370 24716 5646
rect 24676 5364 24728 5370
rect 24676 5306 24728 5312
rect 24780 4729 24808 6151
rect 24490 4720 24546 4729
rect 24490 4655 24492 4664
rect 24544 4655 24546 4664
rect 24766 4720 24822 4729
rect 24766 4655 24822 4664
rect 24492 4626 24544 4632
rect 24676 4480 24728 4486
rect 24676 4422 24728 4428
rect 24768 4480 24820 4486
rect 24768 4422 24820 4428
rect 24289 4380 24585 4400
rect 24345 4378 24369 4380
rect 24425 4378 24449 4380
rect 24505 4378 24529 4380
rect 24367 4326 24369 4378
rect 24431 4326 24443 4378
rect 24505 4326 24507 4378
rect 24345 4324 24369 4326
rect 24425 4324 24449 4326
rect 24505 4324 24529 4326
rect 24289 4304 24585 4324
rect 24306 4040 24362 4049
rect 24306 3975 24362 3984
rect 24490 4040 24546 4049
rect 24490 3975 24546 3984
rect 24320 3670 24348 3975
rect 24504 3738 24532 3975
rect 24492 3732 24544 3738
rect 24492 3674 24544 3680
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 24688 3369 24716 4422
rect 24780 3942 24808 4422
rect 24768 3936 24820 3942
rect 24768 3878 24820 3884
rect 24766 3768 24822 3777
rect 24766 3703 24822 3712
rect 24674 3360 24730 3369
rect 24289 3292 24585 3312
rect 24674 3295 24730 3304
rect 24345 3290 24369 3292
rect 24425 3290 24449 3292
rect 24505 3290 24529 3292
rect 24367 3238 24369 3290
rect 24431 3238 24443 3290
rect 24505 3238 24507 3290
rect 24345 3236 24369 3238
rect 24425 3236 24449 3238
rect 24505 3236 24529 3238
rect 24289 3216 24585 3236
rect 24676 3188 24728 3194
rect 24676 3130 24728 3136
rect 24584 3120 24636 3126
rect 24584 3062 24636 3068
rect 24596 2292 24624 3062
rect 24688 2394 24716 3130
rect 24780 2514 24808 3703
rect 24768 2508 24820 2514
rect 24768 2450 24820 2456
rect 24688 2366 24808 2394
rect 24596 2264 24716 2292
rect 24289 2204 24585 2224
rect 24345 2202 24369 2204
rect 24425 2202 24449 2204
rect 24505 2202 24529 2204
rect 24367 2150 24369 2202
rect 24431 2150 24443 2202
rect 24505 2150 24507 2202
rect 24345 2148 24369 2150
rect 24425 2148 24449 2150
rect 24505 2148 24529 2150
rect 24289 2128 24585 2148
rect 24688 1465 24716 2264
rect 24674 1456 24730 1465
rect 24228 1414 24348 1442
rect 24122 1048 24178 1057
rect 24122 983 24178 992
rect 24320 480 24348 1414
rect 24674 1391 24730 1400
rect 24780 1329 24808 2366
rect 24766 1320 24822 1329
rect 24766 1255 24822 1264
rect 24872 480 24900 6598
rect 25148 6458 25176 9143
rect 25516 8634 25544 12407
rect 25596 12300 25648 12306
rect 25596 12242 25648 12248
rect 25608 11558 25636 12242
rect 25596 11552 25648 11558
rect 25596 11494 25648 11500
rect 25608 11218 25636 11494
rect 25596 11212 25648 11218
rect 25596 11154 25648 11160
rect 25700 10266 25728 17274
rect 25792 11354 25820 17478
rect 25780 11348 25832 11354
rect 25780 11290 25832 11296
rect 25780 11212 25832 11218
rect 25780 11154 25832 11160
rect 25688 10260 25740 10266
rect 25688 10202 25740 10208
rect 25596 9648 25648 9654
rect 25594 9616 25596 9625
rect 25648 9616 25650 9625
rect 25594 9551 25650 9560
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 25226 8120 25282 8129
rect 25226 8055 25282 8064
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25148 6254 25176 6394
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 25044 5024 25096 5030
rect 25044 4966 25096 4972
rect 25136 5024 25188 5030
rect 25136 4966 25188 4972
rect 25056 4865 25084 4966
rect 25042 4856 25098 4865
rect 25042 4791 25098 4800
rect 25044 3936 25096 3942
rect 25042 3904 25044 3913
rect 25096 3904 25098 3913
rect 25042 3839 25098 3848
rect 24952 3596 25004 3602
rect 24952 3538 25004 3544
rect 24964 3194 24992 3538
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24952 3188 25004 3194
rect 24952 3130 25004 3136
rect 25056 3097 25084 3334
rect 25042 3088 25098 3097
rect 25042 3023 25098 3032
rect 25148 2961 25176 4966
rect 25240 4078 25268 8055
rect 25504 7812 25556 7818
rect 25504 7754 25556 7760
rect 25320 7744 25372 7750
rect 25320 7686 25372 7692
rect 25228 4072 25280 4078
rect 25332 4049 25360 7686
rect 25412 6112 25464 6118
rect 25410 6080 25412 6089
rect 25464 6080 25466 6089
rect 25410 6015 25466 6024
rect 25228 4014 25280 4020
rect 25318 4040 25374 4049
rect 25318 3975 25374 3984
rect 25412 3936 25464 3942
rect 25412 3878 25464 3884
rect 25228 3732 25280 3738
rect 25228 3674 25280 3680
rect 25240 3126 25268 3674
rect 25424 3505 25452 3878
rect 25410 3496 25466 3505
rect 25410 3431 25466 3440
rect 25228 3120 25280 3126
rect 25228 3062 25280 3068
rect 25228 2984 25280 2990
rect 25134 2952 25190 2961
rect 25228 2926 25280 2932
rect 25134 2887 25190 2896
rect 25136 2848 25188 2854
rect 25134 2816 25136 2825
rect 25188 2816 25190 2825
rect 25134 2751 25190 2760
rect 24950 2680 25006 2689
rect 24950 2615 24952 2624
rect 25004 2615 25006 2624
rect 24952 2586 25004 2592
rect 25240 1601 25268 2926
rect 25516 2802 25544 7754
rect 25332 2774 25544 2802
rect 25332 2666 25360 2774
rect 25332 2638 25452 2666
rect 25226 1592 25282 1601
rect 25226 1527 25282 1536
rect 25424 480 25452 2638
rect 25608 785 25636 8774
rect 25688 7744 25740 7750
rect 25792 7721 25820 11154
rect 25884 9178 25912 24534
rect 25976 17542 26004 25463
rect 25964 17536 26016 17542
rect 25964 17478 26016 17484
rect 26068 17338 26096 26143
rect 26528 24449 26556 27520
rect 26514 24440 26570 24449
rect 26514 24375 26570 24384
rect 27080 23633 27108 27520
rect 27252 24676 27304 24682
rect 27252 24618 27304 24624
rect 27264 23633 27292 24618
rect 27632 23905 27660 27520
rect 27618 23896 27674 23905
rect 27618 23831 27674 23840
rect 27066 23624 27122 23633
rect 27066 23559 27122 23568
rect 27250 23624 27306 23633
rect 27250 23559 27306 23568
rect 26148 21888 26200 21894
rect 26148 21830 26200 21836
rect 26056 17332 26108 17338
rect 26056 17274 26108 17280
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 25964 15428 26016 15434
rect 25964 15370 26016 15376
rect 25976 15162 26004 15370
rect 25964 15156 26016 15162
rect 25964 15098 26016 15104
rect 25962 13152 26018 13161
rect 25962 13087 26018 13096
rect 25976 9994 26004 13087
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25872 9172 25924 9178
rect 25872 9114 25924 9120
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25870 8256 25926 8265
rect 25870 8191 25926 8200
rect 25688 7686 25740 7692
rect 25778 7712 25834 7721
rect 25700 7449 25728 7686
rect 25778 7647 25834 7656
rect 25778 7576 25834 7585
rect 25884 7546 25912 8191
rect 25778 7511 25780 7520
rect 25832 7511 25834 7520
rect 25872 7540 25924 7546
rect 25780 7482 25832 7488
rect 25872 7482 25924 7488
rect 25686 7440 25742 7449
rect 25976 7426 26004 8910
rect 26068 8634 26096 16458
rect 26160 14657 26188 21830
rect 26240 20868 26292 20874
rect 26240 20810 26292 20816
rect 26252 20602 26280 20810
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26332 19168 26384 19174
rect 26332 19110 26384 19116
rect 26146 14648 26202 14657
rect 26146 14583 26202 14592
rect 26344 14498 26372 19110
rect 26160 14470 26372 14498
rect 26160 8974 26188 14470
rect 26240 13864 26292 13870
rect 26238 13832 26240 13841
rect 26292 13832 26294 13841
rect 26238 13767 26294 13776
rect 26330 13696 26386 13705
rect 26330 13631 26386 13640
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26252 12753 26280 13126
rect 26344 12986 26372 13631
rect 26332 12980 26384 12986
rect 26332 12922 26384 12928
rect 26238 12744 26294 12753
rect 26238 12679 26294 12688
rect 26238 12336 26294 12345
rect 26238 12271 26294 12280
rect 26252 11898 26280 12271
rect 26240 11892 26292 11898
rect 26240 11834 26292 11840
rect 26332 10464 26384 10470
rect 26330 10432 26332 10441
rect 26384 10432 26386 10441
rect 26330 10367 26386 10376
rect 26330 10296 26386 10305
rect 26330 10231 26332 10240
rect 26384 10231 26386 10240
rect 26332 10202 26384 10208
rect 26332 9648 26384 9654
rect 26330 9616 26332 9625
rect 26384 9616 26386 9625
rect 26330 9551 26386 9560
rect 26148 8968 26200 8974
rect 26148 8910 26200 8916
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26056 8628 26108 8634
rect 26056 8570 26108 8576
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 25686 7375 25742 7384
rect 25884 7398 26004 7426
rect 25780 6792 25832 6798
rect 25780 6734 25832 6740
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25700 5137 25728 6598
rect 25792 6458 25820 6734
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 25780 5840 25832 5846
rect 25778 5808 25780 5817
rect 25832 5808 25834 5817
rect 25778 5743 25834 5752
rect 25884 5370 25912 7398
rect 25964 7200 26016 7206
rect 26068 7177 26096 7686
rect 25964 7142 26016 7148
rect 26054 7168 26110 7177
rect 25872 5364 25924 5370
rect 25872 5306 25924 5312
rect 25780 5296 25832 5302
rect 25780 5238 25832 5244
rect 25686 5128 25742 5137
rect 25686 5063 25742 5072
rect 25686 4992 25742 5001
rect 25686 4927 25742 4936
rect 25700 1737 25728 4927
rect 25792 4706 25820 5238
rect 25884 5166 25912 5306
rect 25872 5160 25924 5166
rect 25872 5102 25924 5108
rect 25792 4678 25912 4706
rect 25780 4616 25832 4622
rect 25778 4584 25780 4593
rect 25832 4584 25834 4593
rect 25778 4519 25834 4528
rect 25884 2650 25912 4678
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25686 1728 25742 1737
rect 25686 1663 25742 1672
rect 25594 776 25650 785
rect 25594 711 25650 720
rect 25976 480 26004 7142
rect 26054 7103 26110 7112
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 26068 5778 26096 6598
rect 26056 5772 26108 5778
rect 26056 5714 26108 5720
rect 26068 2514 26096 5714
rect 26056 2508 26108 2514
rect 26056 2450 26108 2456
rect 26160 513 26188 8774
rect 26330 8664 26386 8673
rect 26330 8599 26332 8608
rect 26384 8599 26386 8608
rect 26332 8570 26384 8576
rect 26424 7336 26476 7342
rect 26422 7304 26424 7313
rect 26476 7304 26478 7313
rect 26422 7239 26478 7248
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26252 5953 26280 6054
rect 26238 5944 26294 5953
rect 26238 5879 26294 5888
rect 26424 5568 26476 5574
rect 26424 5510 26476 5516
rect 26332 5092 26384 5098
rect 26332 5034 26384 5040
rect 26240 4480 26292 4486
rect 26240 4422 26292 4428
rect 26252 4185 26280 4422
rect 26238 4176 26294 4185
rect 26238 4111 26294 4120
rect 26240 3664 26292 3670
rect 26238 3632 26240 3641
rect 26292 3632 26294 3641
rect 26238 3567 26294 3576
rect 26344 3233 26372 5034
rect 26330 3224 26386 3233
rect 26330 3159 26386 3168
rect 26240 2848 26292 2854
rect 26240 2790 26292 2796
rect 26252 2417 26280 2790
rect 26238 2408 26294 2417
rect 26238 2343 26294 2352
rect 26436 1873 26464 5510
rect 27066 4040 27122 4049
rect 27066 3975 27122 3984
rect 26514 3360 26570 3369
rect 26514 3295 26570 3304
rect 26422 1864 26478 1873
rect 26422 1799 26478 1808
rect 26146 504 26202 513
rect 20810 96 20866 105
rect 20810 31 20866 40
rect 20994 0 21050 480
rect 21546 0 21602 480
rect 22098 0 22154 480
rect 22650 0 22706 480
rect 23202 0 23258 480
rect 23754 0 23810 480
rect 24306 0 24362 480
rect 24858 0 24914 480
rect 25410 0 25466 480
rect 25962 0 26018 480
rect 26528 480 26556 3295
rect 27080 480 27108 3975
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 27632 480 27660 3431
rect 26146 439 26202 448
rect 26514 0 26570 480
rect 27066 0 27122 480
rect 27618 0 27674 480
<< via2 >>
rect 4250 27648 4306 27704
rect 754 27104 810 27160
rect 1306 26560 1362 26616
rect 1214 25880 1270 25936
rect 1122 24792 1178 24848
rect 938 24112 994 24168
rect 1398 20032 1454 20088
rect 1398 16496 1454 16552
rect 1582 15408 1638 15464
rect 1582 14864 1638 14920
rect 1674 14592 1730 14648
rect 1582 13776 1638 13832
rect 1582 13640 1638 13696
rect 1490 13504 1546 13560
rect 1490 12552 1546 12608
rect 1398 12300 1454 12336
rect 1398 12280 1400 12300
rect 1400 12280 1452 12300
rect 1452 12280 1454 12300
rect 1398 11464 1454 11520
rect 1398 10376 1454 10432
rect 570 8508 572 8528
rect 572 8508 624 8528
rect 624 8508 626 8528
rect 570 8472 626 8508
rect 2870 25336 2926 25392
rect 2226 24112 2282 24168
rect 2134 23976 2190 24032
rect 2502 24692 2504 24712
rect 2504 24692 2556 24712
rect 2556 24692 2558 24712
rect 2502 24656 2558 24692
rect 2410 24404 2466 24440
rect 2410 24384 2412 24404
rect 2412 24384 2464 24404
rect 2464 24384 2466 24404
rect 2410 23316 2466 23352
rect 2410 23296 2412 23316
rect 2412 23296 2464 23316
rect 2464 23296 2466 23316
rect 2410 23160 2466 23216
rect 2318 21936 2374 21992
rect 2410 21664 2466 21720
rect 2502 21528 2558 21584
rect 2318 20576 2374 20632
rect 2410 20304 2466 20360
rect 1950 17856 2006 17912
rect 2134 19252 2136 19272
rect 2136 19252 2188 19272
rect 2188 19252 2190 19272
rect 2134 19216 2190 19252
rect 1858 15428 1914 15464
rect 1858 15408 1860 15428
rect 1860 15408 1912 15428
rect 1912 15408 1914 15428
rect 1766 11328 1822 11384
rect 2042 15000 2098 15056
rect 2226 15308 2228 15328
rect 2228 15308 2280 15328
rect 2280 15308 2282 15328
rect 2226 15272 2282 15308
rect 2410 19352 2466 19408
rect 2686 20712 2742 20768
rect 2410 16088 2466 16144
rect 2870 20032 2926 20088
rect 3146 24792 3202 24848
rect 3422 23180 3478 23216
rect 3422 23160 3424 23180
rect 3424 23160 3476 23180
rect 3476 23160 3478 23180
rect 3330 23024 3386 23080
rect 3330 22344 3386 22400
rect 3238 21256 3294 21312
rect 3146 19760 3202 19816
rect 3054 19252 3056 19272
rect 3056 19252 3108 19272
rect 3108 19252 3110 19272
rect 3054 19216 3110 19252
rect 2962 18944 3018 19000
rect 3146 17856 3202 17912
rect 2778 17720 2834 17776
rect 3054 17040 3110 17096
rect 2962 16904 3018 16960
rect 2410 14612 2466 14648
rect 2410 14592 2412 14612
rect 2412 14592 2464 14612
rect 2464 14592 2466 14612
rect 2042 13912 2098 13968
rect 2042 13776 2098 13832
rect 2042 12980 2098 13016
rect 2042 12960 2044 12980
rect 2044 12960 2096 12980
rect 2096 12960 2098 12980
rect 2410 12588 2412 12608
rect 2412 12588 2464 12608
rect 2464 12588 2466 12608
rect 2410 12552 2466 12588
rect 2962 15000 3018 15056
rect 2870 14492 2872 14512
rect 2872 14492 2924 14512
rect 2924 14492 2926 14512
rect 2870 14456 2926 14492
rect 3054 13640 3110 13696
rect 2226 11600 2282 11656
rect 1766 10376 1822 10432
rect 1766 8880 1822 8936
rect 1582 7792 1638 7848
rect 1398 6976 1454 7032
rect 1674 7248 1730 7304
rect 754 4392 810 4448
rect 2042 9968 2098 10024
rect 2410 10240 2466 10296
rect 3790 24792 3846 24848
rect 3790 23704 3846 23760
rect 3698 23160 3754 23216
rect 3606 23044 3662 23080
rect 3606 23024 3608 23044
rect 3608 23024 3660 23044
rect 3660 23024 3662 23044
rect 3514 22208 3570 22264
rect 3514 21256 3570 21312
rect 3606 20440 3662 20496
rect 3882 23432 3938 23488
rect 3882 22480 3938 22536
rect 23846 27648 23902 27704
rect 4250 22616 4306 22672
rect 3974 21800 4030 21856
rect 4710 26152 4766 26208
rect 4250 20576 4306 20632
rect 4342 20168 4398 20224
rect 4066 19916 4122 19952
rect 4066 19896 4068 19916
rect 4068 19896 4120 19916
rect 4120 19896 4122 19916
rect 3882 18828 3938 18864
rect 3882 18808 3884 18828
rect 3884 18808 3936 18828
rect 3936 18808 3938 18828
rect 3882 17992 3938 18048
rect 3882 16768 3938 16824
rect 3606 15852 3608 15872
rect 3608 15852 3660 15872
rect 3660 15852 3662 15872
rect 3606 15816 3662 15852
rect 4250 17176 4306 17232
rect 4066 16632 4122 16688
rect 2870 12144 2926 12200
rect 2778 12008 2834 12064
rect 2594 10920 2650 10976
rect 2778 10240 2834 10296
rect 2778 9968 2834 10024
rect 2318 9696 2374 9752
rect 1950 9424 2006 9480
rect 1858 8336 1914 8392
rect 2042 6704 2098 6760
rect 2226 7384 2282 7440
rect 2502 9444 2558 9480
rect 2502 9424 2504 9444
rect 2504 9424 2556 9444
rect 2556 9424 2558 9444
rect 2778 9424 2834 9480
rect 2410 8084 2466 8120
rect 2410 8064 2412 8084
rect 2412 8064 2464 8084
rect 2464 8064 2466 8084
rect 2410 7268 2466 7304
rect 2410 7248 2412 7268
rect 2412 7248 2464 7268
rect 2464 7248 2466 7268
rect 2686 8880 2742 8936
rect 3054 9968 3110 10024
rect 3238 9560 3294 9616
rect 3790 13368 3846 13424
rect 4158 13096 4214 13152
rect 3974 12844 4030 12880
rect 3974 12824 3976 12844
rect 3976 12824 4028 12844
rect 4028 12824 4030 12844
rect 3882 12724 3884 12744
rect 3884 12724 3936 12744
rect 3936 12724 3938 12744
rect 3882 12688 3938 12724
rect 3974 12416 4030 12472
rect 4342 15272 4398 15328
rect 4158 12164 4214 12200
rect 4158 12144 4160 12164
rect 4160 12144 4212 12164
rect 4212 12144 4214 12164
rect 3790 11872 3846 11928
rect 3146 9016 3202 9072
rect 3606 9424 3662 9480
rect 3330 8492 3386 8528
rect 3330 8472 3332 8492
rect 3332 8472 3384 8492
rect 3384 8472 3386 8492
rect 3146 7540 3202 7576
rect 3146 7520 3148 7540
rect 3148 7520 3200 7540
rect 3200 7520 3202 7540
rect 1490 5752 1546 5808
rect 1950 5072 2006 5128
rect 1582 4548 1638 4584
rect 1582 4528 1584 4548
rect 1584 4528 1636 4548
rect 1636 4528 1638 4548
rect 1582 3984 1638 4040
rect 1490 3712 1546 3768
rect 662 3440 718 3496
rect 202 1672 258 1728
rect 1766 3712 1822 3768
rect 1398 3032 1454 3088
rect 1950 2896 2006 2952
rect 1214 2760 1270 2816
rect 1582 2080 1638 2136
rect 1950 1672 2006 1728
rect 2318 5888 2374 5944
rect 2318 5772 2374 5808
rect 2318 5752 2320 5772
rect 2320 5752 2372 5772
rect 2372 5752 2374 5772
rect 2870 6704 2926 6760
rect 2686 5752 2742 5808
rect 2594 5616 2650 5672
rect 2410 3168 2466 3224
rect 2226 584 2282 640
rect 2870 3168 2926 3224
rect 3882 11328 3938 11384
rect 3882 10648 3938 10704
rect 4066 10920 4122 10976
rect 3606 6024 3662 6080
rect 3146 1536 3202 1592
rect 3698 5616 3754 5672
rect 4250 10784 4306 10840
rect 4526 21664 4582 21720
rect 4618 19352 4674 19408
rect 4894 22752 4950 22808
rect 4802 17584 4858 17640
rect 4710 17176 4766 17232
rect 4710 14900 4712 14920
rect 4712 14900 4764 14920
rect 4764 14900 4766 14920
rect 4710 14864 4766 14900
rect 4434 12144 4490 12200
rect 4434 11348 4490 11384
rect 4434 11328 4436 11348
rect 4436 11328 4488 11348
rect 4488 11328 4490 11348
rect 4710 12144 4766 12200
rect 5170 23976 5226 24032
rect 5078 23296 5134 23352
rect 5622 25050 5678 25052
rect 5702 25050 5758 25052
rect 5782 25050 5838 25052
rect 5862 25050 5918 25052
rect 5622 24998 5648 25050
rect 5648 24998 5678 25050
rect 5702 24998 5712 25050
rect 5712 24998 5758 25050
rect 5782 24998 5828 25050
rect 5828 24998 5838 25050
rect 5862 24998 5892 25050
rect 5892 24998 5918 25050
rect 5622 24996 5678 24998
rect 5702 24996 5758 24998
rect 5782 24996 5838 24998
rect 5862 24996 5918 24998
rect 5998 24384 6054 24440
rect 5538 24248 5594 24304
rect 5906 24148 5908 24168
rect 5908 24148 5960 24168
rect 5960 24148 5962 24168
rect 5906 24112 5962 24148
rect 5622 23962 5678 23964
rect 5702 23962 5758 23964
rect 5782 23962 5838 23964
rect 5862 23962 5918 23964
rect 5622 23910 5648 23962
rect 5648 23910 5678 23962
rect 5702 23910 5712 23962
rect 5712 23910 5758 23962
rect 5782 23910 5828 23962
rect 5828 23910 5838 23962
rect 5862 23910 5892 23962
rect 5892 23910 5918 23962
rect 5622 23908 5678 23910
rect 5702 23908 5758 23910
rect 5782 23908 5838 23910
rect 5862 23908 5918 23910
rect 6090 23840 6146 23896
rect 5538 23160 5594 23216
rect 5622 22874 5678 22876
rect 5702 22874 5758 22876
rect 5782 22874 5838 22876
rect 5862 22874 5918 22876
rect 5622 22822 5648 22874
rect 5648 22822 5678 22874
rect 5702 22822 5712 22874
rect 5712 22822 5758 22874
rect 5782 22822 5828 22874
rect 5828 22822 5838 22874
rect 5862 22822 5892 22874
rect 5892 22822 5918 22874
rect 5622 22820 5678 22822
rect 5702 22820 5758 22822
rect 5782 22820 5838 22822
rect 5862 22820 5918 22822
rect 5262 22208 5318 22264
rect 5622 21786 5678 21788
rect 5702 21786 5758 21788
rect 5782 21786 5838 21788
rect 5862 21786 5918 21788
rect 5622 21734 5648 21786
rect 5648 21734 5678 21786
rect 5702 21734 5712 21786
rect 5712 21734 5758 21786
rect 5782 21734 5828 21786
rect 5828 21734 5838 21786
rect 5862 21734 5892 21786
rect 5892 21734 5918 21786
rect 5622 21732 5678 21734
rect 5702 21732 5758 21734
rect 5782 21732 5838 21734
rect 5862 21732 5918 21734
rect 5170 21528 5226 21584
rect 5262 20712 5318 20768
rect 5078 17856 5134 17912
rect 5078 17176 5134 17232
rect 4986 16088 5042 16144
rect 4986 15680 5042 15736
rect 4894 14728 4950 14784
rect 4894 13912 4950 13968
rect 5170 17040 5226 17096
rect 5622 20698 5678 20700
rect 5702 20698 5758 20700
rect 5782 20698 5838 20700
rect 5862 20698 5918 20700
rect 5622 20646 5648 20698
rect 5648 20646 5678 20698
rect 5702 20646 5712 20698
rect 5712 20646 5758 20698
rect 5782 20646 5828 20698
rect 5828 20646 5838 20698
rect 5862 20646 5892 20698
rect 5892 20646 5918 20698
rect 5622 20644 5678 20646
rect 5702 20644 5758 20646
rect 5782 20644 5838 20646
rect 5862 20644 5918 20646
rect 5722 20340 5724 20360
rect 5724 20340 5776 20360
rect 5776 20340 5778 20360
rect 5722 20304 5778 20340
rect 5622 19610 5678 19612
rect 5702 19610 5758 19612
rect 5782 19610 5838 19612
rect 5862 19610 5918 19612
rect 5622 19558 5648 19610
rect 5648 19558 5678 19610
rect 5702 19558 5712 19610
rect 5712 19558 5758 19610
rect 5782 19558 5828 19610
rect 5828 19558 5838 19610
rect 5862 19558 5892 19610
rect 5892 19558 5918 19610
rect 5622 19556 5678 19558
rect 5702 19556 5758 19558
rect 5782 19556 5838 19558
rect 5862 19556 5918 19558
rect 5622 18522 5678 18524
rect 5702 18522 5758 18524
rect 5782 18522 5838 18524
rect 5862 18522 5918 18524
rect 5622 18470 5648 18522
rect 5648 18470 5678 18522
rect 5702 18470 5712 18522
rect 5712 18470 5758 18522
rect 5782 18470 5828 18522
rect 5828 18470 5838 18522
rect 5862 18470 5892 18522
rect 5892 18470 5918 18522
rect 5622 18468 5678 18470
rect 5702 18468 5758 18470
rect 5782 18468 5838 18470
rect 5862 18468 5918 18470
rect 5538 18148 5594 18184
rect 5538 18128 5540 18148
rect 5540 18128 5592 18148
rect 5592 18128 5594 18148
rect 5262 16632 5318 16688
rect 4986 13776 5042 13832
rect 5630 17720 5686 17776
rect 5622 17434 5678 17436
rect 5702 17434 5758 17436
rect 5782 17434 5838 17436
rect 5862 17434 5918 17436
rect 5622 17382 5648 17434
rect 5648 17382 5678 17434
rect 5702 17382 5712 17434
rect 5712 17382 5758 17434
rect 5782 17382 5828 17434
rect 5828 17382 5838 17434
rect 5862 17382 5892 17434
rect 5892 17382 5918 17434
rect 5622 17380 5678 17382
rect 5702 17380 5758 17382
rect 5782 17380 5838 17382
rect 5862 17380 5918 17382
rect 5630 17176 5686 17232
rect 5622 16346 5678 16348
rect 5702 16346 5758 16348
rect 5782 16346 5838 16348
rect 5862 16346 5918 16348
rect 5622 16294 5648 16346
rect 5648 16294 5678 16346
rect 5702 16294 5712 16346
rect 5712 16294 5758 16346
rect 5782 16294 5828 16346
rect 5828 16294 5838 16346
rect 5862 16294 5892 16346
rect 5892 16294 5918 16346
rect 5622 16292 5678 16294
rect 5702 16292 5758 16294
rect 5782 16292 5838 16294
rect 5862 16292 5918 16294
rect 5630 16124 5632 16144
rect 5632 16124 5684 16144
rect 5684 16124 5686 16144
rect 5630 16088 5686 16124
rect 5538 15544 5594 15600
rect 5446 15408 5502 15464
rect 5446 15272 5502 15328
rect 5622 15258 5678 15260
rect 5702 15258 5758 15260
rect 5782 15258 5838 15260
rect 5862 15258 5918 15260
rect 5622 15206 5648 15258
rect 5648 15206 5678 15258
rect 5702 15206 5712 15258
rect 5712 15206 5758 15258
rect 5782 15206 5828 15258
rect 5828 15206 5838 15258
rect 5862 15206 5892 15258
rect 5892 15206 5918 15258
rect 5622 15204 5678 15206
rect 5702 15204 5758 15206
rect 5782 15204 5838 15206
rect 5862 15204 5918 15206
rect 5446 14728 5502 14784
rect 4894 12960 4950 13016
rect 4618 9696 4674 9752
rect 4802 10104 4858 10160
rect 4066 8336 4122 8392
rect 4342 7928 4398 7984
rect 4342 6976 4398 7032
rect 4526 6976 4582 7032
rect 3974 6840 4030 6896
rect 4710 7148 4712 7168
rect 4712 7148 4764 7168
rect 4764 7148 4766 7168
rect 4710 7112 4766 7148
rect 4066 5616 4122 5672
rect 4066 4120 4122 4176
rect 4710 5108 4712 5128
rect 4712 5108 4764 5128
rect 4764 5108 4766 5128
rect 4710 5072 4766 5108
rect 4986 9424 5042 9480
rect 5262 13232 5318 13288
rect 5446 13640 5502 13696
rect 5170 12008 5226 12064
rect 5170 11192 5226 11248
rect 4894 8880 4950 8936
rect 5622 14170 5678 14172
rect 5702 14170 5758 14172
rect 5782 14170 5838 14172
rect 5862 14170 5918 14172
rect 5622 14118 5648 14170
rect 5648 14118 5678 14170
rect 5702 14118 5712 14170
rect 5712 14118 5758 14170
rect 5782 14118 5828 14170
rect 5828 14118 5838 14170
rect 5862 14118 5892 14170
rect 5892 14118 5918 14170
rect 5622 14116 5678 14118
rect 5702 14116 5758 14118
rect 5782 14116 5838 14118
rect 5862 14116 5918 14118
rect 5622 13082 5678 13084
rect 5702 13082 5758 13084
rect 5782 13082 5838 13084
rect 5862 13082 5918 13084
rect 5622 13030 5648 13082
rect 5648 13030 5678 13082
rect 5702 13030 5712 13082
rect 5712 13030 5758 13082
rect 5782 13030 5828 13082
rect 5828 13030 5838 13082
rect 5862 13030 5892 13082
rect 5892 13030 5918 13082
rect 5622 13028 5678 13030
rect 5702 13028 5758 13030
rect 5782 13028 5838 13030
rect 5862 13028 5918 13030
rect 5446 11192 5502 11248
rect 5262 9152 5318 9208
rect 5262 8780 5264 8800
rect 5264 8780 5316 8800
rect 5316 8780 5318 8800
rect 5262 8744 5318 8780
rect 5170 6160 5226 6216
rect 5354 6160 5410 6216
rect 4526 3596 4582 3632
rect 4526 3576 4528 3596
rect 4528 3576 4580 3596
rect 4580 3576 4582 3596
rect 3698 856 3754 912
rect 3606 448 3662 504
rect 4986 3440 5042 3496
rect 5170 3168 5226 3224
rect 4066 2796 4068 2816
rect 4068 2796 4120 2816
rect 4120 2796 4122 2816
rect 4066 2760 4122 2796
rect 4802 2644 4858 2680
rect 4802 2624 4804 2644
rect 4804 2624 4856 2644
rect 4856 2624 4858 2644
rect 5622 11994 5678 11996
rect 5702 11994 5758 11996
rect 5782 11994 5838 11996
rect 5862 11994 5918 11996
rect 5622 11942 5648 11994
rect 5648 11942 5678 11994
rect 5702 11942 5712 11994
rect 5712 11942 5758 11994
rect 5782 11942 5828 11994
rect 5828 11942 5838 11994
rect 5862 11942 5892 11994
rect 5892 11942 5918 11994
rect 5622 11940 5678 11942
rect 5702 11940 5758 11942
rect 5782 11940 5838 11942
rect 5862 11940 5918 11942
rect 5622 10906 5678 10908
rect 5702 10906 5758 10908
rect 5782 10906 5838 10908
rect 5862 10906 5918 10908
rect 5622 10854 5648 10906
rect 5648 10854 5678 10906
rect 5702 10854 5712 10906
rect 5712 10854 5758 10906
rect 5782 10854 5828 10906
rect 5828 10854 5838 10906
rect 5862 10854 5892 10906
rect 5892 10854 5918 10906
rect 5622 10852 5678 10854
rect 5702 10852 5758 10854
rect 5782 10852 5838 10854
rect 5862 10852 5918 10854
rect 5814 10512 5870 10568
rect 5906 10376 5962 10432
rect 5622 9818 5678 9820
rect 5702 9818 5758 9820
rect 5782 9818 5838 9820
rect 5862 9818 5918 9820
rect 5622 9766 5648 9818
rect 5648 9766 5678 9818
rect 5702 9766 5712 9818
rect 5712 9766 5758 9818
rect 5782 9766 5828 9818
rect 5828 9766 5838 9818
rect 5862 9766 5892 9818
rect 5892 9766 5918 9818
rect 5622 9764 5678 9766
rect 5702 9764 5758 9766
rect 5782 9764 5838 9766
rect 5862 9764 5918 9766
rect 5622 8730 5678 8732
rect 5702 8730 5758 8732
rect 5782 8730 5838 8732
rect 5862 8730 5918 8732
rect 5622 8678 5648 8730
rect 5648 8678 5678 8730
rect 5702 8678 5712 8730
rect 5712 8678 5758 8730
rect 5782 8678 5828 8730
rect 5828 8678 5838 8730
rect 5862 8678 5892 8730
rect 5892 8678 5918 8730
rect 5622 8676 5678 8678
rect 5702 8676 5758 8678
rect 5782 8676 5838 8678
rect 5862 8676 5918 8678
rect 5622 7642 5678 7644
rect 5702 7642 5758 7644
rect 5782 7642 5838 7644
rect 5862 7642 5918 7644
rect 5622 7590 5648 7642
rect 5648 7590 5678 7642
rect 5702 7590 5712 7642
rect 5712 7590 5758 7642
rect 5782 7590 5828 7642
rect 5828 7590 5838 7642
rect 5862 7590 5892 7642
rect 5892 7590 5918 7642
rect 5622 7588 5678 7590
rect 5702 7588 5758 7590
rect 5782 7588 5838 7590
rect 5862 7588 5918 7590
rect 5814 6860 5870 6896
rect 5814 6840 5816 6860
rect 5816 6840 5868 6860
rect 5868 6840 5870 6860
rect 5630 6724 5686 6760
rect 5630 6704 5632 6724
rect 5632 6704 5684 6724
rect 5684 6704 5686 6724
rect 5622 6554 5678 6556
rect 5702 6554 5758 6556
rect 5782 6554 5838 6556
rect 5862 6554 5918 6556
rect 5622 6502 5648 6554
rect 5648 6502 5678 6554
rect 5702 6502 5712 6554
rect 5712 6502 5758 6554
rect 5782 6502 5828 6554
rect 5828 6502 5838 6554
rect 5862 6502 5892 6554
rect 5892 6502 5918 6554
rect 5622 6500 5678 6502
rect 5702 6500 5758 6502
rect 5782 6500 5838 6502
rect 5862 6500 5918 6502
rect 6458 25064 6514 25120
rect 6366 22480 6422 22536
rect 6366 22092 6422 22128
rect 6366 22072 6368 22092
rect 6368 22072 6420 22092
rect 6420 22072 6422 22092
rect 6734 24112 6790 24168
rect 6550 20712 6606 20768
rect 6366 20032 6422 20088
rect 6642 18808 6698 18864
rect 6458 17484 6460 17504
rect 6460 17484 6512 17504
rect 6512 17484 6514 17504
rect 6458 17448 6514 17484
rect 6550 17312 6606 17368
rect 6458 16768 6514 16824
rect 6274 15272 6330 15328
rect 6274 14612 6330 14648
rect 6274 14592 6276 14612
rect 6276 14592 6328 14612
rect 6328 14592 6330 14612
rect 6550 16360 6606 16416
rect 7378 25336 7434 25392
rect 7286 24792 7342 24848
rect 7286 24656 7342 24712
rect 7010 23468 7012 23488
rect 7012 23468 7064 23488
rect 7064 23468 7066 23488
rect 7010 23432 7066 23468
rect 6918 20848 6974 20904
rect 6826 20576 6882 20632
rect 6826 20460 6882 20496
rect 6826 20440 6828 20460
rect 6828 20440 6880 20460
rect 6880 20440 6882 20460
rect 7194 22072 7250 22128
rect 7102 20440 7158 20496
rect 7194 20032 7250 20088
rect 7010 18672 7066 18728
rect 7102 18400 7158 18456
rect 6918 17176 6974 17232
rect 7010 15952 7066 16008
rect 6182 12688 6238 12744
rect 6734 14728 6790 14784
rect 6918 14728 6974 14784
rect 7010 14340 7066 14376
rect 7010 14320 7012 14340
rect 7012 14320 7064 14340
rect 7064 14320 7066 14340
rect 6366 12824 6422 12880
rect 7470 23724 7526 23760
rect 7470 23704 7472 23724
rect 7472 23704 7524 23724
rect 7524 23704 7526 23724
rect 7654 21684 7710 21720
rect 7654 21664 7656 21684
rect 7656 21664 7708 21684
rect 7708 21664 7710 21684
rect 7654 20884 7656 20904
rect 7656 20884 7708 20904
rect 7708 20884 7710 20904
rect 7654 20848 7710 20884
rect 7470 19760 7526 19816
rect 7746 18808 7802 18864
rect 7470 18672 7526 18728
rect 7470 18028 7472 18048
rect 7472 18028 7524 18048
rect 7524 18028 7526 18048
rect 7470 17992 7526 18028
rect 7470 15408 7526 15464
rect 6458 11600 6514 11656
rect 6458 11192 6514 11248
rect 6274 10784 6330 10840
rect 5622 5466 5678 5468
rect 5702 5466 5758 5468
rect 5782 5466 5838 5468
rect 5862 5466 5918 5468
rect 5622 5414 5648 5466
rect 5648 5414 5678 5466
rect 5702 5414 5712 5466
rect 5712 5414 5758 5466
rect 5782 5414 5828 5466
rect 5828 5414 5838 5466
rect 5862 5414 5892 5466
rect 5892 5414 5918 5466
rect 5622 5412 5678 5414
rect 5702 5412 5758 5414
rect 5782 5412 5838 5414
rect 5862 5412 5918 5414
rect 6090 4800 6146 4856
rect 5622 4378 5678 4380
rect 5702 4378 5758 4380
rect 5782 4378 5838 4380
rect 5862 4378 5918 4380
rect 5622 4326 5648 4378
rect 5648 4326 5678 4378
rect 5702 4326 5712 4378
rect 5712 4326 5758 4378
rect 5782 4326 5828 4378
rect 5828 4326 5838 4378
rect 5862 4326 5892 4378
rect 5892 4326 5918 4378
rect 5622 4324 5678 4326
rect 5702 4324 5758 4326
rect 5782 4324 5838 4326
rect 5862 4324 5918 4326
rect 5622 3290 5678 3292
rect 5702 3290 5758 3292
rect 5782 3290 5838 3292
rect 5862 3290 5918 3292
rect 5622 3238 5648 3290
rect 5648 3238 5678 3290
rect 5702 3238 5712 3290
rect 5712 3238 5758 3290
rect 5782 3238 5828 3290
rect 5828 3238 5838 3290
rect 5862 3238 5892 3290
rect 5892 3238 5918 3290
rect 5622 3236 5678 3238
rect 5702 3236 5758 3238
rect 5782 3236 5838 3238
rect 5862 3236 5918 3238
rect 6274 8336 6330 8392
rect 6550 10124 6606 10160
rect 6550 10104 6552 10124
rect 6552 10104 6604 10124
rect 6604 10104 6606 10124
rect 6734 11600 6790 11656
rect 6826 11464 6882 11520
rect 6642 10004 6644 10024
rect 6644 10004 6696 10024
rect 6696 10004 6698 10024
rect 6642 9968 6698 10004
rect 6458 9832 6514 9888
rect 6642 9696 6698 9752
rect 6274 5908 6330 5944
rect 6274 5888 6276 5908
rect 6276 5888 6328 5908
rect 6328 5888 6330 5908
rect 6366 5072 6422 5128
rect 6366 4120 6422 4176
rect 6550 8336 6606 8392
rect 7102 12180 7104 12200
rect 7104 12180 7156 12200
rect 7156 12180 7158 12200
rect 7102 12144 7158 12180
rect 7010 10920 7066 10976
rect 6734 9560 6790 9616
rect 7286 11872 7342 11928
rect 7102 10104 7158 10160
rect 7010 9288 7066 9344
rect 6734 6296 6790 6352
rect 7194 7928 7250 7984
rect 6642 4664 6698 4720
rect 6826 4392 6882 4448
rect 6734 3304 6790 3360
rect 6274 2252 6276 2272
rect 6276 2252 6328 2272
rect 6328 2252 6330 2272
rect 6274 2216 6330 2252
rect 5622 2202 5678 2204
rect 5702 2202 5758 2204
rect 5782 2202 5838 2204
rect 5862 2202 5918 2204
rect 5622 2150 5648 2202
rect 5648 2150 5678 2202
rect 5702 2150 5712 2202
rect 5712 2150 5758 2202
rect 5782 2150 5828 2202
rect 5828 2150 5838 2202
rect 5862 2150 5892 2202
rect 5892 2150 5918 2202
rect 5622 2148 5678 2150
rect 5702 2148 5758 2150
rect 5782 2148 5838 2150
rect 5862 2148 5918 2150
rect 6550 1556 6606 1592
rect 6550 1536 6552 1556
rect 6552 1536 6604 1556
rect 6604 1536 6606 1556
rect 8022 23044 8078 23080
rect 8022 23024 8024 23044
rect 8024 23024 8076 23044
rect 8076 23024 8078 23044
rect 8482 23296 8538 23352
rect 8482 22208 8538 22264
rect 8390 21120 8446 21176
rect 8574 21664 8630 21720
rect 8574 21528 8630 21584
rect 8206 18284 8262 18320
rect 8206 18264 8208 18284
rect 8208 18264 8260 18284
rect 8260 18264 8262 18284
rect 8206 16940 8208 16960
rect 8208 16940 8260 16960
rect 8260 16940 8262 16960
rect 8206 16904 8262 16940
rect 9034 23976 9090 24032
rect 8758 22616 8814 22672
rect 9494 25916 9496 25936
rect 9496 25916 9548 25936
rect 9548 25916 9550 25936
rect 9494 25880 9550 25916
rect 9494 25780 9496 25800
rect 9496 25780 9548 25800
rect 9548 25780 9550 25800
rect 9494 25744 9550 25780
rect 9494 23568 9550 23624
rect 9494 23180 9550 23216
rect 9494 23160 9496 23180
rect 9496 23160 9548 23180
rect 9548 23160 9550 23180
rect 9678 24792 9734 24848
rect 10289 25594 10345 25596
rect 10369 25594 10425 25596
rect 10449 25594 10505 25596
rect 10529 25594 10585 25596
rect 10289 25542 10315 25594
rect 10315 25542 10345 25594
rect 10369 25542 10379 25594
rect 10379 25542 10425 25594
rect 10449 25542 10495 25594
rect 10495 25542 10505 25594
rect 10529 25542 10559 25594
rect 10559 25542 10585 25594
rect 10289 25540 10345 25542
rect 10369 25540 10425 25542
rect 10449 25540 10505 25542
rect 10529 25540 10585 25542
rect 10874 25472 10930 25528
rect 10138 24792 10194 24848
rect 9678 23296 9734 23352
rect 9678 22344 9734 22400
rect 9126 21392 9182 21448
rect 9218 20848 9274 20904
rect 8666 19624 8722 19680
rect 8850 19624 8906 19680
rect 8482 16652 8538 16688
rect 8482 16632 8484 16652
rect 8484 16632 8536 16652
rect 8536 16632 8538 16652
rect 8666 16360 8722 16416
rect 7838 15544 7894 15600
rect 8114 15700 8170 15736
rect 8114 15680 8116 15700
rect 8116 15680 8168 15700
rect 8168 15680 8170 15700
rect 8022 15428 8078 15464
rect 8022 15408 8024 15428
rect 8024 15408 8076 15428
rect 8076 15408 8078 15428
rect 7930 14592 7986 14648
rect 7746 13504 7802 13560
rect 7746 12688 7802 12744
rect 7838 12280 7894 12336
rect 7562 9696 7618 9752
rect 7746 11192 7802 11248
rect 8022 13504 8078 13560
rect 8022 12416 8078 12472
rect 7930 10920 7986 10976
rect 7838 10648 7894 10704
rect 8482 15952 8538 16008
rect 8298 13776 8354 13832
rect 8942 19488 8998 19544
rect 8850 15156 8906 15192
rect 8850 15136 8852 15156
rect 8852 15136 8904 15156
rect 8904 15136 8906 15156
rect 8666 13912 8722 13968
rect 8574 13640 8630 13696
rect 8390 12980 8446 13016
rect 8390 12960 8392 12980
rect 8392 12960 8444 12980
rect 8444 12960 8446 12980
rect 8206 12144 8262 12200
rect 8114 11328 8170 11384
rect 8114 10260 8170 10296
rect 8114 10240 8116 10260
rect 8116 10240 8168 10260
rect 8168 10240 8170 10260
rect 7470 8744 7526 8800
rect 7470 8336 7526 8392
rect 8206 8336 8262 8392
rect 7470 4936 7526 4992
rect 7746 7964 7748 7984
rect 7748 7964 7800 7984
rect 7800 7964 7802 7984
rect 7746 7928 7802 7964
rect 8758 13368 8814 13424
rect 9218 16632 9274 16688
rect 9218 14184 9274 14240
rect 8850 12280 8906 12336
rect 8850 12008 8906 12064
rect 8758 11600 8814 11656
rect 9218 12588 9220 12608
rect 9220 12588 9272 12608
rect 9272 12588 9274 12608
rect 9218 12552 9274 12588
rect 8850 10512 8906 10568
rect 8482 8608 8538 8664
rect 7654 7540 7710 7576
rect 7654 7520 7656 7540
rect 7656 7520 7708 7540
rect 7708 7520 7710 7540
rect 8114 6704 8170 6760
rect 8022 6432 8078 6488
rect 8390 6296 8446 6352
rect 8206 5752 8262 5808
rect 8206 5480 8262 5536
rect 8114 5092 8170 5128
rect 8114 5072 8116 5092
rect 8116 5072 8168 5092
rect 8168 5072 8170 5092
rect 7838 3460 7894 3496
rect 7838 3440 7840 3460
rect 7840 3440 7892 3460
rect 7892 3440 7894 3460
rect 6918 1536 6974 1592
rect 8666 8472 8722 8528
rect 8666 6840 8722 6896
rect 8850 8472 8906 8528
rect 8574 4820 8630 4856
rect 8574 4800 8576 4820
rect 8576 4800 8628 4820
rect 8628 4800 8630 4820
rect 8574 4120 8630 4176
rect 8390 3168 8446 3224
rect 8390 2896 8446 2952
rect 6918 312 6974 368
rect 8022 448 8078 504
rect 8942 3712 8998 3768
rect 8666 2932 8668 2952
rect 8668 2932 8720 2952
rect 8720 2932 8722 2952
rect 8666 2896 8722 2932
rect 10289 24506 10345 24508
rect 10369 24506 10425 24508
rect 10449 24506 10505 24508
rect 10529 24506 10585 24508
rect 10289 24454 10315 24506
rect 10315 24454 10345 24506
rect 10369 24454 10379 24506
rect 10379 24454 10425 24506
rect 10449 24454 10495 24506
rect 10495 24454 10505 24506
rect 10529 24454 10559 24506
rect 10559 24454 10585 24506
rect 10289 24452 10345 24454
rect 10369 24452 10425 24454
rect 10449 24452 10505 24454
rect 10529 24452 10585 24454
rect 10598 23976 10654 24032
rect 10874 25064 10930 25120
rect 11610 24656 11666 24712
rect 11058 24248 11114 24304
rect 10690 23840 10746 23896
rect 10289 23418 10345 23420
rect 10369 23418 10425 23420
rect 10449 23418 10505 23420
rect 10529 23418 10585 23420
rect 10289 23366 10315 23418
rect 10315 23366 10345 23418
rect 10369 23366 10379 23418
rect 10379 23366 10425 23418
rect 10449 23366 10495 23418
rect 10495 23366 10505 23418
rect 10529 23366 10559 23418
rect 10559 23366 10585 23418
rect 10289 23364 10345 23366
rect 10369 23364 10425 23366
rect 10449 23364 10505 23366
rect 10529 23364 10585 23366
rect 10289 22330 10345 22332
rect 10369 22330 10425 22332
rect 10449 22330 10505 22332
rect 10529 22330 10585 22332
rect 10289 22278 10315 22330
rect 10315 22278 10345 22330
rect 10369 22278 10379 22330
rect 10379 22278 10425 22330
rect 10449 22278 10495 22330
rect 10495 22278 10505 22330
rect 10529 22278 10559 22330
rect 10559 22278 10585 22330
rect 10289 22276 10345 22278
rect 10369 22276 10425 22278
rect 10449 22276 10505 22278
rect 10529 22276 10585 22278
rect 10874 23704 10930 23760
rect 9862 21936 9918 21992
rect 9678 21256 9734 21312
rect 9678 20168 9734 20224
rect 9494 17584 9550 17640
rect 9402 16496 9458 16552
rect 9678 17856 9734 17912
rect 9862 19352 9918 19408
rect 10289 21242 10345 21244
rect 10369 21242 10425 21244
rect 10449 21242 10505 21244
rect 10529 21242 10585 21244
rect 10289 21190 10315 21242
rect 10315 21190 10345 21242
rect 10369 21190 10379 21242
rect 10379 21190 10425 21242
rect 10449 21190 10495 21242
rect 10495 21190 10505 21242
rect 10529 21190 10559 21242
rect 10559 21190 10585 21242
rect 10289 21188 10345 21190
rect 10369 21188 10425 21190
rect 10449 21188 10505 21190
rect 10529 21188 10585 21190
rect 10138 21120 10194 21176
rect 11242 23568 11298 23624
rect 11150 23160 11206 23216
rect 11058 22752 11114 22808
rect 11150 22072 11206 22128
rect 11058 20984 11114 21040
rect 10289 20154 10345 20156
rect 10369 20154 10425 20156
rect 10449 20154 10505 20156
rect 10529 20154 10585 20156
rect 10289 20102 10315 20154
rect 10315 20102 10345 20154
rect 10369 20102 10379 20154
rect 10379 20102 10425 20154
rect 10449 20102 10495 20154
rect 10495 20102 10505 20154
rect 10529 20102 10559 20154
rect 10559 20102 10585 20154
rect 10289 20100 10345 20102
rect 10369 20100 10425 20102
rect 10449 20100 10505 20102
rect 10529 20100 10585 20102
rect 10322 19760 10378 19816
rect 10230 19352 10286 19408
rect 10322 19216 10378 19272
rect 10289 19066 10345 19068
rect 10369 19066 10425 19068
rect 10449 19066 10505 19068
rect 10529 19066 10585 19068
rect 10289 19014 10315 19066
rect 10315 19014 10345 19066
rect 10369 19014 10379 19066
rect 10379 19014 10425 19066
rect 10449 19014 10495 19066
rect 10495 19014 10505 19066
rect 10529 19014 10559 19066
rect 10559 19014 10585 19066
rect 10289 19012 10345 19014
rect 10369 19012 10425 19014
rect 10449 19012 10505 19014
rect 10529 19012 10585 19014
rect 9954 18264 10010 18320
rect 9586 16496 9642 16552
rect 9586 15816 9642 15872
rect 9678 15680 9734 15736
rect 9678 14728 9734 14784
rect 9310 10376 9366 10432
rect 9770 14048 9826 14104
rect 9770 13640 9826 13696
rect 9770 12824 9826 12880
rect 10289 17978 10345 17980
rect 10369 17978 10425 17980
rect 10449 17978 10505 17980
rect 10529 17978 10585 17980
rect 10289 17926 10315 17978
rect 10315 17926 10345 17978
rect 10369 17926 10379 17978
rect 10379 17926 10425 17978
rect 10449 17926 10495 17978
rect 10495 17926 10505 17978
rect 10529 17926 10559 17978
rect 10559 17926 10585 17978
rect 10289 17924 10345 17926
rect 10369 17924 10425 17926
rect 10449 17924 10505 17926
rect 10529 17924 10585 17926
rect 10289 16890 10345 16892
rect 10369 16890 10425 16892
rect 10449 16890 10505 16892
rect 10529 16890 10585 16892
rect 10289 16838 10315 16890
rect 10315 16838 10345 16890
rect 10369 16838 10379 16890
rect 10379 16838 10425 16890
rect 10449 16838 10495 16890
rect 10495 16838 10505 16890
rect 10529 16838 10559 16890
rect 10559 16838 10585 16890
rect 10289 16836 10345 16838
rect 10369 16836 10425 16838
rect 10449 16836 10505 16838
rect 10529 16836 10585 16838
rect 10874 20168 10930 20224
rect 11518 24148 11520 24168
rect 11520 24148 11572 24168
rect 11572 24148 11574 24168
rect 11518 24112 11574 24148
rect 11518 23704 11574 23760
rect 11426 23024 11482 23080
rect 11610 20884 11612 20904
rect 11612 20884 11664 20904
rect 11664 20884 11666 20904
rect 11610 20848 11666 20884
rect 10874 17992 10930 18048
rect 10289 15802 10345 15804
rect 10369 15802 10425 15804
rect 10449 15802 10505 15804
rect 10529 15802 10585 15804
rect 10289 15750 10315 15802
rect 10315 15750 10345 15802
rect 10369 15750 10379 15802
rect 10379 15750 10425 15802
rect 10449 15750 10495 15802
rect 10495 15750 10505 15802
rect 10529 15750 10559 15802
rect 10559 15750 10585 15802
rect 10289 15748 10345 15750
rect 10369 15748 10425 15750
rect 10449 15748 10505 15750
rect 10529 15748 10585 15750
rect 9954 13776 10010 13832
rect 9954 13524 10010 13560
rect 9954 13504 9956 13524
rect 9956 13504 10008 13524
rect 10008 13504 10010 13524
rect 9954 13096 10010 13152
rect 10506 15308 10508 15328
rect 10508 15308 10560 15328
rect 10560 15308 10562 15328
rect 10506 15272 10562 15308
rect 10289 14714 10345 14716
rect 10369 14714 10425 14716
rect 10449 14714 10505 14716
rect 10529 14714 10585 14716
rect 10289 14662 10315 14714
rect 10315 14662 10345 14714
rect 10369 14662 10379 14714
rect 10379 14662 10425 14714
rect 10449 14662 10495 14714
rect 10495 14662 10505 14714
rect 10529 14662 10559 14714
rect 10559 14662 10585 14714
rect 10289 14660 10345 14662
rect 10369 14660 10425 14662
rect 10449 14660 10505 14662
rect 10529 14660 10585 14662
rect 10289 13626 10345 13628
rect 10369 13626 10425 13628
rect 10449 13626 10505 13628
rect 10529 13626 10585 13628
rect 10289 13574 10315 13626
rect 10315 13574 10345 13626
rect 10369 13574 10379 13626
rect 10379 13574 10425 13626
rect 10449 13574 10495 13626
rect 10495 13574 10505 13626
rect 10529 13574 10559 13626
rect 10559 13574 10585 13626
rect 10289 13572 10345 13574
rect 10369 13572 10425 13574
rect 10449 13572 10505 13574
rect 10529 13572 10585 13574
rect 10138 13232 10194 13288
rect 9862 12688 9918 12744
rect 9402 9560 9458 9616
rect 9402 9444 9458 9480
rect 9402 9424 9404 9444
rect 9404 9424 9456 9444
rect 9456 9424 9458 9444
rect 9218 9152 9274 9208
rect 9126 5344 9182 5400
rect 9310 5108 9312 5128
rect 9312 5108 9364 5128
rect 9364 5108 9366 5128
rect 9310 5072 9366 5108
rect 9402 4664 9458 4720
rect 9310 2216 9366 2272
rect 9034 1536 9090 1592
rect 9218 1556 9274 1592
rect 9218 1536 9220 1556
rect 9220 1536 9272 1556
rect 9272 1536 9274 1556
rect 9678 10512 9734 10568
rect 9586 9560 9642 9616
rect 9678 3984 9734 4040
rect 9954 9968 10010 10024
rect 9954 4700 9956 4720
rect 9956 4700 10008 4720
rect 10008 4700 10010 4720
rect 9954 4664 10010 4700
rect 9402 1400 9458 1456
rect 9586 1264 9642 1320
rect 9770 3440 9826 3496
rect 9954 3304 10010 3360
rect 10322 13232 10378 13288
rect 10322 12688 10378 12744
rect 10506 12724 10508 12744
rect 10508 12724 10560 12744
rect 10560 12724 10562 12744
rect 10506 12688 10562 12724
rect 10289 12538 10345 12540
rect 10369 12538 10425 12540
rect 10449 12538 10505 12540
rect 10529 12538 10585 12540
rect 10289 12486 10315 12538
rect 10315 12486 10345 12538
rect 10369 12486 10379 12538
rect 10379 12486 10425 12538
rect 10449 12486 10495 12538
rect 10495 12486 10505 12538
rect 10529 12486 10559 12538
rect 10559 12486 10585 12538
rect 10289 12484 10345 12486
rect 10369 12484 10425 12486
rect 10449 12484 10505 12486
rect 10529 12484 10585 12486
rect 10289 11450 10345 11452
rect 10369 11450 10425 11452
rect 10449 11450 10505 11452
rect 10529 11450 10585 11452
rect 10289 11398 10315 11450
rect 10315 11398 10345 11450
rect 10369 11398 10379 11450
rect 10379 11398 10425 11450
rect 10449 11398 10495 11450
rect 10495 11398 10505 11450
rect 10529 11398 10559 11450
rect 10559 11398 10585 11450
rect 10289 11396 10345 11398
rect 10369 11396 10425 11398
rect 10449 11396 10505 11398
rect 10529 11396 10585 11398
rect 10506 11076 10562 11112
rect 10506 11056 10508 11076
rect 10508 11056 10560 11076
rect 10560 11056 10562 11076
rect 10289 10362 10345 10364
rect 10369 10362 10425 10364
rect 10449 10362 10505 10364
rect 10529 10362 10585 10364
rect 10289 10310 10315 10362
rect 10315 10310 10345 10362
rect 10369 10310 10379 10362
rect 10379 10310 10425 10362
rect 10449 10310 10495 10362
rect 10495 10310 10505 10362
rect 10529 10310 10559 10362
rect 10559 10310 10585 10362
rect 10289 10308 10345 10310
rect 10369 10308 10425 10310
rect 10449 10308 10505 10310
rect 10529 10308 10585 10310
rect 10289 9274 10345 9276
rect 10369 9274 10425 9276
rect 10449 9274 10505 9276
rect 10529 9274 10585 9276
rect 10289 9222 10315 9274
rect 10315 9222 10345 9274
rect 10369 9222 10379 9274
rect 10379 9222 10425 9274
rect 10449 9222 10495 9274
rect 10495 9222 10505 9274
rect 10529 9222 10559 9274
rect 10559 9222 10585 9274
rect 10289 9220 10345 9222
rect 10369 9220 10425 9222
rect 10449 9220 10505 9222
rect 10529 9220 10585 9222
rect 10289 8186 10345 8188
rect 10369 8186 10425 8188
rect 10449 8186 10505 8188
rect 10529 8186 10585 8188
rect 10289 8134 10315 8186
rect 10315 8134 10345 8186
rect 10369 8134 10379 8186
rect 10379 8134 10425 8186
rect 10449 8134 10495 8186
rect 10495 8134 10505 8186
rect 10529 8134 10559 8186
rect 10559 8134 10585 8186
rect 10289 8132 10345 8134
rect 10369 8132 10425 8134
rect 10449 8132 10505 8134
rect 10529 8132 10585 8134
rect 11242 18028 11244 18048
rect 11244 18028 11296 18048
rect 11296 18028 11298 18048
rect 11242 17992 11298 18028
rect 11150 16632 11206 16688
rect 11242 16360 11298 16416
rect 11242 15680 11298 15736
rect 11886 23296 11942 23352
rect 11702 18944 11758 19000
rect 11426 16360 11482 16416
rect 11150 13912 11206 13968
rect 11426 15544 11482 15600
rect 11334 15000 11390 15056
rect 11242 13252 11298 13288
rect 11242 13232 11244 13252
rect 11244 13232 11296 13252
rect 11296 13232 11298 13252
rect 10782 12416 10838 12472
rect 10782 9832 10838 9888
rect 11150 11192 11206 11248
rect 10690 7112 10746 7168
rect 10289 7098 10345 7100
rect 10369 7098 10425 7100
rect 10449 7098 10505 7100
rect 10529 7098 10585 7100
rect 10289 7046 10315 7098
rect 10315 7046 10345 7098
rect 10369 7046 10379 7098
rect 10379 7046 10425 7098
rect 10449 7046 10495 7098
rect 10495 7046 10505 7098
rect 10529 7046 10559 7098
rect 10559 7046 10585 7098
rect 10289 7044 10345 7046
rect 10369 7044 10425 7046
rect 10449 7044 10505 7046
rect 10529 7044 10585 7046
rect 10138 6976 10194 7032
rect 10414 6568 10470 6624
rect 10966 8200 11022 8256
rect 10690 6024 10746 6080
rect 10289 6010 10345 6012
rect 10369 6010 10425 6012
rect 10449 6010 10505 6012
rect 10529 6010 10585 6012
rect 10289 5958 10315 6010
rect 10315 5958 10345 6010
rect 10369 5958 10379 6010
rect 10379 5958 10425 6010
rect 10449 5958 10495 6010
rect 10495 5958 10505 6010
rect 10529 5958 10559 6010
rect 10559 5958 10585 6010
rect 10289 5956 10345 5958
rect 10369 5956 10425 5958
rect 10449 5956 10505 5958
rect 10529 5956 10585 5958
rect 10782 5888 10838 5944
rect 10690 5752 10746 5808
rect 10289 4922 10345 4924
rect 10369 4922 10425 4924
rect 10449 4922 10505 4924
rect 10529 4922 10585 4924
rect 10289 4870 10315 4922
rect 10315 4870 10345 4922
rect 10369 4870 10379 4922
rect 10379 4870 10425 4922
rect 10449 4870 10495 4922
rect 10495 4870 10505 4922
rect 10529 4870 10559 4922
rect 10559 4870 10585 4922
rect 10289 4868 10345 4870
rect 10369 4868 10425 4870
rect 10449 4868 10505 4870
rect 10529 4868 10585 4870
rect 10782 4800 10838 4856
rect 11334 9016 11390 9072
rect 11150 5344 11206 5400
rect 10690 3848 10746 3904
rect 10289 3834 10345 3836
rect 10369 3834 10425 3836
rect 10449 3834 10505 3836
rect 10529 3834 10585 3836
rect 10289 3782 10315 3834
rect 10315 3782 10345 3834
rect 10369 3782 10379 3834
rect 10379 3782 10425 3834
rect 10449 3782 10495 3834
rect 10495 3782 10505 3834
rect 10529 3782 10559 3834
rect 10559 3782 10585 3834
rect 10289 3780 10345 3782
rect 10369 3780 10425 3782
rect 10449 3780 10505 3782
rect 10529 3780 10585 3782
rect 11150 4392 11206 4448
rect 11058 4120 11114 4176
rect 10690 3304 10746 3360
rect 10289 2746 10345 2748
rect 10369 2746 10425 2748
rect 10449 2746 10505 2748
rect 10529 2746 10585 2748
rect 10289 2694 10315 2746
rect 10315 2694 10345 2746
rect 10369 2694 10379 2746
rect 10379 2694 10425 2746
rect 10449 2694 10495 2746
rect 10495 2694 10505 2746
rect 10529 2694 10559 2746
rect 10559 2694 10585 2746
rect 10289 2692 10345 2694
rect 10369 2692 10425 2694
rect 10449 2692 10505 2694
rect 10529 2692 10585 2694
rect 10138 2644 10194 2680
rect 10138 2624 10140 2644
rect 10140 2624 10192 2644
rect 10192 2624 10194 2644
rect 10966 3712 11022 3768
rect 11242 4256 11298 4312
rect 11794 15952 11850 16008
rect 11702 14476 11758 14512
rect 11702 14456 11704 14476
rect 11704 14456 11756 14476
rect 11756 14456 11758 14476
rect 11518 11600 11574 11656
rect 11702 10920 11758 10976
rect 11886 14184 11942 14240
rect 11886 11348 11942 11384
rect 11886 11328 11888 11348
rect 11888 11328 11940 11348
rect 11940 11328 11942 11348
rect 11886 10124 11942 10160
rect 11886 10104 11888 10124
rect 11888 10104 11940 10124
rect 11940 10104 11942 10124
rect 11794 4936 11850 4992
rect 11702 4120 11758 4176
rect 11518 3612 11520 3632
rect 11520 3612 11572 3632
rect 11572 3612 11574 3632
rect 11518 3576 11574 3612
rect 10874 1944 10930 2000
rect 11886 4256 11942 4312
rect 11702 3168 11758 3224
rect 11242 3032 11298 3088
rect 11334 2896 11390 2952
rect 11242 2760 11298 2816
rect 11242 1128 11298 1184
rect 12346 23704 12402 23760
rect 12254 22752 12310 22808
rect 12806 23160 12862 23216
rect 13358 24792 13414 24848
rect 13542 24928 13598 24984
rect 14186 25744 14242 25800
rect 13174 23432 13230 23488
rect 13726 24384 13782 24440
rect 13266 22480 13322 22536
rect 13082 22208 13138 22264
rect 12990 22072 13046 22128
rect 12530 21664 12586 21720
rect 12346 21528 12402 21584
rect 12254 21120 12310 21176
rect 12070 20712 12126 20768
rect 12070 20168 12126 20224
rect 12162 19896 12218 19952
rect 12070 17720 12126 17776
rect 12622 21004 12678 21040
rect 12622 20984 12624 21004
rect 12624 20984 12676 21004
rect 12676 20984 12678 21004
rect 12622 20848 12678 20904
rect 12530 20168 12586 20224
rect 12898 19624 12954 19680
rect 13726 22208 13782 22264
rect 13358 20440 13414 20496
rect 13082 19760 13138 19816
rect 12530 19252 12532 19272
rect 12532 19252 12584 19272
rect 12584 19252 12586 19272
rect 12530 19216 12586 19252
rect 12438 18672 12494 18728
rect 12530 18400 12586 18456
rect 12346 12960 12402 13016
rect 12070 10920 12126 10976
rect 12070 9968 12126 10024
rect 12070 6840 12126 6896
rect 12254 10648 12310 10704
rect 12898 17176 12954 17232
rect 12806 13912 12862 13968
rect 12898 13812 12900 13832
rect 12900 13812 12952 13832
rect 12952 13812 12954 13832
rect 12898 13776 12954 13812
rect 12438 12144 12494 12200
rect 12622 11872 12678 11928
rect 12622 11328 12678 11384
rect 12346 3984 12402 4040
rect 12622 5908 12678 5944
rect 12622 5888 12624 5908
rect 12624 5888 12676 5908
rect 12676 5888 12678 5908
rect 12622 5344 12678 5400
rect 12898 12144 12954 12200
rect 12898 11736 12954 11792
rect 13082 13232 13138 13288
rect 13266 20032 13322 20088
rect 13266 17176 13322 17232
rect 13266 15952 13322 16008
rect 13450 15272 13506 15328
rect 13174 12588 13176 12608
rect 13176 12588 13228 12608
rect 13228 12588 13230 12608
rect 13174 12552 13230 12588
rect 13174 11464 13230 11520
rect 12990 10784 13046 10840
rect 13174 10648 13230 10704
rect 13542 14864 13598 14920
rect 13818 16360 13874 16416
rect 13726 15680 13782 15736
rect 13818 15408 13874 15464
rect 14002 19760 14058 19816
rect 14278 24792 14334 24848
rect 14278 23024 14334 23080
rect 14646 23568 14702 23624
rect 14370 21528 14426 21584
rect 14278 20848 14334 20904
rect 14186 20576 14242 20632
rect 14370 20304 14426 20360
rect 14646 21936 14702 21992
rect 14956 25050 15012 25052
rect 15036 25050 15092 25052
rect 15116 25050 15172 25052
rect 15196 25050 15252 25052
rect 14956 24998 14982 25050
rect 14982 24998 15012 25050
rect 15036 24998 15046 25050
rect 15046 24998 15092 25050
rect 15116 24998 15162 25050
rect 15162 24998 15172 25050
rect 15196 24998 15226 25050
rect 15226 24998 15252 25050
rect 14956 24996 15012 24998
rect 15036 24996 15092 24998
rect 15116 24996 15172 24998
rect 15196 24996 15252 24998
rect 15106 24284 15108 24304
rect 15108 24284 15160 24304
rect 15160 24284 15162 24304
rect 15106 24248 15162 24284
rect 14830 24132 14886 24168
rect 14830 24112 14832 24132
rect 14832 24112 14884 24132
rect 14884 24112 14886 24132
rect 14956 23962 15012 23964
rect 15036 23962 15092 23964
rect 15116 23962 15172 23964
rect 15196 23962 15252 23964
rect 14956 23910 14982 23962
rect 14982 23910 15012 23962
rect 15036 23910 15046 23962
rect 15046 23910 15092 23962
rect 15116 23910 15162 23962
rect 15162 23910 15172 23962
rect 15196 23910 15226 23962
rect 15226 23910 15252 23962
rect 14956 23908 15012 23910
rect 15036 23908 15092 23910
rect 15116 23908 15172 23910
rect 15196 23908 15252 23910
rect 15198 23740 15200 23760
rect 15200 23740 15252 23760
rect 15252 23740 15254 23760
rect 15198 23704 15254 23740
rect 15474 23296 15530 23352
rect 14956 22874 15012 22876
rect 15036 22874 15092 22876
rect 15116 22874 15172 22876
rect 15196 22874 15252 22876
rect 14956 22822 14982 22874
rect 14982 22822 15012 22874
rect 15036 22822 15046 22874
rect 15046 22822 15092 22874
rect 15116 22822 15162 22874
rect 15162 22822 15172 22874
rect 15196 22822 15226 22874
rect 15226 22822 15252 22874
rect 14956 22820 15012 22822
rect 15036 22820 15092 22822
rect 15116 22820 15172 22822
rect 15196 22820 15252 22822
rect 15474 22888 15530 22944
rect 15382 22752 15438 22808
rect 14956 21786 15012 21788
rect 15036 21786 15092 21788
rect 15116 21786 15172 21788
rect 15196 21786 15252 21788
rect 14956 21734 14982 21786
rect 14982 21734 15012 21786
rect 15036 21734 15046 21786
rect 15046 21734 15092 21786
rect 15116 21734 15162 21786
rect 15162 21734 15172 21786
rect 15196 21734 15226 21786
rect 15226 21734 15252 21786
rect 14956 21732 15012 21734
rect 15036 21732 15092 21734
rect 15116 21732 15172 21734
rect 15196 21732 15252 21734
rect 14370 18128 14426 18184
rect 14002 15972 14058 16008
rect 14002 15952 14004 15972
rect 14004 15952 14056 15972
rect 14056 15952 14058 15972
rect 14186 17040 14242 17096
rect 14094 15136 14150 15192
rect 13910 13232 13966 13288
rect 13542 12688 13598 12744
rect 13726 12316 13728 12336
rect 13728 12316 13780 12336
rect 13780 12316 13782 12336
rect 13726 12280 13782 12316
rect 13726 11076 13782 11112
rect 13726 11056 13728 11076
rect 13728 11056 13780 11076
rect 13780 11056 13782 11076
rect 13634 10920 13690 10976
rect 13082 8200 13138 8256
rect 12806 6724 12862 6760
rect 12806 6704 12808 6724
rect 12808 6704 12860 6724
rect 12860 6704 12862 6724
rect 12438 3304 12494 3360
rect 12070 2352 12126 2408
rect 12254 2352 12310 2408
rect 12070 1808 12126 1864
rect 12622 4820 12678 4856
rect 12622 4800 12624 4820
rect 12624 4800 12676 4820
rect 12676 4800 12678 4820
rect 12622 4020 12624 4040
rect 12624 4020 12676 4040
rect 12676 4020 12678 4040
rect 12622 3984 12678 4020
rect 12806 3848 12862 3904
rect 12806 3304 12862 3360
rect 12714 2488 12770 2544
rect 12622 1944 12678 2000
rect 12530 1808 12586 1864
rect 12438 1400 12494 1456
rect 11886 992 11942 1048
rect 13174 5344 13230 5400
rect 13174 4564 13176 4584
rect 13176 4564 13228 4584
rect 13228 4564 13230 4584
rect 13174 4528 13230 4564
rect 13174 3884 13176 3904
rect 13176 3884 13228 3904
rect 13228 3884 13230 3904
rect 13174 3848 13230 3884
rect 13082 3712 13138 3768
rect 13174 2624 13230 2680
rect 13450 9868 13452 9888
rect 13452 9868 13504 9888
rect 13504 9868 13506 9888
rect 13450 9832 13506 9868
rect 13634 10240 13690 10296
rect 13542 9152 13598 9208
rect 13450 5752 13506 5808
rect 14554 17448 14610 17504
rect 14370 16088 14426 16144
rect 14956 20698 15012 20700
rect 15036 20698 15092 20700
rect 15116 20698 15172 20700
rect 15196 20698 15252 20700
rect 14956 20646 14982 20698
rect 14982 20646 15012 20698
rect 15036 20646 15046 20698
rect 15046 20646 15092 20698
rect 15116 20646 15162 20698
rect 15162 20646 15172 20698
rect 15196 20646 15226 20698
rect 15226 20646 15252 20698
rect 14956 20644 15012 20646
rect 15036 20644 15092 20646
rect 15116 20644 15172 20646
rect 15196 20644 15252 20646
rect 14922 20476 14924 20496
rect 14924 20476 14976 20496
rect 14976 20476 14978 20496
rect 14922 20440 14978 20476
rect 15106 20440 15162 20496
rect 15198 20032 15254 20088
rect 14956 19610 15012 19612
rect 15036 19610 15092 19612
rect 15116 19610 15172 19612
rect 15196 19610 15252 19612
rect 14956 19558 14982 19610
rect 14982 19558 15012 19610
rect 15036 19558 15046 19610
rect 15046 19558 15092 19610
rect 15116 19558 15162 19610
rect 15162 19558 15172 19610
rect 15196 19558 15226 19610
rect 15226 19558 15252 19610
rect 14956 19556 15012 19558
rect 15036 19556 15092 19558
rect 15116 19556 15172 19558
rect 15196 19556 15252 19558
rect 14738 18400 14794 18456
rect 14738 18128 14794 18184
rect 14956 18522 15012 18524
rect 15036 18522 15092 18524
rect 15116 18522 15172 18524
rect 15196 18522 15252 18524
rect 14956 18470 14982 18522
rect 14982 18470 15012 18522
rect 15036 18470 15046 18522
rect 15046 18470 15092 18522
rect 15116 18470 15162 18522
rect 15162 18470 15172 18522
rect 15196 18470 15226 18522
rect 15226 18470 15252 18522
rect 14956 18468 15012 18470
rect 15036 18468 15092 18470
rect 15116 18468 15172 18470
rect 15196 18468 15252 18470
rect 14956 17434 15012 17436
rect 15036 17434 15092 17436
rect 15116 17434 15172 17436
rect 15196 17434 15252 17436
rect 14956 17382 14982 17434
rect 14982 17382 15012 17434
rect 15036 17382 15046 17434
rect 15046 17382 15092 17434
rect 15116 17382 15162 17434
rect 15162 17382 15172 17434
rect 15196 17382 15226 17434
rect 15226 17382 15252 17434
rect 14956 17380 15012 17382
rect 15036 17380 15092 17382
rect 15116 17380 15172 17382
rect 15196 17380 15252 17382
rect 14922 16668 14924 16688
rect 14924 16668 14976 16688
rect 14976 16668 14978 16688
rect 14922 16632 14978 16668
rect 14738 16496 14794 16552
rect 15934 24384 15990 24440
rect 15934 23568 15990 23624
rect 16486 24928 16542 24984
rect 15934 22888 15990 22944
rect 15934 22208 15990 22264
rect 15658 20848 15714 20904
rect 15474 20576 15530 20632
rect 15566 19624 15622 19680
rect 15658 19216 15714 19272
rect 15658 18400 15714 18456
rect 15382 17992 15438 18048
rect 15382 17584 15438 17640
rect 14956 16346 15012 16348
rect 15036 16346 15092 16348
rect 15116 16346 15172 16348
rect 15196 16346 15252 16348
rect 14956 16294 14982 16346
rect 14982 16294 15012 16346
rect 15036 16294 15046 16346
rect 15046 16294 15092 16346
rect 15116 16294 15162 16346
rect 15162 16294 15172 16346
rect 15196 16294 15226 16346
rect 15226 16294 15252 16346
rect 14956 16292 15012 16294
rect 15036 16292 15092 16294
rect 15116 16292 15172 16294
rect 15196 16292 15252 16294
rect 14830 15816 14886 15872
rect 15198 15852 15200 15872
rect 15200 15852 15252 15872
rect 15252 15852 15254 15872
rect 14370 13640 14426 13696
rect 14554 14320 14610 14376
rect 14554 13524 14610 13560
rect 14554 13504 14556 13524
rect 14556 13504 14608 13524
rect 14608 13504 14610 13524
rect 14646 13132 14648 13152
rect 14648 13132 14700 13152
rect 14700 13132 14702 13152
rect 14646 13096 14702 13132
rect 14554 12280 14610 12336
rect 14278 12044 14280 12064
rect 14280 12044 14332 12064
rect 14332 12044 14334 12064
rect 14278 12008 14334 12044
rect 14186 11772 14188 11792
rect 14188 11772 14240 11792
rect 14240 11772 14242 11792
rect 14186 11736 14242 11772
rect 15198 15816 15254 15852
rect 15014 15544 15070 15600
rect 14956 15258 15012 15260
rect 15036 15258 15092 15260
rect 15116 15258 15172 15260
rect 15196 15258 15252 15260
rect 14956 15206 14982 15258
rect 14982 15206 15012 15258
rect 15036 15206 15046 15258
rect 15046 15206 15092 15258
rect 15116 15206 15162 15258
rect 15162 15206 15172 15258
rect 15196 15206 15226 15258
rect 15226 15206 15252 15258
rect 14956 15204 15012 15206
rect 15036 15204 15092 15206
rect 15116 15204 15172 15206
rect 15196 15204 15252 15206
rect 15474 16224 15530 16280
rect 14956 14170 15012 14172
rect 15036 14170 15092 14172
rect 15116 14170 15172 14172
rect 15196 14170 15252 14172
rect 14956 14118 14982 14170
rect 14982 14118 15012 14170
rect 15036 14118 15046 14170
rect 15046 14118 15092 14170
rect 15116 14118 15162 14170
rect 15162 14118 15172 14170
rect 15196 14118 15226 14170
rect 15226 14118 15252 14170
rect 14956 14116 15012 14118
rect 15036 14116 15092 14118
rect 15116 14116 15172 14118
rect 15196 14116 15252 14118
rect 14922 13504 14978 13560
rect 14830 13252 14886 13288
rect 14830 13232 14832 13252
rect 14832 13232 14884 13252
rect 14884 13232 14886 13252
rect 14956 13082 15012 13084
rect 15036 13082 15092 13084
rect 15116 13082 15172 13084
rect 15196 13082 15252 13084
rect 14956 13030 14982 13082
rect 14982 13030 15012 13082
rect 15036 13030 15046 13082
rect 15046 13030 15092 13082
rect 15116 13030 15162 13082
rect 15162 13030 15172 13082
rect 15196 13030 15226 13082
rect 15226 13030 15252 13082
rect 14956 13028 15012 13030
rect 15036 13028 15092 13030
rect 15116 13028 15172 13030
rect 15196 13028 15252 13030
rect 15014 12588 15016 12608
rect 15016 12588 15068 12608
rect 15068 12588 15070 12608
rect 15014 12552 15070 12588
rect 14646 11228 14648 11248
rect 14648 11228 14700 11248
rect 14700 11228 14702 11248
rect 14646 11192 14702 11228
rect 14278 9152 14334 9208
rect 13726 5888 13782 5944
rect 13634 5208 13690 5264
rect 13450 3984 13506 4040
rect 13450 2760 13506 2816
rect 13634 3032 13690 3088
rect 13818 2896 13874 2952
rect 13542 2080 13598 2136
rect 14462 10784 14518 10840
rect 14554 10260 14610 10296
rect 14554 10240 14556 10260
rect 14556 10240 14608 10260
rect 14608 10240 14610 10260
rect 14646 8744 14702 8800
rect 14738 7792 14794 7848
rect 14738 7520 14794 7576
rect 14278 4256 14334 4312
rect 14094 4120 14150 4176
rect 14002 2896 14058 2952
rect 14002 1672 14058 1728
rect 14956 11994 15012 11996
rect 15036 11994 15092 11996
rect 15116 11994 15172 11996
rect 15196 11994 15252 11996
rect 14956 11942 14982 11994
rect 14982 11942 15012 11994
rect 15036 11942 15046 11994
rect 15046 11942 15092 11994
rect 15116 11942 15162 11994
rect 15162 11942 15172 11994
rect 15196 11942 15226 11994
rect 15226 11942 15252 11994
rect 14956 11940 15012 11942
rect 15036 11940 15092 11942
rect 15116 11940 15172 11942
rect 15196 11940 15252 11942
rect 15290 11212 15346 11248
rect 15290 11192 15292 11212
rect 15292 11192 15344 11212
rect 15344 11192 15346 11212
rect 14956 10906 15012 10908
rect 15036 10906 15092 10908
rect 15116 10906 15172 10908
rect 15196 10906 15252 10908
rect 14956 10854 14982 10906
rect 14982 10854 15012 10906
rect 15036 10854 15046 10906
rect 15046 10854 15092 10906
rect 15116 10854 15162 10906
rect 15162 10854 15172 10906
rect 15196 10854 15226 10906
rect 15226 10854 15252 10906
rect 14956 10852 15012 10854
rect 15036 10852 15092 10854
rect 15116 10852 15172 10854
rect 15196 10852 15252 10854
rect 15198 10648 15254 10704
rect 15382 10512 15438 10568
rect 14956 9818 15012 9820
rect 15036 9818 15092 9820
rect 15116 9818 15172 9820
rect 15196 9818 15252 9820
rect 14956 9766 14982 9818
rect 14982 9766 15012 9818
rect 15036 9766 15046 9818
rect 15046 9766 15092 9818
rect 15116 9766 15162 9818
rect 15162 9766 15172 9818
rect 15196 9766 15226 9818
rect 15226 9766 15252 9818
rect 14956 9764 15012 9766
rect 15036 9764 15092 9766
rect 15116 9764 15172 9766
rect 15196 9764 15252 9766
rect 15382 9288 15438 9344
rect 14956 8730 15012 8732
rect 15036 8730 15092 8732
rect 15116 8730 15172 8732
rect 15196 8730 15252 8732
rect 14956 8678 14982 8730
rect 14982 8678 15012 8730
rect 15036 8678 15046 8730
rect 15046 8678 15092 8730
rect 15116 8678 15162 8730
rect 15162 8678 15172 8730
rect 15196 8678 15226 8730
rect 15226 8678 15252 8730
rect 14956 8676 15012 8678
rect 15036 8676 15092 8678
rect 15116 8676 15172 8678
rect 15196 8676 15252 8678
rect 15934 19116 15936 19136
rect 15936 19116 15988 19136
rect 15988 19116 15990 19136
rect 15934 19080 15990 19116
rect 15842 18572 15844 18592
rect 15844 18572 15896 18592
rect 15896 18572 15898 18592
rect 15842 18536 15898 18572
rect 16118 17992 16174 18048
rect 15658 15680 15714 15736
rect 15750 14592 15806 14648
rect 15934 14048 15990 14104
rect 15566 13368 15622 13424
rect 15750 11348 15806 11384
rect 15750 11328 15752 11348
rect 15752 11328 15804 11348
rect 15804 11328 15806 11348
rect 15382 9016 15438 9072
rect 15750 9832 15806 9888
rect 15750 9560 15806 9616
rect 15658 8880 15714 8936
rect 15934 13252 15990 13288
rect 15934 13232 15936 13252
rect 15936 13232 15988 13252
rect 15988 13232 15990 13252
rect 16762 24112 16818 24168
rect 16578 23160 16634 23216
rect 16670 22888 16726 22944
rect 16486 22208 16542 22264
rect 16670 21956 16726 21992
rect 16670 21936 16672 21956
rect 16672 21936 16724 21956
rect 16724 21936 16726 21956
rect 16946 24284 16948 24304
rect 16948 24284 17000 24304
rect 17000 24284 17002 24304
rect 16946 24248 17002 24284
rect 17130 24692 17132 24712
rect 17132 24692 17184 24712
rect 17184 24692 17186 24712
rect 17130 24656 17186 24692
rect 17130 24384 17186 24440
rect 17038 23296 17094 23352
rect 16854 22516 16856 22536
rect 16856 22516 16908 22536
rect 16908 22516 16910 22536
rect 16854 22480 16910 22516
rect 17038 22772 17094 22808
rect 17038 22752 17040 22772
rect 17040 22752 17092 22772
rect 17092 22752 17094 22772
rect 16762 20440 16818 20496
rect 16854 19896 16910 19952
rect 16486 19760 16542 19816
rect 16946 19252 16948 19272
rect 16948 19252 17000 19272
rect 17000 19252 17002 19272
rect 16946 19216 17002 19252
rect 16486 18400 16542 18456
rect 16486 18128 16542 18184
rect 16394 16768 16450 16824
rect 16670 16496 16726 16552
rect 16394 16360 16450 16416
rect 16670 16224 16726 16280
rect 16210 14864 16266 14920
rect 16578 15000 16634 15056
rect 16210 13912 16266 13968
rect 16394 12688 16450 12744
rect 16394 12416 16450 12472
rect 16854 14456 16910 14512
rect 16762 12824 16818 12880
rect 16210 11736 16266 11792
rect 17038 13912 17094 13968
rect 16946 13776 17002 13832
rect 16118 10920 16174 10976
rect 16026 10784 16082 10840
rect 15842 9424 15898 9480
rect 15842 9016 15898 9072
rect 15566 8356 15622 8392
rect 15566 8336 15568 8356
rect 15568 8336 15620 8356
rect 15620 8336 15622 8356
rect 14956 7642 15012 7644
rect 15036 7642 15092 7644
rect 15116 7642 15172 7644
rect 15196 7642 15252 7644
rect 14956 7590 14982 7642
rect 14982 7590 15012 7642
rect 15036 7590 15046 7642
rect 15046 7590 15092 7642
rect 15116 7590 15162 7642
rect 15162 7590 15172 7642
rect 15196 7590 15226 7642
rect 15226 7590 15252 7642
rect 14956 7588 15012 7590
rect 15036 7588 15092 7590
rect 15116 7588 15172 7590
rect 15196 7588 15252 7590
rect 14554 6332 14556 6352
rect 14556 6332 14608 6352
rect 14608 6332 14610 6352
rect 14554 6296 14610 6332
rect 14738 6296 14794 6352
rect 14462 6160 14518 6216
rect 14462 4528 14518 4584
rect 14922 6840 14978 6896
rect 15014 6724 15070 6760
rect 15014 6704 15016 6724
rect 15016 6704 15068 6724
rect 15068 6704 15070 6724
rect 14956 6554 15012 6556
rect 15036 6554 15092 6556
rect 15116 6554 15172 6556
rect 15196 6554 15252 6556
rect 14956 6502 14982 6554
rect 14982 6502 15012 6554
rect 15036 6502 15046 6554
rect 15046 6502 15092 6554
rect 15116 6502 15162 6554
rect 15162 6502 15172 6554
rect 15196 6502 15226 6554
rect 15226 6502 15252 6554
rect 14956 6500 15012 6502
rect 15036 6500 15092 6502
rect 15116 6500 15172 6502
rect 15196 6500 15252 6502
rect 15382 6432 15438 6488
rect 15106 6024 15162 6080
rect 15290 6024 15346 6080
rect 15014 5752 15070 5808
rect 15198 5752 15254 5808
rect 14956 5466 15012 5468
rect 15036 5466 15092 5468
rect 15116 5466 15172 5468
rect 15196 5466 15252 5468
rect 14956 5414 14982 5466
rect 14982 5414 15012 5466
rect 15036 5414 15046 5466
rect 15046 5414 15092 5466
rect 15116 5414 15162 5466
rect 15162 5414 15172 5466
rect 15196 5414 15226 5466
rect 15226 5414 15252 5466
rect 14956 5412 15012 5414
rect 15036 5412 15092 5414
rect 15116 5412 15172 5414
rect 15196 5412 15252 5414
rect 14956 4378 15012 4380
rect 15036 4378 15092 4380
rect 15116 4378 15172 4380
rect 15196 4378 15252 4380
rect 14956 4326 14982 4378
rect 14982 4326 15012 4378
rect 15036 4326 15046 4378
rect 15046 4326 15092 4378
rect 15116 4326 15162 4378
rect 15162 4326 15172 4378
rect 15196 4326 15226 4378
rect 15226 4326 15252 4378
rect 14956 4324 15012 4326
rect 15036 4324 15092 4326
rect 15116 4324 15172 4326
rect 15196 4324 15252 4326
rect 14738 3576 14794 3632
rect 15842 7540 15898 7576
rect 15842 7520 15844 7540
rect 15844 7520 15896 7540
rect 15896 7520 15898 7540
rect 14646 3304 14702 3360
rect 14646 2796 14648 2816
rect 14648 2796 14700 2816
rect 14700 2796 14702 2816
rect 14646 2760 14702 2796
rect 14462 2488 14518 2544
rect 15014 3576 15070 3632
rect 14956 3290 15012 3292
rect 15036 3290 15092 3292
rect 15116 3290 15172 3292
rect 15196 3290 15252 3292
rect 14956 3238 14982 3290
rect 14982 3238 15012 3290
rect 15036 3238 15046 3290
rect 15046 3238 15092 3290
rect 15116 3238 15162 3290
rect 15162 3238 15172 3290
rect 15196 3238 15226 3290
rect 15226 3238 15252 3290
rect 14956 3236 15012 3238
rect 15036 3236 15092 3238
rect 15116 3236 15172 3238
rect 15196 3236 15252 3238
rect 15474 3188 15530 3224
rect 15474 3168 15476 3188
rect 15476 3168 15528 3188
rect 15528 3168 15530 3188
rect 15198 2760 15254 2816
rect 14956 2202 15012 2204
rect 15036 2202 15092 2204
rect 15116 2202 15172 2204
rect 15196 2202 15252 2204
rect 14956 2150 14982 2202
rect 14982 2150 15012 2202
rect 15036 2150 15046 2202
rect 15046 2150 15092 2202
rect 15116 2150 15162 2202
rect 15162 2150 15172 2202
rect 15196 2150 15226 2202
rect 15226 2150 15252 2202
rect 14956 2148 15012 2150
rect 15036 2148 15092 2150
rect 15116 2148 15172 2150
rect 15196 2148 15252 2150
rect 15382 2100 15438 2136
rect 15382 2080 15384 2100
rect 15384 2080 15436 2100
rect 15436 2080 15438 2100
rect 15750 3984 15806 4040
rect 15658 3848 15714 3904
rect 15658 2760 15714 2816
rect 16394 10004 16396 10024
rect 16396 10004 16448 10024
rect 16448 10004 16450 10024
rect 16394 9968 16450 10004
rect 16118 8608 16174 8664
rect 16302 8744 16358 8800
rect 17314 21120 17370 21176
rect 17222 20168 17278 20224
rect 17682 24132 17738 24168
rect 17682 24112 17684 24132
rect 17684 24112 17736 24132
rect 17736 24112 17738 24132
rect 17774 23024 17830 23080
rect 18050 23976 18106 24032
rect 18050 21392 18106 21448
rect 17498 20168 17554 20224
rect 17774 20324 17830 20360
rect 17774 20304 17776 20324
rect 17776 20304 17828 20324
rect 17828 20304 17830 20324
rect 17682 20032 17738 20088
rect 17498 19080 17554 19136
rect 17314 18400 17370 18456
rect 17222 17176 17278 17232
rect 17498 17720 17554 17776
rect 17774 18672 17830 18728
rect 17774 18128 17830 18184
rect 18050 19760 18106 19816
rect 17958 16904 18014 16960
rect 17314 15136 17370 15192
rect 17314 13640 17370 13696
rect 18418 21936 18474 21992
rect 18878 24520 18934 24576
rect 18050 16632 18106 16688
rect 18050 16396 18052 16416
rect 18052 16396 18104 16416
rect 18104 16396 18106 16416
rect 18050 16360 18106 16396
rect 18142 15816 18198 15872
rect 18050 15680 18106 15736
rect 18786 23432 18842 23488
rect 18418 18808 18474 18864
rect 18602 18128 18658 18184
rect 18602 17992 18658 18048
rect 18510 17856 18566 17912
rect 18418 16904 18474 16960
rect 18418 16768 18474 16824
rect 18510 15408 18566 15464
rect 20074 26016 20130 26072
rect 20074 25608 20130 25664
rect 19622 25594 19678 25596
rect 19702 25594 19758 25596
rect 19782 25594 19838 25596
rect 19862 25594 19918 25596
rect 19622 25542 19648 25594
rect 19648 25542 19678 25594
rect 19702 25542 19712 25594
rect 19712 25542 19758 25594
rect 19782 25542 19828 25594
rect 19828 25542 19838 25594
rect 19862 25542 19892 25594
rect 19892 25542 19918 25594
rect 19622 25540 19678 25542
rect 19702 25540 19758 25542
rect 19782 25540 19838 25542
rect 19862 25540 19918 25542
rect 19338 23180 19394 23216
rect 19338 23160 19340 23180
rect 19340 23160 19392 23180
rect 19392 23160 19394 23180
rect 19246 22344 19302 22400
rect 19338 21120 19394 21176
rect 18878 20304 18934 20360
rect 19982 24656 20038 24712
rect 19622 24506 19678 24508
rect 19702 24506 19758 24508
rect 19782 24506 19838 24508
rect 19862 24506 19918 24508
rect 19622 24454 19648 24506
rect 19648 24454 19678 24506
rect 19702 24454 19712 24506
rect 19712 24454 19758 24506
rect 19782 24454 19828 24506
rect 19828 24454 19838 24506
rect 19862 24454 19892 24506
rect 19892 24454 19918 24506
rect 19622 24452 19678 24454
rect 19702 24452 19758 24454
rect 19782 24452 19838 24454
rect 19862 24452 19918 24454
rect 19522 24248 19578 24304
rect 19622 23418 19678 23420
rect 19702 23418 19758 23420
rect 19782 23418 19838 23420
rect 19862 23418 19918 23420
rect 19622 23366 19648 23418
rect 19648 23366 19678 23418
rect 19702 23366 19712 23418
rect 19712 23366 19758 23418
rect 19782 23366 19828 23418
rect 19828 23366 19838 23418
rect 19862 23366 19892 23418
rect 19892 23366 19918 23418
rect 19622 23364 19678 23366
rect 19702 23364 19758 23366
rect 19782 23364 19838 23366
rect 19862 23364 19918 23366
rect 20258 24384 20314 24440
rect 20166 24248 20222 24304
rect 20810 25744 20866 25800
rect 20350 23976 20406 24032
rect 20166 22888 20222 22944
rect 20074 22752 20130 22808
rect 20074 22344 20130 22400
rect 19622 22330 19678 22332
rect 19702 22330 19758 22332
rect 19782 22330 19838 22332
rect 19862 22330 19918 22332
rect 19622 22278 19648 22330
rect 19648 22278 19678 22330
rect 19702 22278 19712 22330
rect 19712 22278 19758 22330
rect 19782 22278 19828 22330
rect 19828 22278 19838 22330
rect 19862 22278 19892 22330
rect 19892 22278 19918 22330
rect 19622 22276 19678 22278
rect 19702 22276 19758 22278
rect 19782 22276 19838 22278
rect 19862 22276 19918 22278
rect 19706 21412 19762 21448
rect 19706 21392 19708 21412
rect 19708 21392 19760 21412
rect 19760 21392 19762 21412
rect 19622 21242 19678 21244
rect 19702 21242 19758 21244
rect 19782 21242 19838 21244
rect 19862 21242 19918 21244
rect 19622 21190 19648 21242
rect 19648 21190 19678 21242
rect 19702 21190 19712 21242
rect 19712 21190 19758 21242
rect 19782 21190 19828 21242
rect 19828 21190 19838 21242
rect 19862 21190 19892 21242
rect 19892 21190 19918 21242
rect 19622 21188 19678 21190
rect 19702 21188 19758 21190
rect 19782 21188 19838 21190
rect 19862 21188 19918 21190
rect 19982 20712 20038 20768
rect 19622 20154 19678 20156
rect 19702 20154 19758 20156
rect 19782 20154 19838 20156
rect 19862 20154 19918 20156
rect 19622 20102 19648 20154
rect 19648 20102 19678 20154
rect 19702 20102 19712 20154
rect 19712 20102 19758 20154
rect 19782 20102 19828 20154
rect 19828 20102 19838 20154
rect 19862 20102 19892 20154
rect 19892 20102 19918 20154
rect 19622 20100 19678 20102
rect 19702 20100 19758 20102
rect 19782 20100 19838 20102
rect 19862 20100 19918 20102
rect 19982 19760 20038 19816
rect 18970 17448 19026 17504
rect 18970 16360 19026 16416
rect 17866 13640 17922 13696
rect 17406 12960 17462 13016
rect 17222 12300 17278 12336
rect 17222 12280 17224 12300
rect 17224 12280 17276 12300
rect 17276 12280 17278 12300
rect 16210 6976 16266 7032
rect 16486 6568 16542 6624
rect 16210 856 16266 912
rect 9678 40 9734 96
rect 17130 6704 17186 6760
rect 16854 6296 16910 6352
rect 17130 6432 17186 6488
rect 17314 11328 17370 11384
rect 17498 11192 17554 11248
rect 17406 9324 17408 9344
rect 17408 9324 17460 9344
rect 17460 9324 17462 9344
rect 17406 9288 17462 9324
rect 17682 12280 17738 12336
rect 17774 12144 17830 12200
rect 17590 9152 17646 9208
rect 17038 4392 17094 4448
rect 16946 3884 16948 3904
rect 16948 3884 17000 3904
rect 17000 3884 17002 3904
rect 16946 3848 17002 3884
rect 16854 2644 16910 2680
rect 16854 2624 16856 2644
rect 16856 2624 16908 2644
rect 16908 2624 16910 2644
rect 16670 2488 16726 2544
rect 16670 2216 16726 2272
rect 17498 3984 17554 4040
rect 17038 720 17094 776
rect 17406 1672 17462 1728
rect 17774 11328 17830 11384
rect 17866 10648 17922 10704
rect 18510 14320 18566 14376
rect 18510 13504 18566 13560
rect 18326 13368 18382 13424
rect 18786 14612 18842 14648
rect 18786 14592 18788 14612
rect 18788 14592 18840 14612
rect 18840 14592 18842 14612
rect 18326 10804 18382 10840
rect 18326 10784 18328 10804
rect 18328 10784 18380 10804
rect 18380 10784 18382 10804
rect 17866 10124 17922 10160
rect 17866 10104 17868 10124
rect 17868 10104 17920 10124
rect 17920 10104 17922 10124
rect 17774 9560 17830 9616
rect 17866 8064 17922 8120
rect 18050 8880 18106 8936
rect 18510 10784 18566 10840
rect 18418 10260 18474 10296
rect 18418 10240 18420 10260
rect 18420 10240 18472 10260
rect 18472 10240 18474 10260
rect 18418 9324 18420 9344
rect 18420 9324 18472 9344
rect 18472 9324 18474 9344
rect 18418 9288 18474 9324
rect 18510 8336 18566 8392
rect 18050 3712 18106 3768
rect 18050 2896 18106 2952
rect 18878 11872 18934 11928
rect 18510 6060 18512 6080
rect 18512 6060 18564 6080
rect 18564 6060 18566 6080
rect 18510 6024 18566 6060
rect 18326 5888 18382 5944
rect 18418 5480 18474 5536
rect 18602 5228 18658 5264
rect 18602 5208 18604 5228
rect 18604 5208 18656 5228
rect 18656 5208 18658 5228
rect 18418 4972 18420 4992
rect 18420 4972 18472 4992
rect 18472 4972 18474 4992
rect 18418 4936 18474 4972
rect 18602 4800 18658 4856
rect 18510 4528 18566 4584
rect 18418 3304 18474 3360
rect 19430 19080 19486 19136
rect 19622 19066 19678 19068
rect 19702 19066 19758 19068
rect 19782 19066 19838 19068
rect 19862 19066 19918 19068
rect 19622 19014 19648 19066
rect 19648 19014 19678 19066
rect 19702 19014 19712 19066
rect 19712 19014 19758 19066
rect 19782 19014 19828 19066
rect 19828 19014 19838 19066
rect 19862 19014 19892 19066
rect 19892 19014 19918 19066
rect 19622 19012 19678 19014
rect 19702 19012 19758 19014
rect 19782 19012 19838 19014
rect 19862 19012 19918 19014
rect 19522 18400 19578 18456
rect 19338 18264 19394 18320
rect 19614 18148 19670 18184
rect 19614 18128 19616 18148
rect 19616 18128 19668 18148
rect 19668 18128 19670 18148
rect 19622 17978 19678 17980
rect 19702 17978 19758 17980
rect 19782 17978 19838 17980
rect 19862 17978 19918 17980
rect 19622 17926 19648 17978
rect 19648 17926 19678 17978
rect 19702 17926 19712 17978
rect 19712 17926 19758 17978
rect 19782 17926 19828 17978
rect 19828 17926 19838 17978
rect 19862 17926 19892 17978
rect 19892 17926 19918 17978
rect 19622 17924 19678 17926
rect 19702 17924 19758 17926
rect 19782 17924 19838 17926
rect 19862 17924 19918 17926
rect 19982 17720 20038 17776
rect 19430 17448 19486 17504
rect 19522 17312 19578 17368
rect 19622 16890 19678 16892
rect 19702 16890 19758 16892
rect 19782 16890 19838 16892
rect 19862 16890 19918 16892
rect 19622 16838 19648 16890
rect 19648 16838 19678 16890
rect 19702 16838 19712 16890
rect 19712 16838 19758 16890
rect 19782 16838 19828 16890
rect 19828 16838 19838 16890
rect 19862 16838 19892 16890
rect 19892 16838 19918 16890
rect 19622 16836 19678 16838
rect 19702 16836 19758 16838
rect 19782 16836 19838 16838
rect 19862 16836 19918 16838
rect 19890 16224 19946 16280
rect 19154 15680 19210 15736
rect 19246 14864 19302 14920
rect 19246 14068 19302 14104
rect 19246 14048 19248 14068
rect 19248 14048 19300 14068
rect 19300 14048 19302 14068
rect 19982 16088 20038 16144
rect 19622 15802 19678 15804
rect 19702 15802 19758 15804
rect 19782 15802 19838 15804
rect 19862 15802 19918 15804
rect 19622 15750 19648 15802
rect 19648 15750 19678 15802
rect 19702 15750 19712 15802
rect 19712 15750 19758 15802
rect 19782 15750 19828 15802
rect 19828 15750 19838 15802
rect 19862 15750 19892 15802
rect 19892 15750 19918 15802
rect 19622 15748 19678 15750
rect 19702 15748 19758 15750
rect 19782 15748 19838 15750
rect 19862 15748 19918 15750
rect 19982 15000 20038 15056
rect 19622 14714 19678 14716
rect 19702 14714 19758 14716
rect 19782 14714 19838 14716
rect 19862 14714 19918 14716
rect 19622 14662 19648 14714
rect 19648 14662 19678 14714
rect 19702 14662 19712 14714
rect 19712 14662 19758 14714
rect 19782 14662 19828 14714
rect 19828 14662 19838 14714
rect 19862 14662 19892 14714
rect 19892 14662 19918 14714
rect 19622 14660 19678 14662
rect 19702 14660 19758 14662
rect 19782 14660 19838 14662
rect 19862 14660 19918 14662
rect 19430 13640 19486 13696
rect 19622 13626 19678 13628
rect 19702 13626 19758 13628
rect 19782 13626 19838 13628
rect 19862 13626 19918 13628
rect 19622 13574 19648 13626
rect 19648 13574 19678 13626
rect 19702 13574 19712 13626
rect 19712 13574 19758 13626
rect 19782 13574 19828 13626
rect 19828 13574 19838 13626
rect 19862 13574 19892 13626
rect 19892 13574 19918 13626
rect 19622 13572 19678 13574
rect 19702 13572 19758 13574
rect 19782 13572 19838 13574
rect 19862 13572 19918 13574
rect 20350 22752 20406 22808
rect 19522 12960 19578 13016
rect 19706 12960 19762 13016
rect 19430 12552 19486 12608
rect 19246 11056 19302 11112
rect 18970 9968 19026 10024
rect 19062 9424 19118 9480
rect 19154 9016 19210 9072
rect 19430 11464 19486 11520
rect 19622 12538 19678 12540
rect 19702 12538 19758 12540
rect 19782 12538 19838 12540
rect 19862 12538 19918 12540
rect 19622 12486 19648 12538
rect 19648 12486 19678 12538
rect 19702 12486 19712 12538
rect 19712 12486 19758 12538
rect 19782 12486 19828 12538
rect 19828 12486 19838 12538
rect 19862 12486 19892 12538
rect 19892 12486 19918 12538
rect 19622 12484 19678 12486
rect 19702 12484 19758 12486
rect 19782 12484 19838 12486
rect 19862 12484 19918 12486
rect 19622 11450 19678 11452
rect 19702 11450 19758 11452
rect 19782 11450 19838 11452
rect 19862 11450 19918 11452
rect 19622 11398 19648 11450
rect 19648 11398 19678 11450
rect 19702 11398 19712 11450
rect 19712 11398 19758 11450
rect 19782 11398 19828 11450
rect 19828 11398 19838 11450
rect 19862 11398 19892 11450
rect 19892 11398 19918 11450
rect 19622 11396 19678 11398
rect 19702 11396 19758 11398
rect 19782 11396 19838 11398
rect 19862 11396 19918 11398
rect 19522 10920 19578 10976
rect 20074 11056 20130 11112
rect 19430 9968 19486 10024
rect 19622 10362 19678 10364
rect 19702 10362 19758 10364
rect 19782 10362 19838 10364
rect 19862 10362 19918 10364
rect 19622 10310 19648 10362
rect 19648 10310 19678 10362
rect 19702 10310 19712 10362
rect 19712 10310 19758 10362
rect 19782 10310 19828 10362
rect 19828 10310 19838 10362
rect 19862 10310 19892 10362
rect 19892 10310 19918 10362
rect 19622 10308 19678 10310
rect 19702 10308 19758 10310
rect 19782 10308 19838 10310
rect 19862 10308 19918 10310
rect 20074 10240 20130 10296
rect 19430 9596 19432 9616
rect 19432 9596 19484 9616
rect 19484 9596 19486 9616
rect 19430 9560 19486 9596
rect 19338 9288 19394 9344
rect 19062 8608 19118 8664
rect 19246 7792 19302 7848
rect 19430 8084 19486 8120
rect 19430 8064 19432 8084
rect 19432 8064 19484 8084
rect 19484 8064 19486 8084
rect 19622 9274 19678 9276
rect 19702 9274 19758 9276
rect 19782 9274 19838 9276
rect 19862 9274 19918 9276
rect 19622 9222 19648 9274
rect 19648 9222 19678 9274
rect 19702 9222 19712 9274
rect 19712 9222 19758 9274
rect 19782 9222 19828 9274
rect 19828 9222 19838 9274
rect 19862 9222 19892 9274
rect 19892 9222 19918 9274
rect 19622 9220 19678 9222
rect 19702 9220 19758 9222
rect 19782 9220 19838 9222
rect 19862 9220 19918 9222
rect 19890 8780 19892 8800
rect 19892 8780 19944 8800
rect 19944 8780 19946 8800
rect 19890 8744 19946 8780
rect 19890 8608 19946 8664
rect 20074 8628 20130 8664
rect 20074 8608 20076 8628
rect 20076 8608 20128 8628
rect 20128 8608 20130 8628
rect 19622 8186 19678 8188
rect 19702 8186 19758 8188
rect 19782 8186 19838 8188
rect 19862 8186 19918 8188
rect 19622 8134 19648 8186
rect 19648 8134 19678 8186
rect 19702 8134 19712 8186
rect 19712 8134 19758 8186
rect 19782 8134 19828 8186
rect 19828 8134 19838 8186
rect 19862 8134 19892 8186
rect 19892 8134 19918 8186
rect 19622 8132 19678 8134
rect 19702 8132 19758 8134
rect 19782 8132 19838 8134
rect 19862 8132 19918 8134
rect 20074 8064 20130 8120
rect 19890 7948 19946 7984
rect 19890 7928 19892 7948
rect 19892 7928 19944 7948
rect 19944 7928 19946 7948
rect 20074 7812 20130 7848
rect 20074 7792 20076 7812
rect 20076 7792 20128 7812
rect 20128 7792 20130 7812
rect 19622 7098 19678 7100
rect 19702 7098 19758 7100
rect 19782 7098 19838 7100
rect 19862 7098 19918 7100
rect 19622 7046 19648 7098
rect 19648 7046 19678 7098
rect 19702 7046 19712 7098
rect 19712 7046 19758 7098
rect 19782 7046 19828 7098
rect 19828 7046 19838 7098
rect 19862 7046 19892 7098
rect 19892 7046 19918 7098
rect 19622 7044 19678 7046
rect 19702 7044 19758 7046
rect 19782 7044 19838 7046
rect 19862 7044 19918 7046
rect 19338 6296 19394 6352
rect 19522 6296 19578 6352
rect 19622 6010 19678 6012
rect 19702 6010 19758 6012
rect 19782 6010 19838 6012
rect 19862 6010 19918 6012
rect 19622 5958 19648 6010
rect 19648 5958 19678 6010
rect 19702 5958 19712 6010
rect 19712 5958 19758 6010
rect 19782 5958 19828 6010
rect 19828 5958 19838 6010
rect 19862 5958 19892 6010
rect 19892 5958 19918 6010
rect 19622 5956 19678 5958
rect 19702 5956 19758 5958
rect 19782 5956 19838 5958
rect 19862 5956 19918 5958
rect 19062 4800 19118 4856
rect 19246 3612 19248 3632
rect 19248 3612 19300 3632
rect 19300 3612 19302 3632
rect 19246 3576 19302 3612
rect 18510 3032 18566 3088
rect 18326 1536 18382 1592
rect 17222 856 17278 912
rect 16210 312 16266 368
rect 18234 1400 18290 1456
rect 17222 40 17278 96
rect 18786 2760 18842 2816
rect 18510 2080 18566 2136
rect 18694 2080 18750 2136
rect 18602 1672 18658 1728
rect 18786 1400 18842 1456
rect 19430 5208 19486 5264
rect 19522 5072 19578 5128
rect 19622 4922 19678 4924
rect 19702 4922 19758 4924
rect 19782 4922 19838 4924
rect 19862 4922 19918 4924
rect 19622 4870 19648 4922
rect 19648 4870 19678 4922
rect 19702 4870 19712 4922
rect 19712 4870 19758 4922
rect 19782 4870 19828 4922
rect 19828 4870 19838 4922
rect 19862 4870 19892 4922
rect 19892 4870 19918 4922
rect 19622 4868 19678 4870
rect 19702 4868 19758 4870
rect 19782 4868 19838 4870
rect 19862 4868 19918 4870
rect 19622 3834 19678 3836
rect 19702 3834 19758 3836
rect 19782 3834 19838 3836
rect 19862 3834 19918 3836
rect 19622 3782 19648 3834
rect 19648 3782 19678 3834
rect 19702 3782 19712 3834
rect 19712 3782 19758 3834
rect 19782 3782 19828 3834
rect 19828 3782 19838 3834
rect 19862 3782 19892 3834
rect 19892 3782 19918 3834
rect 19622 3780 19678 3782
rect 19702 3780 19758 3782
rect 19782 3780 19838 3782
rect 19862 3780 19918 3782
rect 19430 3712 19486 3768
rect 19430 2760 19486 2816
rect 19622 2746 19678 2748
rect 19702 2746 19758 2748
rect 19782 2746 19838 2748
rect 19862 2746 19918 2748
rect 19622 2694 19648 2746
rect 19648 2694 19678 2746
rect 19702 2694 19712 2746
rect 19712 2694 19758 2746
rect 19782 2694 19828 2746
rect 19828 2694 19838 2746
rect 19862 2694 19892 2746
rect 19892 2694 19918 2746
rect 19622 2692 19678 2694
rect 19702 2692 19758 2694
rect 19782 2692 19838 2694
rect 19862 2692 19918 2694
rect 19798 2372 19854 2408
rect 19798 2352 19800 2372
rect 19800 2352 19852 2372
rect 19852 2352 19854 2372
rect 18418 176 18474 232
rect 20350 15308 20352 15328
rect 20352 15308 20404 15328
rect 20404 15308 20406 15328
rect 20350 15272 20406 15308
rect 20902 24132 20958 24168
rect 20902 24112 20904 24132
rect 20904 24112 20956 24132
rect 20956 24112 20958 24132
rect 20626 22752 20682 22808
rect 20626 22072 20682 22128
rect 20902 22652 20904 22672
rect 20904 22652 20956 22672
rect 20956 22652 20958 22672
rect 20902 22616 20958 22652
rect 21086 22344 21142 22400
rect 21822 24792 21878 24848
rect 21270 23568 21326 23624
rect 22466 25064 22522 25120
rect 21546 23024 21602 23080
rect 20534 20304 20590 20360
rect 20902 20440 20958 20496
rect 20902 20168 20958 20224
rect 20626 19116 20628 19136
rect 20628 19116 20680 19136
rect 20680 19116 20682 19136
rect 20626 19080 20682 19116
rect 20902 18672 20958 18728
rect 20534 17856 20590 17912
rect 20718 17856 20774 17912
rect 20902 17484 20904 17504
rect 20904 17484 20956 17504
rect 20956 17484 20958 17504
rect 20902 17448 20958 17484
rect 20902 16940 20904 16960
rect 20904 16940 20956 16960
rect 20956 16940 20958 16960
rect 20902 16904 20958 16940
rect 20718 16632 20774 16688
rect 20718 15580 20720 15600
rect 20720 15580 20772 15600
rect 20772 15580 20774 15600
rect 20718 15544 20774 15580
rect 20902 16088 20958 16144
rect 20902 15852 20904 15872
rect 20904 15852 20956 15872
rect 20956 15852 20958 15872
rect 20902 15816 20958 15852
rect 21086 20984 21142 21040
rect 21086 20440 21142 20496
rect 21270 21392 21326 21448
rect 21362 18808 21418 18864
rect 21822 23044 21878 23080
rect 21822 23024 21824 23044
rect 21824 23024 21876 23044
rect 21876 23024 21878 23044
rect 21730 22752 21786 22808
rect 21914 21528 21970 21584
rect 21638 20712 21694 20768
rect 21638 20340 21640 20360
rect 21640 20340 21692 20360
rect 21692 20340 21694 20360
rect 21638 20304 21694 20340
rect 21638 19624 21694 19680
rect 22466 20340 22468 20360
rect 22468 20340 22520 20360
rect 22520 20340 22522 20360
rect 22466 20304 22522 20340
rect 22282 19488 22338 19544
rect 21546 18028 21548 18048
rect 21548 18028 21600 18048
rect 21600 18028 21602 18048
rect 21546 17992 21602 18028
rect 21546 16904 21602 16960
rect 21454 16768 21510 16824
rect 21362 16668 21364 16688
rect 21364 16668 21416 16688
rect 21416 16668 21418 16688
rect 21362 16632 21418 16668
rect 21270 15680 21326 15736
rect 20902 15544 20958 15600
rect 20350 13096 20406 13152
rect 20718 15136 20774 15192
rect 20718 14456 20774 14512
rect 20534 13776 20590 13832
rect 20350 7964 20352 7984
rect 20352 7964 20404 7984
rect 20404 7964 20406 7984
rect 20350 7928 20406 7964
rect 20350 7656 20406 7712
rect 20350 6976 20406 7032
rect 20350 6724 20406 6760
rect 20350 6704 20352 6724
rect 20352 6704 20404 6724
rect 20404 6704 20406 6724
rect 20258 6432 20314 6488
rect 20074 4140 20130 4176
rect 20074 4120 20076 4140
rect 20076 4120 20128 4140
rect 20128 4120 20130 4140
rect 20166 2352 20222 2408
rect 21086 15408 21142 15464
rect 20994 14048 21050 14104
rect 21086 13912 21142 13968
rect 21086 13776 21142 13832
rect 20810 12724 20812 12744
rect 20812 12724 20864 12744
rect 20864 12724 20866 12744
rect 20810 12688 20866 12724
rect 20718 12144 20774 12200
rect 20626 11736 20682 11792
rect 20810 12008 20866 12064
rect 20626 11464 20682 11520
rect 21270 12144 21326 12200
rect 20718 9868 20720 9888
rect 20720 9868 20772 9888
rect 20772 9868 20774 9888
rect 20718 9832 20774 9868
rect 20718 9424 20774 9480
rect 20626 8472 20682 8528
rect 20626 6704 20682 6760
rect 20534 4256 20590 4312
rect 21454 13504 21510 13560
rect 21822 15816 21878 15872
rect 21730 14728 21786 14784
rect 21914 13912 21970 13968
rect 21454 11620 21510 11656
rect 21454 11600 21456 11620
rect 21456 11600 21508 11620
rect 21508 11600 21510 11620
rect 21546 10648 21602 10704
rect 21362 9968 21418 10024
rect 21178 9460 21180 9480
rect 21180 9460 21232 9480
rect 21232 9460 21234 9480
rect 21178 9424 21234 9460
rect 21178 9288 21234 9344
rect 22006 12008 22062 12064
rect 21914 10684 21916 10704
rect 21916 10684 21968 10704
rect 21968 10684 21970 10704
rect 21914 10648 21970 10684
rect 21638 9288 21694 9344
rect 21362 9172 21418 9208
rect 21362 9152 21364 9172
rect 21364 9152 21416 9172
rect 21416 9152 21418 9172
rect 21546 9152 21602 9208
rect 21454 8744 21510 8800
rect 21270 8472 21326 8528
rect 20994 7792 21050 7848
rect 21086 6704 21142 6760
rect 21178 6452 21234 6488
rect 21178 6432 21180 6452
rect 21180 6432 21232 6452
rect 21232 6432 21234 6452
rect 21178 4972 21180 4992
rect 21180 4972 21232 4992
rect 21232 4972 21234 4992
rect 21178 4936 21234 4972
rect 21362 5908 21418 5944
rect 21362 5888 21364 5908
rect 21364 5888 21416 5908
rect 21416 5888 21418 5908
rect 21362 5344 21418 5400
rect 20994 4664 21050 4720
rect 20810 4392 20866 4448
rect 20902 3848 20958 3904
rect 20994 3712 21050 3768
rect 21270 4256 21326 4312
rect 21178 3712 21234 3768
rect 20810 2488 20866 2544
rect 20718 1808 20774 1864
rect 19982 312 20038 368
rect 20902 2252 20904 2272
rect 20904 2252 20956 2272
rect 20956 2252 20958 2272
rect 20902 2216 20958 2252
rect 21086 2760 21142 2816
rect 20994 2080 21050 2136
rect 21178 2488 21234 2544
rect 22374 13232 22430 13288
rect 22282 12552 22338 12608
rect 22374 12008 22430 12064
rect 22282 10376 22338 10432
rect 22466 10376 22522 10432
rect 21822 8744 21878 8800
rect 22006 8744 22062 8800
rect 21638 7792 21694 7848
rect 21546 6432 21602 6488
rect 21914 6840 21970 6896
rect 21730 5616 21786 5672
rect 21546 5344 21602 5400
rect 21638 5092 21694 5128
rect 21638 5072 21640 5092
rect 21640 5072 21692 5092
rect 21692 5072 21694 5092
rect 21546 3168 21602 3224
rect 22006 6160 22062 6216
rect 23018 24656 23074 24712
rect 23570 24792 23626 24848
rect 23202 24248 23258 24304
rect 22926 23704 22982 23760
rect 22834 23024 22890 23080
rect 22650 21800 22706 21856
rect 22742 16360 22798 16416
rect 22834 13504 22890 13560
rect 22834 13096 22890 13152
rect 22650 9560 22706 9616
rect 22282 6296 22338 6352
rect 22558 6568 22614 6624
rect 21914 3984 21970 4040
rect 22558 4256 22614 4312
rect 22006 3168 22062 3224
rect 22098 2896 22154 2952
rect 22374 2352 22430 2408
rect 22558 2216 22614 2272
rect 22374 1808 22430 1864
rect 22558 1128 22614 1184
rect 23110 22752 23166 22808
rect 23478 23196 23480 23216
rect 23480 23196 23532 23216
rect 23532 23196 23534 23216
rect 23478 23160 23534 23196
rect 23386 21664 23442 21720
rect 24030 25880 24086 25936
rect 24030 25472 24086 25528
rect 24214 25880 24270 25936
rect 24766 27104 24822 27160
rect 24766 26560 24822 26616
rect 24858 25372 24860 25392
rect 24860 25372 24912 25392
rect 24912 25372 24914 25392
rect 24858 25336 24914 25372
rect 24289 25050 24345 25052
rect 24369 25050 24425 25052
rect 24449 25050 24505 25052
rect 24529 25050 24585 25052
rect 24289 24998 24315 25050
rect 24315 24998 24345 25050
rect 24369 24998 24379 25050
rect 24379 24998 24425 25050
rect 24449 24998 24495 25050
rect 24495 24998 24505 25050
rect 24529 24998 24559 25050
rect 24559 24998 24585 25050
rect 24289 24996 24345 24998
rect 24369 24996 24425 24998
rect 24449 24996 24505 24998
rect 24529 24996 24585 24998
rect 24766 24792 24822 24848
rect 24214 24656 24270 24712
rect 24674 24404 24730 24440
rect 24674 24384 24676 24404
rect 24676 24384 24728 24404
rect 24728 24384 24730 24404
rect 24122 24112 24178 24168
rect 23938 22888 23994 22944
rect 24289 23962 24345 23964
rect 24369 23962 24425 23964
rect 24449 23962 24505 23964
rect 24529 23962 24585 23964
rect 24289 23910 24315 23962
rect 24315 23910 24345 23962
rect 24369 23910 24379 23962
rect 24379 23910 24425 23962
rect 24449 23910 24495 23962
rect 24495 23910 24505 23962
rect 24529 23910 24559 23962
rect 24559 23910 24585 23962
rect 24289 23908 24345 23910
rect 24369 23908 24425 23910
rect 24449 23908 24505 23910
rect 24529 23908 24585 23910
rect 24766 23860 24822 23896
rect 24766 23840 24768 23860
rect 24768 23840 24820 23860
rect 24820 23840 24822 23860
rect 24766 23568 24822 23624
rect 24306 23432 24362 23488
rect 24490 23468 24492 23488
rect 24492 23468 24544 23488
rect 24544 23468 24546 23488
rect 24490 23432 24546 23468
rect 24289 22874 24345 22876
rect 24369 22874 24425 22876
rect 24449 22874 24505 22876
rect 24529 22874 24585 22876
rect 24289 22822 24315 22874
rect 24315 22822 24345 22874
rect 24369 22822 24379 22874
rect 24379 22822 24425 22874
rect 24449 22822 24495 22874
rect 24495 22822 24505 22874
rect 24529 22822 24559 22874
rect 24559 22822 24585 22874
rect 24289 22820 24345 22822
rect 24369 22820 24425 22822
rect 24449 22820 24505 22822
rect 24529 22820 24585 22822
rect 23662 22616 23718 22672
rect 23478 20596 23534 20632
rect 23478 20576 23480 20596
rect 23480 20576 23532 20596
rect 23532 20576 23534 20596
rect 23202 18536 23258 18592
rect 23662 19216 23718 19272
rect 23018 13640 23074 13696
rect 23018 11056 23074 11112
rect 22926 8916 22928 8936
rect 22928 8916 22980 8936
rect 22980 8916 22982 8936
rect 22926 8880 22982 8916
rect 23018 8372 23020 8392
rect 23020 8372 23072 8392
rect 23072 8372 23074 8392
rect 23018 8336 23074 8372
rect 23570 17856 23626 17912
rect 24766 22480 24822 22536
rect 24030 22208 24086 22264
rect 23938 22092 23994 22128
rect 23938 22072 23940 22092
rect 23940 22072 23992 22092
rect 23992 22072 23994 22092
rect 23938 20712 23994 20768
rect 23938 17992 23994 18048
rect 23754 17312 23810 17368
rect 23386 16496 23442 16552
rect 23662 16768 23718 16824
rect 23570 16224 23626 16280
rect 23478 15952 23534 16008
rect 23386 15308 23388 15328
rect 23388 15308 23440 15328
rect 23440 15308 23442 15328
rect 23386 15272 23442 15308
rect 23294 13912 23350 13968
rect 23662 14864 23718 14920
rect 23570 13912 23626 13968
rect 23570 13404 23572 13424
rect 23572 13404 23624 13424
rect 23624 13404 23626 13424
rect 23570 13368 23626 13404
rect 23570 13232 23626 13288
rect 23478 12980 23534 13016
rect 23478 12960 23480 12980
rect 23480 12960 23532 12980
rect 23532 12960 23534 12980
rect 23478 10804 23534 10840
rect 23478 10784 23480 10804
rect 23480 10784 23532 10804
rect 23532 10784 23534 10804
rect 23478 10260 23534 10296
rect 23478 10240 23480 10260
rect 23480 10240 23532 10260
rect 23532 10240 23534 10260
rect 24289 21786 24345 21788
rect 24369 21786 24425 21788
rect 24449 21786 24505 21788
rect 24529 21786 24585 21788
rect 24289 21734 24315 21786
rect 24315 21734 24345 21786
rect 24369 21734 24379 21786
rect 24379 21734 24425 21786
rect 24449 21734 24495 21786
rect 24495 21734 24505 21786
rect 24529 21734 24559 21786
rect 24559 21734 24585 21786
rect 24289 21732 24345 21734
rect 24369 21732 24425 21734
rect 24449 21732 24505 21734
rect 24529 21732 24585 21734
rect 24674 21256 24730 21312
rect 24289 20698 24345 20700
rect 24369 20698 24425 20700
rect 24449 20698 24505 20700
rect 24529 20698 24585 20700
rect 24289 20646 24315 20698
rect 24315 20646 24345 20698
rect 24369 20646 24379 20698
rect 24379 20646 24425 20698
rect 24449 20646 24495 20698
rect 24495 20646 24505 20698
rect 24529 20646 24559 20698
rect 24559 20646 24585 20698
rect 24289 20644 24345 20646
rect 24369 20644 24425 20646
rect 24449 20644 24505 20646
rect 24529 20644 24585 20646
rect 26054 26152 26110 26208
rect 25962 25472 26018 25528
rect 25870 24656 25926 24712
rect 25318 24112 25374 24168
rect 25410 23024 25466 23080
rect 24766 20032 24822 20088
rect 24289 19610 24345 19612
rect 24369 19610 24425 19612
rect 24449 19610 24505 19612
rect 24529 19610 24585 19612
rect 24289 19558 24315 19610
rect 24315 19558 24345 19610
rect 24369 19558 24379 19610
rect 24379 19558 24425 19610
rect 24449 19558 24495 19610
rect 24495 19558 24505 19610
rect 24529 19558 24559 19610
rect 24559 19558 24585 19610
rect 24289 19556 24345 19558
rect 24369 19556 24425 19558
rect 24449 19556 24505 19558
rect 24529 19556 24585 19558
rect 24674 19488 24730 19544
rect 24289 18522 24345 18524
rect 24369 18522 24425 18524
rect 24449 18522 24505 18524
rect 24529 18522 24585 18524
rect 24289 18470 24315 18522
rect 24315 18470 24345 18522
rect 24369 18470 24379 18522
rect 24379 18470 24425 18522
rect 24449 18470 24495 18522
rect 24495 18470 24505 18522
rect 24529 18470 24559 18522
rect 24559 18470 24585 18522
rect 24289 18468 24345 18470
rect 24369 18468 24425 18470
rect 24449 18468 24505 18470
rect 24529 18468 24585 18470
rect 24214 18264 24270 18320
rect 23754 12552 23810 12608
rect 24030 15580 24032 15600
rect 24032 15580 24084 15600
rect 24084 15580 24086 15600
rect 24030 15544 24086 15580
rect 24289 17434 24345 17436
rect 24369 17434 24425 17436
rect 24449 17434 24505 17436
rect 24529 17434 24585 17436
rect 24289 17382 24315 17434
rect 24315 17382 24345 17434
rect 24369 17382 24379 17434
rect 24379 17382 24425 17434
rect 24449 17382 24495 17434
rect 24495 17382 24505 17434
rect 24529 17382 24559 17434
rect 24559 17382 24585 17434
rect 24289 17380 24345 17382
rect 24369 17380 24425 17382
rect 24449 17380 24505 17382
rect 24529 17380 24585 17382
rect 25318 21936 25374 21992
rect 25502 21800 25558 21856
rect 25042 20204 25044 20224
rect 25044 20204 25096 20224
rect 25096 20204 25098 20224
rect 25042 20168 25098 20204
rect 25042 19352 25098 19408
rect 25410 20712 25466 20768
rect 25226 19896 25282 19952
rect 25594 20440 25650 20496
rect 25594 18944 25650 19000
rect 25042 17856 25098 17912
rect 25042 17756 25044 17776
rect 25044 17756 25096 17776
rect 25096 17756 25098 17776
rect 25042 17720 25098 17756
rect 24950 17584 25006 17640
rect 24289 16346 24345 16348
rect 24369 16346 24425 16348
rect 24449 16346 24505 16348
rect 24529 16346 24585 16348
rect 24289 16294 24315 16346
rect 24315 16294 24345 16346
rect 24369 16294 24379 16346
rect 24379 16294 24425 16346
rect 24449 16294 24495 16346
rect 24495 16294 24505 16346
rect 24529 16294 24559 16346
rect 24559 16294 24585 16346
rect 24289 16292 24345 16294
rect 24369 16292 24425 16294
rect 24449 16292 24505 16294
rect 24529 16292 24585 16294
rect 24306 15952 24362 16008
rect 24490 15700 24546 15736
rect 24490 15680 24492 15700
rect 24492 15680 24544 15700
rect 24544 15680 24546 15700
rect 24306 15544 24362 15600
rect 24289 15258 24345 15260
rect 24369 15258 24425 15260
rect 24449 15258 24505 15260
rect 24529 15258 24585 15260
rect 24289 15206 24315 15258
rect 24315 15206 24345 15258
rect 24369 15206 24379 15258
rect 24379 15206 24425 15258
rect 24449 15206 24495 15258
rect 24495 15206 24505 15258
rect 24529 15206 24559 15258
rect 24559 15206 24585 15258
rect 24289 15204 24345 15206
rect 24369 15204 24425 15206
rect 24449 15204 24505 15206
rect 24529 15204 24585 15206
rect 24122 14764 24124 14784
rect 24124 14764 24176 14784
rect 24176 14764 24178 14784
rect 24122 14728 24178 14764
rect 24122 14592 24178 14648
rect 24030 14184 24086 14240
rect 23938 14048 23994 14104
rect 23938 13912 23994 13968
rect 24030 13504 24086 13560
rect 23386 9152 23442 9208
rect 23294 9016 23350 9072
rect 23202 8356 23258 8392
rect 23202 8336 23204 8356
rect 23204 8336 23256 8356
rect 23256 8336 23258 8356
rect 23110 8064 23166 8120
rect 22926 7928 22982 7984
rect 23662 8472 23718 8528
rect 22742 7148 22744 7168
rect 22744 7148 22796 7168
rect 22796 7148 22798 7168
rect 22742 7112 22798 7148
rect 22742 6180 22798 6216
rect 22742 6160 22744 6180
rect 22744 6160 22796 6180
rect 22796 6160 22798 6180
rect 23018 6024 23074 6080
rect 23386 7520 23442 7576
rect 23478 6976 23534 7032
rect 22834 4800 22890 4856
rect 24858 16496 24914 16552
rect 24858 16088 24914 16144
rect 25226 17076 25228 17096
rect 25228 17076 25280 17096
rect 25280 17076 25282 17096
rect 25226 17040 25282 17076
rect 24766 14864 24822 14920
rect 24289 14170 24345 14172
rect 24369 14170 24425 14172
rect 24449 14170 24505 14172
rect 24529 14170 24585 14172
rect 24289 14118 24315 14170
rect 24315 14118 24345 14170
rect 24369 14118 24379 14170
rect 24379 14118 24425 14170
rect 24449 14118 24495 14170
rect 24495 14118 24505 14170
rect 24529 14118 24559 14170
rect 24559 14118 24585 14170
rect 24289 14116 24345 14118
rect 24369 14116 24425 14118
rect 24449 14116 24505 14118
rect 24529 14116 24585 14118
rect 24950 14728 25006 14784
rect 24674 13640 24730 13696
rect 24289 13082 24345 13084
rect 24369 13082 24425 13084
rect 24449 13082 24505 13084
rect 24529 13082 24585 13084
rect 24289 13030 24315 13082
rect 24315 13030 24345 13082
rect 24369 13030 24379 13082
rect 24379 13030 24425 13082
rect 24449 13030 24495 13082
rect 24495 13030 24505 13082
rect 24529 13030 24559 13082
rect 24559 13030 24585 13082
rect 24289 13028 24345 13030
rect 24369 13028 24425 13030
rect 24449 13028 24505 13030
rect 24529 13028 24585 13030
rect 24122 12552 24178 12608
rect 25410 17720 25466 17776
rect 25502 17176 25558 17232
rect 25410 15952 25466 16008
rect 25318 15544 25374 15600
rect 25318 15272 25374 15328
rect 25318 14864 25374 14920
rect 25226 13912 25282 13968
rect 25134 13368 25190 13424
rect 25042 13232 25098 13288
rect 24674 12552 24730 12608
rect 24582 12416 24638 12472
rect 24122 12008 24178 12064
rect 24289 11994 24345 11996
rect 24369 11994 24425 11996
rect 24449 11994 24505 11996
rect 24529 11994 24585 11996
rect 24289 11942 24315 11994
rect 24315 11942 24345 11994
rect 24369 11942 24379 11994
rect 24379 11942 24425 11994
rect 24449 11942 24495 11994
rect 24495 11942 24505 11994
rect 24529 11942 24559 11994
rect 24559 11942 24585 11994
rect 24289 11940 24345 11942
rect 24369 11940 24425 11942
rect 24449 11940 24505 11942
rect 24529 11940 24585 11942
rect 24122 11872 24178 11928
rect 23938 10648 23994 10704
rect 24582 11464 24638 11520
rect 24030 10140 24032 10160
rect 24032 10140 24084 10160
rect 24084 10140 24086 10160
rect 24030 10104 24086 10140
rect 23938 8200 23994 8256
rect 23570 6704 23626 6760
rect 22742 2488 22798 2544
rect 22926 2624 22982 2680
rect 24289 10906 24345 10908
rect 24369 10906 24425 10908
rect 24449 10906 24505 10908
rect 24529 10906 24585 10908
rect 24289 10854 24315 10906
rect 24315 10854 24345 10906
rect 24369 10854 24379 10906
rect 24379 10854 24425 10906
rect 24449 10854 24495 10906
rect 24495 10854 24505 10906
rect 24529 10854 24559 10906
rect 24559 10854 24585 10906
rect 24289 10852 24345 10854
rect 24369 10852 24425 10854
rect 24449 10852 24505 10854
rect 24529 10852 24585 10854
rect 24289 9818 24345 9820
rect 24369 9818 24425 9820
rect 24449 9818 24505 9820
rect 24529 9818 24585 9820
rect 24289 9766 24315 9818
rect 24315 9766 24345 9818
rect 24369 9766 24379 9818
rect 24379 9766 24425 9818
rect 24449 9766 24495 9818
rect 24495 9766 24505 9818
rect 24529 9766 24559 9818
rect 24559 9766 24585 9818
rect 24289 9764 24345 9766
rect 24369 9764 24425 9766
rect 24449 9764 24505 9766
rect 24529 9764 24585 9766
rect 24858 11736 24914 11792
rect 24950 11636 24952 11656
rect 24952 11636 25004 11656
rect 25004 11636 25006 11656
rect 24950 11600 25006 11636
rect 24858 11464 24914 11520
rect 24950 11328 25006 11384
rect 24582 9560 24638 9616
rect 24398 9288 24454 9344
rect 24858 9460 24860 9480
rect 24860 9460 24912 9480
rect 24912 9460 24914 9480
rect 24858 9424 24914 9460
rect 24858 9036 24914 9072
rect 24858 9016 24860 9036
rect 24860 9016 24912 9036
rect 24912 9016 24914 9036
rect 24674 8744 24730 8800
rect 24289 8730 24345 8732
rect 24369 8730 24425 8732
rect 24449 8730 24505 8732
rect 24529 8730 24585 8732
rect 24289 8678 24315 8730
rect 24315 8678 24345 8730
rect 24369 8678 24379 8730
rect 24379 8678 24425 8730
rect 24449 8678 24495 8730
rect 24495 8678 24505 8730
rect 24529 8678 24559 8730
rect 24559 8678 24585 8730
rect 24289 8676 24345 8678
rect 24369 8676 24425 8678
rect 24449 8676 24505 8678
rect 24529 8676 24585 8678
rect 24858 8508 24860 8528
rect 24860 8508 24912 8528
rect 24912 8508 24914 8528
rect 24858 8472 24914 8508
rect 25594 15272 25650 15328
rect 25502 12824 25558 12880
rect 25502 12416 25558 12472
rect 25134 10920 25190 10976
rect 25410 11228 25412 11248
rect 25412 11228 25464 11248
rect 25464 11228 25466 11248
rect 25410 11192 25466 11228
rect 25410 10920 25466 10976
rect 25318 9968 25374 10024
rect 25134 9152 25190 9208
rect 24289 7642 24345 7644
rect 24369 7642 24425 7644
rect 24449 7642 24505 7644
rect 24529 7642 24585 7644
rect 24289 7590 24315 7642
rect 24315 7590 24345 7642
rect 24369 7590 24379 7642
rect 24379 7590 24425 7642
rect 24449 7590 24495 7642
rect 24495 7590 24505 7642
rect 24529 7590 24559 7642
rect 24559 7590 24585 7642
rect 24289 7588 24345 7590
rect 24369 7588 24425 7590
rect 24449 7588 24505 7590
rect 24529 7588 24585 7590
rect 23754 5244 23756 5264
rect 23756 5244 23808 5264
rect 23808 5244 23810 5264
rect 23754 5208 23810 5244
rect 23662 4936 23718 4992
rect 22834 2352 22890 2408
rect 22926 1400 22982 1456
rect 23478 3440 23534 3496
rect 23478 3340 23480 3360
rect 23480 3340 23532 3360
rect 23532 3340 23534 3360
rect 23478 3304 23534 3340
rect 23478 3188 23534 3224
rect 23478 3168 23480 3188
rect 23480 3168 23532 3188
rect 23532 3168 23534 3188
rect 23662 3304 23718 3360
rect 23938 6024 23994 6080
rect 24030 5636 24086 5672
rect 24030 5616 24032 5636
rect 24032 5616 24084 5636
rect 24084 5616 24086 5636
rect 24030 5480 24086 5536
rect 24122 4664 24178 4720
rect 23938 3712 23994 3768
rect 23846 2252 23848 2272
rect 23848 2252 23900 2272
rect 23900 2252 23902 2272
rect 23846 2216 23902 2252
rect 24950 6976 25006 7032
rect 24766 6840 24822 6896
rect 24289 6554 24345 6556
rect 24369 6554 24425 6556
rect 24449 6554 24505 6556
rect 24529 6554 24585 6556
rect 24289 6502 24315 6554
rect 24315 6502 24345 6554
rect 24369 6502 24379 6554
rect 24379 6502 24425 6554
rect 24449 6502 24495 6554
rect 24495 6502 24505 6554
rect 24529 6502 24559 6554
rect 24559 6502 24585 6554
rect 24289 6500 24345 6502
rect 24369 6500 24425 6502
rect 24449 6500 24505 6502
rect 24529 6500 24585 6502
rect 24766 6432 24822 6488
rect 24766 6160 24822 6216
rect 24289 5466 24345 5468
rect 24369 5466 24425 5468
rect 24449 5466 24505 5468
rect 24529 5466 24585 5468
rect 24289 5414 24315 5466
rect 24315 5414 24345 5466
rect 24369 5414 24379 5466
rect 24379 5414 24425 5466
rect 24449 5414 24495 5466
rect 24495 5414 24505 5466
rect 24529 5414 24559 5466
rect 24559 5414 24585 5466
rect 24289 5412 24345 5414
rect 24369 5412 24425 5414
rect 24449 5412 24505 5414
rect 24529 5412 24585 5414
rect 24490 4684 24546 4720
rect 24490 4664 24492 4684
rect 24492 4664 24544 4684
rect 24544 4664 24546 4684
rect 24766 4664 24822 4720
rect 24289 4378 24345 4380
rect 24369 4378 24425 4380
rect 24449 4378 24505 4380
rect 24529 4378 24585 4380
rect 24289 4326 24315 4378
rect 24315 4326 24345 4378
rect 24369 4326 24379 4378
rect 24379 4326 24425 4378
rect 24449 4326 24495 4378
rect 24495 4326 24505 4378
rect 24529 4326 24559 4378
rect 24559 4326 24585 4378
rect 24289 4324 24345 4326
rect 24369 4324 24425 4326
rect 24449 4324 24505 4326
rect 24529 4324 24585 4326
rect 24306 3984 24362 4040
rect 24490 3984 24546 4040
rect 24766 3712 24822 3768
rect 24674 3304 24730 3360
rect 24289 3290 24345 3292
rect 24369 3290 24425 3292
rect 24449 3290 24505 3292
rect 24529 3290 24585 3292
rect 24289 3238 24315 3290
rect 24315 3238 24345 3290
rect 24369 3238 24379 3290
rect 24379 3238 24425 3290
rect 24449 3238 24495 3290
rect 24495 3238 24505 3290
rect 24529 3238 24559 3290
rect 24559 3238 24585 3290
rect 24289 3236 24345 3238
rect 24369 3236 24425 3238
rect 24449 3236 24505 3238
rect 24529 3236 24585 3238
rect 24289 2202 24345 2204
rect 24369 2202 24425 2204
rect 24449 2202 24505 2204
rect 24529 2202 24585 2204
rect 24289 2150 24315 2202
rect 24315 2150 24345 2202
rect 24369 2150 24379 2202
rect 24379 2150 24425 2202
rect 24449 2150 24495 2202
rect 24495 2150 24505 2202
rect 24529 2150 24559 2202
rect 24559 2150 24585 2202
rect 24289 2148 24345 2150
rect 24369 2148 24425 2150
rect 24449 2148 24505 2150
rect 24529 2148 24585 2150
rect 24122 992 24178 1048
rect 24674 1400 24730 1456
rect 24766 1264 24822 1320
rect 25594 9596 25596 9616
rect 25596 9596 25648 9616
rect 25648 9596 25650 9616
rect 25594 9560 25650 9596
rect 25226 8064 25282 8120
rect 25042 4800 25098 4856
rect 25042 3884 25044 3904
rect 25044 3884 25096 3904
rect 25096 3884 25098 3904
rect 25042 3848 25098 3884
rect 25042 3032 25098 3088
rect 25410 6060 25412 6080
rect 25412 6060 25464 6080
rect 25464 6060 25466 6080
rect 25410 6024 25466 6060
rect 25318 3984 25374 4040
rect 25410 3440 25466 3496
rect 25134 2896 25190 2952
rect 25134 2796 25136 2816
rect 25136 2796 25188 2816
rect 25188 2796 25190 2816
rect 25134 2760 25190 2796
rect 24950 2644 25006 2680
rect 24950 2624 24952 2644
rect 24952 2624 25004 2644
rect 25004 2624 25006 2644
rect 25226 1536 25282 1592
rect 26514 24384 26570 24440
rect 27618 23840 27674 23896
rect 27066 23568 27122 23624
rect 27250 23568 27306 23624
rect 25962 13096 26018 13152
rect 25870 8200 25926 8256
rect 25778 7656 25834 7712
rect 25778 7540 25834 7576
rect 25778 7520 25780 7540
rect 25780 7520 25832 7540
rect 25832 7520 25834 7540
rect 25686 7384 25742 7440
rect 26146 14592 26202 14648
rect 26238 13812 26240 13832
rect 26240 13812 26292 13832
rect 26292 13812 26294 13832
rect 26238 13776 26294 13812
rect 26330 13640 26386 13696
rect 26238 12688 26294 12744
rect 26238 12280 26294 12336
rect 26330 10412 26332 10432
rect 26332 10412 26384 10432
rect 26384 10412 26386 10432
rect 26330 10376 26386 10412
rect 26330 10260 26386 10296
rect 26330 10240 26332 10260
rect 26332 10240 26384 10260
rect 26384 10240 26386 10260
rect 26330 9596 26332 9616
rect 26332 9596 26384 9616
rect 26384 9596 26386 9616
rect 26330 9560 26386 9596
rect 25778 5788 25780 5808
rect 25780 5788 25832 5808
rect 25832 5788 25834 5808
rect 25778 5752 25834 5788
rect 25686 5072 25742 5128
rect 25686 4936 25742 4992
rect 25778 4564 25780 4584
rect 25780 4564 25832 4584
rect 25832 4564 25834 4584
rect 25778 4528 25834 4564
rect 25686 1672 25742 1728
rect 25594 720 25650 776
rect 26054 7112 26110 7168
rect 26330 8628 26386 8664
rect 26330 8608 26332 8628
rect 26332 8608 26384 8628
rect 26384 8608 26386 8628
rect 26422 7284 26424 7304
rect 26424 7284 26476 7304
rect 26476 7284 26478 7304
rect 26422 7248 26478 7284
rect 26238 5888 26294 5944
rect 26238 4120 26294 4176
rect 26238 3612 26240 3632
rect 26240 3612 26292 3632
rect 26292 3612 26294 3632
rect 26238 3576 26294 3612
rect 26330 3168 26386 3224
rect 26238 2352 26294 2408
rect 27066 3984 27122 4040
rect 26514 3304 26570 3360
rect 26422 1808 26478 1864
rect 20810 40 20866 96
rect 26146 448 26202 504
rect 27618 3440 27674 3496
<< metal3 >>
rect 0 27706 480 27736
rect 4245 27706 4311 27709
rect 0 27704 4311 27706
rect 0 27648 4250 27704
rect 4306 27648 4311 27704
rect 0 27646 4311 27648
rect 0 27616 480 27646
rect 4245 27643 4311 27646
rect 23841 27706 23907 27709
rect 27520 27706 28000 27736
rect 23841 27704 28000 27706
rect 23841 27648 23846 27704
rect 23902 27648 28000 27704
rect 23841 27646 28000 27648
rect 23841 27643 23907 27646
rect 27520 27616 28000 27646
rect 0 27162 480 27192
rect 749 27162 815 27165
rect 0 27160 815 27162
rect 0 27104 754 27160
rect 810 27104 815 27160
rect 0 27102 815 27104
rect 0 27072 480 27102
rect 749 27099 815 27102
rect 24761 27162 24827 27165
rect 27520 27162 28000 27192
rect 24761 27160 28000 27162
rect 24761 27104 24766 27160
rect 24822 27104 28000 27160
rect 24761 27102 28000 27104
rect 24761 27099 24827 27102
rect 27520 27072 28000 27102
rect 0 26618 480 26648
rect 1301 26618 1367 26621
rect 0 26616 1367 26618
rect 0 26560 1306 26616
rect 1362 26560 1367 26616
rect 0 26558 1367 26560
rect 0 26528 480 26558
rect 1301 26555 1367 26558
rect 24761 26618 24827 26621
rect 27520 26618 28000 26648
rect 24761 26616 28000 26618
rect 24761 26560 24766 26616
rect 24822 26560 28000 26616
rect 24761 26558 28000 26560
rect 24761 26555 24827 26558
rect 27520 26528 28000 26558
rect 4705 26210 4771 26213
rect 26049 26210 26115 26213
rect 4705 26208 26115 26210
rect 4705 26152 4710 26208
rect 4766 26152 26054 26208
rect 26110 26152 26115 26208
rect 4705 26150 26115 26152
rect 4705 26147 4771 26150
rect 26049 26147 26115 26150
rect 2814 26012 2820 26076
rect 2884 26074 2890 26076
rect 20069 26074 20135 26077
rect 2884 26072 20135 26074
rect 2884 26016 20074 26072
rect 20130 26016 20135 26072
rect 2884 26014 20135 26016
rect 2884 26012 2890 26014
rect 20069 26011 20135 26014
rect 0 25938 480 25968
rect 1209 25938 1275 25941
rect 0 25936 1275 25938
rect 0 25880 1214 25936
rect 1270 25880 1275 25936
rect 0 25878 1275 25880
rect 0 25848 480 25878
rect 1209 25875 1275 25878
rect 9489 25938 9555 25941
rect 24025 25938 24091 25941
rect 9489 25936 24091 25938
rect 9489 25880 9494 25936
rect 9550 25880 24030 25936
rect 24086 25880 24091 25936
rect 9489 25878 24091 25880
rect 9489 25875 9555 25878
rect 24025 25875 24091 25878
rect 24209 25938 24275 25941
rect 27520 25938 28000 25968
rect 24209 25936 28000 25938
rect 24209 25880 24214 25936
rect 24270 25880 28000 25936
rect 24209 25878 28000 25880
rect 24209 25875 24275 25878
rect 27520 25848 28000 25878
rect 9489 25802 9555 25805
rect 14181 25802 14247 25805
rect 20805 25802 20871 25805
rect 9489 25800 14247 25802
rect 9489 25744 9494 25800
rect 9550 25744 14186 25800
rect 14242 25744 14247 25800
rect 9489 25742 14247 25744
rect 9489 25739 9555 25742
rect 14181 25739 14247 25742
rect 19382 25800 20871 25802
rect 19382 25744 20810 25800
rect 20866 25744 20871 25800
rect 19382 25742 20871 25744
rect 10277 25600 10597 25601
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 25535 10597 25536
rect 10869 25530 10935 25533
rect 19382 25530 19442 25742
rect 20805 25739 20871 25742
rect 20069 25666 20135 25669
rect 25814 25666 25820 25668
rect 20069 25664 25820 25666
rect 20069 25608 20074 25664
rect 20130 25608 25820 25664
rect 20069 25606 25820 25608
rect 20069 25603 20135 25606
rect 25814 25604 25820 25606
rect 25884 25604 25890 25668
rect 19610 25600 19930 25601
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 25535 19930 25536
rect 10869 25528 19442 25530
rect 10869 25472 10874 25528
rect 10930 25472 19442 25528
rect 10869 25470 19442 25472
rect 24025 25530 24091 25533
rect 25957 25530 26023 25533
rect 24025 25528 26023 25530
rect 24025 25472 24030 25528
rect 24086 25472 25962 25528
rect 26018 25472 26023 25528
rect 24025 25470 26023 25472
rect 10869 25467 10935 25470
rect 24025 25467 24091 25470
rect 25957 25467 26023 25470
rect 0 25394 480 25424
rect 2865 25394 2931 25397
rect 0 25392 2931 25394
rect 0 25336 2870 25392
rect 2926 25336 2931 25392
rect 0 25334 2931 25336
rect 0 25304 480 25334
rect 2865 25331 2931 25334
rect 7373 25394 7439 25397
rect 23974 25394 23980 25396
rect 7373 25392 23980 25394
rect 7373 25336 7378 25392
rect 7434 25336 23980 25392
rect 7373 25334 23980 25336
rect 7373 25331 7439 25334
rect 23974 25332 23980 25334
rect 24044 25332 24050 25396
rect 24853 25394 24919 25397
rect 27520 25394 28000 25424
rect 24853 25392 28000 25394
rect 24853 25336 24858 25392
rect 24914 25336 28000 25392
rect 24853 25334 28000 25336
rect 24853 25331 24919 25334
rect 27520 25304 28000 25334
rect 10910 25196 10916 25260
rect 10980 25258 10986 25260
rect 21214 25258 21220 25260
rect 10980 25198 21220 25258
rect 10980 25196 10986 25198
rect 21214 25196 21220 25198
rect 21284 25196 21290 25260
rect 6453 25122 6519 25125
rect 10869 25122 10935 25125
rect 22461 25122 22527 25125
rect 6453 25120 10935 25122
rect 6453 25064 6458 25120
rect 6514 25064 10874 25120
rect 10930 25064 10935 25120
rect 6453 25062 10935 25064
rect 6453 25059 6519 25062
rect 10869 25059 10935 25062
rect 15334 25120 22527 25122
rect 15334 25064 22466 25120
rect 22522 25064 22527 25120
rect 15334 25062 22527 25064
rect 5610 25056 5930 25057
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5930 25056
rect 5610 24991 5930 24992
rect 14944 25056 15264 25057
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14944 24991 15264 24992
rect 13537 24986 13603 24989
rect 13537 24984 14842 24986
rect 13537 24928 13542 24984
rect 13598 24928 14842 24984
rect 13537 24926 14842 24928
rect 13537 24923 13603 24926
rect 0 24850 480 24880
rect 1117 24850 1183 24853
rect 0 24848 1183 24850
rect 0 24792 1122 24848
rect 1178 24792 1183 24848
rect 0 24790 1183 24792
rect 0 24760 480 24790
rect 1117 24787 1183 24790
rect 3141 24852 3207 24853
rect 3785 24852 3851 24853
rect 3141 24848 3188 24852
rect 3252 24850 3258 24852
rect 3734 24850 3740 24852
rect 3141 24792 3146 24848
rect 3141 24788 3188 24792
rect 3252 24790 3298 24850
rect 3694 24790 3740 24850
rect 3804 24848 3851 24852
rect 3846 24792 3851 24848
rect 3252 24788 3258 24790
rect 3734 24788 3740 24790
rect 3804 24788 3851 24792
rect 3141 24787 3207 24788
rect 3785 24787 3851 24788
rect 7281 24850 7347 24853
rect 9673 24850 9739 24853
rect 7281 24848 9739 24850
rect 7281 24792 7286 24848
rect 7342 24792 9678 24848
rect 9734 24792 9739 24848
rect 7281 24790 9739 24792
rect 7281 24787 7347 24790
rect 9673 24787 9739 24790
rect 10133 24850 10199 24853
rect 13353 24850 13419 24853
rect 14273 24852 14339 24853
rect 14222 24850 14228 24852
rect 10133 24848 13419 24850
rect 10133 24792 10138 24848
rect 10194 24792 13358 24848
rect 13414 24792 13419 24848
rect 10133 24790 13419 24792
rect 14182 24790 14228 24850
rect 14292 24848 14339 24852
rect 14334 24792 14339 24848
rect 10133 24787 10199 24790
rect 13353 24787 13419 24790
rect 14222 24788 14228 24790
rect 14292 24788 14339 24792
rect 14782 24850 14842 24926
rect 15334 24850 15394 25062
rect 22461 25059 22527 25062
rect 24277 25056 24597 25057
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 24991 24597 24992
rect 16481 24986 16547 24989
rect 23606 24986 23612 24988
rect 16481 24984 23612 24986
rect 16481 24928 16486 24984
rect 16542 24928 23612 24984
rect 16481 24926 23612 24928
rect 16481 24923 16547 24926
rect 23606 24924 23612 24926
rect 23676 24924 23682 24988
rect 14782 24790 15394 24850
rect 21817 24850 21883 24853
rect 23565 24850 23631 24853
rect 21817 24848 23631 24850
rect 21817 24792 21822 24848
rect 21878 24792 23570 24848
rect 23626 24792 23631 24848
rect 21817 24790 23631 24792
rect 14273 24787 14339 24788
rect 21817 24787 21883 24790
rect 23565 24787 23631 24790
rect 24761 24850 24827 24853
rect 27520 24850 28000 24880
rect 24761 24848 28000 24850
rect 24761 24792 24766 24848
rect 24822 24792 28000 24848
rect 24761 24790 28000 24792
rect 24761 24787 24827 24790
rect 27520 24760 28000 24790
rect 2497 24714 2563 24717
rect 2630 24714 2636 24716
rect 2497 24712 2636 24714
rect 2497 24656 2502 24712
rect 2558 24656 2636 24712
rect 2497 24654 2636 24656
rect 2497 24651 2563 24654
rect 2630 24652 2636 24654
rect 2700 24652 2706 24716
rect 7281 24714 7347 24717
rect 11605 24714 11671 24717
rect 17125 24714 17191 24717
rect 7281 24712 10794 24714
rect 7281 24656 7286 24712
rect 7342 24656 10794 24712
rect 7281 24654 10794 24656
rect 7281 24651 7347 24654
rect 10734 24578 10794 24654
rect 11605 24712 17191 24714
rect 11605 24656 11610 24712
rect 11666 24656 17130 24712
rect 17186 24656 17191 24712
rect 11605 24654 17191 24656
rect 11605 24651 11671 24654
rect 17125 24651 17191 24654
rect 19977 24714 20043 24717
rect 23013 24714 23079 24717
rect 19977 24712 23079 24714
rect 19977 24656 19982 24712
rect 20038 24656 23018 24712
rect 23074 24656 23079 24712
rect 19977 24654 23079 24656
rect 19977 24651 20043 24654
rect 23013 24651 23079 24654
rect 24209 24714 24275 24717
rect 25865 24714 25931 24717
rect 24209 24712 25931 24714
rect 24209 24656 24214 24712
rect 24270 24656 25870 24712
rect 25926 24656 25931 24712
rect 24209 24654 25931 24656
rect 24209 24651 24275 24654
rect 25865 24651 25931 24654
rect 18873 24578 18939 24581
rect 10734 24576 18939 24578
rect 10734 24520 18878 24576
rect 18934 24520 18939 24576
rect 10734 24518 18939 24520
rect 18873 24515 18939 24518
rect 10277 24512 10597 24513
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 24447 10597 24448
rect 19610 24512 19930 24513
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 24447 19930 24448
rect 2405 24442 2471 24445
rect 5993 24442 6059 24445
rect 2405 24440 6059 24442
rect 2405 24384 2410 24440
rect 2466 24384 5998 24440
rect 6054 24384 6059 24440
rect 2405 24382 6059 24384
rect 2405 24379 2471 24382
rect 5993 24379 6059 24382
rect 13721 24442 13787 24445
rect 15929 24442 15995 24445
rect 17125 24442 17191 24445
rect 13721 24440 17191 24442
rect 13721 24384 13726 24440
rect 13782 24384 15934 24440
rect 15990 24384 17130 24440
rect 17186 24384 17191 24440
rect 13721 24382 17191 24384
rect 13721 24379 13787 24382
rect 15929 24379 15995 24382
rect 17125 24379 17191 24382
rect 20110 24380 20116 24444
rect 20180 24442 20186 24444
rect 20253 24442 20319 24445
rect 20180 24440 20319 24442
rect 20180 24384 20258 24440
rect 20314 24384 20319 24440
rect 20180 24382 20319 24384
rect 20180 24380 20186 24382
rect 20253 24379 20319 24382
rect 24669 24442 24735 24445
rect 26509 24442 26575 24445
rect 24669 24440 26575 24442
rect 24669 24384 24674 24440
rect 24730 24384 26514 24440
rect 26570 24384 26575 24440
rect 24669 24382 26575 24384
rect 24669 24379 24735 24382
rect 26509 24379 26575 24382
rect 5533 24306 5599 24309
rect 11053 24306 11119 24309
rect 5533 24304 11119 24306
rect 5533 24248 5538 24304
rect 5594 24248 11058 24304
rect 11114 24248 11119 24304
rect 5533 24246 11119 24248
rect 5533 24243 5599 24246
rect 11053 24243 11119 24246
rect 15101 24306 15167 24309
rect 16941 24306 17007 24309
rect 19517 24306 19583 24309
rect 15101 24304 19583 24306
rect 15101 24248 15106 24304
rect 15162 24248 16946 24304
rect 17002 24248 19522 24304
rect 19578 24248 19583 24304
rect 15101 24246 19583 24248
rect 15101 24243 15167 24246
rect 16941 24243 17007 24246
rect 19517 24243 19583 24246
rect 20161 24306 20227 24309
rect 23197 24306 23263 24309
rect 20161 24304 25514 24306
rect 20161 24248 20166 24304
rect 20222 24248 23202 24304
rect 23258 24248 25514 24304
rect 20161 24246 25514 24248
rect 20161 24243 20227 24246
rect 23197 24243 23263 24246
rect 0 24170 480 24200
rect 933 24170 999 24173
rect 0 24168 999 24170
rect 0 24112 938 24168
rect 994 24112 999 24168
rect 0 24110 999 24112
rect 0 24080 480 24110
rect 933 24107 999 24110
rect 2221 24170 2287 24173
rect 5901 24170 5967 24173
rect 2221 24168 5967 24170
rect 2221 24112 2226 24168
rect 2282 24112 5906 24168
rect 5962 24112 5967 24168
rect 2221 24110 5967 24112
rect 2221 24107 2287 24110
rect 5901 24107 5967 24110
rect 6729 24170 6795 24173
rect 11513 24170 11579 24173
rect 6729 24168 11579 24170
rect 6729 24112 6734 24168
rect 6790 24112 11518 24168
rect 11574 24112 11579 24168
rect 6729 24110 11579 24112
rect 6729 24107 6795 24110
rect 11513 24107 11579 24110
rect 14825 24170 14891 24173
rect 16757 24170 16823 24173
rect 14825 24168 16823 24170
rect 14825 24112 14830 24168
rect 14886 24112 16762 24168
rect 16818 24112 16823 24168
rect 14825 24110 16823 24112
rect 14825 24107 14891 24110
rect 16757 24107 16823 24110
rect 17677 24170 17743 24173
rect 20897 24170 20963 24173
rect 17677 24168 20963 24170
rect 17677 24112 17682 24168
rect 17738 24112 20902 24168
rect 20958 24112 20963 24168
rect 17677 24110 20963 24112
rect 17677 24107 17743 24110
rect 20897 24107 20963 24110
rect 24117 24170 24183 24173
rect 25313 24170 25379 24173
rect 24117 24168 25379 24170
rect 24117 24112 24122 24168
rect 24178 24112 25318 24168
rect 25374 24112 25379 24168
rect 24117 24110 25379 24112
rect 25454 24170 25514 24246
rect 27520 24170 28000 24200
rect 25454 24110 28000 24170
rect 24117 24107 24183 24110
rect 25313 24107 25379 24110
rect 27520 24080 28000 24110
rect 2129 24034 2195 24037
rect 5165 24034 5231 24037
rect 2129 24032 5231 24034
rect 2129 23976 2134 24032
rect 2190 23976 5170 24032
rect 5226 23976 5231 24032
rect 2129 23974 5231 23976
rect 2129 23971 2195 23974
rect 5165 23971 5231 23974
rect 9029 24034 9095 24037
rect 10593 24034 10659 24037
rect 9029 24032 10659 24034
rect 9029 23976 9034 24032
rect 9090 23976 10598 24032
rect 10654 23976 10659 24032
rect 9029 23974 10659 23976
rect 9029 23971 9095 23974
rect 10593 23971 10659 23974
rect 18045 24034 18111 24037
rect 20345 24034 20411 24037
rect 18045 24032 20411 24034
rect 18045 23976 18050 24032
rect 18106 23976 20350 24032
rect 20406 23976 20411 24032
rect 18045 23974 20411 23976
rect 18045 23971 18111 23974
rect 20345 23971 20411 23974
rect 5610 23968 5930 23969
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5930 23968
rect 5610 23903 5930 23904
rect 14944 23968 15264 23969
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 23903 15264 23904
rect 24277 23968 24597 23969
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 23903 24597 23904
rect 6085 23898 6151 23901
rect 10685 23898 10751 23901
rect 6085 23896 10751 23898
rect 6085 23840 6090 23896
rect 6146 23840 10690 23896
rect 10746 23840 10751 23896
rect 6085 23838 10751 23840
rect 6085 23835 6151 23838
rect 10685 23835 10751 23838
rect 24761 23898 24827 23901
rect 27613 23898 27679 23901
rect 24761 23896 27679 23898
rect 24761 23840 24766 23896
rect 24822 23840 27618 23896
rect 27674 23840 27679 23896
rect 24761 23838 27679 23840
rect 24761 23835 24827 23838
rect 27613 23835 27679 23838
rect 3785 23762 3851 23765
rect 1350 23760 3851 23762
rect 1350 23704 3790 23760
rect 3846 23704 3851 23760
rect 1350 23702 3851 23704
rect 0 23626 480 23656
rect 1350 23626 1410 23702
rect 3785 23699 3851 23702
rect 7465 23762 7531 23765
rect 10869 23762 10935 23765
rect 7465 23760 10935 23762
rect 7465 23704 7470 23760
rect 7526 23704 10874 23760
rect 10930 23704 10935 23760
rect 7465 23702 10935 23704
rect 7465 23699 7531 23702
rect 10869 23699 10935 23702
rect 11513 23762 11579 23765
rect 12341 23762 12407 23765
rect 15193 23762 15259 23765
rect 22921 23762 22987 23765
rect 11513 23760 15259 23762
rect 11513 23704 11518 23760
rect 11574 23704 12346 23760
rect 12402 23704 15198 23760
rect 15254 23704 15259 23760
rect 11513 23702 15259 23704
rect 11513 23699 11579 23702
rect 12341 23699 12407 23702
rect 15193 23699 15259 23702
rect 15334 23760 22987 23762
rect 15334 23704 22926 23760
rect 22982 23704 22987 23760
rect 15334 23702 22987 23704
rect 0 23566 1410 23626
rect 9489 23626 9555 23629
rect 11237 23626 11303 23629
rect 9489 23624 11303 23626
rect 9489 23568 9494 23624
rect 9550 23568 11242 23624
rect 11298 23568 11303 23624
rect 9489 23566 11303 23568
rect 0 23536 480 23566
rect 9489 23563 9555 23566
rect 11237 23563 11303 23566
rect 14641 23626 14707 23629
rect 15334 23626 15394 23702
rect 22921 23699 22987 23702
rect 14641 23624 15394 23626
rect 14641 23568 14646 23624
rect 14702 23568 15394 23624
rect 14641 23566 15394 23568
rect 15929 23626 15995 23629
rect 21265 23626 21331 23629
rect 15929 23624 21331 23626
rect 15929 23568 15934 23624
rect 15990 23568 21270 23624
rect 21326 23568 21331 23624
rect 15929 23566 21331 23568
rect 14641 23563 14707 23566
rect 15929 23563 15995 23566
rect 21265 23563 21331 23566
rect 24761 23626 24827 23629
rect 27061 23626 27127 23629
rect 24761 23624 27127 23626
rect 24761 23568 24766 23624
rect 24822 23568 27066 23624
rect 27122 23568 27127 23624
rect 24761 23566 27127 23568
rect 24761 23563 24827 23566
rect 27061 23563 27127 23566
rect 27245 23626 27311 23629
rect 27520 23626 28000 23656
rect 27245 23624 28000 23626
rect 27245 23568 27250 23624
rect 27306 23568 28000 23624
rect 27245 23566 28000 23568
rect 27245 23563 27311 23566
rect 27520 23536 28000 23566
rect 3877 23490 3943 23493
rect 7005 23490 7071 23493
rect 3877 23488 7071 23490
rect 3877 23432 3882 23488
rect 3938 23432 7010 23488
rect 7066 23432 7071 23488
rect 3877 23430 7071 23432
rect 3877 23427 3943 23430
rect 7005 23427 7071 23430
rect 13169 23490 13235 23493
rect 18781 23490 18847 23493
rect 13169 23488 18847 23490
rect 13169 23432 13174 23488
rect 13230 23432 18786 23488
rect 18842 23432 18847 23488
rect 13169 23430 18847 23432
rect 13169 23427 13235 23430
rect 18781 23427 18847 23430
rect 20662 23428 20668 23492
rect 20732 23490 20738 23492
rect 24301 23490 24367 23493
rect 20732 23488 24367 23490
rect 20732 23432 24306 23488
rect 24362 23432 24367 23488
rect 20732 23430 24367 23432
rect 20732 23428 20738 23430
rect 24301 23427 24367 23430
rect 24485 23490 24551 23493
rect 24710 23490 24716 23492
rect 24485 23488 24716 23490
rect 24485 23432 24490 23488
rect 24546 23432 24716 23488
rect 24485 23430 24716 23432
rect 24485 23427 24551 23430
rect 24710 23428 24716 23430
rect 24780 23428 24786 23492
rect 10277 23424 10597 23425
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 10277 23359 10597 23360
rect 19610 23424 19930 23425
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 19610 23359 19930 23360
rect 2405 23354 2471 23357
rect 5073 23354 5139 23357
rect 2405 23352 5139 23354
rect 2405 23296 2410 23352
rect 2466 23296 5078 23352
rect 5134 23296 5139 23352
rect 2405 23294 5139 23296
rect 2405 23291 2471 23294
rect 5073 23291 5139 23294
rect 8477 23354 8543 23357
rect 9673 23354 9739 23357
rect 8477 23352 9739 23354
rect 8477 23296 8482 23352
rect 8538 23296 9678 23352
rect 9734 23296 9739 23352
rect 8477 23294 9739 23296
rect 8477 23291 8543 23294
rect 9673 23291 9739 23294
rect 11881 23354 11947 23357
rect 15469 23354 15535 23357
rect 17033 23354 17099 23357
rect 11881 23352 15535 23354
rect 11881 23296 11886 23352
rect 11942 23296 15474 23352
rect 15530 23296 15535 23352
rect 11881 23294 15535 23296
rect 11881 23291 11947 23294
rect 15469 23291 15535 23294
rect 15702 23352 17099 23354
rect 15702 23296 17038 23352
rect 17094 23296 17099 23352
rect 15702 23294 17099 23296
rect 2405 23218 2471 23221
rect 3417 23218 3483 23221
rect 2405 23216 3483 23218
rect 2405 23160 2410 23216
rect 2466 23160 3422 23216
rect 3478 23160 3483 23216
rect 2405 23158 3483 23160
rect 2405 23155 2471 23158
rect 3417 23155 3483 23158
rect 3693 23218 3759 23221
rect 5533 23218 5599 23221
rect 3693 23216 5599 23218
rect 3693 23160 3698 23216
rect 3754 23160 5538 23216
rect 5594 23160 5599 23216
rect 3693 23158 5599 23160
rect 3693 23155 3759 23158
rect 5533 23155 5599 23158
rect 9489 23218 9555 23221
rect 11145 23218 11211 23221
rect 12801 23218 12867 23221
rect 15702 23218 15762 23294
rect 17033 23291 17099 23294
rect 9489 23216 12867 23218
rect 9489 23160 9494 23216
rect 9550 23160 11150 23216
rect 11206 23160 12806 23216
rect 12862 23160 12867 23216
rect 9489 23158 12867 23160
rect 9489 23155 9555 23158
rect 11145 23155 11211 23158
rect 12801 23155 12867 23158
rect 14046 23158 15762 23218
rect 16573 23218 16639 23221
rect 19333 23218 19399 23221
rect 23473 23218 23539 23221
rect 16573 23216 23539 23218
rect 16573 23160 16578 23216
rect 16634 23160 19338 23216
rect 19394 23160 23478 23216
rect 23534 23160 23539 23216
rect 16573 23158 23539 23160
rect 0 23082 480 23112
rect 3325 23082 3391 23085
rect 0 23080 3391 23082
rect 0 23024 3330 23080
rect 3386 23024 3391 23080
rect 0 23022 3391 23024
rect 0 22992 480 23022
rect 3325 23019 3391 23022
rect 3601 23082 3667 23085
rect 8017 23082 8083 23085
rect 3601 23080 8083 23082
rect 3601 23024 3606 23080
rect 3662 23024 8022 23080
rect 8078 23024 8083 23080
rect 3601 23022 8083 23024
rect 3601 23019 3667 23022
rect 8017 23019 8083 23022
rect 11421 23082 11487 23085
rect 14046 23082 14106 23158
rect 16573 23155 16639 23158
rect 19333 23155 19399 23158
rect 23473 23155 23539 23158
rect 11421 23080 14106 23082
rect 11421 23024 11426 23080
rect 11482 23024 14106 23080
rect 11421 23022 14106 23024
rect 14273 23082 14339 23085
rect 17769 23082 17835 23085
rect 21541 23082 21607 23085
rect 14273 23080 17835 23082
rect 14273 23024 14278 23080
rect 14334 23024 17774 23080
rect 17830 23024 17835 23080
rect 14273 23022 17835 23024
rect 11421 23019 11487 23022
rect 14273 23019 14339 23022
rect 17769 23019 17835 23022
rect 17910 23080 21607 23082
rect 17910 23024 21546 23080
rect 21602 23024 21607 23080
rect 17910 23022 21607 23024
rect 15469 22946 15535 22949
rect 15929 22946 15995 22949
rect 15469 22944 15995 22946
rect 15469 22888 15474 22944
rect 15530 22888 15934 22944
rect 15990 22888 15995 22944
rect 15469 22886 15995 22888
rect 15469 22883 15535 22886
rect 15929 22883 15995 22886
rect 16665 22946 16731 22949
rect 17910 22946 17970 23022
rect 21541 23019 21607 23022
rect 21817 23082 21883 23085
rect 22829 23082 22895 23085
rect 21817 23080 22895 23082
rect 21817 23024 21822 23080
rect 21878 23024 22834 23080
rect 22890 23024 22895 23080
rect 21817 23022 22895 23024
rect 21817 23019 21883 23022
rect 22829 23019 22895 23022
rect 25405 23082 25471 23085
rect 27520 23082 28000 23112
rect 25405 23080 28000 23082
rect 25405 23024 25410 23080
rect 25466 23024 28000 23080
rect 25405 23022 28000 23024
rect 25405 23019 25471 23022
rect 27520 22992 28000 23022
rect 16665 22944 17970 22946
rect 16665 22888 16670 22944
rect 16726 22888 17970 22944
rect 16665 22886 17970 22888
rect 20161 22946 20227 22949
rect 23933 22946 23999 22949
rect 20161 22944 23999 22946
rect 20161 22888 20166 22944
rect 20222 22888 23938 22944
rect 23994 22888 23999 22944
rect 20161 22886 23999 22888
rect 16665 22883 16731 22886
rect 20161 22883 20227 22886
rect 23933 22883 23999 22886
rect 5610 22880 5930 22881
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5930 22880
rect 5610 22815 5930 22816
rect 14944 22880 15264 22881
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 22815 15264 22816
rect 24277 22880 24597 22881
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 22815 24597 22816
rect 4889 22810 4955 22813
rect 5022 22810 5028 22812
rect 4889 22808 5028 22810
rect 4889 22752 4894 22808
rect 4950 22752 5028 22808
rect 4889 22750 5028 22752
rect 4889 22747 4955 22750
rect 5022 22748 5028 22750
rect 5092 22748 5098 22812
rect 11053 22810 11119 22813
rect 6318 22808 11119 22810
rect 6318 22752 11058 22808
rect 11114 22752 11119 22808
rect 6318 22750 11119 22752
rect 4245 22674 4311 22677
rect 6318 22674 6378 22750
rect 11053 22747 11119 22750
rect 12249 22810 12315 22813
rect 15377 22810 15443 22813
rect 15510 22810 15516 22812
rect 12249 22808 14842 22810
rect 12249 22752 12254 22808
rect 12310 22752 14842 22808
rect 12249 22750 14842 22752
rect 12249 22747 12315 22750
rect 4245 22672 6378 22674
rect 4245 22616 4250 22672
rect 4306 22616 6378 22672
rect 4245 22614 6378 22616
rect 8753 22674 8819 22677
rect 14782 22674 14842 22750
rect 15377 22808 15516 22810
rect 15377 22752 15382 22808
rect 15438 22752 15516 22808
rect 15377 22750 15516 22752
rect 15377 22747 15443 22750
rect 15510 22748 15516 22750
rect 15580 22748 15586 22812
rect 17033 22810 17099 22813
rect 20069 22810 20135 22813
rect 17033 22808 20135 22810
rect 17033 22752 17038 22808
rect 17094 22752 20074 22808
rect 20130 22752 20135 22808
rect 17033 22750 20135 22752
rect 17033 22747 17099 22750
rect 20069 22747 20135 22750
rect 20345 22810 20411 22813
rect 20621 22810 20687 22813
rect 20345 22808 20687 22810
rect 20345 22752 20350 22808
rect 20406 22752 20626 22808
rect 20682 22752 20687 22808
rect 20345 22750 20687 22752
rect 20345 22747 20411 22750
rect 20621 22747 20687 22750
rect 21725 22810 21791 22813
rect 23105 22810 23171 22813
rect 21725 22808 23171 22810
rect 21725 22752 21730 22808
rect 21786 22752 23110 22808
rect 23166 22752 23171 22808
rect 21725 22750 23171 22752
rect 21725 22747 21791 22750
rect 23105 22747 23171 22750
rect 20897 22674 20963 22677
rect 23657 22674 23723 22677
rect 8753 22672 14704 22674
rect 8753 22616 8758 22672
rect 8814 22616 14704 22672
rect 8753 22614 14704 22616
rect 14782 22672 20963 22674
rect 14782 22616 20902 22672
rect 20958 22616 20963 22672
rect 14782 22614 20963 22616
rect 4245 22611 4311 22614
rect 8753 22611 8819 22614
rect 0 22538 480 22568
rect 3877 22538 3943 22541
rect 0 22536 3943 22538
rect 0 22480 3882 22536
rect 3938 22480 3943 22536
rect 0 22478 3943 22480
rect 0 22448 480 22478
rect 3877 22475 3943 22478
rect 6361 22538 6427 22541
rect 13261 22538 13327 22541
rect 6361 22536 13327 22538
rect 6361 22480 6366 22536
rect 6422 22480 13266 22536
rect 13322 22480 13327 22536
rect 6361 22478 13327 22480
rect 14644 22538 14704 22614
rect 20897 22611 20963 22614
rect 21222 22672 23723 22674
rect 21222 22616 23662 22672
rect 23718 22616 23723 22672
rect 21222 22614 23723 22616
rect 16849 22538 16915 22541
rect 14644 22536 16915 22538
rect 14644 22480 16854 22536
rect 16910 22480 16915 22536
rect 14644 22478 16915 22480
rect 6361 22475 6427 22478
rect 13261 22475 13327 22478
rect 16849 22475 16915 22478
rect 17718 22476 17724 22540
rect 17788 22538 17794 22540
rect 21222 22538 21282 22614
rect 23657 22611 23723 22614
rect 17788 22478 21282 22538
rect 24761 22538 24827 22541
rect 27520 22538 28000 22568
rect 24761 22536 28000 22538
rect 24761 22480 24766 22536
rect 24822 22480 28000 22536
rect 24761 22478 28000 22480
rect 17788 22476 17794 22478
rect 24761 22475 24827 22478
rect 27520 22448 28000 22478
rect 3325 22402 3391 22405
rect 9673 22402 9739 22405
rect 19241 22402 19307 22405
rect 3325 22400 9739 22402
rect 3325 22344 3330 22400
rect 3386 22344 9678 22400
rect 9734 22344 9739 22400
rect 3325 22342 9739 22344
rect 3325 22339 3391 22342
rect 9673 22339 9739 22342
rect 14414 22400 19307 22402
rect 14414 22344 19246 22400
rect 19302 22344 19307 22400
rect 14414 22342 19307 22344
rect 10277 22336 10597 22337
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 22271 10597 22272
rect 3509 22266 3575 22269
rect 5257 22266 5323 22269
rect 8477 22266 8543 22269
rect 3509 22264 5323 22266
rect 3509 22208 3514 22264
rect 3570 22208 5262 22264
rect 5318 22208 5323 22264
rect 3509 22206 5323 22208
rect 3509 22203 3575 22206
rect 5257 22203 5323 22206
rect 7054 22264 8543 22266
rect 7054 22208 8482 22264
rect 8538 22208 8543 22264
rect 7054 22206 8543 22208
rect 6361 22130 6427 22133
rect 7054 22130 7114 22206
rect 8477 22203 8543 22206
rect 13077 22266 13143 22269
rect 13721 22266 13787 22269
rect 14414 22266 14474 22342
rect 19241 22339 19307 22342
rect 20069 22402 20135 22405
rect 21081 22402 21147 22405
rect 20069 22400 21147 22402
rect 20069 22344 20074 22400
rect 20130 22344 21086 22400
rect 21142 22344 21147 22400
rect 20069 22342 21147 22344
rect 20069 22339 20135 22342
rect 21081 22339 21147 22342
rect 19610 22336 19930 22337
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 22271 19930 22272
rect 13077 22264 14474 22266
rect 13077 22208 13082 22264
rect 13138 22208 13726 22264
rect 13782 22208 14474 22264
rect 13077 22206 14474 22208
rect 15929 22266 15995 22269
rect 16481 22266 16547 22269
rect 24025 22266 24091 22269
rect 15929 22264 16547 22266
rect 15929 22208 15934 22264
rect 15990 22208 16486 22264
rect 16542 22208 16547 22264
rect 15929 22206 16547 22208
rect 13077 22203 13143 22206
rect 13721 22203 13787 22206
rect 15929 22203 15995 22206
rect 16481 22203 16547 22206
rect 20118 22264 24091 22266
rect 20118 22208 24030 22264
rect 24086 22208 24091 22264
rect 20118 22206 24091 22208
rect 6361 22128 7114 22130
rect 6361 22072 6366 22128
rect 6422 22072 7114 22128
rect 6361 22070 7114 22072
rect 7189 22130 7255 22133
rect 11145 22130 11211 22133
rect 7189 22128 11211 22130
rect 7189 22072 7194 22128
rect 7250 22072 11150 22128
rect 11206 22072 11211 22128
rect 7189 22070 11211 22072
rect 6361 22067 6427 22070
rect 7189 22067 7255 22070
rect 11145 22067 11211 22070
rect 12985 22130 13051 22133
rect 20118 22130 20178 22206
rect 24025 22203 24091 22206
rect 12985 22128 20178 22130
rect 12985 22072 12990 22128
rect 13046 22072 20178 22128
rect 12985 22070 20178 22072
rect 20621 22130 20687 22133
rect 23933 22130 23999 22133
rect 20621 22128 23999 22130
rect 20621 22072 20626 22128
rect 20682 22072 23938 22128
rect 23994 22072 23999 22128
rect 20621 22070 23999 22072
rect 12985 22067 13051 22070
rect 20621 22067 20687 22070
rect 23933 22067 23999 22070
rect 2313 21994 2379 21997
rect 9857 21994 9923 21997
rect 2313 21992 9923 21994
rect 2313 21936 2318 21992
rect 2374 21936 9862 21992
rect 9918 21936 9923 21992
rect 2313 21934 9923 21936
rect 2313 21931 2379 21934
rect 9857 21931 9923 21934
rect 14641 21994 14707 21997
rect 16665 21994 16731 21997
rect 14641 21992 16731 21994
rect 14641 21936 14646 21992
rect 14702 21936 16670 21992
rect 16726 21936 16731 21992
rect 14641 21934 16731 21936
rect 14641 21931 14707 21934
rect 16665 21931 16731 21934
rect 18413 21994 18479 21997
rect 25313 21994 25379 21997
rect 18413 21992 25379 21994
rect 18413 21936 18418 21992
rect 18474 21936 25318 21992
rect 25374 21936 25379 21992
rect 18413 21934 25379 21936
rect 18413 21931 18479 21934
rect 25313 21931 25379 21934
rect 0 21858 480 21888
rect 3969 21858 4035 21861
rect 0 21856 4035 21858
rect 0 21800 3974 21856
rect 4030 21800 4035 21856
rect 0 21798 4035 21800
rect 0 21768 480 21798
rect 3969 21795 4035 21798
rect 21030 21796 21036 21860
rect 21100 21858 21106 21860
rect 22645 21858 22711 21861
rect 21100 21856 22711 21858
rect 21100 21800 22650 21856
rect 22706 21800 22711 21856
rect 21100 21798 22711 21800
rect 21100 21796 21106 21798
rect 22645 21795 22711 21798
rect 25497 21858 25563 21861
rect 27520 21858 28000 21888
rect 25497 21856 28000 21858
rect 25497 21800 25502 21856
rect 25558 21800 28000 21856
rect 25497 21798 28000 21800
rect 25497 21795 25563 21798
rect 5610 21792 5930 21793
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5930 21792
rect 5610 21727 5930 21728
rect 14944 21792 15264 21793
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 21727 15264 21728
rect 24277 21792 24597 21793
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 27520 21768 28000 21798
rect 24277 21727 24597 21728
rect 2405 21722 2471 21725
rect 4521 21722 4587 21725
rect 2405 21720 4587 21722
rect 2405 21664 2410 21720
rect 2466 21664 4526 21720
rect 4582 21664 4587 21720
rect 2405 21662 4587 21664
rect 2405 21659 2471 21662
rect 4521 21659 4587 21662
rect 7649 21722 7715 21725
rect 8569 21722 8635 21725
rect 12525 21722 12591 21725
rect 23381 21722 23447 21725
rect 7649 21720 12591 21722
rect 7649 21664 7654 21720
rect 7710 21664 8574 21720
rect 8630 21664 12530 21720
rect 12586 21664 12591 21720
rect 7649 21662 12591 21664
rect 7649 21659 7715 21662
rect 8569 21659 8635 21662
rect 12525 21659 12591 21662
rect 15334 21720 23447 21722
rect 15334 21664 23386 21720
rect 23442 21664 23447 21720
rect 15334 21662 23447 21664
rect 2497 21586 2563 21589
rect 2630 21586 2636 21588
rect 2497 21584 2636 21586
rect 2497 21528 2502 21584
rect 2558 21528 2636 21584
rect 2497 21526 2636 21528
rect 2497 21523 2563 21526
rect 2630 21524 2636 21526
rect 2700 21524 2706 21588
rect 5165 21586 5231 21589
rect 8569 21586 8635 21589
rect 12341 21586 12407 21589
rect 5165 21584 12407 21586
rect 5165 21528 5170 21584
rect 5226 21528 8574 21584
rect 8630 21528 12346 21584
rect 12402 21528 12407 21584
rect 5165 21526 12407 21528
rect 2638 21450 2698 21524
rect 5165 21523 5231 21526
rect 8569 21523 8635 21526
rect 12341 21523 12407 21526
rect 14365 21586 14431 21589
rect 15334 21586 15394 21662
rect 23381 21659 23447 21662
rect 21766 21586 21772 21588
rect 14365 21584 15394 21586
rect 14365 21528 14370 21584
rect 14426 21528 15394 21584
rect 14365 21526 15394 21528
rect 16990 21526 21772 21586
rect 14365 21523 14431 21526
rect 9121 21450 9187 21453
rect 9254 21450 9260 21452
rect 2638 21390 3434 21450
rect 0 21314 480 21344
rect 3233 21314 3299 21317
rect 0 21312 3299 21314
rect 0 21256 3238 21312
rect 3294 21256 3299 21312
rect 0 21254 3299 21256
rect 0 21224 480 21254
rect 3233 21251 3299 21254
rect 3374 21042 3434 21390
rect 9121 21448 9260 21450
rect 9121 21392 9126 21448
rect 9182 21392 9260 21448
rect 9121 21390 9260 21392
rect 9121 21387 9187 21390
rect 9254 21388 9260 21390
rect 9324 21388 9330 21452
rect 3509 21314 3575 21317
rect 9673 21314 9739 21317
rect 16990 21314 17050 21526
rect 21766 21524 21772 21526
rect 21836 21524 21842 21588
rect 21909 21586 21975 21589
rect 21909 21584 22018 21586
rect 21909 21528 21914 21584
rect 21970 21528 22018 21584
rect 21909 21523 22018 21528
rect 18045 21450 18111 21453
rect 19701 21450 19767 21453
rect 18045 21448 19767 21450
rect 18045 21392 18050 21448
rect 18106 21392 19706 21448
rect 19762 21392 19767 21448
rect 18045 21390 19767 21392
rect 18045 21387 18111 21390
rect 19701 21387 19767 21390
rect 21265 21450 21331 21453
rect 21958 21450 22018 21523
rect 21265 21448 22018 21450
rect 21265 21392 21270 21448
rect 21326 21392 22018 21448
rect 21265 21390 22018 21392
rect 21265 21387 21331 21390
rect 3509 21312 9739 21314
rect 3509 21256 3514 21312
rect 3570 21256 9678 21312
rect 9734 21256 9739 21312
rect 3509 21254 9739 21256
rect 3509 21251 3575 21254
rect 9673 21251 9739 21254
rect 10734 21254 17050 21314
rect 24669 21314 24735 21317
rect 27520 21314 28000 21344
rect 24669 21312 28000 21314
rect 24669 21256 24674 21312
rect 24730 21256 28000 21312
rect 24669 21254 28000 21256
rect 10277 21248 10597 21249
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 21183 10597 21184
rect 8385 21178 8451 21181
rect 10133 21178 10199 21181
rect 8385 21176 10199 21178
rect 8385 21120 8390 21176
rect 8446 21120 10138 21176
rect 10194 21120 10199 21176
rect 8385 21118 10199 21120
rect 8385 21115 8451 21118
rect 10133 21115 10199 21118
rect 10734 21042 10794 21254
rect 24669 21251 24735 21254
rect 19610 21248 19930 21249
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 27520 21224 28000 21254
rect 19610 21183 19930 21184
rect 12249 21178 12315 21181
rect 17309 21178 17375 21181
rect 19333 21178 19399 21181
rect 12249 21176 19399 21178
rect 12249 21120 12254 21176
rect 12310 21120 17314 21176
rect 17370 21120 19338 21176
rect 19394 21120 19399 21176
rect 12249 21118 19399 21120
rect 12249 21115 12315 21118
rect 17309 21115 17375 21118
rect 19333 21115 19399 21118
rect 3374 20982 10794 21042
rect 11053 21042 11119 21045
rect 12617 21042 12683 21045
rect 21081 21042 21147 21045
rect 11053 21040 12683 21042
rect 11053 20984 11058 21040
rect 11114 20984 12622 21040
rect 12678 20984 12683 21040
rect 11053 20982 12683 20984
rect 11053 20979 11119 20982
rect 12617 20979 12683 20982
rect 14046 21040 21147 21042
rect 14046 20984 21086 21040
rect 21142 20984 21147 21040
rect 14046 20982 21147 20984
rect 2078 20844 2084 20908
rect 2148 20906 2154 20908
rect 6913 20906 6979 20909
rect 2148 20904 6979 20906
rect 2148 20848 6918 20904
rect 6974 20848 6979 20904
rect 2148 20846 6979 20848
rect 2148 20844 2154 20846
rect 6913 20843 6979 20846
rect 7649 20906 7715 20909
rect 9213 20906 9279 20909
rect 11605 20906 11671 20909
rect 7649 20904 11671 20906
rect 7649 20848 7654 20904
rect 7710 20848 9218 20904
rect 9274 20848 11610 20904
rect 11666 20848 11671 20904
rect 7649 20846 11671 20848
rect 7649 20843 7715 20846
rect 9213 20843 9279 20846
rect 11605 20843 11671 20846
rect 12617 20906 12683 20909
rect 14046 20906 14106 20982
rect 21081 20979 21147 20982
rect 12617 20904 14106 20906
rect 12617 20848 12622 20904
rect 12678 20848 14106 20904
rect 12617 20846 14106 20848
rect 14273 20906 14339 20909
rect 15653 20906 15719 20909
rect 14273 20904 15719 20906
rect 14273 20848 14278 20904
rect 14334 20848 15658 20904
rect 15714 20848 15719 20904
rect 14273 20846 15719 20848
rect 12617 20843 12683 20846
rect 14273 20843 14339 20846
rect 15653 20843 15719 20846
rect 0 20770 480 20800
rect 2681 20770 2747 20773
rect 0 20768 2747 20770
rect 0 20712 2686 20768
rect 2742 20712 2747 20768
rect 0 20710 2747 20712
rect 0 20680 480 20710
rect 2681 20707 2747 20710
rect 5257 20770 5323 20773
rect 5390 20770 5396 20772
rect 5257 20768 5396 20770
rect 5257 20712 5262 20768
rect 5318 20712 5396 20768
rect 5257 20710 5396 20712
rect 5257 20707 5323 20710
rect 5390 20708 5396 20710
rect 5460 20708 5466 20772
rect 6545 20770 6611 20773
rect 12065 20770 12131 20773
rect 19977 20770 20043 20773
rect 6545 20768 12131 20770
rect 6545 20712 6550 20768
rect 6606 20712 12070 20768
rect 12126 20712 12131 20768
rect 6545 20710 12131 20712
rect 6545 20707 6611 20710
rect 12065 20707 12131 20710
rect 15334 20768 20043 20770
rect 15334 20712 19982 20768
rect 20038 20712 20043 20768
rect 15334 20710 20043 20712
rect 5610 20704 5930 20705
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5930 20704
rect 5610 20639 5930 20640
rect 14944 20704 15264 20705
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14944 20639 15264 20640
rect 2313 20634 2379 20637
rect 4245 20634 4311 20637
rect 2313 20632 4311 20634
rect 2313 20576 2318 20632
rect 2374 20576 4250 20632
rect 4306 20576 4311 20632
rect 2313 20574 4311 20576
rect 2313 20571 2379 20574
rect 4245 20571 4311 20574
rect 6821 20634 6887 20637
rect 14181 20634 14247 20637
rect 6821 20632 14247 20634
rect 6821 20576 6826 20632
rect 6882 20576 14186 20632
rect 14242 20576 14247 20632
rect 6821 20574 14247 20576
rect 6821 20571 6887 20574
rect 14181 20571 14247 20574
rect 3601 20498 3667 20501
rect 6821 20498 6887 20501
rect 3601 20496 6887 20498
rect 3601 20440 3606 20496
rect 3662 20440 6826 20496
rect 6882 20440 6887 20496
rect 3601 20438 6887 20440
rect 3601 20435 3667 20438
rect 6821 20435 6887 20438
rect 7097 20498 7163 20501
rect 13353 20498 13419 20501
rect 14917 20498 14983 20501
rect 7097 20496 12450 20498
rect 7097 20440 7102 20496
rect 7158 20440 12450 20496
rect 7097 20438 12450 20440
rect 7097 20435 7163 20438
rect 2405 20362 2471 20365
rect 5717 20362 5783 20365
rect 2405 20360 5783 20362
rect 2405 20304 2410 20360
rect 2466 20304 5722 20360
rect 5778 20304 5783 20360
rect 2405 20302 5783 20304
rect 12390 20362 12450 20438
rect 13353 20496 14983 20498
rect 13353 20440 13358 20496
rect 13414 20440 14922 20496
rect 14978 20440 14983 20496
rect 13353 20438 14983 20440
rect 13353 20435 13419 20438
rect 14917 20435 14983 20438
rect 15101 20498 15167 20501
rect 15334 20498 15394 20710
rect 19977 20707 20043 20710
rect 21633 20770 21699 20773
rect 23933 20770 23999 20773
rect 21633 20768 23999 20770
rect 21633 20712 21638 20768
rect 21694 20712 23938 20768
rect 23994 20712 23999 20768
rect 21633 20710 23999 20712
rect 21633 20707 21699 20710
rect 23933 20707 23999 20710
rect 25405 20770 25471 20773
rect 27520 20770 28000 20800
rect 25405 20768 28000 20770
rect 25405 20712 25410 20768
rect 25466 20712 28000 20768
rect 25405 20710 28000 20712
rect 25405 20707 25471 20710
rect 24277 20704 24597 20705
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 27520 20680 28000 20710
rect 24277 20639 24597 20640
rect 15469 20634 15535 20637
rect 23473 20634 23539 20637
rect 15469 20632 23539 20634
rect 15469 20576 15474 20632
rect 15530 20576 23478 20632
rect 23534 20576 23539 20632
rect 15469 20574 23539 20576
rect 15469 20571 15535 20574
rect 23473 20571 23539 20574
rect 15101 20496 15394 20498
rect 15101 20440 15106 20496
rect 15162 20440 15394 20496
rect 15101 20438 15394 20440
rect 16757 20498 16823 20501
rect 20897 20498 20963 20501
rect 16757 20496 20963 20498
rect 16757 20440 16762 20496
rect 16818 20440 20902 20496
rect 20958 20440 20963 20496
rect 16757 20438 20963 20440
rect 15101 20435 15167 20438
rect 16757 20435 16823 20438
rect 20897 20435 20963 20438
rect 21081 20498 21147 20501
rect 25589 20498 25655 20501
rect 21081 20496 25655 20498
rect 21081 20440 21086 20496
rect 21142 20440 25594 20496
rect 25650 20440 25655 20496
rect 21081 20438 25655 20440
rect 21081 20435 21147 20438
rect 25589 20435 25655 20438
rect 14365 20362 14431 20365
rect 12390 20360 14431 20362
rect 12390 20304 14370 20360
rect 14426 20304 14431 20360
rect 12390 20302 14431 20304
rect 2405 20299 2471 20302
rect 5717 20299 5783 20302
rect 14365 20299 14431 20302
rect 14774 20300 14780 20364
rect 14844 20362 14850 20364
rect 17769 20362 17835 20365
rect 18873 20362 18939 20365
rect 20529 20362 20595 20365
rect 14844 20360 18939 20362
rect 14844 20304 17774 20360
rect 17830 20304 18878 20360
rect 18934 20304 18939 20360
rect 14844 20302 18939 20304
rect 14844 20300 14850 20302
rect 17769 20299 17835 20302
rect 18873 20299 18939 20302
rect 19382 20360 20595 20362
rect 19382 20304 20534 20360
rect 20590 20304 20595 20360
rect 19382 20302 20595 20304
rect 4337 20226 4403 20229
rect 9673 20226 9739 20229
rect 10869 20228 10935 20229
rect 10869 20226 10916 20228
rect 4337 20224 9739 20226
rect 4337 20168 4342 20224
rect 4398 20168 9678 20224
rect 9734 20168 9739 20224
rect 4337 20166 9739 20168
rect 10824 20224 10916 20226
rect 10824 20168 10874 20224
rect 10824 20166 10916 20168
rect 4337 20163 4403 20166
rect 9673 20163 9739 20166
rect 10869 20164 10916 20166
rect 10980 20164 10986 20228
rect 12065 20226 12131 20229
rect 12525 20226 12591 20229
rect 17217 20226 17283 20229
rect 12065 20224 17283 20226
rect 12065 20168 12070 20224
rect 12126 20168 12530 20224
rect 12586 20168 17222 20224
rect 17278 20168 17283 20224
rect 12065 20166 17283 20168
rect 10869 20163 10935 20164
rect 12065 20163 12131 20166
rect 12525 20163 12591 20166
rect 17217 20163 17283 20166
rect 17493 20226 17559 20229
rect 19382 20226 19442 20302
rect 20529 20299 20595 20302
rect 21633 20362 21699 20365
rect 22461 20362 22527 20365
rect 21633 20360 22527 20362
rect 21633 20304 21638 20360
rect 21694 20304 22466 20360
rect 22522 20304 22527 20360
rect 21633 20302 22527 20304
rect 21633 20299 21699 20302
rect 22461 20299 22527 20302
rect 17493 20224 19442 20226
rect 17493 20168 17498 20224
rect 17554 20168 19442 20224
rect 17493 20166 19442 20168
rect 20897 20226 20963 20229
rect 25037 20226 25103 20229
rect 20897 20224 25103 20226
rect 20897 20168 20902 20224
rect 20958 20168 25042 20224
rect 25098 20168 25103 20224
rect 20897 20166 25103 20168
rect 17493 20163 17559 20166
rect 20897 20163 20963 20166
rect 25037 20163 25103 20166
rect 10277 20160 10597 20161
rect 0 20090 480 20120
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 10277 20095 10597 20096
rect 19610 20160 19930 20161
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 19610 20095 19930 20096
rect 1393 20090 1459 20093
rect 0 20088 1459 20090
rect 0 20032 1398 20088
rect 1454 20032 1459 20088
rect 0 20030 1459 20032
rect 0 20000 480 20030
rect 1393 20027 1459 20030
rect 2865 20090 2931 20093
rect 6361 20090 6427 20093
rect 7189 20090 7255 20093
rect 2865 20088 7255 20090
rect 2865 20032 2870 20088
rect 2926 20032 6366 20088
rect 6422 20032 7194 20088
rect 7250 20032 7255 20088
rect 2865 20030 7255 20032
rect 2865 20027 2931 20030
rect 6361 20027 6427 20030
rect 7189 20027 7255 20030
rect 13261 20090 13327 20093
rect 15193 20090 15259 20093
rect 13261 20088 15259 20090
rect 13261 20032 13266 20088
rect 13322 20032 15198 20088
rect 15254 20032 15259 20088
rect 13261 20030 15259 20032
rect 13261 20027 13327 20030
rect 15193 20027 15259 20030
rect 17677 20092 17743 20093
rect 17677 20088 17724 20092
rect 17788 20090 17794 20092
rect 24761 20090 24827 20093
rect 27520 20090 28000 20120
rect 17677 20032 17682 20088
rect 17677 20028 17724 20032
rect 17788 20030 17834 20090
rect 24761 20088 28000 20090
rect 24761 20032 24766 20088
rect 24822 20032 28000 20088
rect 24761 20030 28000 20032
rect 17788 20028 17794 20030
rect 17677 20027 17743 20028
rect 24761 20027 24827 20030
rect 27520 20000 28000 20030
rect 4061 19954 4127 19957
rect 12157 19954 12223 19957
rect 4061 19952 12223 19954
rect 4061 19896 4066 19952
rect 4122 19896 12162 19952
rect 12218 19896 12223 19952
rect 4061 19894 12223 19896
rect 4061 19891 4127 19894
rect 12157 19891 12223 19894
rect 16849 19954 16915 19957
rect 25221 19954 25287 19957
rect 16849 19952 25287 19954
rect 16849 19896 16854 19952
rect 16910 19896 25226 19952
rect 25282 19896 25287 19952
rect 16849 19894 25287 19896
rect 16849 19891 16915 19894
rect 25221 19891 25287 19894
rect 3141 19818 3207 19821
rect 7465 19818 7531 19821
rect 3141 19816 7531 19818
rect 3141 19760 3146 19816
rect 3202 19760 7470 19816
rect 7526 19760 7531 19816
rect 3141 19758 7531 19760
rect 3141 19755 3207 19758
rect 7465 19755 7531 19758
rect 10317 19818 10383 19821
rect 13077 19818 13143 19821
rect 10317 19816 13143 19818
rect 10317 19760 10322 19816
rect 10378 19760 13082 19816
rect 13138 19760 13143 19816
rect 10317 19758 13143 19760
rect 10317 19755 10383 19758
rect 13077 19755 13143 19758
rect 13997 19818 14063 19821
rect 16481 19818 16547 19821
rect 18045 19818 18111 19821
rect 13997 19816 15394 19818
rect 13997 19760 14002 19816
rect 14058 19760 15394 19816
rect 13997 19758 15394 19760
rect 13997 19755 14063 19758
rect 8661 19682 8727 19685
rect 8845 19682 8911 19685
rect 8661 19680 10196 19682
rect 8661 19624 8666 19680
rect 8722 19624 8850 19680
rect 8906 19624 10196 19680
rect 8661 19622 10196 19624
rect 8661 19619 8727 19622
rect 8845 19619 8911 19622
rect 5610 19616 5930 19617
rect 0 19546 480 19576
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5930 19616
rect 5610 19551 5930 19552
rect 8937 19546 9003 19549
rect 9070 19546 9076 19548
rect 0 19486 5458 19546
rect 0 19456 480 19486
rect 2405 19410 2471 19413
rect 4613 19410 4679 19413
rect 2405 19408 4679 19410
rect 2405 19352 2410 19408
rect 2466 19352 4618 19408
rect 4674 19352 4679 19408
rect 2405 19350 4679 19352
rect 5398 19410 5458 19486
rect 8937 19544 9076 19546
rect 8937 19488 8942 19544
rect 8998 19488 9076 19544
rect 8937 19486 9076 19488
rect 8937 19483 9003 19486
rect 9070 19484 9076 19486
rect 9140 19484 9146 19548
rect 10136 19546 10196 19622
rect 10726 19620 10732 19684
rect 10796 19682 10802 19684
rect 12893 19682 12959 19685
rect 10796 19680 12959 19682
rect 10796 19624 12898 19680
rect 12954 19624 12959 19680
rect 10796 19622 12959 19624
rect 10796 19620 10802 19622
rect 12893 19619 12959 19622
rect 14944 19616 15264 19617
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14944 19551 15264 19552
rect 14774 19546 14780 19548
rect 10136 19486 14780 19546
rect 14774 19484 14780 19486
rect 14844 19484 14850 19548
rect 15334 19546 15394 19758
rect 16481 19816 18111 19818
rect 16481 19760 16486 19816
rect 16542 19760 18050 19816
rect 18106 19760 18111 19816
rect 16481 19758 18111 19760
rect 16481 19755 16547 19758
rect 18045 19755 18111 19758
rect 19977 19818 20043 19821
rect 20110 19818 20116 19820
rect 19977 19816 20116 19818
rect 19977 19760 19982 19816
rect 20038 19760 20116 19816
rect 19977 19758 20116 19760
rect 19977 19755 20043 19758
rect 20110 19756 20116 19758
rect 20180 19756 20186 19820
rect 15561 19682 15627 19685
rect 21633 19682 21699 19685
rect 15561 19680 21699 19682
rect 15561 19624 15566 19680
rect 15622 19624 21638 19680
rect 21694 19624 21699 19680
rect 15561 19622 21699 19624
rect 15561 19619 15627 19622
rect 21633 19619 21699 19622
rect 24277 19616 24597 19617
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 19551 24597 19552
rect 22277 19546 22343 19549
rect 15334 19544 22343 19546
rect 15334 19488 22282 19544
rect 22338 19488 22343 19544
rect 15334 19486 22343 19488
rect 22277 19483 22343 19486
rect 24669 19546 24735 19549
rect 27520 19546 28000 19576
rect 24669 19544 28000 19546
rect 24669 19488 24674 19544
rect 24730 19488 28000 19544
rect 24669 19486 28000 19488
rect 24669 19483 24735 19486
rect 27520 19456 28000 19486
rect 9857 19410 9923 19413
rect 5398 19408 9923 19410
rect 5398 19352 9862 19408
rect 9918 19352 9923 19408
rect 5398 19350 9923 19352
rect 2405 19347 2471 19350
rect 4613 19347 4679 19350
rect 9857 19347 9923 19350
rect 10225 19410 10291 19413
rect 25037 19410 25103 19413
rect 10225 19408 25103 19410
rect 10225 19352 10230 19408
rect 10286 19352 25042 19408
rect 25098 19352 25103 19408
rect 10225 19350 25103 19352
rect 10225 19347 10291 19350
rect 25037 19347 25103 19350
rect 2129 19274 2195 19277
rect 2262 19274 2268 19276
rect 2129 19272 2268 19274
rect 2129 19216 2134 19272
rect 2190 19216 2268 19272
rect 2129 19214 2268 19216
rect 2129 19211 2195 19214
rect 2262 19212 2268 19214
rect 2332 19212 2338 19276
rect 3049 19274 3115 19277
rect 10317 19274 10383 19277
rect 3049 19272 10383 19274
rect 3049 19216 3054 19272
rect 3110 19216 10322 19272
rect 10378 19216 10383 19272
rect 3049 19214 10383 19216
rect 3049 19211 3115 19214
rect 10317 19211 10383 19214
rect 12525 19274 12591 19277
rect 15653 19274 15719 19277
rect 16941 19274 17007 19277
rect 23657 19274 23723 19277
rect 12525 19272 16866 19274
rect 12525 19216 12530 19272
rect 12586 19216 15658 19272
rect 15714 19216 16866 19272
rect 12525 19214 16866 19216
rect 12525 19211 12591 19214
rect 15653 19211 15719 19214
rect 12934 19076 12940 19140
rect 13004 19138 13010 19140
rect 15929 19138 15995 19141
rect 13004 19136 15995 19138
rect 13004 19080 15934 19136
rect 15990 19080 15995 19136
rect 13004 19078 15995 19080
rect 16806 19138 16866 19214
rect 16941 19272 23723 19274
rect 16941 19216 16946 19272
rect 17002 19216 23662 19272
rect 23718 19216 23723 19272
rect 16941 19214 23723 19216
rect 16941 19211 17007 19214
rect 23657 19211 23723 19214
rect 17493 19138 17559 19141
rect 19425 19140 19491 19141
rect 16806 19136 17559 19138
rect 16806 19080 17498 19136
rect 17554 19080 17559 19136
rect 16806 19078 17559 19080
rect 13004 19076 13010 19078
rect 15929 19075 15995 19078
rect 17493 19075 17559 19078
rect 19374 19076 19380 19140
rect 19444 19138 19491 19140
rect 19444 19136 19536 19138
rect 19486 19080 19536 19136
rect 19444 19078 19536 19080
rect 19444 19076 19491 19078
rect 20294 19076 20300 19140
rect 20364 19138 20370 19140
rect 20621 19138 20687 19141
rect 23790 19138 23796 19140
rect 20364 19136 23796 19138
rect 20364 19080 20626 19136
rect 20682 19080 23796 19136
rect 20364 19078 23796 19080
rect 20364 19076 20370 19078
rect 19425 19075 19491 19076
rect 20621 19075 20687 19078
rect 23790 19076 23796 19078
rect 23860 19076 23866 19140
rect 10277 19072 10597 19073
rect 0 19002 480 19032
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 19007 10597 19008
rect 19610 19072 19930 19073
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 19007 19930 19008
rect 2957 19002 3023 19005
rect 0 19000 3023 19002
rect 0 18944 2962 19000
rect 3018 18944 3023 19000
rect 0 18942 3023 18944
rect 0 18912 480 18942
rect 2957 18939 3023 18942
rect 11697 19002 11763 19005
rect 25589 19002 25655 19005
rect 27520 19002 28000 19032
rect 11697 19000 19442 19002
rect 11697 18944 11702 19000
rect 11758 18944 19442 19000
rect 11697 18942 19442 18944
rect 11697 18939 11763 18942
rect 3877 18866 3943 18869
rect 6637 18866 6703 18869
rect 3877 18864 6703 18866
rect 3877 18808 3882 18864
rect 3938 18808 6642 18864
rect 6698 18808 6703 18864
rect 3877 18806 6703 18808
rect 3877 18803 3943 18806
rect 6637 18803 6703 18806
rect 7741 18866 7807 18869
rect 18413 18866 18479 18869
rect 7741 18864 18479 18866
rect 7741 18808 7746 18864
rect 7802 18808 18418 18864
rect 18474 18808 18479 18864
rect 7741 18806 18479 18808
rect 19382 18866 19442 18942
rect 25589 19000 28000 19002
rect 25589 18944 25594 19000
rect 25650 18944 28000 19000
rect 25589 18942 28000 18944
rect 25589 18939 25655 18942
rect 27520 18912 28000 18942
rect 21357 18866 21423 18869
rect 19382 18864 21423 18866
rect 19382 18808 21362 18864
rect 21418 18808 21423 18864
rect 19382 18806 21423 18808
rect 7741 18803 7807 18806
rect 18413 18803 18479 18806
rect 21357 18803 21423 18806
rect 7005 18730 7071 18733
rect 5352 18728 7071 18730
rect 5352 18672 7010 18728
rect 7066 18672 7071 18728
rect 5352 18670 7071 18672
rect 0 18458 480 18488
rect 5352 18458 5412 18670
rect 7005 18667 7071 18670
rect 7465 18730 7531 18733
rect 12433 18730 12499 18733
rect 7465 18728 12499 18730
rect 7465 18672 7470 18728
rect 7526 18672 12438 18728
rect 12494 18672 12499 18728
rect 7465 18670 12499 18672
rect 7465 18667 7531 18670
rect 12433 18667 12499 18670
rect 17769 18730 17835 18733
rect 20897 18730 20963 18733
rect 17769 18728 20963 18730
rect 17769 18672 17774 18728
rect 17830 18672 20902 18728
rect 20958 18672 20963 18728
rect 17769 18670 20963 18672
rect 17769 18667 17835 18670
rect 20897 18667 20963 18670
rect 15837 18594 15903 18597
rect 23197 18594 23263 18597
rect 15837 18592 23263 18594
rect 15837 18536 15842 18592
rect 15898 18536 23202 18592
rect 23258 18536 23263 18592
rect 15837 18534 23263 18536
rect 15837 18531 15903 18534
rect 23197 18531 23263 18534
rect 5610 18528 5930 18529
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5930 18528
rect 5610 18463 5930 18464
rect 14944 18528 15264 18529
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 18463 15264 18464
rect 24277 18528 24597 18529
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 18463 24597 18464
rect 0 18398 5412 18458
rect 7097 18458 7163 18461
rect 12525 18458 12591 18461
rect 14733 18458 14799 18461
rect 7097 18456 12450 18458
rect 7097 18400 7102 18456
rect 7158 18400 12450 18456
rect 7097 18398 12450 18400
rect 0 18368 480 18398
rect 7097 18395 7163 18398
rect 8201 18322 8267 18325
rect 9949 18322 10015 18325
rect 8201 18320 10015 18322
rect 8201 18264 8206 18320
rect 8262 18264 9954 18320
rect 10010 18264 10015 18320
rect 8201 18262 10015 18264
rect 12390 18322 12450 18398
rect 12525 18456 14799 18458
rect 12525 18400 12530 18456
rect 12586 18400 14738 18456
rect 14794 18400 14799 18456
rect 12525 18398 14799 18400
rect 12525 18395 12591 18398
rect 14733 18395 14799 18398
rect 15653 18458 15719 18461
rect 16481 18458 16547 18461
rect 15653 18456 16547 18458
rect 15653 18400 15658 18456
rect 15714 18400 16486 18456
rect 16542 18400 16547 18456
rect 15653 18398 16547 18400
rect 15653 18395 15719 18398
rect 16481 18395 16547 18398
rect 17309 18458 17375 18461
rect 19517 18458 19583 18461
rect 27520 18458 28000 18488
rect 17309 18456 19583 18458
rect 17309 18400 17314 18456
rect 17370 18400 19522 18456
rect 19578 18400 19583 18456
rect 17309 18398 19583 18400
rect 17309 18395 17375 18398
rect 19517 18395 19583 18398
rect 24718 18398 28000 18458
rect 19333 18322 19399 18325
rect 12390 18320 19399 18322
rect 12390 18264 19338 18320
rect 19394 18264 19399 18320
rect 12390 18262 19399 18264
rect 8201 18259 8267 18262
rect 9949 18259 10015 18262
rect 19333 18259 19399 18262
rect 24209 18322 24275 18325
rect 24718 18322 24778 18398
rect 27520 18368 28000 18398
rect 24209 18320 24778 18322
rect 24209 18264 24214 18320
rect 24270 18264 24778 18320
rect 24209 18262 24778 18264
rect 24209 18259 24275 18262
rect 5533 18186 5599 18189
rect 14365 18186 14431 18189
rect 5533 18184 14431 18186
rect 5533 18128 5538 18184
rect 5594 18128 14370 18184
rect 14426 18128 14431 18184
rect 5533 18126 14431 18128
rect 5533 18123 5599 18126
rect 14365 18123 14431 18126
rect 14733 18186 14799 18189
rect 16481 18186 16547 18189
rect 17769 18186 17835 18189
rect 14733 18184 16314 18186
rect 14733 18128 14738 18184
rect 14794 18128 16314 18184
rect 14733 18126 16314 18128
rect 14733 18123 14799 18126
rect 3877 18050 3943 18053
rect 7465 18050 7531 18053
rect 3877 18048 7531 18050
rect 3877 17992 3882 18048
rect 3938 17992 7470 18048
rect 7526 17992 7531 18048
rect 3877 17990 7531 17992
rect 3877 17987 3943 17990
rect 7465 17987 7531 17990
rect 10869 18050 10935 18053
rect 11237 18050 11303 18053
rect 15377 18050 15443 18053
rect 16113 18050 16179 18053
rect 10869 18048 16179 18050
rect 10869 17992 10874 18048
rect 10930 17992 11242 18048
rect 11298 17992 15382 18048
rect 15438 17992 16118 18048
rect 16174 17992 16179 18048
rect 10869 17990 16179 17992
rect 16254 18050 16314 18126
rect 16481 18184 17835 18186
rect 16481 18128 16486 18184
rect 16542 18128 17774 18184
rect 17830 18128 17835 18184
rect 16481 18126 17835 18128
rect 16481 18123 16547 18126
rect 17769 18123 17835 18126
rect 18597 18186 18663 18189
rect 19609 18186 19675 18189
rect 18597 18184 19488 18186
rect 18597 18128 18602 18184
rect 18658 18152 19488 18184
rect 19566 18184 19675 18186
rect 19566 18152 19614 18184
rect 18658 18128 19614 18152
rect 19670 18128 19675 18184
rect 18597 18126 19675 18128
rect 18597 18123 18663 18126
rect 19428 18123 19675 18126
rect 19428 18092 19626 18123
rect 18597 18050 18663 18053
rect 16254 18048 18663 18050
rect 16254 17992 18602 18048
rect 18658 17992 18663 18048
rect 16254 17990 18663 17992
rect 10869 17987 10935 17990
rect 11237 17987 11303 17990
rect 15377 17987 15443 17990
rect 16113 17987 16179 17990
rect 18597 17987 18663 17990
rect 20294 17988 20300 18052
rect 20364 18050 20370 18052
rect 21030 18050 21036 18052
rect 20364 17990 21036 18050
rect 20364 17988 20370 17990
rect 21030 17988 21036 17990
rect 21100 17988 21106 18052
rect 21541 18050 21607 18053
rect 23933 18050 23999 18053
rect 21541 18048 23999 18050
rect 21541 17992 21546 18048
rect 21602 17992 23938 18048
rect 23994 17992 23999 18048
rect 21541 17990 23999 17992
rect 21541 17987 21607 17990
rect 23933 17987 23999 17990
rect 10277 17984 10597 17985
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 17919 10597 17920
rect 19610 17984 19930 17985
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 17919 19930 17920
rect 1945 17914 2011 17917
rect 3141 17914 3207 17917
rect 1945 17912 3207 17914
rect 1945 17856 1950 17912
rect 2006 17856 3146 17912
rect 3202 17856 3207 17912
rect 1945 17854 3207 17856
rect 1945 17851 2011 17854
rect 3141 17851 3207 17854
rect 5073 17914 5139 17917
rect 9673 17914 9739 17917
rect 5073 17912 9739 17914
rect 5073 17856 5078 17912
rect 5134 17856 9678 17912
rect 9734 17856 9739 17912
rect 5073 17854 9739 17856
rect 5073 17851 5139 17854
rect 9673 17851 9739 17854
rect 10910 17852 10916 17916
rect 10980 17914 10986 17916
rect 18505 17914 18571 17917
rect 10980 17912 18571 17914
rect 10980 17856 18510 17912
rect 18566 17856 18571 17912
rect 10980 17854 18571 17856
rect 10980 17852 10986 17854
rect 18505 17851 18571 17854
rect 20529 17914 20595 17917
rect 20713 17914 20779 17917
rect 22502 17914 22508 17916
rect 20529 17912 22508 17914
rect 20529 17856 20534 17912
rect 20590 17856 20718 17912
rect 20774 17856 22508 17912
rect 20529 17854 22508 17856
rect 20529 17851 20595 17854
rect 20713 17851 20779 17854
rect 22502 17852 22508 17854
rect 22572 17914 22578 17916
rect 23565 17914 23631 17917
rect 22572 17912 23631 17914
rect 22572 17856 23570 17912
rect 23626 17856 23631 17912
rect 22572 17854 23631 17856
rect 22572 17852 22578 17854
rect 23565 17851 23631 17854
rect 25037 17914 25103 17917
rect 25262 17914 25268 17916
rect 25037 17912 25268 17914
rect 25037 17856 25042 17912
rect 25098 17856 25268 17912
rect 25037 17854 25268 17856
rect 25037 17851 25103 17854
rect 25262 17852 25268 17854
rect 25332 17852 25338 17916
rect 0 17778 480 17808
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17688 480 17718
rect 2773 17715 2839 17718
rect 5625 17778 5691 17781
rect 12065 17778 12131 17781
rect 5625 17776 12131 17778
rect 5625 17720 5630 17776
rect 5686 17720 12070 17776
rect 12126 17720 12131 17776
rect 5625 17718 12131 17720
rect 5625 17715 5691 17718
rect 12065 17715 12131 17718
rect 17493 17778 17559 17781
rect 19977 17778 20043 17781
rect 17493 17776 20043 17778
rect 17493 17720 17498 17776
rect 17554 17720 19982 17776
rect 20038 17720 20043 17776
rect 17493 17718 20043 17720
rect 17493 17715 17559 17718
rect 19977 17715 20043 17718
rect 20110 17716 20116 17780
rect 20180 17778 20186 17780
rect 25037 17778 25103 17781
rect 20180 17776 25103 17778
rect 20180 17720 25042 17776
rect 25098 17720 25103 17776
rect 20180 17718 25103 17720
rect 20180 17716 20186 17718
rect 25037 17715 25103 17718
rect 25405 17778 25471 17781
rect 27520 17778 28000 17808
rect 25405 17776 28000 17778
rect 25405 17720 25410 17776
rect 25466 17720 28000 17776
rect 25405 17718 28000 17720
rect 25405 17715 25471 17718
rect 27520 17688 28000 17718
rect 4797 17642 4863 17645
rect 9489 17642 9555 17645
rect 4797 17640 9555 17642
rect 4797 17584 4802 17640
rect 4858 17584 9494 17640
rect 9550 17584 9555 17640
rect 4797 17582 9555 17584
rect 4797 17579 4863 17582
rect 9489 17579 9555 17582
rect 15377 17642 15443 17645
rect 24945 17642 25011 17645
rect 15377 17640 25011 17642
rect 15377 17584 15382 17640
rect 15438 17584 24950 17640
rect 25006 17584 25011 17640
rect 15377 17582 25011 17584
rect 15377 17579 15443 17582
rect 24945 17579 25011 17582
rect 6453 17506 6519 17509
rect 14549 17506 14615 17509
rect 6453 17504 14615 17506
rect 6453 17448 6458 17504
rect 6514 17448 14554 17504
rect 14610 17448 14615 17504
rect 6453 17446 14615 17448
rect 6453 17443 6519 17446
rect 14549 17443 14615 17446
rect 18965 17506 19031 17509
rect 19425 17506 19491 17509
rect 20897 17506 20963 17509
rect 18965 17504 19304 17506
rect 18965 17448 18970 17504
rect 19026 17448 19304 17504
rect 18965 17446 19304 17448
rect 18965 17443 19031 17446
rect 5610 17440 5930 17441
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5930 17440
rect 5610 17375 5930 17376
rect 14944 17440 15264 17441
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 17375 15264 17376
rect 6545 17370 6611 17373
rect 10910 17370 10916 17372
rect 6545 17368 10916 17370
rect 6545 17312 6550 17368
rect 6606 17312 10916 17368
rect 6545 17310 10916 17312
rect 6545 17307 6611 17310
rect 10910 17308 10916 17310
rect 10980 17308 10986 17372
rect 19244 17370 19304 17446
rect 19425 17504 20963 17506
rect 19425 17448 19430 17504
rect 19486 17448 20902 17504
rect 20958 17448 20963 17504
rect 19425 17446 20963 17448
rect 19425 17443 19491 17446
rect 20897 17443 20963 17446
rect 24277 17440 24597 17441
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 17375 24597 17376
rect 19517 17370 19583 17373
rect 23749 17370 23815 17373
rect 19244 17368 23815 17370
rect 19244 17312 19522 17368
rect 19578 17312 23754 17368
rect 23810 17312 23815 17368
rect 19244 17310 23815 17312
rect 19517 17307 19583 17310
rect 23749 17307 23815 17310
rect 0 17234 480 17264
rect 4245 17234 4311 17237
rect 0 17232 4311 17234
rect 0 17176 4250 17232
rect 4306 17176 4311 17232
rect 0 17174 4311 17176
rect 0 17144 480 17174
rect 4245 17171 4311 17174
rect 4705 17234 4771 17237
rect 5073 17234 5139 17237
rect 4705 17232 5139 17234
rect 4705 17176 4710 17232
rect 4766 17176 5078 17232
rect 5134 17176 5139 17232
rect 4705 17174 5139 17176
rect 4705 17171 4771 17174
rect 5073 17171 5139 17174
rect 5625 17234 5691 17237
rect 6126 17234 6132 17236
rect 5625 17232 6132 17234
rect 5625 17176 5630 17232
rect 5686 17176 6132 17232
rect 5625 17174 6132 17176
rect 5625 17171 5691 17174
rect 6126 17172 6132 17174
rect 6196 17172 6202 17236
rect 6913 17234 6979 17237
rect 12893 17234 12959 17237
rect 13261 17234 13327 17237
rect 17217 17234 17283 17237
rect 22870 17234 22876 17236
rect 6913 17232 11944 17234
rect 6913 17176 6918 17232
rect 6974 17176 11944 17232
rect 6913 17174 11944 17176
rect 6913 17171 6979 17174
rect 3049 17098 3115 17101
rect 5165 17098 5231 17101
rect 11884 17098 11944 17174
rect 12893 17232 14428 17234
rect 12893 17176 12898 17232
rect 12954 17176 13266 17232
rect 13322 17176 14428 17232
rect 12893 17174 14428 17176
rect 12893 17171 12959 17174
rect 13261 17171 13327 17174
rect 14181 17098 14247 17101
rect 3049 17096 11346 17098
rect 3049 17040 3054 17096
rect 3110 17040 5170 17096
rect 5226 17040 11346 17096
rect 3049 17038 11346 17040
rect 11884 17096 14247 17098
rect 11884 17040 14186 17096
rect 14242 17040 14247 17096
rect 11884 17038 14247 17040
rect 14368 17098 14428 17174
rect 17217 17232 22876 17234
rect 17217 17176 17222 17232
rect 17278 17176 22876 17232
rect 17217 17174 22876 17176
rect 17217 17171 17283 17174
rect 22870 17172 22876 17174
rect 22940 17172 22946 17236
rect 25497 17234 25563 17237
rect 27520 17234 28000 17264
rect 25497 17232 28000 17234
rect 25497 17176 25502 17232
rect 25558 17176 28000 17232
rect 25497 17174 28000 17176
rect 25497 17171 25563 17174
rect 27520 17144 28000 17174
rect 20110 17098 20116 17100
rect 14368 17038 20116 17098
rect 3049 17035 3115 17038
rect 5165 17035 5231 17038
rect 2957 16962 3023 16965
rect 8201 16962 8267 16965
rect 2957 16960 8267 16962
rect 2957 16904 2962 16960
rect 3018 16904 8206 16960
rect 8262 16904 8267 16960
rect 2957 16902 8267 16904
rect 2957 16899 3023 16902
rect 8201 16899 8267 16902
rect 10277 16896 10597 16897
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 10277 16831 10597 16832
rect 3877 16826 3943 16829
rect 6453 16826 6519 16829
rect 3877 16824 6519 16826
rect 3877 16768 3882 16824
rect 3938 16768 6458 16824
rect 6514 16768 6519 16824
rect 3877 16766 6519 16768
rect 3877 16763 3943 16766
rect 6453 16763 6519 16766
rect 0 16690 480 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 480 16630
rect 4061 16627 4127 16630
rect 5257 16690 5323 16693
rect 8477 16690 8543 16693
rect 5257 16688 8543 16690
rect 5257 16632 5262 16688
rect 5318 16632 8482 16688
rect 8538 16632 8543 16688
rect 5257 16630 8543 16632
rect 5257 16627 5323 16630
rect 8477 16627 8543 16630
rect 9213 16690 9279 16693
rect 11145 16690 11211 16693
rect 9213 16688 11211 16690
rect 9213 16632 9218 16688
rect 9274 16632 11150 16688
rect 11206 16632 11211 16688
rect 9213 16630 11211 16632
rect 11286 16690 11346 17038
rect 14181 17035 14247 17038
rect 20110 17036 20116 17038
rect 20180 17036 20186 17100
rect 20478 17036 20484 17100
rect 20548 17098 20554 17100
rect 25221 17098 25287 17101
rect 20548 17096 25287 17098
rect 20548 17040 25226 17096
rect 25282 17040 25287 17096
rect 20548 17038 25287 17040
rect 20548 17036 20554 17038
rect 25221 17035 25287 17038
rect 17953 16962 18019 16965
rect 18413 16962 18479 16965
rect 17953 16960 18479 16962
rect 17953 16904 17958 16960
rect 18014 16904 18418 16960
rect 18474 16904 18479 16960
rect 17953 16902 18479 16904
rect 17953 16899 18019 16902
rect 18413 16899 18479 16902
rect 20662 16900 20668 16964
rect 20732 16962 20738 16964
rect 20897 16962 20963 16965
rect 20732 16960 20963 16962
rect 20732 16904 20902 16960
rect 20958 16904 20963 16960
rect 20732 16902 20963 16904
rect 20732 16900 20738 16902
rect 20897 16899 20963 16902
rect 21541 16962 21607 16965
rect 21541 16960 24962 16962
rect 21541 16904 21546 16960
rect 21602 16904 24962 16960
rect 21541 16902 24962 16904
rect 21541 16899 21607 16902
rect 19610 16896 19930 16897
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 16831 19930 16832
rect 16389 16826 16455 16829
rect 18413 16826 18479 16829
rect 16389 16824 18479 16826
rect 16389 16768 16394 16824
rect 16450 16768 18418 16824
rect 18474 16768 18479 16824
rect 16389 16766 18479 16768
rect 16389 16763 16455 16766
rect 18413 16763 18479 16766
rect 21449 16826 21515 16829
rect 23657 16826 23723 16829
rect 21449 16824 23723 16826
rect 21449 16768 21454 16824
rect 21510 16768 23662 16824
rect 23718 16768 23723 16824
rect 21449 16766 23723 16768
rect 21449 16763 21515 16766
rect 23657 16763 23723 16766
rect 14917 16690 14983 16693
rect 11286 16688 14983 16690
rect 11286 16632 14922 16688
rect 14978 16632 14983 16688
rect 11286 16630 14983 16632
rect 9213 16627 9279 16630
rect 11145 16627 11211 16630
rect 14917 16627 14983 16630
rect 18045 16690 18111 16693
rect 20713 16690 20779 16693
rect 18045 16688 20779 16690
rect 18045 16632 18050 16688
rect 18106 16632 20718 16688
rect 20774 16632 20779 16688
rect 18045 16630 20779 16632
rect 18045 16627 18111 16630
rect 20713 16627 20779 16630
rect 21357 16690 21423 16693
rect 24902 16690 24962 16902
rect 27520 16690 28000 16720
rect 21357 16688 24778 16690
rect 21357 16632 21362 16688
rect 21418 16632 24778 16688
rect 21357 16630 24778 16632
rect 24902 16630 28000 16690
rect 21357 16627 21423 16630
rect 1393 16554 1459 16557
rect 9397 16554 9463 16557
rect 1393 16552 9463 16554
rect 1393 16496 1398 16552
rect 1454 16496 9402 16552
rect 9458 16496 9463 16552
rect 1393 16494 9463 16496
rect 1393 16491 1459 16494
rect 9397 16491 9463 16494
rect 9581 16554 9647 16557
rect 14733 16554 14799 16557
rect 9581 16552 14799 16554
rect 9581 16496 9586 16552
rect 9642 16496 14738 16552
rect 14794 16496 14799 16552
rect 9581 16494 14799 16496
rect 9581 16491 9647 16494
rect 14733 16491 14799 16494
rect 16665 16554 16731 16557
rect 23381 16554 23447 16557
rect 16665 16552 23447 16554
rect 16665 16496 16670 16552
rect 16726 16496 23386 16552
rect 23442 16496 23447 16552
rect 16665 16494 23447 16496
rect 24718 16554 24778 16630
rect 27520 16600 28000 16630
rect 24853 16554 24919 16557
rect 24718 16552 24919 16554
rect 24718 16496 24858 16552
rect 24914 16496 24919 16552
rect 24718 16494 24919 16496
rect 16665 16491 16731 16494
rect 23381 16491 23447 16494
rect 24853 16491 24919 16494
rect 6545 16418 6611 16421
rect 6678 16418 6684 16420
rect 6545 16416 6684 16418
rect 6545 16360 6550 16416
rect 6606 16360 6684 16416
rect 6545 16358 6684 16360
rect 6545 16355 6611 16358
rect 6678 16356 6684 16358
rect 6748 16356 6754 16420
rect 8661 16418 8727 16421
rect 11237 16418 11303 16421
rect 8661 16416 11303 16418
rect 8661 16360 8666 16416
rect 8722 16360 11242 16416
rect 11298 16360 11303 16416
rect 8661 16358 11303 16360
rect 8661 16355 8727 16358
rect 11237 16355 11303 16358
rect 11421 16418 11487 16421
rect 13813 16418 13879 16421
rect 11421 16416 13879 16418
rect 11421 16360 11426 16416
rect 11482 16360 13818 16416
rect 13874 16360 13879 16416
rect 11421 16358 13879 16360
rect 11421 16355 11487 16358
rect 13813 16355 13879 16358
rect 16389 16418 16455 16421
rect 18045 16418 18111 16421
rect 16389 16416 18111 16418
rect 16389 16360 16394 16416
rect 16450 16360 18050 16416
rect 18106 16360 18111 16416
rect 16389 16358 18111 16360
rect 16389 16355 16455 16358
rect 18045 16355 18111 16358
rect 18965 16418 19031 16421
rect 22737 16418 22803 16421
rect 18965 16416 22803 16418
rect 18965 16360 18970 16416
rect 19026 16360 22742 16416
rect 22798 16360 22803 16416
rect 18965 16358 22803 16360
rect 18965 16355 19031 16358
rect 22737 16355 22803 16358
rect 5610 16352 5930 16353
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5930 16352
rect 5610 16287 5930 16288
rect 14944 16352 15264 16353
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14944 16287 15264 16288
rect 24277 16352 24597 16353
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 16287 24597 16288
rect 9990 16220 9996 16284
rect 10060 16282 10066 16284
rect 14590 16282 14596 16284
rect 10060 16222 14596 16282
rect 10060 16220 10066 16222
rect 14590 16220 14596 16222
rect 14660 16220 14666 16284
rect 15469 16282 15535 16285
rect 16665 16282 16731 16285
rect 15469 16280 16731 16282
rect 15469 16224 15474 16280
rect 15530 16224 16670 16280
rect 16726 16224 16731 16280
rect 15469 16222 16731 16224
rect 15469 16219 15535 16222
rect 16665 16219 16731 16222
rect 19885 16282 19951 16285
rect 23565 16282 23631 16285
rect 19885 16280 23631 16282
rect 19885 16224 19890 16280
rect 19946 16224 23570 16280
rect 23626 16224 23631 16280
rect 19885 16222 23631 16224
rect 19885 16219 19951 16222
rect 23565 16219 23631 16222
rect 2405 16146 2471 16149
rect 4981 16146 5047 16149
rect 2405 16144 5047 16146
rect 2405 16088 2410 16144
rect 2466 16088 4986 16144
rect 5042 16088 5047 16144
rect 2405 16086 5047 16088
rect 2405 16083 2471 16086
rect 4981 16083 5047 16086
rect 5625 16146 5691 16149
rect 14365 16146 14431 16149
rect 5625 16144 14431 16146
rect 5625 16088 5630 16144
rect 5686 16088 14370 16144
rect 14426 16088 14431 16144
rect 5625 16086 14431 16088
rect 5625 16083 5691 16086
rect 14365 16083 14431 16086
rect 19977 16146 20043 16149
rect 20897 16146 20963 16149
rect 24853 16146 24919 16149
rect 19977 16144 24919 16146
rect 19977 16088 19982 16144
rect 20038 16088 20902 16144
rect 20958 16088 24858 16144
rect 24914 16088 24919 16144
rect 19977 16086 24919 16088
rect 19977 16083 20043 16086
rect 20897 16083 20963 16086
rect 24853 16083 24919 16086
rect 0 16010 480 16040
rect 7005 16010 7071 16013
rect 0 16008 7071 16010
rect 0 15952 7010 16008
rect 7066 15952 7071 16008
rect 0 15950 7071 15952
rect 0 15920 480 15950
rect 7005 15947 7071 15950
rect 8477 16010 8543 16013
rect 11789 16010 11855 16013
rect 13261 16012 13327 16013
rect 13261 16010 13308 16012
rect 8477 16008 11855 16010
rect 8477 15952 8482 16008
rect 8538 15952 11794 16008
rect 11850 15952 11855 16008
rect 8477 15950 11855 15952
rect 13216 16008 13308 16010
rect 13216 15952 13266 16008
rect 13216 15950 13308 15952
rect 8477 15947 8543 15950
rect 11789 15947 11855 15950
rect 13261 15948 13308 15950
rect 13372 15948 13378 16012
rect 13997 16010 14063 16013
rect 21030 16010 21036 16012
rect 13997 16008 21036 16010
rect 13997 15952 14002 16008
rect 14058 15952 21036 16008
rect 13997 15950 21036 15952
rect 13261 15947 13327 15948
rect 13997 15947 14063 15950
rect 21030 15948 21036 15950
rect 21100 15948 21106 16012
rect 23473 16010 23539 16013
rect 24301 16010 24367 16013
rect 23473 16008 24367 16010
rect 23473 15952 23478 16008
rect 23534 15952 24306 16008
rect 24362 15952 24367 16008
rect 23473 15950 24367 15952
rect 23473 15947 23539 15950
rect 24301 15947 24367 15950
rect 25405 16010 25471 16013
rect 27520 16010 28000 16040
rect 25405 16008 28000 16010
rect 25405 15952 25410 16008
rect 25466 15952 28000 16008
rect 25405 15950 28000 15952
rect 25405 15947 25471 15950
rect 27520 15920 28000 15950
rect 3601 15874 3667 15877
rect 9581 15874 9647 15877
rect 3601 15872 9647 15874
rect 3601 15816 3606 15872
rect 3662 15816 9586 15872
rect 9642 15816 9647 15872
rect 3601 15814 9647 15816
rect 3601 15811 3667 15814
rect 9581 15811 9647 15814
rect 14825 15874 14891 15877
rect 15193 15874 15259 15877
rect 18137 15874 18203 15877
rect 20897 15876 20963 15877
rect 14825 15872 18203 15874
rect 14825 15816 14830 15872
rect 14886 15816 15198 15872
rect 15254 15816 18142 15872
rect 18198 15816 18203 15872
rect 14825 15814 18203 15816
rect 14825 15811 14891 15814
rect 15193 15811 15259 15814
rect 18137 15811 18203 15814
rect 20846 15812 20852 15876
rect 20916 15874 20963 15876
rect 21817 15874 21883 15877
rect 20916 15872 21883 15874
rect 20958 15816 21822 15872
rect 21878 15816 21883 15872
rect 20916 15814 21883 15816
rect 20916 15812 20963 15814
rect 20897 15811 20963 15812
rect 21817 15811 21883 15814
rect 10277 15808 10597 15809
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 15743 10597 15744
rect 19610 15808 19930 15809
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 15743 19930 15744
rect 4981 15738 5047 15741
rect 6126 15738 6132 15740
rect 4981 15736 6132 15738
rect 4981 15680 4986 15736
rect 5042 15680 6132 15736
rect 4981 15678 6132 15680
rect 4981 15675 5047 15678
rect 6126 15676 6132 15678
rect 6196 15676 6202 15740
rect 8109 15738 8175 15741
rect 9673 15738 9739 15741
rect 8109 15736 9739 15738
rect 8109 15680 8114 15736
rect 8170 15680 9678 15736
rect 9734 15680 9739 15736
rect 8109 15678 9739 15680
rect 8109 15675 8175 15678
rect 9673 15675 9739 15678
rect 11237 15738 11303 15741
rect 13721 15738 13787 15741
rect 15653 15738 15719 15741
rect 11237 15736 15719 15738
rect 11237 15680 11242 15736
rect 11298 15680 13726 15736
rect 13782 15680 15658 15736
rect 15714 15680 15719 15736
rect 11237 15678 15719 15680
rect 11237 15675 11303 15678
rect 13721 15675 13787 15678
rect 15653 15675 15719 15678
rect 18045 15738 18111 15741
rect 19149 15738 19215 15741
rect 18045 15736 19215 15738
rect 18045 15680 18050 15736
rect 18106 15680 19154 15736
rect 19210 15680 19215 15736
rect 18045 15678 19215 15680
rect 18045 15675 18111 15678
rect 19149 15675 19215 15678
rect 21265 15738 21331 15741
rect 24485 15738 24551 15741
rect 21265 15736 24551 15738
rect 21265 15680 21270 15736
rect 21326 15680 24490 15736
rect 24546 15680 24551 15736
rect 21265 15678 24551 15680
rect 21265 15675 21331 15678
rect 24485 15675 24551 15678
rect 5533 15602 5599 15605
rect 7833 15602 7899 15605
rect 11421 15602 11487 15605
rect 5533 15600 11487 15602
rect 5533 15544 5538 15600
rect 5594 15544 7838 15600
rect 7894 15544 11426 15600
rect 11482 15544 11487 15600
rect 5533 15542 11487 15544
rect 5533 15539 5599 15542
rect 7833 15539 7899 15542
rect 11421 15539 11487 15542
rect 15009 15602 15075 15605
rect 20713 15602 20779 15605
rect 15009 15600 20779 15602
rect 15009 15544 15014 15600
rect 15070 15544 20718 15600
rect 20774 15544 20779 15600
rect 15009 15542 20779 15544
rect 15009 15539 15075 15542
rect 20713 15539 20779 15542
rect 20897 15602 20963 15605
rect 24025 15602 24091 15605
rect 20897 15600 24091 15602
rect 20897 15544 20902 15600
rect 20958 15544 24030 15600
rect 24086 15544 24091 15600
rect 20897 15542 24091 15544
rect 20897 15539 20963 15542
rect 24025 15539 24091 15542
rect 24301 15602 24367 15605
rect 25313 15602 25379 15605
rect 24301 15600 25379 15602
rect 24301 15544 24306 15600
rect 24362 15544 25318 15600
rect 25374 15544 25379 15600
rect 24301 15542 25379 15544
rect 24301 15539 24367 15542
rect 25313 15539 25379 15542
rect 0 15466 480 15496
rect 1577 15466 1643 15469
rect 0 15464 1643 15466
rect 0 15408 1582 15464
rect 1638 15408 1643 15464
rect 0 15406 1643 15408
rect 0 15376 480 15406
rect 1577 15403 1643 15406
rect 1853 15466 1919 15469
rect 5441 15466 5507 15469
rect 7465 15466 7531 15469
rect 1853 15464 5320 15466
rect 1853 15408 1858 15464
rect 1914 15408 5320 15464
rect 1853 15406 5320 15408
rect 1853 15403 1919 15406
rect 2221 15330 2287 15333
rect 4337 15330 4403 15333
rect 2221 15328 4403 15330
rect 2221 15272 2226 15328
rect 2282 15272 4342 15328
rect 4398 15272 4403 15328
rect 2221 15270 4403 15272
rect 5260 15330 5320 15406
rect 5441 15464 7531 15466
rect 5441 15408 5446 15464
rect 5502 15408 7470 15464
rect 7526 15408 7531 15464
rect 5441 15406 7531 15408
rect 5441 15403 5507 15406
rect 7465 15403 7531 15406
rect 8017 15466 8083 15469
rect 13813 15466 13879 15469
rect 18505 15466 18571 15469
rect 8017 15464 13879 15466
rect 8017 15408 8022 15464
rect 8078 15408 13818 15464
rect 13874 15408 13879 15464
rect 8017 15406 13879 15408
rect 8017 15403 8083 15406
rect 13813 15403 13879 15406
rect 14414 15464 18571 15466
rect 14414 15408 18510 15464
rect 18566 15408 18571 15464
rect 14414 15406 18571 15408
rect 5441 15330 5507 15333
rect 5260 15328 5507 15330
rect 5260 15272 5446 15328
rect 5502 15272 5507 15328
rect 5260 15270 5507 15272
rect 2221 15267 2287 15270
rect 4337 15267 4403 15270
rect 5441 15267 5507 15270
rect 6269 15330 6335 15333
rect 10501 15330 10567 15333
rect 6269 15328 10567 15330
rect 6269 15272 6274 15328
rect 6330 15272 10506 15328
rect 10562 15272 10567 15328
rect 6269 15270 10567 15272
rect 6269 15267 6335 15270
rect 10501 15267 10567 15270
rect 13445 15330 13511 15333
rect 14414 15330 14474 15406
rect 18505 15403 18571 15406
rect 21081 15466 21147 15469
rect 27520 15466 28000 15496
rect 21081 15464 28000 15466
rect 21081 15408 21086 15464
rect 21142 15408 28000 15464
rect 21081 15406 28000 15408
rect 21081 15403 21147 15406
rect 27520 15376 28000 15406
rect 13445 15328 14474 15330
rect 13445 15272 13450 15328
rect 13506 15272 14474 15328
rect 13445 15270 14474 15272
rect 20345 15330 20411 15333
rect 23381 15330 23447 15333
rect 20345 15328 23447 15330
rect 20345 15272 20350 15328
rect 20406 15272 23386 15328
rect 23442 15272 23447 15328
rect 20345 15270 23447 15272
rect 13445 15267 13511 15270
rect 20345 15267 20411 15270
rect 23381 15267 23447 15270
rect 25313 15330 25379 15333
rect 25589 15330 25655 15333
rect 25313 15328 25655 15330
rect 25313 15272 25318 15328
rect 25374 15272 25594 15328
rect 25650 15272 25655 15328
rect 25313 15270 25655 15272
rect 25313 15267 25379 15270
rect 25589 15267 25655 15270
rect 5610 15264 5930 15265
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5930 15264
rect 5610 15199 5930 15200
rect 14944 15264 15264 15265
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14944 15199 15264 15200
rect 24277 15264 24597 15265
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 15199 24597 15200
rect 8845 15194 8911 15197
rect 8845 15192 13508 15194
rect 8845 15136 8850 15192
rect 8906 15136 13508 15192
rect 8845 15134 13508 15136
rect 8845 15131 8911 15134
rect 2037 15058 2103 15061
rect 2957 15058 3023 15061
rect 11329 15058 11395 15061
rect 2037 15056 11395 15058
rect 2037 15000 2042 15056
rect 2098 15000 2962 15056
rect 3018 15000 11334 15056
rect 11390 15000 11395 15056
rect 2037 14998 11395 15000
rect 13448 15058 13508 15134
rect 13854 15132 13860 15196
rect 13924 15194 13930 15196
rect 14089 15194 14155 15197
rect 13924 15192 14155 15194
rect 13924 15136 14094 15192
rect 14150 15136 14155 15192
rect 13924 15134 14155 15136
rect 13924 15132 13930 15134
rect 14089 15131 14155 15134
rect 17309 15194 17375 15197
rect 20713 15194 20779 15197
rect 17309 15192 20779 15194
rect 17309 15136 17314 15192
rect 17370 15136 20718 15192
rect 20774 15136 20779 15192
rect 17309 15134 20779 15136
rect 17309 15131 17375 15134
rect 20713 15131 20779 15134
rect 16573 15058 16639 15061
rect 19977 15058 20043 15061
rect 20294 15058 20300 15060
rect 13448 15056 16639 15058
rect 13448 15000 16578 15056
rect 16634 15000 16639 15056
rect 13448 14998 16639 15000
rect 2037 14995 2103 14998
rect 2957 14995 3023 14998
rect 11329 14995 11395 14998
rect 16573 14995 16639 14998
rect 17772 15056 20300 15058
rect 17772 15000 19982 15056
rect 20038 15000 20300 15056
rect 17772 14998 20300 15000
rect 0 14922 480 14952
rect 1577 14922 1643 14925
rect 0 14920 1643 14922
rect 0 14864 1582 14920
rect 1638 14864 1643 14920
rect 0 14862 1643 14864
rect 0 14832 480 14862
rect 1577 14859 1643 14862
rect 4705 14922 4771 14925
rect 13537 14922 13603 14925
rect 4705 14920 13603 14922
rect 4705 14864 4710 14920
rect 4766 14864 13542 14920
rect 13598 14864 13603 14920
rect 4705 14862 13603 14864
rect 4705 14859 4771 14862
rect 13537 14859 13603 14862
rect 16205 14922 16271 14925
rect 17772 14922 17832 14998
rect 19977 14995 20043 14998
rect 20294 14996 20300 14998
rect 20364 14996 20370 15060
rect 23238 14996 23244 15060
rect 23308 15058 23314 15060
rect 24894 15058 24900 15060
rect 23308 14998 24900 15058
rect 23308 14996 23314 14998
rect 24894 14996 24900 14998
rect 24964 14996 24970 15060
rect 16205 14920 17832 14922
rect 16205 14864 16210 14920
rect 16266 14864 17832 14920
rect 16205 14862 17832 14864
rect 19241 14922 19307 14925
rect 20478 14922 20484 14924
rect 19241 14920 20484 14922
rect 19241 14864 19246 14920
rect 19302 14864 20484 14920
rect 19241 14862 20484 14864
rect 16205 14859 16271 14862
rect 19241 14859 19307 14862
rect 20478 14860 20484 14862
rect 20548 14860 20554 14924
rect 23657 14922 23723 14925
rect 24761 14922 24827 14925
rect 23657 14920 24827 14922
rect 23657 14864 23662 14920
rect 23718 14864 24766 14920
rect 24822 14864 24827 14920
rect 23657 14862 24827 14864
rect 23657 14859 23723 14862
rect 24761 14859 24827 14862
rect 25313 14922 25379 14925
rect 27520 14922 28000 14952
rect 25313 14920 28000 14922
rect 25313 14864 25318 14920
rect 25374 14864 28000 14920
rect 25313 14862 28000 14864
rect 25313 14859 25379 14862
rect 27520 14832 28000 14862
rect 4889 14786 4955 14789
rect 1718 14784 4955 14786
rect 1718 14728 4894 14784
rect 4950 14728 4955 14784
rect 1718 14726 4955 14728
rect 1718 14653 1778 14726
rect 4889 14723 4955 14726
rect 5441 14786 5507 14789
rect 6310 14786 6316 14788
rect 5441 14784 6316 14786
rect 5441 14728 5446 14784
rect 5502 14728 6316 14784
rect 5441 14726 6316 14728
rect 5441 14723 5507 14726
rect 6310 14724 6316 14726
rect 6380 14786 6386 14788
rect 6729 14786 6795 14789
rect 6380 14784 6795 14786
rect 6380 14728 6734 14784
rect 6790 14728 6795 14784
rect 6380 14726 6795 14728
rect 6380 14724 6386 14726
rect 6729 14723 6795 14726
rect 6913 14786 6979 14789
rect 9673 14786 9739 14789
rect 6913 14784 9739 14786
rect 6913 14728 6918 14784
rect 6974 14728 9678 14784
rect 9734 14728 9739 14784
rect 6913 14726 9739 14728
rect 6913 14723 6979 14726
rect 9673 14723 9739 14726
rect 21725 14786 21791 14789
rect 24117 14786 24183 14789
rect 21725 14784 24183 14786
rect 21725 14728 21730 14784
rect 21786 14728 24122 14784
rect 24178 14728 24183 14784
rect 21725 14726 24183 14728
rect 21725 14723 21791 14726
rect 24117 14723 24183 14726
rect 24710 14724 24716 14788
rect 24780 14786 24786 14788
rect 24945 14786 25011 14789
rect 24780 14784 25011 14786
rect 24780 14728 24950 14784
rect 25006 14728 25011 14784
rect 24780 14726 25011 14728
rect 24780 14724 24786 14726
rect 24945 14723 25011 14726
rect 10277 14720 10597 14721
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 14655 10597 14656
rect 19610 14720 19930 14721
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 14655 19930 14656
rect 1669 14648 1778 14653
rect 1669 14592 1674 14648
rect 1730 14592 1778 14648
rect 1669 14590 1778 14592
rect 2405 14650 2471 14653
rect 6269 14650 6335 14653
rect 2405 14648 6335 14650
rect 2405 14592 2410 14648
rect 2466 14592 6274 14648
rect 6330 14592 6335 14648
rect 2405 14590 6335 14592
rect 1669 14587 1735 14590
rect 2405 14587 2471 14590
rect 6269 14587 6335 14590
rect 7925 14650 7991 14653
rect 9622 14650 9628 14652
rect 7925 14648 9628 14650
rect 7925 14592 7930 14648
rect 7986 14592 9628 14648
rect 7925 14590 9628 14592
rect 7925 14587 7991 14590
rect 9622 14588 9628 14590
rect 9692 14588 9698 14652
rect 15745 14650 15811 14653
rect 18781 14650 18847 14653
rect 15745 14648 18847 14650
rect 15745 14592 15750 14648
rect 15806 14592 18786 14648
rect 18842 14592 18847 14648
rect 15745 14590 18847 14592
rect 15745 14587 15811 14590
rect 18781 14587 18847 14590
rect 24117 14650 24183 14653
rect 26141 14650 26207 14653
rect 24117 14648 26207 14650
rect 24117 14592 24122 14648
rect 24178 14592 26146 14648
rect 26202 14592 26207 14648
rect 24117 14590 26207 14592
rect 24117 14587 24183 14590
rect 26141 14587 26207 14590
rect 2865 14514 2931 14517
rect 11697 14514 11763 14517
rect 2865 14512 11763 14514
rect 2865 14456 2870 14512
rect 2926 14456 11702 14512
rect 11758 14456 11763 14512
rect 2865 14454 11763 14456
rect 2865 14451 2931 14454
rect 11697 14451 11763 14454
rect 16849 14514 16915 14517
rect 20713 14514 20779 14517
rect 16849 14512 20779 14514
rect 16849 14456 16854 14512
rect 16910 14456 20718 14512
rect 20774 14456 20779 14512
rect 16849 14454 20779 14456
rect 16849 14451 16915 14454
rect 20713 14451 20779 14454
rect 0 14378 480 14408
rect 7005 14378 7071 14381
rect 14549 14378 14615 14381
rect 0 14376 7071 14378
rect 0 14320 7010 14376
rect 7066 14320 7071 14376
rect 0 14318 7071 14320
rect 0 14288 480 14318
rect 7005 14315 7071 14318
rect 7238 14376 14615 14378
rect 7238 14320 14554 14376
rect 14610 14320 14615 14376
rect 7238 14318 14615 14320
rect 5610 14176 5930 14177
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5930 14176
rect 5610 14111 5930 14112
rect 2037 13970 2103 13973
rect 2446 13970 2452 13972
rect 2037 13968 2452 13970
rect 2037 13912 2042 13968
rect 2098 13912 2452 13968
rect 2037 13910 2452 13912
rect 2037 13907 2103 13910
rect 2446 13908 2452 13910
rect 2516 13908 2522 13972
rect 4889 13970 4955 13973
rect 7238 13970 7298 14318
rect 14549 14315 14615 14318
rect 18505 14378 18571 14381
rect 27520 14378 28000 14408
rect 18505 14376 28000 14378
rect 18505 14320 18510 14376
rect 18566 14320 28000 14376
rect 18505 14318 28000 14320
rect 18505 14315 18571 14318
rect 27520 14288 28000 14318
rect 9213 14242 9279 14245
rect 11881 14242 11947 14245
rect 14222 14242 14228 14244
rect 9213 14240 14228 14242
rect 9213 14184 9218 14240
rect 9274 14184 11886 14240
rect 11942 14184 14228 14240
rect 9213 14182 14228 14184
rect 9213 14179 9279 14182
rect 11881 14179 11947 14182
rect 14222 14180 14228 14182
rect 14292 14180 14298 14244
rect 22318 14180 22324 14244
rect 22388 14242 22394 14244
rect 24025 14242 24091 14245
rect 22388 14240 24091 14242
rect 22388 14184 24030 14240
rect 24086 14184 24091 14240
rect 22388 14182 24091 14184
rect 22388 14180 22394 14182
rect 24025 14179 24091 14182
rect 14944 14176 15264 14177
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 14111 15264 14112
rect 24277 14176 24597 14177
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 14111 24597 14112
rect 9765 14106 9831 14109
rect 11094 14106 11100 14108
rect 9765 14104 11100 14106
rect 9765 14048 9770 14104
rect 9826 14048 11100 14104
rect 9765 14046 11100 14048
rect 9765 14043 9831 14046
rect 11094 14044 11100 14046
rect 11164 14044 11170 14108
rect 15929 14106 15995 14109
rect 19241 14106 19307 14109
rect 15929 14104 19307 14106
rect 15929 14048 15934 14104
rect 15990 14048 19246 14104
rect 19302 14048 19307 14104
rect 15929 14046 19307 14048
rect 15929 14043 15995 14046
rect 19241 14043 19307 14046
rect 20989 14106 21055 14109
rect 23933 14106 23999 14109
rect 20989 14104 23999 14106
rect 20989 14048 20994 14104
rect 21050 14048 23938 14104
rect 23994 14048 23999 14104
rect 20989 14046 23999 14048
rect 20989 14043 21055 14046
rect 23933 14043 23999 14046
rect 4889 13968 7298 13970
rect 4889 13912 4894 13968
rect 4950 13912 7298 13968
rect 4889 13910 7298 13912
rect 8661 13970 8727 13973
rect 11145 13970 11211 13973
rect 8661 13968 11211 13970
rect 8661 13912 8666 13968
rect 8722 13912 11150 13968
rect 11206 13912 11211 13968
rect 8661 13910 11211 13912
rect 4889 13907 4955 13910
rect 8661 13907 8727 13910
rect 11145 13907 11211 13910
rect 12801 13970 12867 13973
rect 16205 13970 16271 13973
rect 12801 13968 16271 13970
rect 12801 13912 12806 13968
rect 12862 13912 16210 13968
rect 16266 13912 16271 13968
rect 12801 13910 16271 13912
rect 12801 13907 12867 13910
rect 16205 13907 16271 13910
rect 17033 13970 17099 13973
rect 21081 13970 21147 13973
rect 17033 13968 21147 13970
rect 17033 13912 17038 13968
rect 17094 13912 21086 13968
rect 21142 13912 21147 13968
rect 17033 13910 21147 13912
rect 17033 13907 17099 13910
rect 21081 13907 21147 13910
rect 21909 13970 21975 13973
rect 23289 13970 23355 13973
rect 21909 13968 23355 13970
rect 21909 13912 21914 13968
rect 21970 13912 23294 13968
rect 23350 13912 23355 13968
rect 21909 13910 23355 13912
rect 21909 13907 21975 13910
rect 23289 13907 23355 13910
rect 23565 13970 23631 13973
rect 23933 13970 23999 13973
rect 25221 13970 25287 13973
rect 23565 13968 25287 13970
rect 23565 13912 23570 13968
rect 23626 13912 23938 13968
rect 23994 13912 25226 13968
rect 25282 13912 25287 13968
rect 23565 13910 25287 13912
rect 23565 13907 23631 13910
rect 23933 13907 23999 13910
rect 25221 13907 25287 13910
rect 1577 13834 1643 13837
rect 2037 13834 2103 13837
rect 1577 13832 2103 13834
rect 1577 13776 1582 13832
rect 1638 13776 2042 13832
rect 2098 13776 2103 13832
rect 1577 13774 2103 13776
rect 1577 13771 1643 13774
rect 2037 13771 2103 13774
rect 4981 13834 5047 13837
rect 8293 13834 8359 13837
rect 4981 13832 8359 13834
rect 4981 13776 4986 13832
rect 5042 13776 8298 13832
rect 8354 13776 8359 13832
rect 4981 13774 8359 13776
rect 4981 13771 5047 13774
rect 8293 13771 8359 13774
rect 9949 13834 10015 13837
rect 12893 13834 12959 13837
rect 16941 13834 17007 13837
rect 9949 13832 17007 13834
rect 9949 13776 9954 13832
rect 10010 13776 12898 13832
rect 12954 13776 16946 13832
rect 17002 13776 17007 13832
rect 9949 13774 17007 13776
rect 9949 13771 10015 13774
rect 12893 13771 12959 13774
rect 16941 13771 17007 13774
rect 20529 13834 20595 13837
rect 21081 13836 21147 13837
rect 20846 13834 20852 13836
rect 20529 13832 20852 13834
rect 20529 13776 20534 13832
rect 20590 13776 20852 13832
rect 20529 13774 20852 13776
rect 20529 13771 20595 13774
rect 20846 13772 20852 13774
rect 20916 13772 20922 13836
rect 21030 13834 21036 13836
rect 20990 13774 21036 13834
rect 21100 13832 21147 13836
rect 26233 13834 26299 13837
rect 21142 13776 21147 13832
rect 21030 13772 21036 13774
rect 21100 13772 21147 13776
rect 21081 13771 21147 13772
rect 22326 13832 26299 13834
rect 22326 13776 26238 13832
rect 26294 13776 26299 13832
rect 22326 13774 26299 13776
rect 0 13698 480 13728
rect 1577 13698 1643 13701
rect 0 13696 1643 13698
rect 0 13640 1582 13696
rect 1638 13640 1643 13696
rect 0 13638 1643 13640
rect 0 13608 480 13638
rect 1577 13635 1643 13638
rect 3049 13698 3115 13701
rect 5206 13698 5212 13700
rect 3049 13696 5212 13698
rect 3049 13640 3054 13696
rect 3110 13640 5212 13696
rect 3049 13638 5212 13640
rect 3049 13635 3115 13638
rect 5206 13636 5212 13638
rect 5276 13636 5282 13700
rect 5441 13698 5507 13701
rect 8569 13698 8635 13701
rect 5441 13696 8635 13698
rect 5441 13640 5446 13696
rect 5502 13640 8574 13696
rect 8630 13640 8635 13696
rect 5441 13638 8635 13640
rect 5441 13635 5507 13638
rect 8569 13635 8635 13638
rect 9765 13700 9831 13701
rect 9765 13696 9812 13700
rect 9876 13698 9882 13700
rect 14365 13698 14431 13701
rect 17309 13698 17375 13701
rect 9765 13640 9770 13696
rect 9765 13636 9812 13640
rect 9876 13638 9922 13698
rect 14365 13696 17375 13698
rect 14365 13640 14370 13696
rect 14426 13640 17314 13696
rect 17370 13640 17375 13696
rect 14365 13638 17375 13640
rect 9876 13636 9882 13638
rect 9765 13635 9831 13636
rect 14365 13635 14431 13638
rect 17309 13635 17375 13638
rect 17861 13698 17927 13701
rect 19425 13698 19491 13701
rect 17861 13696 19491 13698
rect 17861 13640 17866 13696
rect 17922 13640 19430 13696
rect 19486 13640 19491 13696
rect 17861 13638 19491 13640
rect 17861 13635 17927 13638
rect 19425 13635 19491 13638
rect 20662 13636 20668 13700
rect 20732 13698 20738 13700
rect 22326 13698 22386 13774
rect 26233 13771 26299 13774
rect 20732 13638 22386 13698
rect 23013 13698 23079 13701
rect 24669 13698 24735 13701
rect 26325 13698 26391 13701
rect 27520 13698 28000 13728
rect 23013 13696 26391 13698
rect 23013 13640 23018 13696
rect 23074 13640 24674 13696
rect 24730 13640 26330 13696
rect 26386 13640 26391 13696
rect 23013 13638 26391 13640
rect 20732 13636 20738 13638
rect 23013 13635 23079 13638
rect 24669 13635 24735 13638
rect 26325 13635 26391 13638
rect 26558 13638 28000 13698
rect 10277 13632 10597 13633
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 13567 10597 13568
rect 19610 13632 19930 13633
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 19610 13567 19930 13568
rect 1485 13562 1551 13565
rect 7741 13562 7807 13565
rect 1485 13560 7807 13562
rect 1485 13504 1490 13560
rect 1546 13504 7746 13560
rect 7802 13504 7807 13560
rect 1485 13502 7807 13504
rect 1485 13499 1551 13502
rect 7741 13499 7807 13502
rect 8017 13562 8083 13565
rect 8017 13560 8954 13562
rect 8017 13504 8022 13560
rect 8078 13504 8954 13560
rect 8017 13502 8954 13504
rect 8017 13499 8083 13502
rect 3785 13426 3851 13429
rect 8753 13426 8819 13429
rect 3785 13424 8819 13426
rect 3785 13368 3790 13424
rect 3846 13368 8758 13424
rect 8814 13368 8819 13424
rect 3785 13366 8819 13368
rect 8894 13426 8954 13502
rect 9622 13500 9628 13564
rect 9692 13562 9698 13564
rect 9949 13562 10015 13565
rect 14549 13562 14615 13565
rect 9692 13560 10015 13562
rect 9692 13504 9954 13560
rect 10010 13504 10015 13560
rect 9692 13502 10015 13504
rect 9692 13500 9698 13502
rect 9949 13499 10015 13502
rect 10734 13560 14615 13562
rect 10734 13504 14554 13560
rect 14610 13504 14615 13560
rect 10734 13502 14615 13504
rect 10734 13426 10794 13502
rect 14549 13499 14615 13502
rect 14917 13562 14983 13565
rect 18505 13562 18571 13565
rect 14917 13560 18571 13562
rect 14917 13504 14922 13560
rect 14978 13504 18510 13560
rect 18566 13504 18571 13560
rect 14917 13502 18571 13504
rect 14917 13499 14983 13502
rect 18505 13499 18571 13502
rect 21449 13562 21515 13565
rect 22829 13562 22895 13565
rect 21449 13560 22895 13562
rect 21449 13504 21454 13560
rect 21510 13504 22834 13560
rect 22890 13504 22895 13560
rect 21449 13502 22895 13504
rect 21449 13499 21515 13502
rect 22829 13499 22895 13502
rect 24025 13562 24091 13565
rect 26558 13562 26618 13638
rect 27520 13608 28000 13638
rect 24025 13560 26618 13562
rect 24025 13504 24030 13560
rect 24086 13504 26618 13560
rect 24025 13502 26618 13504
rect 24025 13499 24091 13502
rect 15561 13426 15627 13429
rect 8894 13366 10794 13426
rect 10918 13424 15627 13426
rect 10918 13368 15566 13424
rect 15622 13368 15627 13424
rect 10918 13366 15627 13368
rect 3785 13363 3851 13366
rect 8753 13363 8819 13366
rect 5257 13290 5323 13293
rect 10133 13290 10199 13293
rect 5257 13288 10199 13290
rect 5257 13232 5262 13288
rect 5318 13232 10138 13288
rect 10194 13232 10199 13288
rect 5257 13230 10199 13232
rect 5257 13227 5323 13230
rect 10133 13227 10199 13230
rect 10317 13290 10383 13293
rect 10918 13290 10978 13366
rect 15561 13363 15627 13366
rect 18321 13426 18387 13429
rect 23565 13426 23631 13429
rect 18321 13424 23631 13426
rect 18321 13368 18326 13424
rect 18382 13368 23570 13424
rect 23626 13368 23631 13424
rect 18321 13366 23631 13368
rect 18321 13363 18387 13366
rect 23565 13363 23631 13366
rect 24710 13364 24716 13428
rect 24780 13426 24786 13428
rect 25129 13426 25195 13429
rect 24780 13424 25195 13426
rect 24780 13368 25134 13424
rect 25190 13368 25195 13424
rect 24780 13366 25195 13368
rect 24780 13364 24786 13366
rect 25129 13363 25195 13366
rect 10317 13288 10978 13290
rect 10317 13232 10322 13288
rect 10378 13232 10978 13288
rect 10317 13230 10978 13232
rect 11237 13290 11303 13293
rect 13077 13290 13143 13293
rect 11237 13288 13143 13290
rect 11237 13232 11242 13288
rect 11298 13232 13082 13288
rect 13138 13232 13143 13288
rect 11237 13230 13143 13232
rect 10317 13227 10383 13230
rect 11237 13227 11303 13230
rect 13077 13227 13143 13230
rect 13670 13228 13676 13292
rect 13740 13290 13746 13292
rect 13905 13290 13971 13293
rect 13740 13288 13971 13290
rect 13740 13232 13910 13288
rect 13966 13232 13971 13288
rect 13740 13230 13971 13232
rect 13740 13228 13746 13230
rect 13905 13227 13971 13230
rect 14825 13290 14891 13293
rect 15929 13290 15995 13293
rect 22369 13290 22435 13293
rect 14825 13288 15394 13290
rect 14825 13232 14830 13288
rect 14886 13232 15394 13288
rect 14825 13230 15394 13232
rect 14825 13227 14891 13230
rect 0 13154 480 13184
rect 4153 13154 4219 13157
rect 0 13152 4219 13154
rect 0 13096 4158 13152
rect 4214 13096 4219 13152
rect 0 13094 4219 13096
rect 0 13064 480 13094
rect 4153 13091 4219 13094
rect 9949 13154 10015 13157
rect 14641 13154 14707 13157
rect 9949 13152 14707 13154
rect 9949 13096 9954 13152
rect 10010 13096 14646 13152
rect 14702 13096 14707 13152
rect 9949 13094 14707 13096
rect 15334 13154 15394 13230
rect 15929 13288 22435 13290
rect 15929 13232 15934 13288
rect 15990 13232 22374 13288
rect 22430 13232 22435 13288
rect 15929 13230 22435 13232
rect 15929 13227 15995 13230
rect 22369 13227 22435 13230
rect 23565 13290 23631 13293
rect 25037 13290 25103 13293
rect 23565 13288 25103 13290
rect 23565 13232 23570 13288
rect 23626 13232 25042 13288
rect 25098 13232 25103 13288
rect 23565 13230 25103 13232
rect 23565 13227 23631 13230
rect 25037 13227 25103 13230
rect 20110 13154 20116 13156
rect 15334 13094 20116 13154
rect 9949 13091 10015 13094
rect 14641 13091 14707 13094
rect 20110 13092 20116 13094
rect 20180 13092 20186 13156
rect 20345 13154 20411 13157
rect 22829 13154 22895 13157
rect 20345 13152 22895 13154
rect 20345 13096 20350 13152
rect 20406 13096 22834 13152
rect 22890 13096 22895 13152
rect 20345 13094 22895 13096
rect 20345 13091 20411 13094
rect 22829 13091 22895 13094
rect 25957 13154 26023 13157
rect 27520 13154 28000 13184
rect 25957 13152 28000 13154
rect 25957 13096 25962 13152
rect 26018 13096 28000 13152
rect 25957 13094 28000 13096
rect 25957 13091 26023 13094
rect 5610 13088 5930 13089
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5930 13088
rect 5610 13023 5930 13024
rect 14944 13088 15264 13089
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 14944 13023 15264 13024
rect 24277 13088 24597 13089
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 27520 13064 28000 13094
rect 24277 13023 24597 13024
rect 2037 13020 2103 13021
rect 4889 13020 4955 13021
rect 2037 13018 2084 13020
rect 1992 13016 2084 13018
rect 1992 12960 2042 13016
rect 1992 12958 2084 12960
rect 2037 12956 2084 12958
rect 2148 12956 2154 13020
rect 4838 13018 4844 13020
rect 4798 12958 4844 13018
rect 4908 13016 4955 13020
rect 8385 13018 8451 13021
rect 12341 13018 12407 13021
rect 4950 12960 4955 13016
rect 4838 12956 4844 12958
rect 4908 12956 4955 12960
rect 2037 12955 2103 12956
rect 4889 12955 4955 12956
rect 5996 13016 12407 13018
rect 5996 12960 8390 13016
rect 8446 12960 12346 13016
rect 12402 12960 12407 13016
rect 5996 12958 12407 12960
rect 3969 12882 4035 12885
rect 5996 12882 6056 12958
rect 8385 12955 8451 12958
rect 12341 12955 12407 12958
rect 15878 12956 15884 13020
rect 15948 13018 15954 13020
rect 17401 13018 17467 13021
rect 17718 13018 17724 13020
rect 15948 12958 17050 13018
rect 15948 12956 15954 12958
rect 3969 12880 6056 12882
rect 3969 12824 3974 12880
rect 4030 12824 6056 12880
rect 3969 12822 6056 12824
rect 3969 12819 4035 12822
rect 6126 12820 6132 12884
rect 6196 12882 6202 12884
rect 6361 12882 6427 12885
rect 6196 12880 6427 12882
rect 6196 12824 6366 12880
rect 6422 12824 6427 12880
rect 6196 12822 6427 12824
rect 6196 12820 6202 12822
rect 6361 12819 6427 12822
rect 9765 12882 9831 12885
rect 16757 12882 16823 12885
rect 9765 12880 16823 12882
rect 9765 12824 9770 12880
rect 9826 12824 16762 12880
rect 16818 12824 16823 12880
rect 9765 12822 16823 12824
rect 16990 12882 17050 12958
rect 17401 13016 17724 13018
rect 17401 12960 17406 13016
rect 17462 12960 17724 13016
rect 17401 12958 17724 12960
rect 17401 12955 17467 12958
rect 17718 12956 17724 12958
rect 17788 12956 17794 13020
rect 19374 12956 19380 13020
rect 19444 13018 19450 13020
rect 19517 13018 19583 13021
rect 19444 13016 19583 13018
rect 19444 12960 19522 13016
rect 19578 12960 19583 13016
rect 19444 12958 19583 12960
rect 19444 12956 19450 12958
rect 19517 12955 19583 12958
rect 19701 13018 19767 13021
rect 23473 13018 23539 13021
rect 19701 13016 23539 13018
rect 19701 12960 19706 13016
rect 19762 12960 23478 13016
rect 23534 12960 23539 13016
rect 19701 12958 23539 12960
rect 19701 12955 19767 12958
rect 23473 12955 23539 12958
rect 21030 12882 21036 12884
rect 16990 12822 21036 12882
rect 9765 12819 9831 12822
rect 16757 12819 16823 12822
rect 21030 12820 21036 12822
rect 21100 12820 21106 12884
rect 25497 12882 25563 12885
rect 21222 12880 25563 12882
rect 21222 12824 25502 12880
rect 25558 12824 25563 12880
rect 21222 12822 25563 12824
rect 3877 12746 3943 12749
rect 6177 12746 6243 12749
rect 3877 12744 6243 12746
rect 3877 12688 3882 12744
rect 3938 12688 6182 12744
rect 6238 12688 6243 12744
rect 3877 12686 6243 12688
rect 3877 12683 3943 12686
rect 6177 12683 6243 12686
rect 7741 12746 7807 12749
rect 9857 12746 9923 12749
rect 10317 12746 10383 12749
rect 7741 12744 10383 12746
rect 7741 12688 7746 12744
rect 7802 12688 9862 12744
rect 9918 12688 10322 12744
rect 10378 12688 10383 12744
rect 7741 12686 10383 12688
rect 7741 12683 7807 12686
rect 9857 12683 9923 12686
rect 10317 12683 10383 12686
rect 10501 12746 10567 12749
rect 13537 12746 13603 12749
rect 10501 12744 13603 12746
rect 10501 12688 10506 12744
rect 10562 12688 13542 12744
rect 13598 12688 13603 12744
rect 10501 12686 13603 12688
rect 10501 12683 10567 12686
rect 13537 12683 13603 12686
rect 16389 12746 16455 12749
rect 20805 12746 20871 12749
rect 21222 12746 21282 12822
rect 25497 12819 25563 12822
rect 16389 12744 20132 12746
rect 16389 12688 16394 12744
rect 16450 12688 20132 12744
rect 16389 12686 20132 12688
rect 16389 12683 16455 12686
rect 0 12610 480 12640
rect 1485 12610 1551 12613
rect 0 12608 1551 12610
rect 0 12552 1490 12608
rect 1546 12552 1551 12608
rect 0 12550 1551 12552
rect 0 12520 480 12550
rect 1485 12547 1551 12550
rect 2405 12610 2471 12613
rect 9213 12610 9279 12613
rect 2405 12608 9279 12610
rect 2405 12552 2410 12608
rect 2466 12552 9218 12608
rect 9274 12552 9279 12608
rect 2405 12550 9279 12552
rect 2405 12547 2471 12550
rect 9213 12547 9279 12550
rect 12934 12548 12940 12612
rect 13004 12610 13010 12612
rect 13169 12610 13235 12613
rect 13004 12608 13235 12610
rect 13004 12552 13174 12608
rect 13230 12552 13235 12608
rect 13004 12550 13235 12552
rect 13004 12548 13010 12550
rect 13169 12547 13235 12550
rect 15009 12610 15075 12613
rect 19425 12610 19491 12613
rect 15009 12608 19491 12610
rect 15009 12552 15014 12608
rect 15070 12552 19430 12608
rect 19486 12552 19491 12608
rect 15009 12550 19491 12552
rect 15009 12547 15075 12550
rect 19425 12547 19491 12550
rect 10277 12544 10597 12545
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 12479 10597 12480
rect 19610 12544 19930 12545
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 19610 12479 19930 12480
rect 3969 12474 4035 12477
rect 8017 12474 8083 12477
rect 3969 12472 8083 12474
rect 3969 12416 3974 12472
rect 4030 12416 8022 12472
rect 8078 12416 8083 12472
rect 3969 12414 8083 12416
rect 3969 12411 4035 12414
rect 8017 12411 8083 12414
rect 10777 12474 10843 12477
rect 16389 12474 16455 12477
rect 10777 12472 16455 12474
rect 10777 12416 10782 12472
rect 10838 12416 16394 12472
rect 16450 12416 16455 12472
rect 10777 12414 16455 12416
rect 20072 12474 20132 12686
rect 20805 12744 21282 12746
rect 20805 12688 20810 12744
rect 20866 12688 21282 12744
rect 20805 12686 21282 12688
rect 20805 12683 20871 12686
rect 21950 12684 21956 12748
rect 22020 12746 22026 12748
rect 26233 12746 26299 12749
rect 22020 12744 26299 12746
rect 22020 12688 26238 12744
rect 26294 12688 26299 12744
rect 22020 12686 26299 12688
rect 22020 12684 22026 12686
rect 26233 12683 26299 12686
rect 22277 12610 22343 12613
rect 22502 12610 22508 12612
rect 22277 12608 22508 12610
rect 22277 12552 22282 12608
rect 22338 12552 22508 12608
rect 22277 12550 22508 12552
rect 22277 12547 22343 12550
rect 22502 12548 22508 12550
rect 22572 12548 22578 12612
rect 23749 12610 23815 12613
rect 24117 12610 24183 12613
rect 23749 12608 24183 12610
rect 23749 12552 23754 12608
rect 23810 12552 24122 12608
rect 24178 12552 24183 12608
rect 23749 12550 24183 12552
rect 23749 12547 23815 12550
rect 24117 12547 24183 12550
rect 24669 12610 24735 12613
rect 27520 12610 28000 12640
rect 24669 12608 28000 12610
rect 24669 12552 24674 12608
rect 24730 12552 28000 12608
rect 24669 12550 28000 12552
rect 24669 12547 24735 12550
rect 27520 12520 28000 12550
rect 24577 12474 24643 12477
rect 20072 12472 24643 12474
rect 20072 12416 24582 12472
rect 24638 12416 24643 12472
rect 20072 12414 24643 12416
rect 10777 12411 10843 12414
rect 16389 12411 16455 12414
rect 24577 12411 24643 12414
rect 25262 12412 25268 12476
rect 25332 12474 25338 12476
rect 25497 12474 25563 12477
rect 25332 12472 25563 12474
rect 25332 12416 25502 12472
rect 25558 12416 25563 12472
rect 25332 12414 25563 12416
rect 25332 12412 25338 12414
rect 25497 12411 25563 12414
rect 1393 12338 1459 12341
rect 7598 12338 7604 12340
rect 1393 12336 7604 12338
rect 1393 12280 1398 12336
rect 1454 12280 7604 12336
rect 1393 12278 7604 12280
rect 1393 12275 1459 12278
rect 7598 12276 7604 12278
rect 7668 12276 7674 12340
rect 7833 12338 7899 12341
rect 8845 12338 8911 12341
rect 13721 12338 13787 12341
rect 7833 12336 13787 12338
rect 7833 12280 7838 12336
rect 7894 12280 8850 12336
rect 8906 12280 13726 12336
rect 13782 12280 13787 12336
rect 7833 12278 13787 12280
rect 7833 12275 7899 12278
rect 8845 12275 8911 12278
rect 13721 12275 13787 12278
rect 14549 12338 14615 12341
rect 17217 12338 17283 12341
rect 14549 12336 17283 12338
rect 14549 12280 14554 12336
rect 14610 12280 17222 12336
rect 17278 12280 17283 12336
rect 14549 12278 17283 12280
rect 14549 12275 14615 12278
rect 17217 12275 17283 12278
rect 17677 12338 17743 12341
rect 26233 12338 26299 12341
rect 17677 12336 26299 12338
rect 17677 12280 17682 12336
rect 17738 12280 26238 12336
rect 26294 12280 26299 12336
rect 17677 12278 26299 12280
rect 17677 12275 17743 12278
rect 26233 12275 26299 12278
rect 2865 12202 2931 12205
rect 3182 12202 3188 12204
rect 2865 12200 3188 12202
rect 2865 12144 2870 12200
rect 2926 12144 3188 12200
rect 2865 12142 3188 12144
rect 2865 12139 2931 12142
rect 3182 12140 3188 12142
rect 3252 12202 3258 12204
rect 4153 12202 4219 12205
rect 3252 12200 4219 12202
rect 3252 12144 4158 12200
rect 4214 12144 4219 12200
rect 3252 12142 4219 12144
rect 3252 12140 3258 12142
rect 4153 12139 4219 12142
rect 4429 12202 4495 12205
rect 4705 12202 4771 12205
rect 7097 12202 7163 12205
rect 4429 12200 7163 12202
rect 4429 12144 4434 12200
rect 4490 12144 4710 12200
rect 4766 12144 7102 12200
rect 7158 12144 7163 12200
rect 4429 12142 7163 12144
rect 4429 12139 4495 12142
rect 4705 12139 4771 12142
rect 7097 12139 7163 12142
rect 8201 12202 8267 12205
rect 12433 12202 12499 12205
rect 8201 12200 12499 12202
rect 8201 12144 8206 12200
rect 8262 12144 12438 12200
rect 12494 12144 12499 12200
rect 8201 12142 12499 12144
rect 8201 12139 8267 12142
rect 12433 12139 12499 12142
rect 12893 12202 12959 12205
rect 15510 12202 15516 12204
rect 12893 12200 15516 12202
rect 12893 12144 12898 12200
rect 12954 12144 15516 12200
rect 12893 12142 15516 12144
rect 12893 12139 12959 12142
rect 15510 12140 15516 12142
rect 15580 12140 15586 12204
rect 17769 12202 17835 12205
rect 20713 12202 20779 12205
rect 17769 12200 20779 12202
rect 17769 12144 17774 12200
rect 17830 12144 20718 12200
rect 20774 12144 20779 12200
rect 17769 12142 20779 12144
rect 17769 12139 17835 12142
rect 20713 12139 20779 12142
rect 21265 12202 21331 12205
rect 21265 12200 23490 12202
rect 21265 12144 21270 12200
rect 21326 12144 23490 12200
rect 21265 12142 23490 12144
rect 21265 12139 21331 12142
rect 2773 12066 2839 12069
rect 3734 12066 3740 12068
rect 2773 12064 3740 12066
rect 2773 12008 2778 12064
rect 2834 12008 3740 12064
rect 2773 12006 3740 12008
rect 2773 12003 2839 12006
rect 3734 12004 3740 12006
rect 3804 12066 3810 12068
rect 5165 12066 5231 12069
rect 3804 12064 5231 12066
rect 3804 12008 5170 12064
rect 5226 12008 5231 12064
rect 3804 12006 5231 12008
rect 3804 12004 3810 12006
rect 5165 12003 5231 12006
rect 8845 12066 8911 12069
rect 14273 12066 14339 12069
rect 8845 12064 14339 12066
rect 8845 12008 8850 12064
rect 8906 12008 14278 12064
rect 14334 12008 14339 12064
rect 8845 12006 14339 12008
rect 8845 12003 8911 12006
rect 14273 12003 14339 12006
rect 20805 12066 20871 12069
rect 22001 12066 22067 12069
rect 20805 12064 22067 12066
rect 20805 12008 20810 12064
rect 20866 12008 22006 12064
rect 22062 12008 22067 12064
rect 20805 12006 22067 12008
rect 20805 12003 20871 12006
rect 22001 12003 22067 12006
rect 22134 12004 22140 12068
rect 22204 12066 22210 12068
rect 22369 12066 22435 12069
rect 22204 12064 22435 12066
rect 22204 12008 22374 12064
rect 22430 12008 22435 12064
rect 22204 12006 22435 12008
rect 23430 12066 23490 12142
rect 23606 12140 23612 12204
rect 23676 12202 23682 12204
rect 23974 12202 23980 12204
rect 23676 12142 23980 12202
rect 23676 12140 23682 12142
rect 23974 12140 23980 12142
rect 24044 12140 24050 12204
rect 24117 12066 24183 12069
rect 23430 12064 24183 12066
rect 23430 12008 24122 12064
rect 24178 12008 24183 12064
rect 23430 12006 24183 12008
rect 22204 12004 22210 12006
rect 22369 12003 22435 12006
rect 24117 12003 24183 12006
rect 5610 12000 5930 12001
rect 0 11930 480 11960
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5930 12000
rect 5610 11935 5930 11936
rect 14944 12000 15264 12001
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14944 11935 15264 11936
rect 24277 12000 24597 12001
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 24277 11935 24597 11936
rect 3785 11930 3851 11933
rect 7281 11932 7347 11933
rect 0 11928 3851 11930
rect 0 11872 3790 11928
rect 3846 11872 3851 11928
rect 0 11870 3851 11872
rect 0 11840 480 11870
rect 3785 11867 3851 11870
rect 7230 11868 7236 11932
rect 7300 11930 7347 11932
rect 7300 11928 7392 11930
rect 7342 11872 7392 11928
rect 7300 11870 7392 11872
rect 7300 11868 7347 11870
rect 7598 11868 7604 11932
rect 7668 11930 7674 11932
rect 12617 11930 12683 11933
rect 7668 11928 12683 11930
rect 7668 11872 12622 11928
rect 12678 11872 12683 11928
rect 7668 11870 12683 11872
rect 7668 11868 7674 11870
rect 7281 11867 7347 11868
rect 12617 11867 12683 11870
rect 18873 11930 18939 11933
rect 24117 11930 24183 11933
rect 27520 11930 28000 11960
rect 18873 11928 24183 11930
rect 18873 11872 18878 11928
rect 18934 11872 24122 11928
rect 24178 11872 24183 11928
rect 18873 11870 24183 11872
rect 18873 11867 18939 11870
rect 24117 11867 24183 11870
rect 25086 11870 28000 11930
rect 12893 11794 12959 11797
rect 1166 11792 12959 11794
rect 1166 11736 12898 11792
rect 12954 11736 12959 11792
rect 1166 11734 12959 11736
rect 0 11386 480 11416
rect 1166 11386 1226 11734
rect 12893 11731 12959 11734
rect 14038 11732 14044 11796
rect 14108 11794 14114 11796
rect 14181 11794 14247 11797
rect 14108 11792 14247 11794
rect 14108 11736 14186 11792
rect 14242 11736 14247 11792
rect 14108 11734 14247 11736
rect 14108 11732 14114 11734
rect 14181 11731 14247 11734
rect 16205 11794 16271 11797
rect 20621 11794 20687 11797
rect 24853 11794 24919 11797
rect 16205 11792 24919 11794
rect 16205 11736 16210 11792
rect 16266 11736 20626 11792
rect 20682 11736 24858 11792
rect 24914 11736 24919 11792
rect 16205 11734 24919 11736
rect 16205 11731 16271 11734
rect 20621 11731 20687 11734
rect 24853 11731 24919 11734
rect 2221 11658 2287 11661
rect 6453 11658 6519 11661
rect 2221 11656 6519 11658
rect 2221 11600 2226 11656
rect 2282 11600 6458 11656
rect 6514 11600 6519 11656
rect 2221 11598 6519 11600
rect 2221 11595 2287 11598
rect 6453 11595 6519 11598
rect 6729 11658 6795 11661
rect 8753 11658 8819 11661
rect 11513 11658 11579 11661
rect 6729 11656 8819 11658
rect 6729 11600 6734 11656
rect 6790 11600 8758 11656
rect 8814 11600 8819 11656
rect 6729 11598 8819 11600
rect 6729 11595 6795 11598
rect 8753 11595 8819 11598
rect 8894 11656 11579 11658
rect 8894 11600 11518 11656
rect 11574 11600 11579 11656
rect 8894 11598 11579 11600
rect 1393 11522 1459 11525
rect 6821 11522 6887 11525
rect 8894 11522 8954 11598
rect 11513 11595 11579 11598
rect 14590 11596 14596 11660
rect 14660 11658 14666 11660
rect 21449 11658 21515 11661
rect 14660 11656 21515 11658
rect 14660 11600 21454 11656
rect 21510 11600 21515 11656
rect 14660 11598 21515 11600
rect 14660 11596 14666 11598
rect 21449 11595 21515 11598
rect 23974 11596 23980 11660
rect 24044 11658 24050 11660
rect 24945 11658 25011 11661
rect 24044 11656 25011 11658
rect 24044 11600 24950 11656
rect 25006 11600 25011 11656
rect 24044 11598 25011 11600
rect 24044 11596 24050 11598
rect 24945 11595 25011 11598
rect 1393 11520 4354 11522
rect 1393 11464 1398 11520
rect 1454 11464 4354 11520
rect 1393 11462 4354 11464
rect 1393 11459 1459 11462
rect 0 11326 1226 11386
rect 1761 11386 1827 11389
rect 3877 11386 3943 11389
rect 1761 11384 3943 11386
rect 1761 11328 1766 11384
rect 1822 11328 3882 11384
rect 3938 11328 3943 11384
rect 1761 11326 3943 11328
rect 4294 11386 4354 11462
rect 6821 11520 8954 11522
rect 6821 11464 6826 11520
rect 6882 11464 8954 11520
rect 6821 11462 8954 11464
rect 13169 11522 13235 11525
rect 19425 11522 19491 11525
rect 13169 11520 19491 11522
rect 13169 11464 13174 11520
rect 13230 11464 19430 11520
rect 19486 11464 19491 11520
rect 13169 11462 19491 11464
rect 6821 11459 6887 11462
rect 13169 11459 13235 11462
rect 19425 11459 19491 11462
rect 20621 11522 20687 11525
rect 22318 11522 22324 11524
rect 20621 11520 22324 11522
rect 20621 11464 20626 11520
rect 20682 11464 22324 11520
rect 20621 11462 22324 11464
rect 20621 11459 20687 11462
rect 22318 11460 22324 11462
rect 22388 11460 22394 11524
rect 23422 11460 23428 11524
rect 23492 11522 23498 11524
rect 24577 11522 24643 11525
rect 23492 11520 24643 11522
rect 23492 11464 24582 11520
rect 24638 11464 24643 11520
rect 23492 11462 24643 11464
rect 23492 11460 23498 11462
rect 24577 11459 24643 11462
rect 24853 11522 24919 11525
rect 25086 11522 25146 11870
rect 27520 11840 28000 11870
rect 24853 11520 25146 11522
rect 24853 11464 24858 11520
rect 24914 11464 25146 11520
rect 24853 11462 25146 11464
rect 24853 11459 24919 11462
rect 10277 11456 10597 11457
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 11391 10597 11392
rect 19610 11456 19930 11457
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 11391 19930 11392
rect 4429 11386 4495 11389
rect 8109 11386 8175 11389
rect 11881 11386 11947 11389
rect 4294 11384 8175 11386
rect 4294 11328 4434 11384
rect 4490 11328 8114 11384
rect 8170 11328 8175 11384
rect 4294 11326 8175 11328
rect 0 11296 480 11326
rect 1761 11323 1827 11326
rect 3877 11323 3943 11326
rect 4429 11323 4495 11326
rect 8109 11323 8175 11326
rect 10734 11384 11947 11386
rect 10734 11328 11886 11384
rect 11942 11328 11947 11384
rect 10734 11326 11947 11328
rect 5165 11252 5231 11253
rect 5165 11250 5212 11252
rect 5120 11248 5212 11250
rect 5120 11192 5170 11248
rect 5120 11190 5212 11192
rect 5165 11188 5212 11190
rect 5276 11188 5282 11252
rect 5441 11250 5507 11253
rect 6453 11250 6519 11253
rect 5441 11248 6519 11250
rect 5441 11192 5446 11248
rect 5502 11192 6458 11248
rect 6514 11192 6519 11248
rect 5441 11190 6519 11192
rect 5165 11187 5231 11188
rect 5441 11187 5507 11190
rect 6453 11187 6519 11190
rect 7741 11250 7807 11253
rect 10734 11250 10794 11326
rect 11881 11323 11947 11326
rect 12617 11386 12683 11389
rect 15745 11386 15811 11389
rect 12617 11384 15811 11386
rect 12617 11328 12622 11384
rect 12678 11328 15750 11384
rect 15806 11328 15811 11384
rect 12617 11326 15811 11328
rect 12617 11323 12683 11326
rect 15745 11323 15811 11326
rect 17309 11386 17375 11389
rect 17769 11386 17835 11389
rect 17309 11384 17835 11386
rect 17309 11328 17314 11384
rect 17370 11328 17774 11384
rect 17830 11328 17835 11384
rect 17309 11326 17835 11328
rect 17309 11323 17375 11326
rect 17769 11323 17835 11326
rect 21030 11324 21036 11388
rect 21100 11386 21106 11388
rect 24945 11386 25011 11389
rect 27520 11386 28000 11416
rect 21100 11384 25011 11386
rect 21100 11328 24950 11384
rect 25006 11328 25011 11384
rect 21100 11326 25011 11328
rect 21100 11324 21106 11326
rect 24945 11323 25011 11326
rect 25638 11326 28000 11386
rect 7741 11248 10794 11250
rect 7741 11192 7746 11248
rect 7802 11192 10794 11248
rect 7741 11190 10794 11192
rect 11145 11250 11211 11253
rect 14641 11250 14707 11253
rect 11145 11248 14707 11250
rect 11145 11192 11150 11248
rect 11206 11192 14646 11248
rect 14702 11192 14707 11248
rect 11145 11190 14707 11192
rect 7741 11187 7807 11190
rect 11145 11187 11211 11190
rect 14641 11187 14707 11190
rect 15285 11250 15351 11253
rect 15878 11250 15884 11252
rect 15285 11248 15884 11250
rect 15285 11192 15290 11248
rect 15346 11192 15884 11248
rect 15285 11190 15884 11192
rect 15285 11187 15351 11190
rect 15878 11188 15884 11190
rect 15948 11188 15954 11252
rect 17493 11250 17559 11253
rect 25405 11250 25471 11253
rect 17493 11248 25471 11250
rect 17493 11192 17498 11248
rect 17554 11192 25410 11248
rect 25466 11192 25471 11248
rect 17493 11190 25471 11192
rect 17493 11187 17559 11190
rect 25405 11187 25471 11190
rect 7230 11052 7236 11116
rect 7300 11052 7306 11116
rect 10501 11114 10567 11117
rect 13721 11114 13787 11117
rect 10501 11112 13787 11114
rect 10501 11056 10506 11112
rect 10562 11056 13726 11112
rect 13782 11056 13787 11112
rect 10501 11054 13787 11056
rect 2589 10978 2655 10981
rect 4061 10978 4127 10981
rect 2589 10976 4127 10978
rect 2589 10920 2594 10976
rect 2650 10920 4066 10976
rect 4122 10920 4127 10976
rect 2589 10918 4127 10920
rect 2589 10915 2655 10918
rect 4061 10915 4127 10918
rect 7005 10978 7071 10981
rect 7238 10978 7298 11052
rect 10501 11051 10567 11054
rect 13721 11051 13787 11054
rect 13854 11052 13860 11116
rect 13924 11114 13930 11116
rect 19241 11114 19307 11117
rect 13924 11112 19307 11114
rect 13924 11056 19246 11112
rect 19302 11056 19307 11112
rect 13924 11054 19307 11056
rect 13924 11052 13930 11054
rect 19241 11051 19307 11054
rect 20069 11114 20135 11117
rect 23013 11114 23079 11117
rect 25638 11114 25698 11326
rect 27520 11296 28000 11326
rect 20069 11112 23079 11114
rect 20069 11056 20074 11112
rect 20130 11056 23018 11112
rect 23074 11056 23079 11112
rect 20069 11054 23079 11056
rect 20069 11051 20135 11054
rect 23013 11051 23079 11054
rect 25454 11054 25698 11114
rect 25454 10981 25514 11054
rect 7005 10976 7298 10978
rect 7005 10920 7010 10976
rect 7066 10920 7298 10976
rect 7005 10918 7298 10920
rect 7925 10978 7991 10981
rect 11697 10978 11763 10981
rect 7925 10976 11763 10978
rect 7925 10920 7930 10976
rect 7986 10920 11702 10976
rect 11758 10920 11763 10976
rect 7925 10918 11763 10920
rect 7005 10915 7071 10918
rect 7925 10915 7991 10918
rect 11697 10915 11763 10918
rect 12065 10978 12131 10981
rect 13629 10978 13695 10981
rect 12065 10976 13695 10978
rect 12065 10920 12070 10976
rect 12126 10920 13634 10976
rect 13690 10920 13695 10976
rect 12065 10918 13695 10920
rect 12065 10915 12131 10918
rect 13629 10915 13695 10918
rect 16113 10978 16179 10981
rect 19517 10978 19583 10981
rect 25129 10980 25195 10981
rect 25078 10978 25084 10980
rect 16113 10976 24180 10978
rect 16113 10920 16118 10976
rect 16174 10920 19522 10976
rect 19578 10920 24180 10976
rect 16113 10918 24180 10920
rect 25038 10918 25084 10978
rect 25148 10976 25195 10980
rect 25190 10920 25195 10976
rect 16113 10915 16179 10918
rect 19517 10915 19583 10918
rect 5610 10912 5930 10913
rect 0 10842 480 10872
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5930 10912
rect 5610 10847 5930 10848
rect 14944 10912 15264 10913
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 10847 15264 10848
rect 4245 10842 4311 10845
rect 0 10840 4311 10842
rect 0 10784 4250 10840
rect 4306 10784 4311 10840
rect 0 10782 4311 10784
rect 0 10752 480 10782
rect 4245 10779 4311 10782
rect 6269 10842 6335 10845
rect 12985 10842 13051 10845
rect 14457 10842 14523 10845
rect 6269 10840 14523 10842
rect 6269 10784 6274 10840
rect 6330 10784 12990 10840
rect 13046 10784 14462 10840
rect 14518 10784 14523 10840
rect 6269 10782 14523 10784
rect 6269 10779 6335 10782
rect 12985 10779 13051 10782
rect 14457 10779 14523 10782
rect 16021 10842 16087 10845
rect 18321 10842 18387 10845
rect 16021 10840 18387 10842
rect 16021 10784 16026 10840
rect 16082 10784 18326 10840
rect 18382 10784 18387 10840
rect 16021 10782 18387 10784
rect 16021 10779 16087 10782
rect 18321 10779 18387 10782
rect 18505 10842 18571 10845
rect 23473 10842 23539 10845
rect 18505 10840 23539 10842
rect 18505 10784 18510 10840
rect 18566 10784 23478 10840
rect 23534 10784 23539 10840
rect 18505 10782 23539 10784
rect 18505 10779 18571 10782
rect 23473 10779 23539 10782
rect 3877 10706 3943 10709
rect 6494 10706 6500 10708
rect 3877 10704 6500 10706
rect 3877 10648 3882 10704
rect 3938 10648 6500 10704
rect 3877 10646 6500 10648
rect 3877 10643 3943 10646
rect 6494 10644 6500 10646
rect 6564 10644 6570 10708
rect 7833 10706 7899 10709
rect 12249 10706 12315 10709
rect 7833 10704 12315 10706
rect 7833 10648 7838 10704
rect 7894 10648 12254 10704
rect 12310 10648 12315 10704
rect 7833 10646 12315 10648
rect 7833 10643 7899 10646
rect 12249 10643 12315 10646
rect 13169 10706 13235 10709
rect 15193 10706 15259 10709
rect 13169 10704 15259 10706
rect 13169 10648 13174 10704
rect 13230 10648 15198 10704
rect 15254 10648 15259 10704
rect 13169 10646 15259 10648
rect 13169 10643 13235 10646
rect 15193 10643 15259 10646
rect 17861 10706 17927 10709
rect 21541 10706 21607 10709
rect 17861 10704 21607 10706
rect 17861 10648 17866 10704
rect 17922 10648 21546 10704
rect 21602 10648 21607 10704
rect 17861 10646 21607 10648
rect 17861 10643 17927 10646
rect 21541 10643 21607 10646
rect 21909 10706 21975 10709
rect 23933 10706 23999 10709
rect 21909 10704 23999 10706
rect 21909 10648 21914 10704
rect 21970 10648 23938 10704
rect 23994 10648 23999 10704
rect 21909 10646 23999 10648
rect 24120 10706 24180 10918
rect 25078 10916 25084 10918
rect 25148 10916 25195 10920
rect 25129 10915 25195 10916
rect 25405 10976 25514 10981
rect 25405 10920 25410 10976
rect 25466 10920 25514 10976
rect 25405 10918 25514 10920
rect 25405 10915 25471 10918
rect 24277 10912 24597 10913
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 10847 24597 10848
rect 27520 10842 28000 10872
rect 24672 10782 28000 10842
rect 24672 10706 24732 10782
rect 27520 10752 28000 10782
rect 24120 10646 24732 10706
rect 21909 10643 21975 10646
rect 23933 10643 23999 10646
rect 4838 10508 4844 10572
rect 4908 10570 4914 10572
rect 5809 10570 5875 10573
rect 8845 10570 8911 10573
rect 4908 10568 8911 10570
rect 4908 10512 5814 10568
rect 5870 10512 8850 10568
rect 8906 10512 8911 10568
rect 4908 10510 8911 10512
rect 4908 10508 4914 10510
rect 5809 10507 5875 10510
rect 8845 10507 8911 10510
rect 9673 10570 9739 10573
rect 10910 10570 10916 10572
rect 9673 10568 10916 10570
rect 9673 10512 9678 10568
rect 9734 10512 10916 10568
rect 9673 10510 10916 10512
rect 9673 10507 9739 10510
rect 10910 10508 10916 10510
rect 10980 10508 10986 10572
rect 15377 10570 15443 10573
rect 15377 10568 26986 10570
rect 15377 10512 15382 10568
rect 15438 10512 26986 10568
rect 15377 10510 26986 10512
rect 15377 10507 15443 10510
rect 1393 10434 1459 10437
rect 1761 10434 1827 10437
rect 5901 10434 5967 10437
rect 1393 10432 5967 10434
rect 1393 10376 1398 10432
rect 1454 10376 1766 10432
rect 1822 10376 5906 10432
rect 5962 10376 5967 10432
rect 1393 10374 5967 10376
rect 1393 10371 1459 10374
rect 1761 10371 1827 10374
rect 5901 10371 5967 10374
rect 6494 10372 6500 10436
rect 6564 10434 6570 10436
rect 9305 10434 9371 10437
rect 6564 10432 9371 10434
rect 6564 10376 9310 10432
rect 9366 10376 9371 10432
rect 6564 10374 9371 10376
rect 6564 10372 6570 10374
rect 9305 10371 9371 10374
rect 20110 10372 20116 10436
rect 20180 10434 20186 10436
rect 22277 10434 22343 10437
rect 20180 10432 22343 10434
rect 20180 10376 22282 10432
rect 22338 10376 22343 10432
rect 20180 10374 22343 10376
rect 20180 10372 20186 10374
rect 22277 10371 22343 10374
rect 22461 10434 22527 10437
rect 26325 10434 26391 10437
rect 22461 10432 26391 10434
rect 22461 10376 22466 10432
rect 22522 10376 26330 10432
rect 26386 10376 26391 10432
rect 22461 10374 26391 10376
rect 22461 10371 22527 10374
rect 26325 10371 26391 10374
rect 10277 10368 10597 10369
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 10303 10597 10304
rect 19610 10368 19930 10369
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19610 10303 19930 10304
rect 1710 10236 1716 10300
rect 1780 10298 1786 10300
rect 2405 10298 2471 10301
rect 1780 10296 2471 10298
rect 1780 10240 2410 10296
rect 2466 10240 2471 10296
rect 1780 10238 2471 10240
rect 1780 10236 1786 10238
rect 2405 10235 2471 10238
rect 2773 10298 2839 10301
rect 8109 10298 8175 10301
rect 2773 10296 8175 10298
rect 2773 10240 2778 10296
rect 2834 10240 8114 10296
rect 8170 10240 8175 10296
rect 2773 10238 8175 10240
rect 2773 10235 2839 10238
rect 8109 10235 8175 10238
rect 10910 10236 10916 10300
rect 10980 10298 10986 10300
rect 13629 10298 13695 10301
rect 10980 10296 13695 10298
rect 10980 10240 13634 10296
rect 13690 10240 13695 10296
rect 10980 10238 13695 10240
rect 10980 10236 10986 10238
rect 13629 10235 13695 10238
rect 14549 10298 14615 10301
rect 18413 10298 18479 10301
rect 14549 10296 18479 10298
rect 14549 10240 14554 10296
rect 14610 10240 18418 10296
rect 18474 10240 18479 10296
rect 14549 10238 18479 10240
rect 14549 10235 14615 10238
rect 18413 10235 18479 10238
rect 20069 10298 20135 10301
rect 23473 10298 23539 10301
rect 20069 10296 23539 10298
rect 20069 10240 20074 10296
rect 20130 10240 23478 10296
rect 23534 10240 23539 10296
rect 20069 10238 23539 10240
rect 20069 10235 20135 10238
rect 23473 10235 23539 10238
rect 26325 10298 26391 10301
rect 26734 10298 26740 10300
rect 26325 10296 26740 10298
rect 26325 10240 26330 10296
rect 26386 10240 26740 10296
rect 26325 10238 26740 10240
rect 26325 10235 26391 10238
rect 26734 10236 26740 10238
rect 26804 10236 26810 10300
rect 0 10162 480 10192
rect 4797 10162 4863 10165
rect 6126 10162 6132 10164
rect 0 10102 4354 10162
rect 0 10072 480 10102
rect 2037 10026 2103 10029
rect 2773 10026 2839 10029
rect 3049 10028 3115 10029
rect 2037 10024 2839 10026
rect 2037 9968 2042 10024
rect 2098 9968 2778 10024
rect 2834 9968 2839 10024
rect 2037 9966 2839 9968
rect 2037 9963 2103 9966
rect 2773 9963 2839 9966
rect 2998 9964 3004 10028
rect 3068 10026 3115 10028
rect 4294 10026 4354 10102
rect 4797 10160 6132 10162
rect 4797 10104 4802 10160
rect 4858 10104 6132 10160
rect 4797 10102 6132 10104
rect 4797 10099 4863 10102
rect 6126 10100 6132 10102
rect 6196 10100 6202 10164
rect 6545 10162 6611 10165
rect 7097 10162 7163 10165
rect 11881 10162 11947 10165
rect 6545 10160 11947 10162
rect 6545 10104 6550 10160
rect 6606 10104 7102 10160
rect 7158 10104 11886 10160
rect 11942 10104 11947 10160
rect 6545 10102 11947 10104
rect 6545 10099 6611 10102
rect 7097 10099 7163 10102
rect 11881 10099 11947 10102
rect 17861 10162 17927 10165
rect 24025 10162 24091 10165
rect 17861 10160 24091 10162
rect 17861 10104 17866 10160
rect 17922 10104 24030 10160
rect 24086 10104 24091 10160
rect 17861 10102 24091 10104
rect 26926 10162 26986 10510
rect 27520 10162 28000 10192
rect 26926 10102 28000 10162
rect 17861 10099 17927 10102
rect 24025 10099 24091 10102
rect 27520 10072 28000 10102
rect 6494 10026 6500 10028
rect 3068 10024 3160 10026
rect 3110 9968 3160 10024
rect 3068 9966 3160 9968
rect 4294 9966 6500 10026
rect 3068 9964 3115 9966
rect 6494 9964 6500 9966
rect 6564 9964 6570 10028
rect 6637 10026 6703 10029
rect 9949 10026 10015 10029
rect 12065 10026 12131 10029
rect 16389 10026 16455 10029
rect 18965 10026 19031 10029
rect 19425 10026 19491 10029
rect 6637 10024 10015 10026
rect 6637 9968 6642 10024
rect 6698 9968 9954 10024
rect 10010 9968 10015 10024
rect 6637 9966 10015 9968
rect 3049 9963 3115 9964
rect 6637 9963 6703 9966
rect 9949 9963 10015 9966
rect 10136 10024 12131 10026
rect 10136 9968 12070 10024
rect 12126 9968 12131 10024
rect 10136 9966 12131 9968
rect 6453 9890 6519 9893
rect 10136 9890 10196 9966
rect 12065 9963 12131 9966
rect 14782 10024 19491 10026
rect 14782 9968 16394 10024
rect 16450 9968 18970 10024
rect 19026 9968 19430 10024
rect 19486 9968 19491 10024
rect 14782 9966 19491 9968
rect 6453 9888 10196 9890
rect 6453 9832 6458 9888
rect 6514 9832 10196 9888
rect 6453 9830 10196 9832
rect 10777 9890 10843 9893
rect 13445 9890 13511 9893
rect 10777 9888 13511 9890
rect 10777 9832 10782 9888
rect 10838 9832 13450 9888
rect 13506 9832 13511 9888
rect 10777 9830 13511 9832
rect 6453 9827 6519 9830
rect 10777 9827 10843 9830
rect 13445 9827 13511 9830
rect 5610 9824 5930 9825
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5930 9824
rect 5610 9759 5930 9760
rect 2313 9754 2379 9757
rect 4613 9754 4679 9757
rect 2313 9752 4679 9754
rect 2313 9696 2318 9752
rect 2374 9696 4618 9752
rect 4674 9696 4679 9752
rect 2313 9694 4679 9696
rect 2313 9691 2379 9694
rect 4613 9691 4679 9694
rect 6637 9756 6703 9757
rect 6637 9752 6684 9756
rect 6748 9754 6754 9756
rect 7557 9754 7623 9757
rect 14782 9754 14842 9966
rect 16389 9963 16455 9966
rect 18965 9963 19031 9966
rect 19425 9963 19491 9966
rect 21357 10026 21423 10029
rect 25313 10026 25379 10029
rect 21357 10024 25379 10026
rect 21357 9968 21362 10024
rect 21418 9968 25318 10024
rect 25374 9968 25379 10024
rect 21357 9966 25379 9968
rect 21357 9963 21423 9966
rect 25313 9963 25379 9966
rect 15745 9890 15811 9893
rect 20713 9890 20779 9893
rect 15745 9888 20779 9890
rect 15745 9832 15750 9888
rect 15806 9832 20718 9888
rect 20774 9832 20779 9888
rect 15745 9830 20779 9832
rect 15745 9827 15811 9830
rect 20713 9827 20779 9830
rect 14944 9824 15264 9825
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 14944 9759 15264 9760
rect 24277 9824 24597 9825
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 24277 9759 24597 9760
rect 6637 9696 6642 9752
rect 6637 9692 6684 9696
rect 6748 9694 6794 9754
rect 7557 9752 14842 9754
rect 7557 9696 7562 9752
rect 7618 9696 14842 9752
rect 7557 9694 14842 9696
rect 19198 9694 19810 9754
rect 6748 9692 6754 9694
rect 6637 9691 6703 9692
rect 7557 9691 7623 9694
rect 0 9618 480 9648
rect 3233 9618 3299 9621
rect 6729 9618 6795 9621
rect 0 9558 2698 9618
rect 0 9528 480 9558
rect 1945 9482 2011 9485
rect 2497 9482 2563 9485
rect 1945 9480 2563 9482
rect 1945 9424 1950 9480
rect 2006 9424 2502 9480
rect 2558 9424 2563 9480
rect 1945 9422 2563 9424
rect 1945 9419 2011 9422
rect 2497 9419 2563 9422
rect 2638 9210 2698 9558
rect 3233 9616 6795 9618
rect 3233 9560 3238 9616
rect 3294 9560 6734 9616
rect 6790 9560 6795 9616
rect 3233 9558 6795 9560
rect 3233 9555 3299 9558
rect 6729 9555 6795 9558
rect 9254 9556 9260 9620
rect 9324 9618 9330 9620
rect 9397 9618 9463 9621
rect 9324 9616 9463 9618
rect 9324 9560 9402 9616
rect 9458 9560 9463 9616
rect 9324 9558 9463 9560
rect 9324 9556 9330 9558
rect 9397 9555 9463 9558
rect 9581 9618 9647 9621
rect 15745 9618 15811 9621
rect 17769 9618 17835 9621
rect 19198 9618 19258 9694
rect 19425 9620 19491 9621
rect 9581 9616 15624 9618
rect 9581 9560 9586 9616
rect 9642 9560 15624 9616
rect 9581 9558 15624 9560
rect 9581 9555 9647 9558
rect 2773 9482 2839 9485
rect 3601 9482 3667 9485
rect 4981 9482 5047 9485
rect 2773 9480 5047 9482
rect 2773 9424 2778 9480
rect 2834 9424 3606 9480
rect 3662 9424 4986 9480
rect 5042 9424 5047 9480
rect 2773 9422 5047 9424
rect 2773 9419 2839 9422
rect 3601 9419 3667 9422
rect 4981 9419 5047 9422
rect 9397 9482 9463 9485
rect 15564 9482 15624 9558
rect 15745 9616 19258 9618
rect 15745 9560 15750 9616
rect 15806 9560 17774 9616
rect 17830 9560 19258 9616
rect 15745 9558 19258 9560
rect 15745 9555 15811 9558
rect 17769 9555 17835 9558
rect 19374 9556 19380 9620
rect 19444 9618 19491 9620
rect 19750 9618 19810 9694
rect 22645 9618 22711 9621
rect 19444 9616 19536 9618
rect 19486 9560 19536 9616
rect 19444 9558 19536 9560
rect 19750 9616 22711 9618
rect 19750 9560 22650 9616
rect 22706 9560 22711 9616
rect 19750 9558 22711 9560
rect 19444 9556 19491 9558
rect 19425 9555 19491 9556
rect 22645 9555 22711 9558
rect 22870 9556 22876 9620
rect 22940 9618 22946 9620
rect 24577 9618 24643 9621
rect 22940 9616 24643 9618
rect 22940 9560 24582 9616
rect 24638 9560 24643 9616
rect 22940 9558 24643 9560
rect 22940 9556 22946 9558
rect 24577 9555 24643 9558
rect 25446 9556 25452 9620
rect 25516 9618 25522 9620
rect 25589 9618 25655 9621
rect 26325 9620 26391 9621
rect 26325 9618 26372 9620
rect 25516 9616 25655 9618
rect 25516 9560 25594 9616
rect 25650 9560 25655 9616
rect 25516 9558 25655 9560
rect 26280 9616 26372 9618
rect 26280 9560 26330 9616
rect 26280 9558 26372 9560
rect 25516 9556 25522 9558
rect 25589 9555 25655 9558
rect 26325 9556 26372 9558
rect 26436 9556 26442 9620
rect 27520 9618 28000 9648
rect 26558 9558 28000 9618
rect 26325 9555 26391 9556
rect 15837 9482 15903 9485
rect 9397 9480 10794 9482
rect 9397 9424 9402 9480
rect 9458 9424 10794 9480
rect 9397 9422 10794 9424
rect 15564 9480 15903 9482
rect 15564 9424 15842 9480
rect 15898 9424 15903 9480
rect 15564 9422 15903 9424
rect 9397 9419 9463 9422
rect 7005 9346 7071 9349
rect 5030 9344 7071 9346
rect 5030 9288 7010 9344
rect 7066 9288 7071 9344
rect 5030 9286 7071 9288
rect 10734 9346 10794 9422
rect 15837 9419 15903 9422
rect 19057 9482 19123 9485
rect 20713 9482 20779 9485
rect 19057 9480 20779 9482
rect 19057 9424 19062 9480
rect 19118 9424 20718 9480
rect 20774 9424 20779 9480
rect 19057 9422 20779 9424
rect 19057 9419 19123 9422
rect 20713 9419 20779 9422
rect 21173 9482 21239 9485
rect 24853 9482 24919 9485
rect 21173 9480 24919 9482
rect 21173 9424 21178 9480
rect 21234 9424 24858 9480
rect 24914 9424 24919 9480
rect 21173 9422 24919 9424
rect 21173 9419 21239 9422
rect 24853 9419 24919 9422
rect 13854 9346 13860 9348
rect 10734 9286 13860 9346
rect 5030 9210 5090 9286
rect 7005 9283 7071 9286
rect 13854 9284 13860 9286
rect 13924 9284 13930 9348
rect 15377 9346 15443 9349
rect 17401 9346 17467 9349
rect 15377 9344 17467 9346
rect 15377 9288 15382 9344
rect 15438 9288 17406 9344
rect 17462 9288 17467 9344
rect 15377 9286 17467 9288
rect 15377 9283 15443 9286
rect 17401 9283 17467 9286
rect 18413 9346 18479 9349
rect 19333 9346 19399 9349
rect 18413 9344 19399 9346
rect 18413 9288 18418 9344
rect 18474 9288 19338 9344
rect 19394 9288 19399 9344
rect 18413 9286 19399 9288
rect 18413 9283 18479 9286
rect 19333 9283 19399 9286
rect 20662 9284 20668 9348
rect 20732 9346 20738 9348
rect 21173 9346 21239 9349
rect 20732 9344 21239 9346
rect 20732 9288 21178 9344
rect 21234 9288 21239 9344
rect 20732 9286 21239 9288
rect 20732 9284 20738 9286
rect 21173 9283 21239 9286
rect 21633 9346 21699 9349
rect 24393 9346 24459 9349
rect 21633 9344 24459 9346
rect 21633 9288 21638 9344
rect 21694 9288 24398 9344
rect 24454 9288 24459 9344
rect 21633 9286 24459 9288
rect 21633 9283 21699 9286
rect 24393 9283 24459 9286
rect 10277 9280 10597 9281
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 9215 10597 9216
rect 19610 9280 19930 9281
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 9215 19930 9216
rect 2638 9150 5090 9210
rect 5257 9210 5323 9213
rect 9213 9210 9279 9213
rect 5257 9208 9279 9210
rect 5257 9152 5262 9208
rect 5318 9152 9218 9208
rect 9274 9152 9279 9208
rect 5257 9150 9279 9152
rect 5257 9147 5323 9150
rect 9213 9147 9279 9150
rect 13537 9210 13603 9213
rect 14273 9210 14339 9213
rect 17585 9210 17651 9213
rect 13537 9208 17651 9210
rect 13537 9152 13542 9208
rect 13598 9152 14278 9208
rect 14334 9152 17590 9208
rect 17646 9152 17651 9208
rect 13537 9150 17651 9152
rect 13537 9147 13603 9150
rect 14273 9147 14339 9150
rect 17585 9147 17651 9150
rect 21214 9148 21220 9212
rect 21284 9210 21290 9212
rect 21357 9210 21423 9213
rect 21284 9208 21423 9210
rect 21284 9152 21362 9208
rect 21418 9152 21423 9208
rect 21284 9150 21423 9152
rect 21284 9148 21290 9150
rect 21357 9147 21423 9150
rect 21541 9210 21607 9213
rect 21950 9210 21956 9212
rect 21541 9208 21956 9210
rect 21541 9152 21546 9208
rect 21602 9152 21956 9208
rect 21541 9150 21956 9152
rect 21541 9147 21607 9150
rect 21950 9148 21956 9150
rect 22020 9148 22026 9212
rect 23381 9210 23447 9213
rect 25129 9210 25195 9213
rect 23381 9208 25195 9210
rect 23381 9152 23386 9208
rect 23442 9152 25134 9208
rect 25190 9152 25195 9208
rect 23381 9150 25195 9152
rect 23381 9147 23447 9150
rect 25129 9147 25195 9150
rect 0 9074 480 9104
rect 3141 9074 3207 9077
rect 0 9072 3207 9074
rect 0 9016 3146 9072
rect 3202 9016 3207 9072
rect 0 9014 3207 9016
rect 0 8984 480 9014
rect 3141 9011 3207 9014
rect 11329 9074 11395 9077
rect 15377 9074 15443 9077
rect 11329 9072 15443 9074
rect 11329 9016 11334 9072
rect 11390 9016 15382 9072
rect 15438 9016 15443 9072
rect 11329 9014 15443 9016
rect 11329 9011 11395 9014
rect 15377 9011 15443 9014
rect 15837 9074 15903 9077
rect 19149 9074 19215 9077
rect 23289 9074 23355 9077
rect 15837 9072 23355 9074
rect 15837 9016 15842 9072
rect 15898 9016 19154 9072
rect 19210 9016 23294 9072
rect 23350 9016 23355 9072
rect 15837 9014 23355 9016
rect 15837 9011 15903 9014
rect 19149 9011 19215 9014
rect 23289 9011 23355 9014
rect 23974 9012 23980 9076
rect 24044 9074 24050 9076
rect 24853 9074 24919 9077
rect 24044 9072 24919 9074
rect 24044 9016 24858 9072
rect 24914 9016 24919 9072
rect 24044 9014 24919 9016
rect 24044 9012 24050 9014
rect 24853 9011 24919 9014
rect 1761 8938 1827 8941
rect 2446 8938 2452 8940
rect 1761 8936 2452 8938
rect 1761 8880 1766 8936
rect 1822 8880 2452 8936
rect 1761 8878 2452 8880
rect 1761 8875 1827 8878
rect 2446 8876 2452 8878
rect 2516 8938 2522 8940
rect 2681 8938 2747 8941
rect 2516 8936 2747 8938
rect 2516 8880 2686 8936
rect 2742 8880 2747 8936
rect 2516 8878 2747 8880
rect 2516 8876 2522 8878
rect 2681 8875 2747 8878
rect 4889 8938 4955 8941
rect 15653 8938 15719 8941
rect 18045 8938 18111 8941
rect 22921 8938 22987 8941
rect 26558 8938 26618 9558
rect 27520 9528 28000 9558
rect 27520 9074 28000 9104
rect 4889 8936 15578 8938
rect 4889 8880 4894 8936
rect 4950 8880 15578 8936
rect 4889 8878 15578 8880
rect 4889 8875 4955 8878
rect 5257 8802 5323 8805
rect 5390 8802 5396 8804
rect 5257 8800 5396 8802
rect 5257 8744 5262 8800
rect 5318 8744 5396 8800
rect 5257 8742 5396 8744
rect 5257 8739 5323 8742
rect 5390 8740 5396 8742
rect 5460 8740 5466 8804
rect 7465 8802 7531 8805
rect 14641 8802 14707 8805
rect 7465 8800 14707 8802
rect 7465 8744 7470 8800
rect 7526 8744 14646 8800
rect 14702 8744 14707 8800
rect 7465 8742 14707 8744
rect 15518 8802 15578 8878
rect 15653 8936 22987 8938
rect 15653 8880 15658 8936
rect 15714 8880 18050 8936
rect 18106 8880 22926 8936
rect 22982 8880 22987 8936
rect 15653 8878 22987 8880
rect 15653 8875 15719 8878
rect 18045 8875 18111 8878
rect 22921 8875 22987 8878
rect 24120 8878 26618 8938
rect 26742 9014 28000 9074
rect 16297 8802 16363 8805
rect 15518 8800 16363 8802
rect 15518 8744 16302 8800
rect 16358 8744 16363 8800
rect 15518 8742 16363 8744
rect 7465 8739 7531 8742
rect 14641 8739 14707 8742
rect 16297 8739 16363 8742
rect 19885 8802 19951 8805
rect 21449 8802 21515 8805
rect 21817 8804 21883 8805
rect 19885 8800 21515 8802
rect 19885 8744 19890 8800
rect 19946 8744 21454 8800
rect 21510 8744 21515 8800
rect 19885 8742 21515 8744
rect 19885 8739 19951 8742
rect 21449 8739 21515 8742
rect 21766 8740 21772 8804
rect 21836 8802 21883 8804
rect 22001 8802 22067 8805
rect 24120 8802 24180 8878
rect 21836 8800 21928 8802
rect 21878 8744 21928 8800
rect 21836 8742 21928 8744
rect 22001 8800 24180 8802
rect 22001 8744 22006 8800
rect 22062 8744 24180 8800
rect 22001 8742 24180 8744
rect 24669 8802 24735 8805
rect 26742 8802 26802 9014
rect 27520 8984 28000 9014
rect 24669 8800 26802 8802
rect 24669 8744 24674 8800
rect 24730 8744 26802 8800
rect 24669 8742 26802 8744
rect 21836 8740 21883 8742
rect 21817 8739 21883 8740
rect 22001 8739 22067 8742
rect 24669 8739 24735 8742
rect 5610 8736 5930 8737
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5930 8736
rect 5610 8671 5930 8672
rect 14944 8736 15264 8737
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 8671 15264 8672
rect 24277 8736 24597 8737
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 8671 24597 8672
rect 8477 8666 8543 8669
rect 16113 8666 16179 8669
rect 19057 8666 19123 8669
rect 19885 8666 19951 8669
rect 8477 8664 14520 8666
rect 8477 8608 8482 8664
rect 8538 8608 14520 8664
rect 8477 8606 14520 8608
rect 8477 8603 8543 8606
rect 0 8530 480 8560
rect 565 8530 631 8533
rect 0 8528 631 8530
rect 0 8472 570 8528
rect 626 8472 631 8528
rect 0 8470 631 8472
rect 0 8440 480 8470
rect 565 8467 631 8470
rect 3325 8530 3391 8533
rect 8661 8530 8727 8533
rect 3325 8528 8727 8530
rect 3325 8472 3330 8528
rect 3386 8472 8666 8528
rect 8722 8472 8727 8528
rect 3325 8470 8727 8472
rect 3325 8467 3391 8470
rect 8661 8467 8727 8470
rect 8845 8530 8911 8533
rect 14460 8530 14520 8606
rect 16113 8664 19123 8666
rect 16113 8608 16118 8664
rect 16174 8608 19062 8664
rect 19118 8608 19123 8664
rect 19382 8664 19951 8666
rect 19382 8632 19890 8664
rect 16113 8606 19123 8608
rect 16113 8603 16179 8606
rect 19057 8603 19123 8606
rect 19336 8608 19890 8632
rect 19946 8608 19951 8664
rect 19336 8606 19951 8608
rect 19336 8572 19442 8606
rect 19885 8603 19951 8606
rect 20069 8666 20135 8669
rect 26325 8666 26391 8669
rect 27286 8666 27292 8668
rect 20069 8664 23858 8666
rect 20069 8608 20074 8664
rect 20130 8608 23858 8664
rect 20069 8606 23858 8608
rect 20069 8603 20135 8606
rect 19336 8564 19396 8572
rect 19244 8530 19396 8564
rect 8845 8528 11162 8530
rect 8845 8472 8850 8528
rect 8906 8472 11162 8528
rect 8845 8470 11162 8472
rect 14460 8504 19396 8530
rect 20621 8532 20687 8533
rect 20621 8528 20668 8532
rect 20732 8530 20738 8532
rect 21265 8530 21331 8533
rect 23657 8530 23723 8533
rect 14460 8470 19304 8504
rect 20621 8472 20626 8528
rect 8845 8467 8911 8470
rect 1853 8394 1919 8397
rect 4061 8394 4127 8397
rect 6269 8394 6335 8397
rect 1853 8392 6335 8394
rect 1853 8336 1858 8392
rect 1914 8336 4066 8392
rect 4122 8336 6274 8392
rect 6330 8336 6335 8392
rect 1853 8334 6335 8336
rect 1853 8331 1919 8334
rect 4061 8331 4127 8334
rect 6269 8331 6335 8334
rect 6545 8394 6611 8397
rect 7465 8394 7531 8397
rect 6545 8392 7531 8394
rect 6545 8336 6550 8392
rect 6606 8336 7470 8392
rect 7526 8336 7531 8392
rect 6545 8334 7531 8336
rect 6545 8331 6611 8334
rect 7465 8331 7531 8334
rect 8201 8394 8267 8397
rect 8201 8392 10978 8394
rect 8201 8336 8206 8392
rect 8262 8336 10978 8392
rect 8201 8334 10978 8336
rect 8201 8331 8267 8334
rect 10918 8261 10978 8334
rect 8150 8258 8156 8260
rect 1350 8198 8156 8258
rect 0 7850 480 7880
rect 1350 7850 1410 8198
rect 8150 8196 8156 8198
rect 8220 8196 8226 8260
rect 10918 8256 11027 8261
rect 10918 8200 10966 8256
rect 11022 8200 11027 8256
rect 10918 8198 11027 8200
rect 11102 8258 11162 8470
rect 20621 8468 20668 8472
rect 20732 8470 20778 8530
rect 21265 8528 23723 8530
rect 21265 8472 21270 8528
rect 21326 8472 23662 8528
rect 23718 8472 23723 8528
rect 21265 8470 23723 8472
rect 23798 8530 23858 8606
rect 26325 8664 27292 8666
rect 26325 8608 26330 8664
rect 26386 8608 27292 8664
rect 26325 8606 27292 8608
rect 26325 8603 26391 8606
rect 27286 8604 27292 8606
rect 27356 8604 27362 8668
rect 24853 8530 24919 8533
rect 27520 8530 28000 8560
rect 23798 8528 24919 8530
rect 23798 8472 24858 8528
rect 24914 8472 24919 8528
rect 23798 8470 24919 8472
rect 20732 8468 20738 8470
rect 20621 8467 20687 8468
rect 21265 8467 21331 8470
rect 23657 8467 23723 8470
rect 24853 8467 24919 8470
rect 25086 8470 28000 8530
rect 15561 8396 15627 8397
rect 15510 8332 15516 8396
rect 15580 8394 15627 8396
rect 18505 8394 18571 8397
rect 15580 8392 15672 8394
rect 15622 8336 15672 8392
rect 15580 8334 15672 8336
rect 18505 8392 21834 8394
rect 18505 8336 18510 8392
rect 18566 8336 21834 8392
rect 18505 8334 21834 8336
rect 15580 8332 15627 8334
rect 15561 8331 15627 8332
rect 18505 8331 18571 8334
rect 13077 8258 13143 8261
rect 11102 8256 13143 8258
rect 11102 8200 13082 8256
rect 13138 8200 13143 8256
rect 11102 8198 13143 8200
rect 21774 8258 21834 8334
rect 21950 8332 21956 8396
rect 22020 8394 22026 8396
rect 23013 8394 23079 8397
rect 22020 8392 23079 8394
rect 22020 8336 23018 8392
rect 23074 8336 23079 8392
rect 22020 8334 23079 8336
rect 22020 8332 22026 8334
rect 23013 8331 23079 8334
rect 23197 8394 23263 8397
rect 25086 8394 25146 8470
rect 27520 8440 28000 8470
rect 23197 8392 25146 8394
rect 23197 8336 23202 8392
rect 23258 8336 25146 8392
rect 23197 8334 25146 8336
rect 23197 8331 23263 8334
rect 23933 8258 23999 8261
rect 21774 8256 23999 8258
rect 21774 8200 23938 8256
rect 23994 8200 23999 8256
rect 21774 8198 23999 8200
rect 10961 8195 11027 8198
rect 13077 8195 13143 8198
rect 23933 8195 23999 8198
rect 24894 8196 24900 8260
rect 24964 8258 24970 8260
rect 25865 8258 25931 8261
rect 24964 8256 25931 8258
rect 24964 8200 25870 8256
rect 25926 8200 25931 8256
rect 24964 8198 25931 8200
rect 24964 8196 24970 8198
rect 25865 8195 25931 8198
rect 10277 8192 10597 8193
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 10277 8127 10597 8128
rect 19610 8192 19930 8193
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 19610 8127 19930 8128
rect 2405 8122 2471 8125
rect 9990 8122 9996 8124
rect 2405 8120 9996 8122
rect 2405 8064 2410 8120
rect 2466 8064 9996 8120
rect 2405 8062 9996 8064
rect 2405 8059 2471 8062
rect 9990 8060 9996 8062
rect 10060 8060 10066 8124
rect 17861 8122 17927 8125
rect 19425 8122 19491 8125
rect 17861 8120 19491 8122
rect 17861 8064 17866 8120
rect 17922 8064 19430 8120
rect 19486 8064 19491 8120
rect 17861 8062 19491 8064
rect 17861 8059 17927 8062
rect 19425 8059 19491 8062
rect 20069 8122 20135 8125
rect 22870 8122 22876 8124
rect 20069 8120 22876 8122
rect 20069 8064 20074 8120
rect 20130 8064 22876 8120
rect 20069 8062 22876 8064
rect 20069 8059 20135 8062
rect 22870 8060 22876 8062
rect 22940 8060 22946 8124
rect 23105 8122 23171 8125
rect 25221 8122 25287 8125
rect 23105 8120 25287 8122
rect 23105 8064 23110 8120
rect 23166 8064 25226 8120
rect 25282 8064 25287 8120
rect 23105 8062 25287 8064
rect 23105 8059 23171 8062
rect 25221 8059 25287 8062
rect 4337 7986 4403 7989
rect 7189 7986 7255 7989
rect 4337 7984 7255 7986
rect 4337 7928 4342 7984
rect 4398 7928 7194 7984
rect 7250 7928 7255 7984
rect 4337 7926 7255 7928
rect 4337 7923 4403 7926
rect 7189 7923 7255 7926
rect 7741 7986 7807 7989
rect 19885 7986 19951 7989
rect 7741 7984 19951 7986
rect 7741 7928 7746 7984
rect 7802 7928 19890 7984
rect 19946 7928 19951 7984
rect 7741 7926 19951 7928
rect 7741 7923 7807 7926
rect 19885 7923 19951 7926
rect 20345 7986 20411 7989
rect 22921 7986 22987 7989
rect 20345 7984 22987 7986
rect 20345 7928 20350 7984
rect 20406 7928 22926 7984
rect 22982 7928 22987 7984
rect 20345 7926 22987 7928
rect 20345 7923 20411 7926
rect 22921 7923 22987 7926
rect 0 7790 1410 7850
rect 1577 7850 1643 7853
rect 14733 7850 14799 7853
rect 19241 7850 19307 7853
rect 1577 7848 14799 7850
rect 1577 7792 1582 7848
rect 1638 7792 14738 7848
rect 14794 7792 14799 7848
rect 1577 7790 14799 7792
rect 0 7760 480 7790
rect 1577 7787 1643 7790
rect 14733 7787 14799 7790
rect 15702 7848 19307 7850
rect 15702 7792 19246 7848
rect 19302 7792 19307 7848
rect 15702 7790 19307 7792
rect 5610 7648 5930 7649
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5930 7648
rect 5610 7583 5930 7584
rect 14944 7648 15264 7649
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 7583 15264 7584
rect 2814 7516 2820 7580
rect 2884 7578 2890 7580
rect 3141 7578 3207 7581
rect 2884 7576 3207 7578
rect 2884 7520 3146 7576
rect 3202 7520 3207 7576
rect 2884 7518 3207 7520
rect 2884 7516 2890 7518
rect 3141 7515 3207 7518
rect 7649 7578 7715 7581
rect 14733 7578 14799 7581
rect 7649 7576 14799 7578
rect 7649 7520 7654 7576
rect 7710 7520 14738 7576
rect 14794 7520 14799 7576
rect 7649 7518 14799 7520
rect 7649 7515 7715 7518
rect 14733 7515 14799 7518
rect 2221 7442 2287 7445
rect 15702 7442 15762 7790
rect 19241 7787 19307 7790
rect 19374 7788 19380 7852
rect 19444 7850 19450 7852
rect 20069 7850 20135 7853
rect 19444 7848 20135 7850
rect 19444 7792 20074 7848
rect 20130 7792 20135 7848
rect 19444 7790 20135 7792
rect 19444 7788 19450 7790
rect 20069 7787 20135 7790
rect 20989 7850 21055 7853
rect 21633 7850 21699 7853
rect 27520 7850 28000 7880
rect 20989 7848 28000 7850
rect 20989 7792 20994 7848
rect 21050 7792 21638 7848
rect 21694 7792 28000 7848
rect 20989 7790 28000 7792
rect 20989 7787 21055 7790
rect 21633 7787 21699 7790
rect 27520 7760 28000 7790
rect 17718 7652 17724 7716
rect 17788 7714 17794 7716
rect 20345 7714 20411 7717
rect 17788 7712 20411 7714
rect 17788 7656 20350 7712
rect 20406 7656 20411 7712
rect 17788 7654 20411 7656
rect 17788 7652 17794 7654
rect 20345 7651 20411 7654
rect 25773 7714 25839 7717
rect 25773 7712 26618 7714
rect 25773 7656 25778 7712
rect 25834 7656 26618 7712
rect 25773 7654 26618 7656
rect 25773 7651 25839 7654
rect 24277 7648 24597 7649
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 7583 24597 7584
rect 15837 7578 15903 7581
rect 23381 7578 23447 7581
rect 25773 7580 25839 7581
rect 25773 7578 25820 7580
rect 15837 7576 23447 7578
rect 15837 7520 15842 7576
rect 15898 7520 23386 7576
rect 23442 7520 23447 7576
rect 15837 7518 23447 7520
rect 25728 7576 25820 7578
rect 25728 7520 25778 7576
rect 25728 7518 25820 7520
rect 15837 7515 15903 7518
rect 23381 7515 23447 7518
rect 25773 7516 25820 7518
rect 25884 7516 25890 7580
rect 25773 7515 25839 7516
rect 25681 7442 25747 7445
rect 2221 7440 15762 7442
rect 2221 7384 2226 7440
rect 2282 7384 15762 7440
rect 2221 7382 15762 7384
rect 17174 7440 25747 7442
rect 17174 7384 25686 7440
rect 25742 7384 25747 7440
rect 17174 7382 25747 7384
rect 2221 7379 2287 7382
rect 0 7306 480 7336
rect 1669 7306 1735 7309
rect 0 7304 1735 7306
rect 0 7248 1674 7304
rect 1730 7248 1735 7304
rect 0 7246 1735 7248
rect 0 7216 480 7246
rect 1669 7243 1735 7246
rect 2405 7306 2471 7309
rect 17174 7306 17234 7382
rect 25681 7379 25747 7382
rect 26417 7306 26483 7309
rect 2405 7304 17234 7306
rect 2405 7248 2410 7304
rect 2466 7248 17234 7304
rect 2405 7246 17234 7248
rect 17358 7304 26483 7306
rect 17358 7248 26422 7304
rect 26478 7248 26483 7304
rect 17358 7246 26483 7248
rect 26558 7306 26618 7654
rect 27520 7306 28000 7336
rect 26558 7246 28000 7306
rect 2405 7243 2471 7246
rect 4705 7170 4771 7173
rect 5390 7170 5396 7172
rect 4705 7168 5396 7170
rect 4705 7112 4710 7168
rect 4766 7112 5396 7168
rect 4705 7110 5396 7112
rect 4705 7107 4771 7110
rect 5390 7108 5396 7110
rect 5460 7108 5466 7172
rect 10685 7170 10751 7173
rect 17358 7170 17418 7246
rect 26417 7243 26483 7246
rect 27520 7216 28000 7246
rect 10685 7168 17418 7170
rect 10685 7112 10690 7168
rect 10746 7112 17418 7168
rect 10685 7110 17418 7112
rect 22737 7170 22803 7173
rect 22737 7168 23674 7170
rect 22737 7112 22742 7168
rect 22798 7112 23674 7168
rect 22737 7110 23674 7112
rect 10685 7107 10751 7110
rect 22737 7107 22803 7110
rect 10277 7104 10597 7105
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 10277 7039 10597 7040
rect 19610 7104 19930 7105
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 7039 19930 7040
rect 1393 7034 1459 7037
rect 4337 7034 4403 7037
rect 1393 7032 4403 7034
rect 1393 6976 1398 7032
rect 1454 6976 4342 7032
rect 4398 6976 4403 7032
rect 1393 6974 4403 6976
rect 1393 6971 1459 6974
rect 4337 6971 4403 6974
rect 4521 7034 4587 7037
rect 10133 7034 10199 7037
rect 16205 7034 16271 7037
rect 4521 7032 10199 7034
rect 4521 6976 4526 7032
rect 4582 6976 10138 7032
rect 10194 6976 10199 7032
rect 4521 6974 10199 6976
rect 4521 6971 4587 6974
rect 10133 6971 10199 6974
rect 14782 7032 16271 7034
rect 14782 6976 16210 7032
rect 16266 6976 16271 7032
rect 14782 6974 16271 6976
rect 3969 6898 4035 6901
rect 5809 6898 5875 6901
rect 3969 6896 5875 6898
rect 3969 6840 3974 6896
rect 4030 6840 5814 6896
rect 5870 6840 5875 6896
rect 3969 6838 5875 6840
rect 3969 6835 4035 6838
rect 5809 6835 5875 6838
rect 8661 6898 8727 6901
rect 12065 6898 12131 6901
rect 8661 6896 12131 6898
rect 8661 6840 8666 6896
rect 8722 6840 12070 6896
rect 12126 6840 12131 6896
rect 8661 6838 12131 6840
rect 8661 6835 8727 6838
rect 12065 6835 12131 6838
rect 0 6762 480 6792
rect 2037 6762 2103 6765
rect 0 6760 2103 6762
rect 0 6704 2042 6760
rect 2098 6704 2103 6760
rect 0 6702 2103 6704
rect 0 6672 480 6702
rect 2037 6699 2103 6702
rect 2865 6762 2931 6765
rect 5625 6762 5691 6765
rect 2865 6760 5691 6762
rect 2865 6704 2870 6760
rect 2926 6704 5630 6760
rect 5686 6704 5691 6760
rect 2865 6702 5691 6704
rect 2865 6699 2931 6702
rect 5625 6699 5691 6702
rect 8109 6762 8175 6765
rect 12801 6762 12867 6765
rect 8109 6760 12867 6762
rect 8109 6704 8114 6760
rect 8170 6704 12806 6760
rect 12862 6704 12867 6760
rect 8109 6702 12867 6704
rect 8109 6699 8175 6702
rect 12801 6699 12867 6702
rect 10409 6626 10475 6629
rect 10726 6626 10732 6628
rect 10409 6624 10732 6626
rect 10409 6568 10414 6624
rect 10470 6568 10732 6624
rect 10409 6566 10732 6568
rect 10409 6563 10475 6566
rect 10726 6564 10732 6566
rect 10796 6564 10802 6628
rect 5610 6560 5930 6561
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5930 6560
rect 5610 6495 5930 6496
rect 8017 6490 8083 6493
rect 14782 6490 14842 6974
rect 16205 6971 16271 6974
rect 20345 7034 20411 7037
rect 23473 7034 23539 7037
rect 20345 7032 23539 7034
rect 20345 6976 20350 7032
rect 20406 6976 23478 7032
rect 23534 6976 23539 7032
rect 20345 6974 23539 6976
rect 20345 6971 20411 6974
rect 23473 6971 23539 6974
rect 14917 6898 14983 6901
rect 21909 6898 21975 6901
rect 14917 6896 21975 6898
rect 14917 6840 14922 6896
rect 14978 6840 21914 6896
rect 21970 6840 21975 6896
rect 14917 6838 21975 6840
rect 23614 6898 23674 7110
rect 25262 7108 25268 7172
rect 25332 7170 25338 7172
rect 26049 7170 26115 7173
rect 25332 7168 26115 7170
rect 25332 7112 26054 7168
rect 26110 7112 26115 7168
rect 25332 7110 26115 7112
rect 25332 7108 25338 7110
rect 26049 7107 26115 7110
rect 24945 7036 25011 7037
rect 24894 7034 24900 7036
rect 24854 6974 24900 7034
rect 24964 7032 25011 7036
rect 25006 6976 25011 7032
rect 24894 6972 24900 6974
rect 24964 6972 25011 6976
rect 24945 6971 25011 6972
rect 24761 6898 24827 6901
rect 23614 6896 24827 6898
rect 23614 6840 24766 6896
rect 24822 6840 24827 6896
rect 23614 6838 24827 6840
rect 14917 6835 14983 6838
rect 21909 6835 21975 6838
rect 24761 6835 24827 6838
rect 15009 6762 15075 6765
rect 17125 6762 17191 6765
rect 20345 6764 20411 6765
rect 15009 6760 17191 6762
rect 15009 6704 15014 6760
rect 15070 6704 17130 6760
rect 17186 6704 17191 6760
rect 15009 6702 17191 6704
rect 15009 6699 15075 6702
rect 17125 6699 17191 6702
rect 20294 6700 20300 6764
rect 20364 6762 20411 6764
rect 20621 6764 20687 6765
rect 20621 6762 20668 6764
rect 20364 6760 20456 6762
rect 20406 6704 20456 6760
rect 20364 6702 20456 6704
rect 20576 6760 20668 6762
rect 20576 6704 20626 6760
rect 20576 6702 20668 6704
rect 20364 6700 20411 6702
rect 20345 6699 20411 6700
rect 20621 6700 20668 6702
rect 20732 6700 20738 6764
rect 21081 6762 21147 6765
rect 23565 6762 23631 6765
rect 27520 6762 28000 6792
rect 21081 6760 23631 6762
rect 21081 6704 21086 6760
rect 21142 6704 23570 6760
rect 23626 6704 23631 6760
rect 21081 6702 23631 6704
rect 20621 6699 20687 6700
rect 21081 6699 21147 6702
rect 23565 6699 23631 6702
rect 23798 6702 28000 6762
rect 16481 6626 16547 6629
rect 21950 6626 21956 6628
rect 16481 6624 21956 6626
rect 16481 6568 16486 6624
rect 16542 6568 21956 6624
rect 16481 6566 21956 6568
rect 16481 6563 16547 6566
rect 21950 6564 21956 6566
rect 22020 6564 22026 6628
rect 22553 6626 22619 6629
rect 23798 6626 23858 6702
rect 27520 6672 28000 6702
rect 22553 6624 23858 6626
rect 22553 6568 22558 6624
rect 22614 6568 23858 6624
rect 22553 6566 23858 6568
rect 22553 6563 22619 6566
rect 14944 6560 15264 6561
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 6495 15264 6496
rect 24277 6560 24597 6561
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 6495 24597 6496
rect 8017 6488 14842 6490
rect 8017 6432 8022 6488
rect 8078 6432 14842 6488
rect 8017 6430 14842 6432
rect 15377 6490 15443 6493
rect 17125 6490 17191 6493
rect 20253 6490 20319 6493
rect 15377 6488 17050 6490
rect 15377 6432 15382 6488
rect 15438 6432 17050 6488
rect 15377 6430 17050 6432
rect 8017 6427 8083 6430
rect 15377 6427 15443 6430
rect 6729 6354 6795 6357
rect 8385 6354 8451 6357
rect 14549 6354 14615 6357
rect 6729 6352 8451 6354
rect 6729 6296 6734 6352
rect 6790 6296 8390 6352
rect 8446 6296 8451 6352
rect 6729 6294 8451 6296
rect 6729 6291 6795 6294
rect 8385 6291 8451 6294
rect 14230 6352 14615 6354
rect 14230 6296 14554 6352
rect 14610 6296 14615 6352
rect 14230 6294 14615 6296
rect 5165 6218 5231 6221
rect 5349 6218 5415 6221
rect 9990 6218 9996 6220
rect 5165 6216 9996 6218
rect 5165 6160 5170 6216
rect 5226 6160 5354 6216
rect 5410 6160 9996 6216
rect 5165 6158 9996 6160
rect 5165 6155 5231 6158
rect 5349 6155 5415 6158
rect 9990 6156 9996 6158
rect 10060 6156 10066 6220
rect 14230 6218 14290 6294
rect 14549 6291 14615 6294
rect 14733 6354 14799 6357
rect 16849 6354 16915 6357
rect 14733 6352 16915 6354
rect 14733 6296 14738 6352
rect 14794 6296 16854 6352
rect 16910 6296 16915 6352
rect 14733 6294 16915 6296
rect 16990 6354 17050 6430
rect 17125 6488 20319 6490
rect 17125 6432 17130 6488
rect 17186 6432 20258 6488
rect 20314 6432 20319 6488
rect 17125 6430 20319 6432
rect 17125 6427 17191 6430
rect 20253 6427 20319 6430
rect 20662 6428 20668 6492
rect 20732 6490 20738 6492
rect 21173 6490 21239 6493
rect 20732 6488 21239 6490
rect 20732 6432 21178 6488
rect 21234 6432 21239 6488
rect 20732 6430 21239 6432
rect 20732 6428 20738 6430
rect 21173 6427 21239 6430
rect 21541 6492 21607 6493
rect 21541 6488 21588 6492
rect 21652 6490 21658 6492
rect 24761 6490 24827 6493
rect 21541 6432 21546 6488
rect 21541 6428 21588 6432
rect 21652 6430 21698 6490
rect 24761 6488 25698 6490
rect 24761 6432 24766 6488
rect 24822 6432 25698 6488
rect 24761 6430 25698 6432
rect 21652 6428 21658 6430
rect 21541 6427 21607 6428
rect 24761 6427 24827 6430
rect 19333 6354 19399 6357
rect 16990 6352 19399 6354
rect 16990 6296 19338 6352
rect 19394 6296 19399 6352
rect 16990 6294 19399 6296
rect 14733 6291 14799 6294
rect 16849 6291 16915 6294
rect 19333 6291 19399 6294
rect 19517 6354 19583 6357
rect 22277 6354 22343 6357
rect 19517 6352 22343 6354
rect 19517 6296 19522 6352
rect 19578 6296 22282 6352
rect 22338 6296 22343 6352
rect 19517 6294 22343 6296
rect 19517 6291 19583 6294
rect 22277 6291 22343 6294
rect 10136 6158 14290 6218
rect 14457 6218 14523 6221
rect 22001 6218 22067 6221
rect 14457 6216 22067 6218
rect 14457 6160 14462 6216
rect 14518 6160 22006 6216
rect 22062 6160 22067 6216
rect 14457 6158 22067 6160
rect 0 6082 480 6112
rect 3601 6082 3667 6085
rect 0 6080 3667 6082
rect 0 6024 3606 6080
rect 3662 6024 3667 6080
rect 0 6022 3667 6024
rect 0 5992 480 6022
rect 3601 6019 3667 6022
rect 2313 5946 2379 5949
rect 6269 5946 6335 5949
rect 10136 5946 10196 6158
rect 14457 6155 14523 6158
rect 22001 6155 22067 6158
rect 22737 6218 22803 6221
rect 24761 6218 24827 6221
rect 22737 6216 24827 6218
rect 22737 6160 22742 6216
rect 22798 6160 24766 6216
rect 24822 6160 24827 6216
rect 22737 6158 24827 6160
rect 22737 6155 22803 6158
rect 24761 6155 24827 6158
rect 10685 6082 10751 6085
rect 15101 6082 15167 6085
rect 10685 6080 15167 6082
rect 10685 6024 10690 6080
rect 10746 6024 15106 6080
rect 15162 6024 15167 6080
rect 10685 6022 15167 6024
rect 10685 6019 10751 6022
rect 15101 6019 15167 6022
rect 15285 6082 15351 6085
rect 18505 6082 18571 6085
rect 15285 6080 18571 6082
rect 15285 6024 15290 6080
rect 15346 6024 18510 6080
rect 18566 6024 18571 6080
rect 15285 6022 18571 6024
rect 15285 6019 15351 6022
rect 18505 6019 18571 6022
rect 22870 6020 22876 6084
rect 22940 6082 22946 6084
rect 23013 6082 23079 6085
rect 22940 6080 23079 6082
rect 22940 6024 23018 6080
rect 23074 6024 23079 6080
rect 22940 6022 23079 6024
rect 22940 6020 22946 6022
rect 23013 6019 23079 6022
rect 23933 6082 23999 6085
rect 25405 6082 25471 6085
rect 23933 6080 25471 6082
rect 23933 6024 23938 6080
rect 23994 6024 25410 6080
rect 25466 6024 25471 6080
rect 23933 6022 25471 6024
rect 25638 6082 25698 6430
rect 27520 6082 28000 6112
rect 25638 6022 28000 6082
rect 23933 6019 23999 6022
rect 25405 6019 25471 6022
rect 10277 6016 10597 6017
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 5951 10597 5952
rect 19610 6016 19930 6017
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 27520 5992 28000 6022
rect 19610 5951 19930 5952
rect 2313 5944 6335 5946
rect 2313 5888 2318 5944
rect 2374 5888 6274 5944
rect 6330 5888 6335 5944
rect 2313 5886 6335 5888
rect 2313 5883 2379 5886
rect 6269 5883 6335 5886
rect 7606 5886 10196 5946
rect 10777 5946 10843 5949
rect 12617 5946 12683 5949
rect 10777 5944 12683 5946
rect 10777 5888 10782 5944
rect 10838 5888 12622 5944
rect 12678 5888 12683 5944
rect 10777 5886 12683 5888
rect 1485 5810 1551 5813
rect 2313 5810 2379 5813
rect 2681 5810 2747 5813
rect 7606 5810 7666 5886
rect 10777 5883 10843 5886
rect 12617 5883 12683 5886
rect 13721 5946 13787 5949
rect 18321 5946 18387 5949
rect 13721 5944 18387 5946
rect 13721 5888 13726 5944
rect 13782 5888 18326 5944
rect 18382 5888 18387 5944
rect 13721 5886 18387 5888
rect 13721 5883 13787 5886
rect 18321 5883 18387 5886
rect 21357 5946 21423 5949
rect 26233 5946 26299 5949
rect 21357 5944 26299 5946
rect 21357 5888 21362 5944
rect 21418 5888 26238 5944
rect 26294 5888 26299 5944
rect 21357 5886 26299 5888
rect 21357 5883 21423 5886
rect 26233 5883 26299 5886
rect 1485 5808 7666 5810
rect 1485 5752 1490 5808
rect 1546 5752 2318 5808
rect 2374 5752 2686 5808
rect 2742 5752 7666 5808
rect 1485 5750 7666 5752
rect 8201 5810 8267 5813
rect 10685 5810 10751 5813
rect 8201 5808 10751 5810
rect 8201 5752 8206 5808
rect 8262 5752 10690 5808
rect 10746 5752 10751 5808
rect 8201 5750 10751 5752
rect 1485 5747 1551 5750
rect 2313 5747 2379 5750
rect 2681 5747 2747 5750
rect 8201 5747 8267 5750
rect 10685 5747 10751 5750
rect 13445 5810 13511 5813
rect 15009 5810 15075 5813
rect 13445 5808 15075 5810
rect 13445 5752 13450 5808
rect 13506 5752 15014 5808
rect 15070 5752 15075 5808
rect 13445 5750 15075 5752
rect 13445 5747 13511 5750
rect 15009 5747 15075 5750
rect 15193 5810 15259 5813
rect 25773 5810 25839 5813
rect 15193 5808 17786 5810
rect 15193 5752 15198 5808
rect 15254 5752 17786 5808
rect 15193 5750 17786 5752
rect 15193 5747 15259 5750
rect 2589 5674 2655 5677
rect 3693 5674 3759 5677
rect 4061 5676 4127 5677
rect 4061 5674 4108 5676
rect 2589 5672 3759 5674
rect 2589 5616 2594 5672
rect 2650 5616 3698 5672
rect 3754 5616 3759 5672
rect 2589 5614 3759 5616
rect 4016 5672 4108 5674
rect 4016 5616 4066 5672
rect 4016 5614 4108 5616
rect 2589 5611 2655 5614
rect 3693 5611 3759 5614
rect 4061 5612 4108 5614
rect 4172 5612 4178 5676
rect 4061 5611 4127 5612
rect 0 5538 480 5568
rect 8201 5538 8267 5541
rect 0 5478 4906 5538
rect 0 5448 480 5478
rect 4846 5266 4906 5478
rect 8201 5536 14842 5538
rect 8201 5480 8206 5536
rect 8262 5480 14842 5536
rect 8201 5478 14842 5480
rect 8201 5475 8267 5478
rect 5610 5472 5930 5473
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5930 5472
rect 5610 5407 5930 5408
rect 9121 5402 9187 5405
rect 11145 5402 11211 5405
rect 9121 5400 11211 5402
rect 9121 5344 9126 5400
rect 9182 5344 11150 5400
rect 11206 5344 11211 5400
rect 9121 5342 11211 5344
rect 9121 5339 9187 5342
rect 11145 5339 11211 5342
rect 12382 5340 12388 5404
rect 12452 5402 12458 5404
rect 12617 5402 12683 5405
rect 13169 5402 13235 5405
rect 12452 5400 13235 5402
rect 12452 5344 12622 5400
rect 12678 5344 13174 5400
rect 13230 5344 13235 5400
rect 12452 5342 13235 5344
rect 12452 5340 12458 5342
rect 12617 5339 12683 5342
rect 13169 5339 13235 5342
rect 13629 5266 13695 5269
rect 4846 5264 13695 5266
rect 4846 5208 13634 5264
rect 13690 5208 13695 5264
rect 4846 5206 13695 5208
rect 14782 5266 14842 5478
rect 14944 5472 15264 5473
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 14944 5407 15264 5408
rect 17726 5402 17786 5750
rect 19382 5808 25839 5810
rect 19382 5752 25778 5808
rect 25834 5752 25839 5808
rect 19382 5750 25839 5752
rect 18413 5538 18479 5541
rect 19382 5538 19442 5750
rect 25773 5747 25839 5750
rect 21725 5674 21791 5677
rect 24025 5674 24091 5677
rect 21725 5672 24091 5674
rect 21725 5616 21730 5672
rect 21786 5616 24030 5672
rect 24086 5616 24091 5672
rect 21725 5614 24091 5616
rect 21725 5611 21791 5614
rect 24025 5611 24091 5614
rect 18413 5536 19442 5538
rect 18413 5480 18418 5536
rect 18474 5480 19442 5536
rect 18413 5478 19442 5480
rect 18413 5475 18479 5478
rect 23606 5476 23612 5540
rect 23676 5538 23682 5540
rect 24025 5538 24091 5541
rect 27520 5538 28000 5568
rect 23676 5536 24091 5538
rect 23676 5480 24030 5536
rect 24086 5480 24091 5536
rect 23676 5478 24091 5480
rect 23676 5476 23682 5478
rect 24025 5475 24091 5478
rect 24902 5478 28000 5538
rect 24277 5472 24597 5473
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 5407 24597 5408
rect 21357 5402 21423 5405
rect 17726 5400 21423 5402
rect 17726 5344 21362 5400
rect 21418 5344 21423 5400
rect 17726 5342 21423 5344
rect 21357 5339 21423 5342
rect 21541 5402 21607 5405
rect 21541 5400 24180 5402
rect 21541 5344 21546 5400
rect 21602 5344 24180 5400
rect 21541 5342 24180 5344
rect 21541 5339 21607 5342
rect 18597 5266 18663 5269
rect 14782 5264 18663 5266
rect 14782 5208 18602 5264
rect 18658 5208 18663 5264
rect 14782 5206 18663 5208
rect 13629 5203 13695 5206
rect 18597 5203 18663 5206
rect 19425 5266 19491 5269
rect 23749 5266 23815 5269
rect 19425 5264 23815 5266
rect 19425 5208 19430 5264
rect 19486 5208 23754 5264
rect 23810 5208 23815 5264
rect 19425 5206 23815 5208
rect 24120 5266 24180 5342
rect 24902 5266 24962 5478
rect 27520 5448 28000 5478
rect 24120 5206 24962 5266
rect 19425 5203 19491 5206
rect 23749 5203 23815 5206
rect 1945 5130 2011 5133
rect 2078 5130 2084 5132
rect 1945 5128 2084 5130
rect 1945 5072 1950 5128
rect 2006 5072 2084 5128
rect 1945 5070 2084 5072
rect 1945 5067 2011 5070
rect 2078 5068 2084 5070
rect 2148 5068 2154 5132
rect 4705 5130 4771 5133
rect 6361 5130 6427 5133
rect 8109 5132 8175 5133
rect 8109 5130 8156 5132
rect 4705 5128 6427 5130
rect 4705 5072 4710 5128
rect 4766 5072 6366 5128
rect 6422 5072 6427 5128
rect 4705 5070 6427 5072
rect 8064 5128 8156 5130
rect 8064 5072 8114 5128
rect 8064 5070 8156 5072
rect 4705 5067 4771 5070
rect 6361 5067 6427 5070
rect 8109 5068 8156 5070
rect 8220 5068 8226 5132
rect 9305 5130 9371 5133
rect 19517 5130 19583 5133
rect 9305 5128 19583 5130
rect 9305 5072 9310 5128
rect 9366 5072 19522 5128
rect 19578 5072 19583 5128
rect 9305 5070 19583 5072
rect 8109 5067 8175 5068
rect 9305 5067 9371 5070
rect 19517 5067 19583 5070
rect 21633 5130 21699 5133
rect 25681 5130 25747 5133
rect 21633 5128 25747 5130
rect 21633 5072 21638 5128
rect 21694 5072 25686 5128
rect 25742 5072 25747 5128
rect 21633 5070 25747 5072
rect 21633 5067 21699 5070
rect 25681 5067 25747 5070
rect 0 4994 480 5024
rect 7465 4994 7531 4997
rect 0 4992 7531 4994
rect 0 4936 7470 4992
rect 7526 4936 7531 4992
rect 0 4934 7531 4936
rect 0 4904 480 4934
rect 7465 4931 7531 4934
rect 11789 4994 11855 4997
rect 18413 4994 18479 4997
rect 11789 4992 18479 4994
rect 11789 4936 11794 4992
rect 11850 4936 18418 4992
rect 18474 4936 18479 4992
rect 11789 4934 18479 4936
rect 11789 4931 11855 4934
rect 18413 4931 18479 4934
rect 21173 4994 21239 4997
rect 23657 4994 23723 4997
rect 21173 4992 23723 4994
rect 21173 4936 21178 4992
rect 21234 4936 23662 4992
rect 23718 4936 23723 4992
rect 21173 4934 23723 4936
rect 21173 4931 21239 4934
rect 23657 4931 23723 4934
rect 25681 4994 25747 4997
rect 27520 4994 28000 5024
rect 25681 4992 28000 4994
rect 25681 4936 25686 4992
rect 25742 4936 28000 4992
rect 25681 4934 28000 4936
rect 25681 4931 25747 4934
rect 10277 4928 10597 4929
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 10277 4863 10597 4864
rect 19610 4928 19930 4929
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 27520 4904 28000 4934
rect 19610 4863 19930 4864
rect 6085 4858 6151 4861
rect 8569 4858 8635 4861
rect 9622 4858 9628 4860
rect 6085 4856 9628 4858
rect 6085 4800 6090 4856
rect 6146 4800 8574 4856
rect 8630 4800 9628 4856
rect 6085 4798 9628 4800
rect 6085 4795 6151 4798
rect 8569 4795 8635 4798
rect 9622 4796 9628 4798
rect 9692 4796 9698 4860
rect 10777 4858 10843 4861
rect 12382 4858 12388 4860
rect 10777 4856 12388 4858
rect 10777 4800 10782 4856
rect 10838 4800 12388 4856
rect 10777 4798 12388 4800
rect 10777 4795 10843 4798
rect 12382 4796 12388 4798
rect 12452 4796 12458 4860
rect 12617 4858 12683 4861
rect 18597 4858 18663 4861
rect 19057 4858 19123 4861
rect 12617 4856 19123 4858
rect 12617 4800 12622 4856
rect 12678 4800 18602 4856
rect 18658 4800 19062 4856
rect 19118 4800 19123 4856
rect 12617 4798 19123 4800
rect 12617 4795 12683 4798
rect 18597 4795 18663 4798
rect 19057 4795 19123 4798
rect 22829 4858 22895 4861
rect 25037 4858 25103 4861
rect 22829 4856 25103 4858
rect 22829 4800 22834 4856
rect 22890 4800 25042 4856
rect 25098 4800 25103 4856
rect 22829 4798 25103 4800
rect 22829 4795 22895 4798
rect 25037 4795 25103 4798
rect 6637 4724 6703 4725
rect 6637 4722 6684 4724
rect 6592 4720 6684 4722
rect 6592 4664 6642 4720
rect 6592 4662 6684 4664
rect 6637 4660 6684 4662
rect 6748 4660 6754 4724
rect 9254 4660 9260 4724
rect 9324 4722 9330 4724
rect 9397 4722 9463 4725
rect 9324 4720 9463 4722
rect 9324 4664 9402 4720
rect 9458 4664 9463 4720
rect 9324 4662 9463 4664
rect 9324 4660 9330 4662
rect 6637 4659 6703 4660
rect 9397 4659 9463 4662
rect 9949 4722 10015 4725
rect 20989 4722 21055 4725
rect 9949 4720 21055 4722
rect 9949 4664 9954 4720
rect 10010 4664 20994 4720
rect 21050 4664 21055 4720
rect 9949 4662 21055 4664
rect 9949 4659 10015 4662
rect 20989 4659 21055 4662
rect 23790 4660 23796 4724
rect 23860 4722 23866 4724
rect 24117 4722 24183 4725
rect 24485 4722 24551 4725
rect 23860 4720 24551 4722
rect 23860 4664 24122 4720
rect 24178 4664 24490 4720
rect 24546 4664 24551 4720
rect 23860 4662 24551 4664
rect 23860 4660 23866 4662
rect 24117 4659 24183 4662
rect 24485 4659 24551 4662
rect 24761 4722 24827 4725
rect 24761 4720 26066 4722
rect 24761 4664 24766 4720
rect 24822 4664 26066 4720
rect 24761 4662 26066 4664
rect 24761 4659 24827 4662
rect 1577 4586 1643 4589
rect 13169 4586 13235 4589
rect 1577 4584 13235 4586
rect 1577 4528 1582 4584
rect 1638 4528 13174 4584
rect 13230 4528 13235 4584
rect 1577 4526 13235 4528
rect 1577 4523 1643 4526
rect 13169 4523 13235 4526
rect 14457 4586 14523 4589
rect 18505 4586 18571 4589
rect 25773 4586 25839 4589
rect 14457 4584 15394 4586
rect 14457 4528 14462 4584
rect 14518 4528 15394 4584
rect 14457 4526 15394 4528
rect 14457 4523 14523 4526
rect 0 4450 480 4480
rect 749 4450 815 4453
rect 0 4448 815 4450
rect 0 4392 754 4448
rect 810 4392 815 4448
rect 0 4390 815 4392
rect 0 4360 480 4390
rect 749 4387 815 4390
rect 6821 4450 6887 4453
rect 11145 4450 11211 4453
rect 6821 4448 11211 4450
rect 6821 4392 6826 4448
rect 6882 4392 11150 4448
rect 11206 4392 11211 4448
rect 6821 4390 11211 4392
rect 6821 4387 6887 4390
rect 11145 4387 11211 4390
rect 5610 4384 5930 4385
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5930 4384
rect 5610 4319 5930 4320
rect 14944 4384 15264 4385
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 14944 4319 15264 4320
rect 11237 4314 11303 4317
rect 6134 4312 11303 4314
rect 6134 4256 11242 4312
rect 11298 4256 11303 4312
rect 6134 4254 11303 4256
rect 4061 4178 4127 4181
rect 6134 4178 6194 4254
rect 11237 4251 11303 4254
rect 11881 4314 11947 4317
rect 14273 4314 14339 4317
rect 11881 4312 14339 4314
rect 11881 4256 11886 4312
rect 11942 4256 14278 4312
rect 14334 4256 14339 4312
rect 11881 4254 14339 4256
rect 15334 4314 15394 4526
rect 18505 4584 25839 4586
rect 18505 4528 18510 4584
rect 18566 4528 25778 4584
rect 25834 4528 25839 4584
rect 18505 4526 25839 4528
rect 18505 4523 18571 4526
rect 25773 4523 25839 4526
rect 17033 4450 17099 4453
rect 20805 4450 20871 4453
rect 17033 4448 20871 4450
rect 17033 4392 17038 4448
rect 17094 4392 20810 4448
rect 20866 4392 20871 4448
rect 17033 4390 20871 4392
rect 26006 4450 26066 4662
rect 27520 4450 28000 4480
rect 26006 4390 28000 4450
rect 17033 4387 17099 4390
rect 20805 4387 20871 4390
rect 24277 4384 24597 4385
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 27520 4360 28000 4390
rect 24277 4319 24597 4320
rect 20529 4314 20595 4317
rect 15334 4312 20595 4314
rect 15334 4256 20534 4312
rect 20590 4256 20595 4312
rect 15334 4254 20595 4256
rect 11881 4251 11947 4254
rect 14273 4251 14339 4254
rect 20529 4251 20595 4254
rect 20662 4252 20668 4316
rect 20732 4314 20738 4316
rect 21265 4314 21331 4317
rect 22553 4314 22619 4317
rect 20732 4312 22619 4314
rect 20732 4256 21270 4312
rect 21326 4256 22558 4312
rect 22614 4256 22619 4312
rect 20732 4254 22619 4256
rect 20732 4252 20738 4254
rect 21265 4251 21331 4254
rect 22553 4251 22619 4254
rect 4061 4176 6194 4178
rect 4061 4120 4066 4176
rect 4122 4120 6194 4176
rect 4061 4118 6194 4120
rect 6361 4178 6427 4181
rect 8569 4178 8635 4181
rect 11053 4178 11119 4181
rect 6361 4176 8635 4178
rect 6361 4120 6366 4176
rect 6422 4120 8574 4176
rect 8630 4120 8635 4176
rect 6361 4118 8635 4120
rect 4061 4115 4127 4118
rect 6361 4115 6427 4118
rect 8569 4115 8635 4118
rect 8710 4176 11119 4178
rect 8710 4120 11058 4176
rect 11114 4120 11119 4176
rect 8710 4118 11119 4120
rect 1577 4042 1643 4045
rect 8710 4042 8770 4118
rect 11053 4115 11119 4118
rect 11697 4178 11763 4181
rect 14089 4178 14155 4181
rect 11697 4176 14155 4178
rect 11697 4120 11702 4176
rect 11758 4120 14094 4176
rect 14150 4120 14155 4176
rect 11697 4118 14155 4120
rect 11697 4115 11763 4118
rect 14089 4115 14155 4118
rect 20069 4178 20135 4181
rect 26233 4178 26299 4181
rect 20069 4176 26299 4178
rect 20069 4120 20074 4176
rect 20130 4120 26238 4176
rect 26294 4120 26299 4176
rect 20069 4118 26299 4120
rect 20069 4115 20135 4118
rect 26233 4115 26299 4118
rect 1577 4040 8770 4042
rect 1577 3984 1582 4040
rect 1638 3984 8770 4040
rect 1577 3982 8770 3984
rect 9673 4042 9739 4045
rect 12341 4042 12407 4045
rect 9673 4040 12407 4042
rect 9673 3984 9678 4040
rect 9734 3984 12346 4040
rect 12402 3984 12407 4040
rect 9673 3982 12407 3984
rect 1577 3979 1643 3982
rect 9673 3979 9739 3982
rect 12341 3979 12407 3982
rect 12617 4042 12683 4045
rect 13445 4042 13511 4045
rect 12617 4040 13511 4042
rect 12617 3984 12622 4040
rect 12678 3984 13450 4040
rect 13506 3984 13511 4040
rect 12617 3982 13511 3984
rect 12617 3979 12683 3982
rect 13445 3979 13511 3982
rect 15745 4042 15811 4045
rect 17493 4042 17559 4045
rect 15745 4040 17559 4042
rect 15745 3984 15750 4040
rect 15806 3984 17498 4040
rect 17554 3984 17559 4040
rect 15745 3982 17559 3984
rect 15745 3979 15811 3982
rect 17493 3979 17559 3982
rect 21909 4042 21975 4045
rect 24301 4042 24367 4045
rect 21909 4040 24367 4042
rect 21909 3984 21914 4040
rect 21970 3984 24306 4040
rect 24362 3984 24367 4040
rect 21909 3982 24367 3984
rect 21909 3979 21975 3982
rect 24301 3979 24367 3982
rect 24485 4042 24551 4045
rect 24710 4042 24716 4044
rect 24485 4040 24716 4042
rect 24485 3984 24490 4040
rect 24546 3984 24716 4040
rect 24485 3982 24716 3984
rect 24485 3979 24551 3982
rect 24710 3980 24716 3982
rect 24780 3980 24786 4044
rect 25313 4042 25379 4045
rect 27061 4042 27127 4045
rect 25313 4040 27127 4042
rect 25313 3984 25318 4040
rect 25374 3984 27066 4040
rect 27122 3984 27127 4040
rect 25313 3982 27127 3984
rect 25313 3979 25379 3982
rect 27061 3979 27127 3982
rect 10685 3906 10751 3909
rect 12801 3906 12867 3909
rect 10685 3904 12867 3906
rect 10685 3848 10690 3904
rect 10746 3848 12806 3904
rect 12862 3848 12867 3904
rect 10685 3846 12867 3848
rect 10685 3843 10751 3846
rect 12801 3843 12867 3846
rect 13169 3906 13235 3909
rect 15653 3906 15719 3909
rect 13169 3904 15719 3906
rect 13169 3848 13174 3904
rect 13230 3848 15658 3904
rect 15714 3848 15719 3904
rect 13169 3846 15719 3848
rect 13169 3843 13235 3846
rect 15653 3843 15719 3846
rect 16430 3844 16436 3908
rect 16500 3906 16506 3908
rect 16941 3906 17007 3909
rect 16500 3904 17007 3906
rect 16500 3848 16946 3904
rect 17002 3848 17007 3904
rect 16500 3846 17007 3848
rect 16500 3844 16506 3846
rect 16941 3843 17007 3846
rect 20897 3906 20963 3909
rect 25037 3906 25103 3909
rect 20897 3904 25103 3906
rect 20897 3848 20902 3904
rect 20958 3848 25042 3904
rect 25098 3848 25103 3904
rect 20897 3846 25103 3848
rect 20897 3843 20963 3846
rect 25037 3843 25103 3846
rect 10277 3840 10597 3841
rect 0 3770 480 3800
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 10277 3775 10597 3776
rect 19610 3840 19930 3841
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 3775 19930 3776
rect 1485 3770 1551 3773
rect 0 3768 1551 3770
rect 0 3712 1490 3768
rect 1546 3712 1551 3768
rect 0 3710 1551 3712
rect 0 3680 480 3710
rect 1485 3707 1551 3710
rect 1761 3770 1827 3773
rect 8937 3770 9003 3773
rect 10961 3770 11027 3773
rect 13077 3770 13143 3773
rect 18045 3770 18111 3773
rect 19425 3770 19491 3773
rect 20989 3772 21055 3773
rect 20989 3770 21036 3772
rect 1761 3768 9138 3770
rect 1761 3712 1766 3768
rect 1822 3712 8942 3768
rect 8998 3712 9138 3768
rect 1761 3710 9138 3712
rect 1761 3707 1827 3710
rect 8937 3707 9003 3710
rect 4521 3634 4587 3637
rect 4654 3634 4660 3636
rect 4521 3632 4660 3634
rect 4521 3576 4526 3632
rect 4582 3576 4660 3632
rect 4521 3574 4660 3576
rect 4521 3571 4587 3574
rect 4654 3572 4660 3574
rect 4724 3572 4730 3636
rect 9078 3634 9138 3710
rect 10961 3768 11898 3770
rect 10961 3712 10966 3768
rect 11022 3712 11898 3768
rect 10961 3710 11898 3712
rect 10961 3707 11027 3710
rect 11513 3634 11579 3637
rect 11838 3636 11898 3710
rect 13077 3768 18111 3770
rect 13077 3712 13082 3768
rect 13138 3712 18050 3768
rect 18106 3712 18111 3768
rect 13077 3710 18111 3712
rect 13077 3707 13143 3710
rect 18045 3707 18111 3710
rect 19014 3768 19491 3770
rect 19014 3712 19430 3768
rect 19486 3712 19491 3768
rect 19014 3710 19491 3712
rect 20944 3768 21036 3770
rect 20944 3712 20994 3768
rect 20944 3710 21036 3712
rect 4846 3574 7666 3634
rect 9078 3632 11579 3634
rect 9078 3576 11518 3632
rect 11574 3576 11579 3632
rect 9078 3574 11579 3576
rect 657 3498 723 3501
rect 4846 3498 4906 3574
rect 657 3496 4906 3498
rect 657 3440 662 3496
rect 718 3440 4906 3496
rect 657 3438 4906 3440
rect 4981 3498 5047 3501
rect 6678 3498 6684 3500
rect 4981 3496 6684 3498
rect 4981 3440 4986 3496
rect 5042 3440 6684 3496
rect 4981 3438 6684 3440
rect 657 3435 723 3438
rect 4981 3435 5047 3438
rect 6678 3436 6684 3438
rect 6748 3436 6754 3500
rect 6310 3300 6316 3364
rect 6380 3362 6386 3364
rect 6729 3362 6795 3365
rect 6380 3360 6795 3362
rect 6380 3304 6734 3360
rect 6790 3304 6795 3360
rect 6380 3302 6795 3304
rect 7606 3362 7666 3574
rect 11513 3571 11579 3574
rect 11830 3572 11836 3636
rect 11900 3634 11906 3636
rect 14733 3634 14799 3637
rect 11900 3632 14799 3634
rect 11900 3576 14738 3632
rect 14794 3576 14799 3632
rect 11900 3574 14799 3576
rect 11900 3572 11906 3574
rect 14733 3571 14799 3574
rect 15009 3634 15075 3637
rect 19014 3634 19074 3710
rect 19425 3707 19491 3710
rect 20989 3708 21036 3710
rect 21100 3708 21106 3772
rect 21173 3770 21239 3773
rect 23933 3770 23999 3773
rect 21173 3768 23999 3770
rect 21173 3712 21178 3768
rect 21234 3712 23938 3768
rect 23994 3712 23999 3768
rect 21173 3710 23999 3712
rect 20989 3707 21055 3708
rect 21173 3707 21239 3710
rect 23933 3707 23999 3710
rect 24761 3770 24827 3773
rect 27520 3770 28000 3800
rect 24761 3768 28000 3770
rect 24761 3712 24766 3768
rect 24822 3712 28000 3768
rect 24761 3710 28000 3712
rect 24761 3707 24827 3710
rect 27520 3680 28000 3710
rect 15009 3632 19074 3634
rect 15009 3576 15014 3632
rect 15070 3576 19074 3632
rect 15009 3574 19074 3576
rect 19241 3634 19307 3637
rect 26233 3634 26299 3637
rect 19241 3632 26299 3634
rect 19241 3576 19246 3632
rect 19302 3576 26238 3632
rect 26294 3576 26299 3632
rect 19241 3574 26299 3576
rect 15009 3571 15075 3574
rect 19241 3571 19307 3574
rect 26233 3571 26299 3574
rect 7833 3498 7899 3501
rect 9765 3498 9831 3501
rect 23473 3498 23539 3501
rect 7833 3496 23539 3498
rect 7833 3440 7838 3496
rect 7894 3440 9770 3496
rect 9826 3440 23478 3496
rect 23534 3440 23539 3496
rect 7833 3438 23539 3440
rect 7833 3435 7899 3438
rect 9765 3435 9831 3438
rect 23473 3435 23539 3438
rect 25405 3498 25471 3501
rect 27613 3498 27679 3501
rect 25405 3496 27679 3498
rect 25405 3440 25410 3496
rect 25466 3440 27618 3496
rect 27674 3440 27679 3496
rect 25405 3438 27679 3440
rect 25405 3435 25471 3438
rect 27613 3435 27679 3438
rect 9949 3362 10015 3365
rect 7606 3360 10015 3362
rect 7606 3304 9954 3360
rect 10010 3304 10015 3360
rect 7606 3302 10015 3304
rect 6380 3300 6386 3302
rect 6729 3299 6795 3302
rect 9949 3299 10015 3302
rect 10685 3362 10751 3365
rect 12433 3362 12499 3365
rect 10685 3360 12499 3362
rect 10685 3304 10690 3360
rect 10746 3304 12438 3360
rect 12494 3304 12499 3360
rect 10685 3302 12499 3304
rect 10685 3299 10751 3302
rect 12433 3299 12499 3302
rect 12801 3362 12867 3365
rect 14641 3362 14707 3365
rect 12801 3360 14707 3362
rect 12801 3304 12806 3360
rect 12862 3304 14646 3360
rect 14702 3304 14707 3360
rect 12801 3302 14707 3304
rect 12801 3299 12867 3302
rect 14641 3299 14707 3302
rect 18413 3362 18479 3365
rect 23473 3362 23539 3365
rect 23657 3364 23723 3365
rect 18413 3360 23539 3362
rect 18413 3304 18418 3360
rect 18474 3304 23478 3360
rect 23534 3304 23539 3360
rect 18413 3302 23539 3304
rect 18413 3299 18479 3302
rect 23473 3299 23539 3302
rect 23606 3300 23612 3364
rect 23676 3362 23723 3364
rect 24669 3362 24735 3365
rect 26509 3362 26575 3365
rect 23676 3360 23768 3362
rect 23718 3304 23768 3360
rect 23676 3302 23768 3304
rect 24669 3360 26575 3362
rect 24669 3304 24674 3360
rect 24730 3304 26514 3360
rect 26570 3304 26575 3360
rect 24669 3302 26575 3304
rect 23676 3300 23723 3302
rect 23657 3299 23723 3300
rect 24669 3299 24735 3302
rect 26509 3299 26575 3302
rect 5610 3296 5930 3297
rect 0 3226 480 3256
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5930 3296
rect 5610 3231 5930 3232
rect 14944 3296 15264 3297
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 14944 3231 15264 3232
rect 24277 3296 24597 3297
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 3231 24597 3232
rect 2405 3226 2471 3229
rect 0 3224 2471 3226
rect 0 3168 2410 3224
rect 2466 3168 2471 3224
rect 0 3166 2471 3168
rect 0 3136 480 3166
rect 2405 3163 2471 3166
rect 2865 3226 2931 3229
rect 5165 3226 5231 3229
rect 2865 3224 5231 3226
rect 2865 3168 2870 3224
rect 2926 3168 5170 3224
rect 5226 3168 5231 3224
rect 2865 3166 5231 3168
rect 2865 3163 2931 3166
rect 5165 3163 5231 3166
rect 8385 3226 8451 3229
rect 11697 3226 11763 3229
rect 8385 3224 11763 3226
rect 8385 3168 8390 3224
rect 8446 3168 11702 3224
rect 11758 3168 11763 3224
rect 8385 3166 11763 3168
rect 8385 3163 8451 3166
rect 11697 3163 11763 3166
rect 15469 3226 15535 3229
rect 21541 3226 21607 3229
rect 22001 3226 22067 3229
rect 23473 3228 23539 3229
rect 15469 3224 22067 3226
rect 15469 3168 15474 3224
rect 15530 3168 21546 3224
rect 21602 3168 22006 3224
rect 22062 3168 22067 3224
rect 15469 3166 22067 3168
rect 15469 3163 15535 3166
rect 21541 3163 21607 3166
rect 22001 3163 22067 3166
rect 23422 3164 23428 3228
rect 23492 3226 23539 3228
rect 26325 3226 26391 3229
rect 27520 3226 28000 3256
rect 23492 3224 23584 3226
rect 23534 3168 23584 3224
rect 23492 3166 23584 3168
rect 26325 3224 28000 3226
rect 26325 3168 26330 3224
rect 26386 3168 28000 3224
rect 26325 3166 28000 3168
rect 23492 3164 23539 3166
rect 23473 3163 23539 3164
rect 26325 3163 26391 3166
rect 27520 3136 28000 3166
rect 1393 3090 1459 3093
rect 11237 3090 11303 3093
rect 1393 3088 11303 3090
rect 1393 3032 1398 3088
rect 1454 3032 11242 3088
rect 11298 3032 11303 3088
rect 1393 3030 11303 3032
rect 1393 3027 1459 3030
rect 11237 3027 11303 3030
rect 13629 3090 13695 3093
rect 18505 3090 18571 3093
rect 25037 3090 25103 3093
rect 13629 3088 25103 3090
rect 13629 3032 13634 3088
rect 13690 3032 18510 3088
rect 18566 3032 25042 3088
rect 25098 3032 25103 3088
rect 13629 3030 25103 3032
rect 13629 3027 13695 3030
rect 18505 3027 18571 3030
rect 25037 3027 25103 3030
rect 1945 2954 2011 2957
rect 8385 2954 8451 2957
rect 1945 2952 8451 2954
rect 1945 2896 1950 2952
rect 2006 2896 8390 2952
rect 8446 2896 8451 2952
rect 1945 2894 8451 2896
rect 1945 2891 2011 2894
rect 8385 2891 8451 2894
rect 8661 2954 8727 2957
rect 11329 2954 11395 2957
rect 13813 2954 13879 2957
rect 8661 2952 10794 2954
rect 8661 2896 8666 2952
rect 8722 2896 10794 2952
rect 8661 2894 10794 2896
rect 8661 2891 8727 2894
rect 1209 2818 1275 2821
rect 4061 2818 4127 2821
rect 10734 2818 10794 2894
rect 11329 2952 13879 2954
rect 11329 2896 11334 2952
rect 11390 2896 13818 2952
rect 13874 2896 13879 2952
rect 11329 2894 13879 2896
rect 11329 2891 11395 2894
rect 13813 2891 13879 2894
rect 13997 2954 14063 2957
rect 18045 2954 18111 2957
rect 13997 2952 18111 2954
rect 13997 2896 14002 2952
rect 14058 2896 18050 2952
rect 18106 2896 18111 2952
rect 13997 2894 18111 2896
rect 13997 2891 14063 2894
rect 18045 2891 18111 2894
rect 22093 2954 22159 2957
rect 25129 2954 25195 2957
rect 22093 2952 25195 2954
rect 22093 2896 22098 2952
rect 22154 2896 25134 2952
rect 25190 2896 25195 2952
rect 22093 2894 25195 2896
rect 22093 2891 22159 2894
rect 25129 2891 25195 2894
rect 11237 2818 11303 2821
rect 1209 2816 4722 2818
rect 1209 2760 1214 2816
rect 1270 2760 4066 2816
rect 4122 2760 4722 2816
rect 1209 2758 4722 2760
rect 10734 2816 11303 2818
rect 10734 2760 11242 2816
rect 11298 2760 11303 2816
rect 10734 2758 11303 2760
rect 1209 2755 1275 2758
rect 4061 2755 4127 2758
rect 0 2682 480 2712
rect 0 2622 3802 2682
rect 0 2592 480 2622
rect 3742 2410 3802 2622
rect 4662 2546 4722 2758
rect 11237 2755 11303 2758
rect 13445 2818 13511 2821
rect 14641 2818 14707 2821
rect 15193 2818 15259 2821
rect 13445 2816 15259 2818
rect 13445 2760 13450 2816
rect 13506 2760 14646 2816
rect 14702 2760 15198 2816
rect 15254 2760 15259 2816
rect 13445 2758 15259 2760
rect 13445 2755 13511 2758
rect 14641 2755 14707 2758
rect 15193 2755 15259 2758
rect 15653 2818 15719 2821
rect 18781 2818 18847 2821
rect 19425 2818 19491 2821
rect 15653 2816 19491 2818
rect 15653 2760 15658 2816
rect 15714 2760 18786 2816
rect 18842 2760 19430 2816
rect 19486 2760 19491 2816
rect 15653 2758 19491 2760
rect 15653 2755 15719 2758
rect 18781 2755 18847 2758
rect 19425 2755 19491 2758
rect 21081 2818 21147 2821
rect 25129 2818 25195 2821
rect 21081 2816 25195 2818
rect 21081 2760 21086 2816
rect 21142 2760 25134 2816
rect 25190 2760 25195 2816
rect 21081 2758 25195 2760
rect 21081 2755 21147 2758
rect 25129 2755 25195 2758
rect 10277 2752 10597 2753
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2687 10597 2688
rect 19610 2752 19930 2753
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 19610 2687 19930 2688
rect 4797 2682 4863 2685
rect 10133 2682 10199 2685
rect 4797 2680 10199 2682
rect 4797 2624 4802 2680
rect 4858 2624 10138 2680
rect 10194 2624 10199 2680
rect 4797 2622 10199 2624
rect 4797 2619 4863 2622
rect 10133 2619 10199 2622
rect 12382 2620 12388 2684
rect 12452 2682 12458 2684
rect 13169 2682 13235 2685
rect 16849 2682 16915 2685
rect 12452 2622 13002 2682
rect 12452 2620 12458 2622
rect 12709 2546 12775 2549
rect 4662 2544 12775 2546
rect 4662 2488 12714 2544
rect 12770 2488 12775 2544
rect 4662 2486 12775 2488
rect 12942 2546 13002 2622
rect 13169 2680 16915 2682
rect 13169 2624 13174 2680
rect 13230 2624 16854 2680
rect 16910 2624 16915 2680
rect 13169 2622 16915 2624
rect 13169 2619 13235 2622
rect 16849 2619 16915 2622
rect 22921 2682 22987 2685
rect 24945 2682 25011 2685
rect 27520 2682 28000 2712
rect 22921 2680 25011 2682
rect 22921 2624 22926 2680
rect 22982 2624 24950 2680
rect 25006 2624 25011 2680
rect 22921 2622 25011 2624
rect 22921 2619 22987 2622
rect 24945 2619 25011 2622
rect 25086 2622 28000 2682
rect 14457 2546 14523 2549
rect 16665 2546 16731 2549
rect 12942 2544 14523 2546
rect 12942 2488 14462 2544
rect 14518 2488 14523 2544
rect 12942 2486 14523 2488
rect 12709 2483 12775 2486
rect 14457 2483 14523 2486
rect 14598 2544 16731 2546
rect 14598 2488 16670 2544
rect 16726 2488 16731 2544
rect 14598 2486 16731 2488
rect 12065 2410 12131 2413
rect 3742 2408 12131 2410
rect 3742 2352 12070 2408
rect 12126 2352 12131 2408
rect 3742 2350 12131 2352
rect 12065 2347 12131 2350
rect 12249 2410 12315 2413
rect 14598 2410 14658 2486
rect 16665 2483 16731 2486
rect 16798 2484 16804 2548
rect 16868 2546 16874 2548
rect 20805 2546 20871 2549
rect 16868 2544 20871 2546
rect 16868 2488 20810 2544
rect 20866 2488 20871 2544
rect 16868 2486 20871 2488
rect 16868 2484 16874 2486
rect 20805 2483 20871 2486
rect 21173 2546 21239 2549
rect 22737 2546 22803 2549
rect 25086 2546 25146 2622
rect 27520 2592 28000 2622
rect 21173 2544 22570 2546
rect 21173 2488 21178 2544
rect 21234 2488 22570 2544
rect 21173 2486 22570 2488
rect 21173 2483 21239 2486
rect 19793 2410 19859 2413
rect 12249 2408 14658 2410
rect 12249 2352 12254 2408
rect 12310 2352 14658 2408
rect 12249 2350 14658 2352
rect 14782 2408 19859 2410
rect 14782 2352 19798 2408
rect 19854 2352 19859 2408
rect 14782 2350 19859 2352
rect 12249 2347 12315 2350
rect 6269 2274 6335 2277
rect 9305 2274 9371 2277
rect 14782 2274 14842 2350
rect 19793 2347 19859 2350
rect 20161 2410 20227 2413
rect 22369 2410 22435 2413
rect 20161 2408 22435 2410
rect 20161 2352 20166 2408
rect 20222 2352 22374 2408
rect 22430 2352 22435 2408
rect 20161 2350 22435 2352
rect 22510 2410 22570 2486
rect 22737 2544 25146 2546
rect 22737 2488 22742 2544
rect 22798 2488 25146 2544
rect 22737 2486 25146 2488
rect 22737 2483 22803 2486
rect 22829 2410 22895 2413
rect 26233 2410 26299 2413
rect 22510 2408 26299 2410
rect 22510 2352 22834 2408
rect 22890 2352 26238 2408
rect 26294 2352 26299 2408
rect 22510 2350 26299 2352
rect 20161 2347 20227 2350
rect 22369 2347 22435 2350
rect 22829 2347 22895 2350
rect 26233 2347 26299 2350
rect 6269 2272 14842 2274
rect 6269 2216 6274 2272
rect 6330 2216 9310 2272
rect 9366 2216 14842 2272
rect 6269 2214 14842 2216
rect 16665 2274 16731 2277
rect 20897 2274 20963 2277
rect 16665 2272 20963 2274
rect 16665 2216 16670 2272
rect 16726 2216 20902 2272
rect 20958 2216 20963 2272
rect 16665 2214 20963 2216
rect 6269 2211 6335 2214
rect 9305 2211 9371 2214
rect 16665 2211 16731 2214
rect 20897 2211 20963 2214
rect 22553 2274 22619 2277
rect 23841 2274 23907 2277
rect 22553 2272 23907 2274
rect 22553 2216 22558 2272
rect 22614 2216 23846 2272
rect 23902 2216 23907 2272
rect 22553 2214 23907 2216
rect 22553 2211 22619 2214
rect 23841 2211 23907 2214
rect 5610 2208 5930 2209
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5930 2208
rect 5610 2143 5930 2144
rect 14944 2208 15264 2209
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2143 15264 2144
rect 24277 2208 24597 2209
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2143 24597 2144
rect 1577 2138 1643 2141
rect 13537 2138 13603 2141
rect 1577 2136 5458 2138
rect 1577 2080 1582 2136
rect 1638 2080 5458 2136
rect 1577 2078 5458 2080
rect 1577 2075 1643 2078
rect 0 2002 480 2032
rect 5398 2002 5458 2078
rect 6870 2136 13603 2138
rect 6870 2080 13542 2136
rect 13598 2080 13603 2136
rect 6870 2078 13603 2080
rect 6870 2002 6930 2078
rect 13537 2075 13603 2078
rect 15377 2138 15443 2141
rect 18505 2138 18571 2141
rect 15377 2136 18571 2138
rect 15377 2080 15382 2136
rect 15438 2080 18510 2136
rect 18566 2080 18571 2136
rect 15377 2078 18571 2080
rect 15377 2075 15443 2078
rect 18505 2075 18571 2078
rect 18689 2138 18755 2141
rect 20989 2138 21055 2141
rect 18689 2136 21055 2138
rect 18689 2080 18694 2136
rect 18750 2080 20994 2136
rect 21050 2080 21055 2136
rect 18689 2078 21055 2080
rect 18689 2075 18755 2078
rect 20989 2075 21055 2078
rect 0 1942 5274 2002
rect 5398 1942 6930 2002
rect 10869 2002 10935 2005
rect 12617 2002 12683 2005
rect 27520 2002 28000 2032
rect 10869 2000 12266 2002
rect 10869 1944 10874 2000
rect 10930 1944 12266 2000
rect 10869 1942 12266 1944
rect 0 1912 480 1942
rect 5214 1866 5274 1942
rect 10869 1939 10935 1942
rect 12065 1866 12131 1869
rect 5214 1864 12131 1866
rect 5214 1808 12070 1864
rect 12126 1808 12131 1864
rect 5214 1806 12131 1808
rect 12206 1866 12266 1942
rect 12617 2000 28000 2002
rect 12617 1944 12622 2000
rect 12678 1944 28000 2000
rect 12617 1942 28000 1944
rect 12617 1939 12683 1942
rect 27520 1912 28000 1942
rect 12382 1866 12388 1868
rect 12206 1806 12388 1866
rect 12065 1803 12131 1806
rect 12382 1804 12388 1806
rect 12452 1804 12458 1868
rect 12525 1866 12591 1869
rect 15510 1866 15516 1868
rect 12525 1864 15516 1866
rect 12525 1808 12530 1864
rect 12586 1808 15516 1864
rect 12525 1806 15516 1808
rect 12525 1803 12591 1806
rect 15510 1804 15516 1806
rect 15580 1866 15586 1868
rect 20713 1866 20779 1869
rect 15580 1864 20779 1866
rect 15580 1808 20718 1864
rect 20774 1808 20779 1864
rect 15580 1806 20779 1808
rect 15580 1804 15586 1806
rect 20713 1803 20779 1806
rect 22369 1866 22435 1869
rect 26417 1866 26483 1869
rect 22369 1864 26483 1866
rect 22369 1808 22374 1864
rect 22430 1808 26422 1864
rect 26478 1808 26483 1864
rect 22369 1806 26483 1808
rect 22369 1803 22435 1806
rect 26417 1803 26483 1806
rect 197 1730 263 1733
rect 1945 1730 2011 1733
rect 2078 1730 2084 1732
rect 197 1728 674 1730
rect 197 1672 202 1728
rect 258 1672 674 1728
rect 197 1670 674 1672
rect 197 1667 263 1670
rect 614 1594 674 1670
rect 1945 1728 2084 1730
rect 1945 1672 1950 1728
rect 2006 1672 2084 1728
rect 1945 1670 2084 1672
rect 1945 1667 2011 1670
rect 2078 1668 2084 1670
rect 2148 1668 2154 1732
rect 13997 1730 14063 1733
rect 2270 1728 14063 1730
rect 2270 1672 14002 1728
rect 14058 1672 14063 1728
rect 2270 1670 14063 1672
rect 2270 1594 2330 1670
rect 13997 1667 14063 1670
rect 17401 1730 17467 1733
rect 18597 1730 18663 1733
rect 25681 1730 25747 1733
rect 17401 1728 18522 1730
rect 17401 1672 17406 1728
rect 17462 1672 18522 1728
rect 17401 1670 18522 1672
rect 17401 1667 17467 1670
rect 614 1534 2330 1594
rect 3141 1594 3207 1597
rect 6545 1594 6611 1597
rect 3141 1592 6611 1594
rect 3141 1536 3146 1592
rect 3202 1536 6550 1592
rect 6606 1536 6611 1592
rect 3141 1534 6611 1536
rect 3141 1531 3207 1534
rect 6545 1531 6611 1534
rect 6913 1594 6979 1597
rect 9029 1594 9095 1597
rect 6913 1592 9095 1594
rect 6913 1536 6918 1592
rect 6974 1536 9034 1592
rect 9090 1536 9095 1592
rect 6913 1534 9095 1536
rect 6913 1531 6979 1534
rect 9029 1531 9095 1534
rect 9213 1594 9279 1597
rect 18321 1594 18387 1597
rect 9213 1592 18387 1594
rect 9213 1536 9218 1592
rect 9274 1536 18326 1592
rect 18382 1536 18387 1592
rect 9213 1534 18387 1536
rect 18462 1594 18522 1670
rect 18597 1728 25747 1730
rect 18597 1672 18602 1728
rect 18658 1672 25686 1728
rect 25742 1672 25747 1728
rect 18597 1670 25747 1672
rect 18597 1667 18663 1670
rect 25681 1667 25747 1670
rect 25221 1594 25287 1597
rect 18462 1592 25287 1594
rect 18462 1536 25226 1592
rect 25282 1536 25287 1592
rect 18462 1534 25287 1536
rect 9213 1531 9279 1534
rect 18321 1531 18387 1534
rect 25221 1531 25287 1534
rect 0 1458 480 1488
rect 9397 1458 9463 1461
rect 0 1456 9463 1458
rect 0 1400 9402 1456
rect 9458 1400 9463 1456
rect 0 1398 9463 1400
rect 0 1368 480 1398
rect 9397 1395 9463 1398
rect 12433 1458 12499 1461
rect 18229 1458 18295 1461
rect 12433 1456 18295 1458
rect 12433 1400 12438 1456
rect 12494 1400 18234 1456
rect 18290 1400 18295 1456
rect 12433 1398 18295 1400
rect 12433 1395 12499 1398
rect 18229 1395 18295 1398
rect 18781 1458 18847 1461
rect 22921 1458 22987 1461
rect 18781 1456 22987 1458
rect 18781 1400 18786 1456
rect 18842 1400 22926 1456
rect 22982 1400 22987 1456
rect 18781 1398 22987 1400
rect 18781 1395 18847 1398
rect 22921 1395 22987 1398
rect 24669 1458 24735 1461
rect 27520 1458 28000 1488
rect 24669 1456 28000 1458
rect 24669 1400 24674 1456
rect 24730 1400 28000 1456
rect 24669 1398 28000 1400
rect 24669 1395 24735 1398
rect 27520 1368 28000 1398
rect 9581 1322 9647 1325
rect 24761 1322 24827 1325
rect 9581 1320 24827 1322
rect 9581 1264 9586 1320
rect 9642 1264 24766 1320
rect 24822 1264 24827 1320
rect 9581 1262 24827 1264
rect 9581 1259 9647 1262
rect 24761 1259 24827 1262
rect 11237 1186 11303 1189
rect 22553 1186 22619 1189
rect 11237 1184 22619 1186
rect 11237 1128 11242 1184
rect 11298 1128 22558 1184
rect 22614 1128 22619 1184
rect 11237 1126 22619 1128
rect 11237 1123 11303 1126
rect 22553 1123 22619 1126
rect 11881 1050 11947 1053
rect 24117 1050 24183 1053
rect 11881 1048 24183 1050
rect 11881 992 11886 1048
rect 11942 992 24122 1048
rect 24178 992 24183 1048
rect 11881 990 24183 992
rect 11881 987 11947 990
rect 24117 987 24183 990
rect 0 914 480 944
rect 3693 914 3759 917
rect 16205 914 16271 917
rect 0 854 3618 914
rect 0 824 480 854
rect 3558 778 3618 854
rect 3693 912 16271 914
rect 3693 856 3698 912
rect 3754 856 16210 912
rect 16266 856 16271 912
rect 3693 854 16271 856
rect 3693 851 3759 854
rect 16205 851 16271 854
rect 17217 914 17283 917
rect 27520 914 28000 944
rect 17217 912 28000 914
rect 17217 856 17222 912
rect 17278 856 28000 912
rect 17217 854 28000 856
rect 17217 851 17283 854
rect 27520 824 28000 854
rect 17033 778 17099 781
rect 25589 778 25655 781
rect 3558 776 17099 778
rect 3558 720 17038 776
rect 17094 720 17099 776
rect 3558 718 17099 720
rect 17033 715 17099 718
rect 17174 776 25655 778
rect 17174 720 25594 776
rect 25650 720 25655 776
rect 17174 718 25655 720
rect 2221 642 2287 645
rect 17174 642 17234 718
rect 25589 715 25655 718
rect 2221 640 17234 642
rect 2221 584 2226 640
rect 2282 584 17234 640
rect 2221 582 17234 584
rect 2221 579 2287 582
rect 3601 506 3667 509
rect 8017 506 8083 509
rect 26141 506 26207 509
rect 3601 504 7114 506
rect 3601 448 3606 504
rect 3662 448 7114 504
rect 3601 446 7114 448
rect 3601 443 3667 446
rect 0 370 480 400
rect 6913 370 6979 373
rect 0 368 6979 370
rect 0 312 6918 368
rect 6974 312 6979 368
rect 0 310 6979 312
rect 7054 370 7114 446
rect 8017 504 26207 506
rect 8017 448 8022 504
rect 8078 448 26146 504
rect 26202 448 26207 504
rect 8017 446 26207 448
rect 8017 443 8083 446
rect 26141 443 26207 446
rect 16205 370 16271 373
rect 19977 370 20043 373
rect 27520 370 28000 400
rect 7054 310 16130 370
rect 0 280 480 310
rect 6913 307 6979 310
rect 16070 234 16130 310
rect 16205 368 20043 370
rect 16205 312 16210 368
rect 16266 312 19982 368
rect 20038 312 20043 368
rect 16205 310 20043 312
rect 16205 307 16271 310
rect 19977 307 20043 310
rect 27478 280 28000 370
rect 18413 234 18479 237
rect 27478 234 27538 280
rect 16070 174 17418 234
rect 9673 98 9739 101
rect 17217 98 17283 101
rect 9673 96 17283 98
rect 9673 40 9678 96
rect 9734 40 17222 96
rect 17278 40 17283 96
rect 9673 38 17283 40
rect 17358 98 17418 174
rect 18413 232 27538 234
rect 18413 176 18418 232
rect 18474 176 27538 232
rect 18413 174 27538 176
rect 18413 171 18479 174
rect 20805 98 20871 101
rect 17358 96 20871 98
rect 17358 40 20810 96
rect 20866 40 20871 96
rect 17358 38 20871 40
rect 9673 35 9739 38
rect 17217 35 17283 38
rect 20805 35 20871 38
<< via3 >>
rect 2820 26012 2884 26076
rect 10285 25596 10349 25600
rect 10285 25540 10289 25596
rect 10289 25540 10345 25596
rect 10345 25540 10349 25596
rect 10285 25536 10349 25540
rect 10365 25596 10429 25600
rect 10365 25540 10369 25596
rect 10369 25540 10425 25596
rect 10425 25540 10429 25596
rect 10365 25536 10429 25540
rect 10445 25596 10509 25600
rect 10445 25540 10449 25596
rect 10449 25540 10505 25596
rect 10505 25540 10509 25596
rect 10445 25536 10509 25540
rect 10525 25596 10589 25600
rect 10525 25540 10529 25596
rect 10529 25540 10585 25596
rect 10585 25540 10589 25596
rect 10525 25536 10589 25540
rect 25820 25604 25884 25668
rect 19618 25596 19682 25600
rect 19618 25540 19622 25596
rect 19622 25540 19678 25596
rect 19678 25540 19682 25596
rect 19618 25536 19682 25540
rect 19698 25596 19762 25600
rect 19698 25540 19702 25596
rect 19702 25540 19758 25596
rect 19758 25540 19762 25596
rect 19698 25536 19762 25540
rect 19778 25596 19842 25600
rect 19778 25540 19782 25596
rect 19782 25540 19838 25596
rect 19838 25540 19842 25596
rect 19778 25536 19842 25540
rect 19858 25596 19922 25600
rect 19858 25540 19862 25596
rect 19862 25540 19918 25596
rect 19918 25540 19922 25596
rect 19858 25536 19922 25540
rect 23980 25332 24044 25396
rect 10916 25196 10980 25260
rect 21220 25196 21284 25260
rect 5618 25052 5682 25056
rect 5618 24996 5622 25052
rect 5622 24996 5678 25052
rect 5678 24996 5682 25052
rect 5618 24992 5682 24996
rect 5698 25052 5762 25056
rect 5698 24996 5702 25052
rect 5702 24996 5758 25052
rect 5758 24996 5762 25052
rect 5698 24992 5762 24996
rect 5778 25052 5842 25056
rect 5778 24996 5782 25052
rect 5782 24996 5838 25052
rect 5838 24996 5842 25052
rect 5778 24992 5842 24996
rect 5858 25052 5922 25056
rect 5858 24996 5862 25052
rect 5862 24996 5918 25052
rect 5918 24996 5922 25052
rect 5858 24992 5922 24996
rect 14952 25052 15016 25056
rect 14952 24996 14956 25052
rect 14956 24996 15012 25052
rect 15012 24996 15016 25052
rect 14952 24992 15016 24996
rect 15032 25052 15096 25056
rect 15032 24996 15036 25052
rect 15036 24996 15092 25052
rect 15092 24996 15096 25052
rect 15032 24992 15096 24996
rect 15112 25052 15176 25056
rect 15112 24996 15116 25052
rect 15116 24996 15172 25052
rect 15172 24996 15176 25052
rect 15112 24992 15176 24996
rect 15192 25052 15256 25056
rect 15192 24996 15196 25052
rect 15196 24996 15252 25052
rect 15252 24996 15256 25052
rect 15192 24992 15256 24996
rect 3188 24848 3252 24852
rect 3188 24792 3202 24848
rect 3202 24792 3252 24848
rect 3188 24788 3252 24792
rect 3740 24848 3804 24852
rect 3740 24792 3790 24848
rect 3790 24792 3804 24848
rect 3740 24788 3804 24792
rect 14228 24848 14292 24852
rect 14228 24792 14278 24848
rect 14278 24792 14292 24848
rect 14228 24788 14292 24792
rect 24285 25052 24349 25056
rect 24285 24996 24289 25052
rect 24289 24996 24345 25052
rect 24345 24996 24349 25052
rect 24285 24992 24349 24996
rect 24365 25052 24429 25056
rect 24365 24996 24369 25052
rect 24369 24996 24425 25052
rect 24425 24996 24429 25052
rect 24365 24992 24429 24996
rect 24445 25052 24509 25056
rect 24445 24996 24449 25052
rect 24449 24996 24505 25052
rect 24505 24996 24509 25052
rect 24445 24992 24509 24996
rect 24525 25052 24589 25056
rect 24525 24996 24529 25052
rect 24529 24996 24585 25052
rect 24585 24996 24589 25052
rect 24525 24992 24589 24996
rect 23612 24924 23676 24988
rect 2636 24652 2700 24716
rect 10285 24508 10349 24512
rect 10285 24452 10289 24508
rect 10289 24452 10345 24508
rect 10345 24452 10349 24508
rect 10285 24448 10349 24452
rect 10365 24508 10429 24512
rect 10365 24452 10369 24508
rect 10369 24452 10425 24508
rect 10425 24452 10429 24508
rect 10365 24448 10429 24452
rect 10445 24508 10509 24512
rect 10445 24452 10449 24508
rect 10449 24452 10505 24508
rect 10505 24452 10509 24508
rect 10445 24448 10509 24452
rect 10525 24508 10589 24512
rect 10525 24452 10529 24508
rect 10529 24452 10585 24508
rect 10585 24452 10589 24508
rect 10525 24448 10589 24452
rect 19618 24508 19682 24512
rect 19618 24452 19622 24508
rect 19622 24452 19678 24508
rect 19678 24452 19682 24508
rect 19618 24448 19682 24452
rect 19698 24508 19762 24512
rect 19698 24452 19702 24508
rect 19702 24452 19758 24508
rect 19758 24452 19762 24508
rect 19698 24448 19762 24452
rect 19778 24508 19842 24512
rect 19778 24452 19782 24508
rect 19782 24452 19838 24508
rect 19838 24452 19842 24508
rect 19778 24448 19842 24452
rect 19858 24508 19922 24512
rect 19858 24452 19862 24508
rect 19862 24452 19918 24508
rect 19918 24452 19922 24508
rect 19858 24448 19922 24452
rect 20116 24380 20180 24444
rect 5618 23964 5682 23968
rect 5618 23908 5622 23964
rect 5622 23908 5678 23964
rect 5678 23908 5682 23964
rect 5618 23904 5682 23908
rect 5698 23964 5762 23968
rect 5698 23908 5702 23964
rect 5702 23908 5758 23964
rect 5758 23908 5762 23964
rect 5698 23904 5762 23908
rect 5778 23964 5842 23968
rect 5778 23908 5782 23964
rect 5782 23908 5838 23964
rect 5838 23908 5842 23964
rect 5778 23904 5842 23908
rect 5858 23964 5922 23968
rect 5858 23908 5862 23964
rect 5862 23908 5918 23964
rect 5918 23908 5922 23964
rect 5858 23904 5922 23908
rect 14952 23964 15016 23968
rect 14952 23908 14956 23964
rect 14956 23908 15012 23964
rect 15012 23908 15016 23964
rect 14952 23904 15016 23908
rect 15032 23964 15096 23968
rect 15032 23908 15036 23964
rect 15036 23908 15092 23964
rect 15092 23908 15096 23964
rect 15032 23904 15096 23908
rect 15112 23964 15176 23968
rect 15112 23908 15116 23964
rect 15116 23908 15172 23964
rect 15172 23908 15176 23964
rect 15112 23904 15176 23908
rect 15192 23964 15256 23968
rect 15192 23908 15196 23964
rect 15196 23908 15252 23964
rect 15252 23908 15256 23964
rect 15192 23904 15256 23908
rect 24285 23964 24349 23968
rect 24285 23908 24289 23964
rect 24289 23908 24345 23964
rect 24345 23908 24349 23964
rect 24285 23904 24349 23908
rect 24365 23964 24429 23968
rect 24365 23908 24369 23964
rect 24369 23908 24425 23964
rect 24425 23908 24429 23964
rect 24365 23904 24429 23908
rect 24445 23964 24509 23968
rect 24445 23908 24449 23964
rect 24449 23908 24505 23964
rect 24505 23908 24509 23964
rect 24445 23904 24509 23908
rect 24525 23964 24589 23968
rect 24525 23908 24529 23964
rect 24529 23908 24585 23964
rect 24585 23908 24589 23964
rect 24525 23904 24589 23908
rect 20668 23428 20732 23492
rect 24716 23428 24780 23492
rect 10285 23420 10349 23424
rect 10285 23364 10289 23420
rect 10289 23364 10345 23420
rect 10345 23364 10349 23420
rect 10285 23360 10349 23364
rect 10365 23420 10429 23424
rect 10365 23364 10369 23420
rect 10369 23364 10425 23420
rect 10425 23364 10429 23420
rect 10365 23360 10429 23364
rect 10445 23420 10509 23424
rect 10445 23364 10449 23420
rect 10449 23364 10505 23420
rect 10505 23364 10509 23420
rect 10445 23360 10509 23364
rect 10525 23420 10589 23424
rect 10525 23364 10529 23420
rect 10529 23364 10585 23420
rect 10585 23364 10589 23420
rect 10525 23360 10589 23364
rect 19618 23420 19682 23424
rect 19618 23364 19622 23420
rect 19622 23364 19678 23420
rect 19678 23364 19682 23420
rect 19618 23360 19682 23364
rect 19698 23420 19762 23424
rect 19698 23364 19702 23420
rect 19702 23364 19758 23420
rect 19758 23364 19762 23420
rect 19698 23360 19762 23364
rect 19778 23420 19842 23424
rect 19778 23364 19782 23420
rect 19782 23364 19838 23420
rect 19838 23364 19842 23420
rect 19778 23360 19842 23364
rect 19858 23420 19922 23424
rect 19858 23364 19862 23420
rect 19862 23364 19918 23420
rect 19918 23364 19922 23420
rect 19858 23360 19922 23364
rect 5618 22876 5682 22880
rect 5618 22820 5622 22876
rect 5622 22820 5678 22876
rect 5678 22820 5682 22876
rect 5618 22816 5682 22820
rect 5698 22876 5762 22880
rect 5698 22820 5702 22876
rect 5702 22820 5758 22876
rect 5758 22820 5762 22876
rect 5698 22816 5762 22820
rect 5778 22876 5842 22880
rect 5778 22820 5782 22876
rect 5782 22820 5838 22876
rect 5838 22820 5842 22876
rect 5778 22816 5842 22820
rect 5858 22876 5922 22880
rect 5858 22820 5862 22876
rect 5862 22820 5918 22876
rect 5918 22820 5922 22876
rect 5858 22816 5922 22820
rect 14952 22876 15016 22880
rect 14952 22820 14956 22876
rect 14956 22820 15012 22876
rect 15012 22820 15016 22876
rect 14952 22816 15016 22820
rect 15032 22876 15096 22880
rect 15032 22820 15036 22876
rect 15036 22820 15092 22876
rect 15092 22820 15096 22876
rect 15032 22816 15096 22820
rect 15112 22876 15176 22880
rect 15112 22820 15116 22876
rect 15116 22820 15172 22876
rect 15172 22820 15176 22876
rect 15112 22816 15176 22820
rect 15192 22876 15256 22880
rect 15192 22820 15196 22876
rect 15196 22820 15252 22876
rect 15252 22820 15256 22876
rect 15192 22816 15256 22820
rect 24285 22876 24349 22880
rect 24285 22820 24289 22876
rect 24289 22820 24345 22876
rect 24345 22820 24349 22876
rect 24285 22816 24349 22820
rect 24365 22876 24429 22880
rect 24365 22820 24369 22876
rect 24369 22820 24425 22876
rect 24425 22820 24429 22876
rect 24365 22816 24429 22820
rect 24445 22876 24509 22880
rect 24445 22820 24449 22876
rect 24449 22820 24505 22876
rect 24505 22820 24509 22876
rect 24445 22816 24509 22820
rect 24525 22876 24589 22880
rect 24525 22820 24529 22876
rect 24529 22820 24585 22876
rect 24585 22820 24589 22876
rect 24525 22816 24589 22820
rect 5028 22748 5092 22812
rect 15516 22748 15580 22812
rect 17724 22476 17788 22540
rect 10285 22332 10349 22336
rect 10285 22276 10289 22332
rect 10289 22276 10345 22332
rect 10345 22276 10349 22332
rect 10285 22272 10349 22276
rect 10365 22332 10429 22336
rect 10365 22276 10369 22332
rect 10369 22276 10425 22332
rect 10425 22276 10429 22332
rect 10365 22272 10429 22276
rect 10445 22332 10509 22336
rect 10445 22276 10449 22332
rect 10449 22276 10505 22332
rect 10505 22276 10509 22332
rect 10445 22272 10509 22276
rect 10525 22332 10589 22336
rect 10525 22276 10529 22332
rect 10529 22276 10585 22332
rect 10585 22276 10589 22332
rect 10525 22272 10589 22276
rect 19618 22332 19682 22336
rect 19618 22276 19622 22332
rect 19622 22276 19678 22332
rect 19678 22276 19682 22332
rect 19618 22272 19682 22276
rect 19698 22332 19762 22336
rect 19698 22276 19702 22332
rect 19702 22276 19758 22332
rect 19758 22276 19762 22332
rect 19698 22272 19762 22276
rect 19778 22332 19842 22336
rect 19778 22276 19782 22332
rect 19782 22276 19838 22332
rect 19838 22276 19842 22332
rect 19778 22272 19842 22276
rect 19858 22332 19922 22336
rect 19858 22276 19862 22332
rect 19862 22276 19918 22332
rect 19918 22276 19922 22332
rect 19858 22272 19922 22276
rect 21036 21796 21100 21860
rect 5618 21788 5682 21792
rect 5618 21732 5622 21788
rect 5622 21732 5678 21788
rect 5678 21732 5682 21788
rect 5618 21728 5682 21732
rect 5698 21788 5762 21792
rect 5698 21732 5702 21788
rect 5702 21732 5758 21788
rect 5758 21732 5762 21788
rect 5698 21728 5762 21732
rect 5778 21788 5842 21792
rect 5778 21732 5782 21788
rect 5782 21732 5838 21788
rect 5838 21732 5842 21788
rect 5778 21728 5842 21732
rect 5858 21788 5922 21792
rect 5858 21732 5862 21788
rect 5862 21732 5918 21788
rect 5918 21732 5922 21788
rect 5858 21728 5922 21732
rect 14952 21788 15016 21792
rect 14952 21732 14956 21788
rect 14956 21732 15012 21788
rect 15012 21732 15016 21788
rect 14952 21728 15016 21732
rect 15032 21788 15096 21792
rect 15032 21732 15036 21788
rect 15036 21732 15092 21788
rect 15092 21732 15096 21788
rect 15032 21728 15096 21732
rect 15112 21788 15176 21792
rect 15112 21732 15116 21788
rect 15116 21732 15172 21788
rect 15172 21732 15176 21788
rect 15112 21728 15176 21732
rect 15192 21788 15256 21792
rect 15192 21732 15196 21788
rect 15196 21732 15252 21788
rect 15252 21732 15256 21788
rect 15192 21728 15256 21732
rect 24285 21788 24349 21792
rect 24285 21732 24289 21788
rect 24289 21732 24345 21788
rect 24345 21732 24349 21788
rect 24285 21728 24349 21732
rect 24365 21788 24429 21792
rect 24365 21732 24369 21788
rect 24369 21732 24425 21788
rect 24425 21732 24429 21788
rect 24365 21728 24429 21732
rect 24445 21788 24509 21792
rect 24445 21732 24449 21788
rect 24449 21732 24505 21788
rect 24505 21732 24509 21788
rect 24445 21728 24509 21732
rect 24525 21788 24589 21792
rect 24525 21732 24529 21788
rect 24529 21732 24585 21788
rect 24585 21732 24589 21788
rect 24525 21728 24589 21732
rect 2636 21524 2700 21588
rect 9260 21388 9324 21452
rect 21772 21524 21836 21588
rect 10285 21244 10349 21248
rect 10285 21188 10289 21244
rect 10289 21188 10345 21244
rect 10345 21188 10349 21244
rect 10285 21184 10349 21188
rect 10365 21244 10429 21248
rect 10365 21188 10369 21244
rect 10369 21188 10425 21244
rect 10425 21188 10429 21244
rect 10365 21184 10429 21188
rect 10445 21244 10509 21248
rect 10445 21188 10449 21244
rect 10449 21188 10505 21244
rect 10505 21188 10509 21244
rect 10445 21184 10509 21188
rect 10525 21244 10589 21248
rect 10525 21188 10529 21244
rect 10529 21188 10585 21244
rect 10585 21188 10589 21244
rect 10525 21184 10589 21188
rect 19618 21244 19682 21248
rect 19618 21188 19622 21244
rect 19622 21188 19678 21244
rect 19678 21188 19682 21244
rect 19618 21184 19682 21188
rect 19698 21244 19762 21248
rect 19698 21188 19702 21244
rect 19702 21188 19758 21244
rect 19758 21188 19762 21244
rect 19698 21184 19762 21188
rect 19778 21244 19842 21248
rect 19778 21188 19782 21244
rect 19782 21188 19838 21244
rect 19838 21188 19842 21244
rect 19778 21184 19842 21188
rect 19858 21244 19922 21248
rect 19858 21188 19862 21244
rect 19862 21188 19918 21244
rect 19918 21188 19922 21244
rect 19858 21184 19922 21188
rect 2084 20844 2148 20908
rect 5396 20708 5460 20772
rect 5618 20700 5682 20704
rect 5618 20644 5622 20700
rect 5622 20644 5678 20700
rect 5678 20644 5682 20700
rect 5618 20640 5682 20644
rect 5698 20700 5762 20704
rect 5698 20644 5702 20700
rect 5702 20644 5758 20700
rect 5758 20644 5762 20700
rect 5698 20640 5762 20644
rect 5778 20700 5842 20704
rect 5778 20644 5782 20700
rect 5782 20644 5838 20700
rect 5838 20644 5842 20700
rect 5778 20640 5842 20644
rect 5858 20700 5922 20704
rect 5858 20644 5862 20700
rect 5862 20644 5918 20700
rect 5918 20644 5922 20700
rect 5858 20640 5922 20644
rect 14952 20700 15016 20704
rect 14952 20644 14956 20700
rect 14956 20644 15012 20700
rect 15012 20644 15016 20700
rect 14952 20640 15016 20644
rect 15032 20700 15096 20704
rect 15032 20644 15036 20700
rect 15036 20644 15092 20700
rect 15092 20644 15096 20700
rect 15032 20640 15096 20644
rect 15112 20700 15176 20704
rect 15112 20644 15116 20700
rect 15116 20644 15172 20700
rect 15172 20644 15176 20700
rect 15112 20640 15176 20644
rect 15192 20700 15256 20704
rect 15192 20644 15196 20700
rect 15196 20644 15252 20700
rect 15252 20644 15256 20700
rect 15192 20640 15256 20644
rect 24285 20700 24349 20704
rect 24285 20644 24289 20700
rect 24289 20644 24345 20700
rect 24345 20644 24349 20700
rect 24285 20640 24349 20644
rect 24365 20700 24429 20704
rect 24365 20644 24369 20700
rect 24369 20644 24425 20700
rect 24425 20644 24429 20700
rect 24365 20640 24429 20644
rect 24445 20700 24509 20704
rect 24445 20644 24449 20700
rect 24449 20644 24505 20700
rect 24505 20644 24509 20700
rect 24445 20640 24509 20644
rect 24525 20700 24589 20704
rect 24525 20644 24529 20700
rect 24529 20644 24585 20700
rect 24585 20644 24589 20700
rect 24525 20640 24589 20644
rect 14780 20300 14844 20364
rect 10916 20224 10980 20228
rect 10916 20168 10930 20224
rect 10930 20168 10980 20224
rect 10916 20164 10980 20168
rect 10285 20156 10349 20160
rect 10285 20100 10289 20156
rect 10289 20100 10345 20156
rect 10345 20100 10349 20156
rect 10285 20096 10349 20100
rect 10365 20156 10429 20160
rect 10365 20100 10369 20156
rect 10369 20100 10425 20156
rect 10425 20100 10429 20156
rect 10365 20096 10429 20100
rect 10445 20156 10509 20160
rect 10445 20100 10449 20156
rect 10449 20100 10505 20156
rect 10505 20100 10509 20156
rect 10445 20096 10509 20100
rect 10525 20156 10589 20160
rect 10525 20100 10529 20156
rect 10529 20100 10585 20156
rect 10585 20100 10589 20156
rect 10525 20096 10589 20100
rect 19618 20156 19682 20160
rect 19618 20100 19622 20156
rect 19622 20100 19678 20156
rect 19678 20100 19682 20156
rect 19618 20096 19682 20100
rect 19698 20156 19762 20160
rect 19698 20100 19702 20156
rect 19702 20100 19758 20156
rect 19758 20100 19762 20156
rect 19698 20096 19762 20100
rect 19778 20156 19842 20160
rect 19778 20100 19782 20156
rect 19782 20100 19838 20156
rect 19838 20100 19842 20156
rect 19778 20096 19842 20100
rect 19858 20156 19922 20160
rect 19858 20100 19862 20156
rect 19862 20100 19918 20156
rect 19918 20100 19922 20156
rect 19858 20096 19922 20100
rect 17724 20088 17788 20092
rect 17724 20032 17738 20088
rect 17738 20032 17788 20088
rect 17724 20028 17788 20032
rect 5618 19612 5682 19616
rect 5618 19556 5622 19612
rect 5622 19556 5678 19612
rect 5678 19556 5682 19612
rect 5618 19552 5682 19556
rect 5698 19612 5762 19616
rect 5698 19556 5702 19612
rect 5702 19556 5758 19612
rect 5758 19556 5762 19612
rect 5698 19552 5762 19556
rect 5778 19612 5842 19616
rect 5778 19556 5782 19612
rect 5782 19556 5838 19612
rect 5838 19556 5842 19612
rect 5778 19552 5842 19556
rect 5858 19612 5922 19616
rect 5858 19556 5862 19612
rect 5862 19556 5918 19612
rect 5918 19556 5922 19612
rect 5858 19552 5922 19556
rect 9076 19484 9140 19548
rect 10732 19620 10796 19684
rect 14952 19612 15016 19616
rect 14952 19556 14956 19612
rect 14956 19556 15012 19612
rect 15012 19556 15016 19612
rect 14952 19552 15016 19556
rect 15032 19612 15096 19616
rect 15032 19556 15036 19612
rect 15036 19556 15092 19612
rect 15092 19556 15096 19612
rect 15032 19552 15096 19556
rect 15112 19612 15176 19616
rect 15112 19556 15116 19612
rect 15116 19556 15172 19612
rect 15172 19556 15176 19612
rect 15112 19552 15176 19556
rect 15192 19612 15256 19616
rect 15192 19556 15196 19612
rect 15196 19556 15252 19612
rect 15252 19556 15256 19612
rect 15192 19552 15256 19556
rect 14780 19484 14844 19548
rect 20116 19756 20180 19820
rect 24285 19612 24349 19616
rect 24285 19556 24289 19612
rect 24289 19556 24345 19612
rect 24345 19556 24349 19612
rect 24285 19552 24349 19556
rect 24365 19612 24429 19616
rect 24365 19556 24369 19612
rect 24369 19556 24425 19612
rect 24425 19556 24429 19612
rect 24365 19552 24429 19556
rect 24445 19612 24509 19616
rect 24445 19556 24449 19612
rect 24449 19556 24505 19612
rect 24505 19556 24509 19612
rect 24445 19552 24509 19556
rect 24525 19612 24589 19616
rect 24525 19556 24529 19612
rect 24529 19556 24585 19612
rect 24585 19556 24589 19612
rect 24525 19552 24589 19556
rect 2268 19212 2332 19276
rect 12940 19076 13004 19140
rect 19380 19136 19444 19140
rect 19380 19080 19430 19136
rect 19430 19080 19444 19136
rect 19380 19076 19444 19080
rect 20300 19076 20364 19140
rect 23796 19076 23860 19140
rect 10285 19068 10349 19072
rect 10285 19012 10289 19068
rect 10289 19012 10345 19068
rect 10345 19012 10349 19068
rect 10285 19008 10349 19012
rect 10365 19068 10429 19072
rect 10365 19012 10369 19068
rect 10369 19012 10425 19068
rect 10425 19012 10429 19068
rect 10365 19008 10429 19012
rect 10445 19068 10509 19072
rect 10445 19012 10449 19068
rect 10449 19012 10505 19068
rect 10505 19012 10509 19068
rect 10445 19008 10509 19012
rect 10525 19068 10589 19072
rect 10525 19012 10529 19068
rect 10529 19012 10585 19068
rect 10585 19012 10589 19068
rect 10525 19008 10589 19012
rect 19618 19068 19682 19072
rect 19618 19012 19622 19068
rect 19622 19012 19678 19068
rect 19678 19012 19682 19068
rect 19618 19008 19682 19012
rect 19698 19068 19762 19072
rect 19698 19012 19702 19068
rect 19702 19012 19758 19068
rect 19758 19012 19762 19068
rect 19698 19008 19762 19012
rect 19778 19068 19842 19072
rect 19778 19012 19782 19068
rect 19782 19012 19838 19068
rect 19838 19012 19842 19068
rect 19778 19008 19842 19012
rect 19858 19068 19922 19072
rect 19858 19012 19862 19068
rect 19862 19012 19918 19068
rect 19918 19012 19922 19068
rect 19858 19008 19922 19012
rect 5618 18524 5682 18528
rect 5618 18468 5622 18524
rect 5622 18468 5678 18524
rect 5678 18468 5682 18524
rect 5618 18464 5682 18468
rect 5698 18524 5762 18528
rect 5698 18468 5702 18524
rect 5702 18468 5758 18524
rect 5758 18468 5762 18524
rect 5698 18464 5762 18468
rect 5778 18524 5842 18528
rect 5778 18468 5782 18524
rect 5782 18468 5838 18524
rect 5838 18468 5842 18524
rect 5778 18464 5842 18468
rect 5858 18524 5922 18528
rect 5858 18468 5862 18524
rect 5862 18468 5918 18524
rect 5918 18468 5922 18524
rect 5858 18464 5922 18468
rect 14952 18524 15016 18528
rect 14952 18468 14956 18524
rect 14956 18468 15012 18524
rect 15012 18468 15016 18524
rect 14952 18464 15016 18468
rect 15032 18524 15096 18528
rect 15032 18468 15036 18524
rect 15036 18468 15092 18524
rect 15092 18468 15096 18524
rect 15032 18464 15096 18468
rect 15112 18524 15176 18528
rect 15112 18468 15116 18524
rect 15116 18468 15172 18524
rect 15172 18468 15176 18524
rect 15112 18464 15176 18468
rect 15192 18524 15256 18528
rect 15192 18468 15196 18524
rect 15196 18468 15252 18524
rect 15252 18468 15256 18524
rect 15192 18464 15256 18468
rect 24285 18524 24349 18528
rect 24285 18468 24289 18524
rect 24289 18468 24345 18524
rect 24345 18468 24349 18524
rect 24285 18464 24349 18468
rect 24365 18524 24429 18528
rect 24365 18468 24369 18524
rect 24369 18468 24425 18524
rect 24425 18468 24429 18524
rect 24365 18464 24429 18468
rect 24445 18524 24509 18528
rect 24445 18468 24449 18524
rect 24449 18468 24505 18524
rect 24505 18468 24509 18524
rect 24445 18464 24509 18468
rect 24525 18524 24589 18528
rect 24525 18468 24529 18524
rect 24529 18468 24585 18524
rect 24585 18468 24589 18524
rect 24525 18464 24589 18468
rect 20300 17988 20364 18052
rect 21036 17988 21100 18052
rect 10285 17980 10349 17984
rect 10285 17924 10289 17980
rect 10289 17924 10345 17980
rect 10345 17924 10349 17980
rect 10285 17920 10349 17924
rect 10365 17980 10429 17984
rect 10365 17924 10369 17980
rect 10369 17924 10425 17980
rect 10425 17924 10429 17980
rect 10365 17920 10429 17924
rect 10445 17980 10509 17984
rect 10445 17924 10449 17980
rect 10449 17924 10505 17980
rect 10505 17924 10509 17980
rect 10445 17920 10509 17924
rect 10525 17980 10589 17984
rect 10525 17924 10529 17980
rect 10529 17924 10585 17980
rect 10585 17924 10589 17980
rect 10525 17920 10589 17924
rect 19618 17980 19682 17984
rect 19618 17924 19622 17980
rect 19622 17924 19678 17980
rect 19678 17924 19682 17980
rect 19618 17920 19682 17924
rect 19698 17980 19762 17984
rect 19698 17924 19702 17980
rect 19702 17924 19758 17980
rect 19758 17924 19762 17980
rect 19698 17920 19762 17924
rect 19778 17980 19842 17984
rect 19778 17924 19782 17980
rect 19782 17924 19838 17980
rect 19838 17924 19842 17980
rect 19778 17920 19842 17924
rect 19858 17980 19922 17984
rect 19858 17924 19862 17980
rect 19862 17924 19918 17980
rect 19918 17924 19922 17980
rect 19858 17920 19922 17924
rect 10916 17852 10980 17916
rect 22508 17852 22572 17916
rect 25268 17852 25332 17916
rect 20116 17716 20180 17780
rect 5618 17436 5682 17440
rect 5618 17380 5622 17436
rect 5622 17380 5678 17436
rect 5678 17380 5682 17436
rect 5618 17376 5682 17380
rect 5698 17436 5762 17440
rect 5698 17380 5702 17436
rect 5702 17380 5758 17436
rect 5758 17380 5762 17436
rect 5698 17376 5762 17380
rect 5778 17436 5842 17440
rect 5778 17380 5782 17436
rect 5782 17380 5838 17436
rect 5838 17380 5842 17436
rect 5778 17376 5842 17380
rect 5858 17436 5922 17440
rect 5858 17380 5862 17436
rect 5862 17380 5918 17436
rect 5918 17380 5922 17436
rect 5858 17376 5922 17380
rect 14952 17436 15016 17440
rect 14952 17380 14956 17436
rect 14956 17380 15012 17436
rect 15012 17380 15016 17436
rect 14952 17376 15016 17380
rect 15032 17436 15096 17440
rect 15032 17380 15036 17436
rect 15036 17380 15092 17436
rect 15092 17380 15096 17436
rect 15032 17376 15096 17380
rect 15112 17436 15176 17440
rect 15112 17380 15116 17436
rect 15116 17380 15172 17436
rect 15172 17380 15176 17436
rect 15112 17376 15176 17380
rect 15192 17436 15256 17440
rect 15192 17380 15196 17436
rect 15196 17380 15252 17436
rect 15252 17380 15256 17436
rect 15192 17376 15256 17380
rect 10916 17308 10980 17372
rect 24285 17436 24349 17440
rect 24285 17380 24289 17436
rect 24289 17380 24345 17436
rect 24345 17380 24349 17436
rect 24285 17376 24349 17380
rect 24365 17436 24429 17440
rect 24365 17380 24369 17436
rect 24369 17380 24425 17436
rect 24425 17380 24429 17436
rect 24365 17376 24429 17380
rect 24445 17436 24509 17440
rect 24445 17380 24449 17436
rect 24449 17380 24505 17436
rect 24505 17380 24509 17436
rect 24445 17376 24509 17380
rect 24525 17436 24589 17440
rect 24525 17380 24529 17436
rect 24529 17380 24585 17436
rect 24585 17380 24589 17436
rect 24525 17376 24589 17380
rect 6132 17172 6196 17236
rect 22876 17172 22940 17236
rect 10285 16892 10349 16896
rect 10285 16836 10289 16892
rect 10289 16836 10345 16892
rect 10345 16836 10349 16892
rect 10285 16832 10349 16836
rect 10365 16892 10429 16896
rect 10365 16836 10369 16892
rect 10369 16836 10425 16892
rect 10425 16836 10429 16892
rect 10365 16832 10429 16836
rect 10445 16892 10509 16896
rect 10445 16836 10449 16892
rect 10449 16836 10505 16892
rect 10505 16836 10509 16892
rect 10445 16832 10509 16836
rect 10525 16892 10589 16896
rect 10525 16836 10529 16892
rect 10529 16836 10585 16892
rect 10585 16836 10589 16892
rect 10525 16832 10589 16836
rect 20116 17036 20180 17100
rect 20484 17036 20548 17100
rect 20668 16900 20732 16964
rect 19618 16892 19682 16896
rect 19618 16836 19622 16892
rect 19622 16836 19678 16892
rect 19678 16836 19682 16892
rect 19618 16832 19682 16836
rect 19698 16892 19762 16896
rect 19698 16836 19702 16892
rect 19702 16836 19758 16892
rect 19758 16836 19762 16892
rect 19698 16832 19762 16836
rect 19778 16892 19842 16896
rect 19778 16836 19782 16892
rect 19782 16836 19838 16892
rect 19838 16836 19842 16892
rect 19778 16832 19842 16836
rect 19858 16892 19922 16896
rect 19858 16836 19862 16892
rect 19862 16836 19918 16892
rect 19918 16836 19922 16892
rect 19858 16832 19922 16836
rect 6684 16356 6748 16420
rect 5618 16348 5682 16352
rect 5618 16292 5622 16348
rect 5622 16292 5678 16348
rect 5678 16292 5682 16348
rect 5618 16288 5682 16292
rect 5698 16348 5762 16352
rect 5698 16292 5702 16348
rect 5702 16292 5758 16348
rect 5758 16292 5762 16348
rect 5698 16288 5762 16292
rect 5778 16348 5842 16352
rect 5778 16292 5782 16348
rect 5782 16292 5838 16348
rect 5838 16292 5842 16348
rect 5778 16288 5842 16292
rect 5858 16348 5922 16352
rect 5858 16292 5862 16348
rect 5862 16292 5918 16348
rect 5918 16292 5922 16348
rect 5858 16288 5922 16292
rect 14952 16348 15016 16352
rect 14952 16292 14956 16348
rect 14956 16292 15012 16348
rect 15012 16292 15016 16348
rect 14952 16288 15016 16292
rect 15032 16348 15096 16352
rect 15032 16292 15036 16348
rect 15036 16292 15092 16348
rect 15092 16292 15096 16348
rect 15032 16288 15096 16292
rect 15112 16348 15176 16352
rect 15112 16292 15116 16348
rect 15116 16292 15172 16348
rect 15172 16292 15176 16348
rect 15112 16288 15176 16292
rect 15192 16348 15256 16352
rect 15192 16292 15196 16348
rect 15196 16292 15252 16348
rect 15252 16292 15256 16348
rect 15192 16288 15256 16292
rect 24285 16348 24349 16352
rect 24285 16292 24289 16348
rect 24289 16292 24345 16348
rect 24345 16292 24349 16348
rect 24285 16288 24349 16292
rect 24365 16348 24429 16352
rect 24365 16292 24369 16348
rect 24369 16292 24425 16348
rect 24425 16292 24429 16348
rect 24365 16288 24429 16292
rect 24445 16348 24509 16352
rect 24445 16292 24449 16348
rect 24449 16292 24505 16348
rect 24505 16292 24509 16348
rect 24445 16288 24509 16292
rect 24525 16348 24589 16352
rect 24525 16292 24529 16348
rect 24529 16292 24585 16348
rect 24585 16292 24589 16348
rect 24525 16288 24589 16292
rect 9996 16220 10060 16284
rect 14596 16220 14660 16284
rect 13308 16008 13372 16012
rect 13308 15952 13322 16008
rect 13322 15952 13372 16008
rect 13308 15948 13372 15952
rect 21036 15948 21100 16012
rect 20852 15872 20916 15876
rect 20852 15816 20902 15872
rect 20902 15816 20916 15872
rect 20852 15812 20916 15816
rect 10285 15804 10349 15808
rect 10285 15748 10289 15804
rect 10289 15748 10345 15804
rect 10345 15748 10349 15804
rect 10285 15744 10349 15748
rect 10365 15804 10429 15808
rect 10365 15748 10369 15804
rect 10369 15748 10425 15804
rect 10425 15748 10429 15804
rect 10365 15744 10429 15748
rect 10445 15804 10509 15808
rect 10445 15748 10449 15804
rect 10449 15748 10505 15804
rect 10505 15748 10509 15804
rect 10445 15744 10509 15748
rect 10525 15804 10589 15808
rect 10525 15748 10529 15804
rect 10529 15748 10585 15804
rect 10585 15748 10589 15804
rect 10525 15744 10589 15748
rect 19618 15804 19682 15808
rect 19618 15748 19622 15804
rect 19622 15748 19678 15804
rect 19678 15748 19682 15804
rect 19618 15744 19682 15748
rect 19698 15804 19762 15808
rect 19698 15748 19702 15804
rect 19702 15748 19758 15804
rect 19758 15748 19762 15804
rect 19698 15744 19762 15748
rect 19778 15804 19842 15808
rect 19778 15748 19782 15804
rect 19782 15748 19838 15804
rect 19838 15748 19842 15804
rect 19778 15744 19842 15748
rect 19858 15804 19922 15808
rect 19858 15748 19862 15804
rect 19862 15748 19918 15804
rect 19918 15748 19922 15804
rect 19858 15744 19922 15748
rect 6132 15676 6196 15740
rect 5618 15260 5682 15264
rect 5618 15204 5622 15260
rect 5622 15204 5678 15260
rect 5678 15204 5682 15260
rect 5618 15200 5682 15204
rect 5698 15260 5762 15264
rect 5698 15204 5702 15260
rect 5702 15204 5758 15260
rect 5758 15204 5762 15260
rect 5698 15200 5762 15204
rect 5778 15260 5842 15264
rect 5778 15204 5782 15260
rect 5782 15204 5838 15260
rect 5838 15204 5842 15260
rect 5778 15200 5842 15204
rect 5858 15260 5922 15264
rect 5858 15204 5862 15260
rect 5862 15204 5918 15260
rect 5918 15204 5922 15260
rect 5858 15200 5922 15204
rect 14952 15260 15016 15264
rect 14952 15204 14956 15260
rect 14956 15204 15012 15260
rect 15012 15204 15016 15260
rect 14952 15200 15016 15204
rect 15032 15260 15096 15264
rect 15032 15204 15036 15260
rect 15036 15204 15092 15260
rect 15092 15204 15096 15260
rect 15032 15200 15096 15204
rect 15112 15260 15176 15264
rect 15112 15204 15116 15260
rect 15116 15204 15172 15260
rect 15172 15204 15176 15260
rect 15112 15200 15176 15204
rect 15192 15260 15256 15264
rect 15192 15204 15196 15260
rect 15196 15204 15252 15260
rect 15252 15204 15256 15260
rect 15192 15200 15256 15204
rect 24285 15260 24349 15264
rect 24285 15204 24289 15260
rect 24289 15204 24345 15260
rect 24345 15204 24349 15260
rect 24285 15200 24349 15204
rect 24365 15260 24429 15264
rect 24365 15204 24369 15260
rect 24369 15204 24425 15260
rect 24425 15204 24429 15260
rect 24365 15200 24429 15204
rect 24445 15260 24509 15264
rect 24445 15204 24449 15260
rect 24449 15204 24505 15260
rect 24505 15204 24509 15260
rect 24445 15200 24509 15204
rect 24525 15260 24589 15264
rect 24525 15204 24529 15260
rect 24529 15204 24585 15260
rect 24585 15204 24589 15260
rect 24525 15200 24589 15204
rect 13860 15132 13924 15196
rect 20300 14996 20364 15060
rect 23244 14996 23308 15060
rect 24900 14996 24964 15060
rect 20484 14860 20548 14924
rect 6316 14724 6380 14788
rect 24716 14724 24780 14788
rect 10285 14716 10349 14720
rect 10285 14660 10289 14716
rect 10289 14660 10345 14716
rect 10345 14660 10349 14716
rect 10285 14656 10349 14660
rect 10365 14716 10429 14720
rect 10365 14660 10369 14716
rect 10369 14660 10425 14716
rect 10425 14660 10429 14716
rect 10365 14656 10429 14660
rect 10445 14716 10509 14720
rect 10445 14660 10449 14716
rect 10449 14660 10505 14716
rect 10505 14660 10509 14716
rect 10445 14656 10509 14660
rect 10525 14716 10589 14720
rect 10525 14660 10529 14716
rect 10529 14660 10585 14716
rect 10585 14660 10589 14716
rect 10525 14656 10589 14660
rect 19618 14716 19682 14720
rect 19618 14660 19622 14716
rect 19622 14660 19678 14716
rect 19678 14660 19682 14716
rect 19618 14656 19682 14660
rect 19698 14716 19762 14720
rect 19698 14660 19702 14716
rect 19702 14660 19758 14716
rect 19758 14660 19762 14716
rect 19698 14656 19762 14660
rect 19778 14716 19842 14720
rect 19778 14660 19782 14716
rect 19782 14660 19838 14716
rect 19838 14660 19842 14716
rect 19778 14656 19842 14660
rect 19858 14716 19922 14720
rect 19858 14660 19862 14716
rect 19862 14660 19918 14716
rect 19918 14660 19922 14716
rect 19858 14656 19922 14660
rect 9628 14588 9692 14652
rect 5618 14172 5682 14176
rect 5618 14116 5622 14172
rect 5622 14116 5678 14172
rect 5678 14116 5682 14172
rect 5618 14112 5682 14116
rect 5698 14172 5762 14176
rect 5698 14116 5702 14172
rect 5702 14116 5758 14172
rect 5758 14116 5762 14172
rect 5698 14112 5762 14116
rect 5778 14172 5842 14176
rect 5778 14116 5782 14172
rect 5782 14116 5838 14172
rect 5838 14116 5842 14172
rect 5778 14112 5842 14116
rect 5858 14172 5922 14176
rect 5858 14116 5862 14172
rect 5862 14116 5918 14172
rect 5918 14116 5922 14172
rect 5858 14112 5922 14116
rect 2452 13908 2516 13972
rect 14228 14180 14292 14244
rect 22324 14180 22388 14244
rect 14952 14172 15016 14176
rect 14952 14116 14956 14172
rect 14956 14116 15012 14172
rect 15012 14116 15016 14172
rect 14952 14112 15016 14116
rect 15032 14172 15096 14176
rect 15032 14116 15036 14172
rect 15036 14116 15092 14172
rect 15092 14116 15096 14172
rect 15032 14112 15096 14116
rect 15112 14172 15176 14176
rect 15112 14116 15116 14172
rect 15116 14116 15172 14172
rect 15172 14116 15176 14172
rect 15112 14112 15176 14116
rect 15192 14172 15256 14176
rect 15192 14116 15196 14172
rect 15196 14116 15252 14172
rect 15252 14116 15256 14172
rect 15192 14112 15256 14116
rect 24285 14172 24349 14176
rect 24285 14116 24289 14172
rect 24289 14116 24345 14172
rect 24345 14116 24349 14172
rect 24285 14112 24349 14116
rect 24365 14172 24429 14176
rect 24365 14116 24369 14172
rect 24369 14116 24425 14172
rect 24425 14116 24429 14172
rect 24365 14112 24429 14116
rect 24445 14172 24509 14176
rect 24445 14116 24449 14172
rect 24449 14116 24505 14172
rect 24505 14116 24509 14172
rect 24445 14112 24509 14116
rect 24525 14172 24589 14176
rect 24525 14116 24529 14172
rect 24529 14116 24585 14172
rect 24585 14116 24589 14172
rect 24525 14112 24589 14116
rect 11100 14044 11164 14108
rect 20852 13772 20916 13836
rect 21036 13832 21100 13836
rect 21036 13776 21086 13832
rect 21086 13776 21100 13832
rect 21036 13772 21100 13776
rect 5212 13636 5276 13700
rect 9812 13696 9876 13700
rect 9812 13640 9826 13696
rect 9826 13640 9876 13696
rect 9812 13636 9876 13640
rect 20668 13636 20732 13700
rect 10285 13628 10349 13632
rect 10285 13572 10289 13628
rect 10289 13572 10345 13628
rect 10345 13572 10349 13628
rect 10285 13568 10349 13572
rect 10365 13628 10429 13632
rect 10365 13572 10369 13628
rect 10369 13572 10425 13628
rect 10425 13572 10429 13628
rect 10365 13568 10429 13572
rect 10445 13628 10509 13632
rect 10445 13572 10449 13628
rect 10449 13572 10505 13628
rect 10505 13572 10509 13628
rect 10445 13568 10509 13572
rect 10525 13628 10589 13632
rect 10525 13572 10529 13628
rect 10529 13572 10585 13628
rect 10585 13572 10589 13628
rect 10525 13568 10589 13572
rect 19618 13628 19682 13632
rect 19618 13572 19622 13628
rect 19622 13572 19678 13628
rect 19678 13572 19682 13628
rect 19618 13568 19682 13572
rect 19698 13628 19762 13632
rect 19698 13572 19702 13628
rect 19702 13572 19758 13628
rect 19758 13572 19762 13628
rect 19698 13568 19762 13572
rect 19778 13628 19842 13632
rect 19778 13572 19782 13628
rect 19782 13572 19838 13628
rect 19838 13572 19842 13628
rect 19778 13568 19842 13572
rect 19858 13628 19922 13632
rect 19858 13572 19862 13628
rect 19862 13572 19918 13628
rect 19918 13572 19922 13628
rect 19858 13568 19922 13572
rect 9628 13500 9692 13564
rect 24716 13364 24780 13428
rect 13676 13228 13740 13292
rect 20116 13092 20180 13156
rect 5618 13084 5682 13088
rect 5618 13028 5622 13084
rect 5622 13028 5678 13084
rect 5678 13028 5682 13084
rect 5618 13024 5682 13028
rect 5698 13084 5762 13088
rect 5698 13028 5702 13084
rect 5702 13028 5758 13084
rect 5758 13028 5762 13084
rect 5698 13024 5762 13028
rect 5778 13084 5842 13088
rect 5778 13028 5782 13084
rect 5782 13028 5838 13084
rect 5838 13028 5842 13084
rect 5778 13024 5842 13028
rect 5858 13084 5922 13088
rect 5858 13028 5862 13084
rect 5862 13028 5918 13084
rect 5918 13028 5922 13084
rect 5858 13024 5922 13028
rect 14952 13084 15016 13088
rect 14952 13028 14956 13084
rect 14956 13028 15012 13084
rect 15012 13028 15016 13084
rect 14952 13024 15016 13028
rect 15032 13084 15096 13088
rect 15032 13028 15036 13084
rect 15036 13028 15092 13084
rect 15092 13028 15096 13084
rect 15032 13024 15096 13028
rect 15112 13084 15176 13088
rect 15112 13028 15116 13084
rect 15116 13028 15172 13084
rect 15172 13028 15176 13084
rect 15112 13024 15176 13028
rect 15192 13084 15256 13088
rect 15192 13028 15196 13084
rect 15196 13028 15252 13084
rect 15252 13028 15256 13084
rect 15192 13024 15256 13028
rect 24285 13084 24349 13088
rect 24285 13028 24289 13084
rect 24289 13028 24345 13084
rect 24345 13028 24349 13084
rect 24285 13024 24349 13028
rect 24365 13084 24429 13088
rect 24365 13028 24369 13084
rect 24369 13028 24425 13084
rect 24425 13028 24429 13084
rect 24365 13024 24429 13028
rect 24445 13084 24509 13088
rect 24445 13028 24449 13084
rect 24449 13028 24505 13084
rect 24505 13028 24509 13084
rect 24445 13024 24509 13028
rect 24525 13084 24589 13088
rect 24525 13028 24529 13084
rect 24529 13028 24585 13084
rect 24585 13028 24589 13084
rect 24525 13024 24589 13028
rect 2084 13016 2148 13020
rect 2084 12960 2098 13016
rect 2098 12960 2148 13016
rect 2084 12956 2148 12960
rect 4844 13016 4908 13020
rect 4844 12960 4894 13016
rect 4894 12960 4908 13016
rect 4844 12956 4908 12960
rect 15884 12956 15948 13020
rect 6132 12820 6196 12884
rect 17724 12956 17788 13020
rect 19380 12956 19444 13020
rect 21036 12820 21100 12884
rect 12940 12548 13004 12612
rect 10285 12540 10349 12544
rect 10285 12484 10289 12540
rect 10289 12484 10345 12540
rect 10345 12484 10349 12540
rect 10285 12480 10349 12484
rect 10365 12540 10429 12544
rect 10365 12484 10369 12540
rect 10369 12484 10425 12540
rect 10425 12484 10429 12540
rect 10365 12480 10429 12484
rect 10445 12540 10509 12544
rect 10445 12484 10449 12540
rect 10449 12484 10505 12540
rect 10505 12484 10509 12540
rect 10445 12480 10509 12484
rect 10525 12540 10589 12544
rect 10525 12484 10529 12540
rect 10529 12484 10585 12540
rect 10585 12484 10589 12540
rect 10525 12480 10589 12484
rect 19618 12540 19682 12544
rect 19618 12484 19622 12540
rect 19622 12484 19678 12540
rect 19678 12484 19682 12540
rect 19618 12480 19682 12484
rect 19698 12540 19762 12544
rect 19698 12484 19702 12540
rect 19702 12484 19758 12540
rect 19758 12484 19762 12540
rect 19698 12480 19762 12484
rect 19778 12540 19842 12544
rect 19778 12484 19782 12540
rect 19782 12484 19838 12540
rect 19838 12484 19842 12540
rect 19778 12480 19842 12484
rect 19858 12540 19922 12544
rect 19858 12484 19862 12540
rect 19862 12484 19918 12540
rect 19918 12484 19922 12540
rect 19858 12480 19922 12484
rect 21956 12684 22020 12748
rect 22508 12548 22572 12612
rect 25268 12412 25332 12476
rect 7604 12276 7668 12340
rect 3188 12140 3252 12204
rect 15516 12140 15580 12204
rect 3740 12004 3804 12068
rect 22140 12004 22204 12068
rect 23612 12140 23676 12204
rect 23980 12140 24044 12204
rect 5618 11996 5682 12000
rect 5618 11940 5622 11996
rect 5622 11940 5678 11996
rect 5678 11940 5682 11996
rect 5618 11936 5682 11940
rect 5698 11996 5762 12000
rect 5698 11940 5702 11996
rect 5702 11940 5758 11996
rect 5758 11940 5762 11996
rect 5698 11936 5762 11940
rect 5778 11996 5842 12000
rect 5778 11940 5782 11996
rect 5782 11940 5838 11996
rect 5838 11940 5842 11996
rect 5778 11936 5842 11940
rect 5858 11996 5922 12000
rect 5858 11940 5862 11996
rect 5862 11940 5918 11996
rect 5918 11940 5922 11996
rect 5858 11936 5922 11940
rect 14952 11996 15016 12000
rect 14952 11940 14956 11996
rect 14956 11940 15012 11996
rect 15012 11940 15016 11996
rect 14952 11936 15016 11940
rect 15032 11996 15096 12000
rect 15032 11940 15036 11996
rect 15036 11940 15092 11996
rect 15092 11940 15096 11996
rect 15032 11936 15096 11940
rect 15112 11996 15176 12000
rect 15112 11940 15116 11996
rect 15116 11940 15172 11996
rect 15172 11940 15176 11996
rect 15112 11936 15176 11940
rect 15192 11996 15256 12000
rect 15192 11940 15196 11996
rect 15196 11940 15252 11996
rect 15252 11940 15256 11996
rect 15192 11936 15256 11940
rect 24285 11996 24349 12000
rect 24285 11940 24289 11996
rect 24289 11940 24345 11996
rect 24345 11940 24349 11996
rect 24285 11936 24349 11940
rect 24365 11996 24429 12000
rect 24365 11940 24369 11996
rect 24369 11940 24425 11996
rect 24425 11940 24429 11996
rect 24365 11936 24429 11940
rect 24445 11996 24509 12000
rect 24445 11940 24449 11996
rect 24449 11940 24505 11996
rect 24505 11940 24509 11996
rect 24445 11936 24509 11940
rect 24525 11996 24589 12000
rect 24525 11940 24529 11996
rect 24529 11940 24585 11996
rect 24585 11940 24589 11996
rect 24525 11936 24589 11940
rect 7236 11928 7300 11932
rect 7236 11872 7286 11928
rect 7286 11872 7300 11928
rect 7236 11868 7300 11872
rect 7604 11868 7668 11932
rect 14044 11732 14108 11796
rect 14596 11596 14660 11660
rect 23980 11596 24044 11660
rect 22324 11460 22388 11524
rect 23428 11460 23492 11524
rect 10285 11452 10349 11456
rect 10285 11396 10289 11452
rect 10289 11396 10345 11452
rect 10345 11396 10349 11452
rect 10285 11392 10349 11396
rect 10365 11452 10429 11456
rect 10365 11396 10369 11452
rect 10369 11396 10425 11452
rect 10425 11396 10429 11452
rect 10365 11392 10429 11396
rect 10445 11452 10509 11456
rect 10445 11396 10449 11452
rect 10449 11396 10505 11452
rect 10505 11396 10509 11452
rect 10445 11392 10509 11396
rect 10525 11452 10589 11456
rect 10525 11396 10529 11452
rect 10529 11396 10585 11452
rect 10585 11396 10589 11452
rect 10525 11392 10589 11396
rect 19618 11452 19682 11456
rect 19618 11396 19622 11452
rect 19622 11396 19678 11452
rect 19678 11396 19682 11452
rect 19618 11392 19682 11396
rect 19698 11452 19762 11456
rect 19698 11396 19702 11452
rect 19702 11396 19758 11452
rect 19758 11396 19762 11452
rect 19698 11392 19762 11396
rect 19778 11452 19842 11456
rect 19778 11396 19782 11452
rect 19782 11396 19838 11452
rect 19838 11396 19842 11452
rect 19778 11392 19842 11396
rect 19858 11452 19922 11456
rect 19858 11396 19862 11452
rect 19862 11396 19918 11452
rect 19918 11396 19922 11452
rect 19858 11392 19922 11396
rect 5212 11248 5276 11252
rect 5212 11192 5226 11248
rect 5226 11192 5276 11248
rect 5212 11188 5276 11192
rect 21036 11324 21100 11388
rect 15884 11188 15948 11252
rect 7236 11052 7300 11116
rect 13860 11052 13924 11116
rect 25084 10976 25148 10980
rect 25084 10920 25134 10976
rect 25134 10920 25148 10976
rect 5618 10908 5682 10912
rect 5618 10852 5622 10908
rect 5622 10852 5678 10908
rect 5678 10852 5682 10908
rect 5618 10848 5682 10852
rect 5698 10908 5762 10912
rect 5698 10852 5702 10908
rect 5702 10852 5758 10908
rect 5758 10852 5762 10908
rect 5698 10848 5762 10852
rect 5778 10908 5842 10912
rect 5778 10852 5782 10908
rect 5782 10852 5838 10908
rect 5838 10852 5842 10908
rect 5778 10848 5842 10852
rect 5858 10908 5922 10912
rect 5858 10852 5862 10908
rect 5862 10852 5918 10908
rect 5918 10852 5922 10908
rect 5858 10848 5922 10852
rect 14952 10908 15016 10912
rect 14952 10852 14956 10908
rect 14956 10852 15012 10908
rect 15012 10852 15016 10908
rect 14952 10848 15016 10852
rect 15032 10908 15096 10912
rect 15032 10852 15036 10908
rect 15036 10852 15092 10908
rect 15092 10852 15096 10908
rect 15032 10848 15096 10852
rect 15112 10908 15176 10912
rect 15112 10852 15116 10908
rect 15116 10852 15172 10908
rect 15172 10852 15176 10908
rect 15112 10848 15176 10852
rect 15192 10908 15256 10912
rect 15192 10852 15196 10908
rect 15196 10852 15252 10908
rect 15252 10852 15256 10908
rect 15192 10848 15256 10852
rect 6500 10644 6564 10708
rect 25084 10916 25148 10920
rect 24285 10908 24349 10912
rect 24285 10852 24289 10908
rect 24289 10852 24345 10908
rect 24345 10852 24349 10908
rect 24285 10848 24349 10852
rect 24365 10908 24429 10912
rect 24365 10852 24369 10908
rect 24369 10852 24425 10908
rect 24425 10852 24429 10908
rect 24365 10848 24429 10852
rect 24445 10908 24509 10912
rect 24445 10852 24449 10908
rect 24449 10852 24505 10908
rect 24505 10852 24509 10908
rect 24445 10848 24509 10852
rect 24525 10908 24589 10912
rect 24525 10852 24529 10908
rect 24529 10852 24585 10908
rect 24585 10852 24589 10908
rect 24525 10848 24589 10852
rect 4844 10508 4908 10572
rect 10916 10508 10980 10572
rect 6500 10372 6564 10436
rect 20116 10372 20180 10436
rect 10285 10364 10349 10368
rect 10285 10308 10289 10364
rect 10289 10308 10345 10364
rect 10345 10308 10349 10364
rect 10285 10304 10349 10308
rect 10365 10364 10429 10368
rect 10365 10308 10369 10364
rect 10369 10308 10425 10364
rect 10425 10308 10429 10364
rect 10365 10304 10429 10308
rect 10445 10364 10509 10368
rect 10445 10308 10449 10364
rect 10449 10308 10505 10364
rect 10505 10308 10509 10364
rect 10445 10304 10509 10308
rect 10525 10364 10589 10368
rect 10525 10308 10529 10364
rect 10529 10308 10585 10364
rect 10585 10308 10589 10364
rect 10525 10304 10589 10308
rect 19618 10364 19682 10368
rect 19618 10308 19622 10364
rect 19622 10308 19678 10364
rect 19678 10308 19682 10364
rect 19618 10304 19682 10308
rect 19698 10364 19762 10368
rect 19698 10308 19702 10364
rect 19702 10308 19758 10364
rect 19758 10308 19762 10364
rect 19698 10304 19762 10308
rect 19778 10364 19842 10368
rect 19778 10308 19782 10364
rect 19782 10308 19838 10364
rect 19838 10308 19842 10364
rect 19778 10304 19842 10308
rect 19858 10364 19922 10368
rect 19858 10308 19862 10364
rect 19862 10308 19918 10364
rect 19918 10308 19922 10364
rect 19858 10304 19922 10308
rect 1716 10236 1780 10300
rect 10916 10236 10980 10300
rect 26740 10236 26804 10300
rect 3004 10024 3068 10028
rect 6132 10100 6196 10164
rect 3004 9968 3054 10024
rect 3054 9968 3068 10024
rect 3004 9964 3068 9968
rect 6500 9964 6564 10028
rect 5618 9820 5682 9824
rect 5618 9764 5622 9820
rect 5622 9764 5678 9820
rect 5678 9764 5682 9820
rect 5618 9760 5682 9764
rect 5698 9820 5762 9824
rect 5698 9764 5702 9820
rect 5702 9764 5758 9820
rect 5758 9764 5762 9820
rect 5698 9760 5762 9764
rect 5778 9820 5842 9824
rect 5778 9764 5782 9820
rect 5782 9764 5838 9820
rect 5838 9764 5842 9820
rect 5778 9760 5842 9764
rect 5858 9820 5922 9824
rect 5858 9764 5862 9820
rect 5862 9764 5918 9820
rect 5918 9764 5922 9820
rect 5858 9760 5922 9764
rect 6684 9752 6748 9756
rect 14952 9820 15016 9824
rect 14952 9764 14956 9820
rect 14956 9764 15012 9820
rect 15012 9764 15016 9820
rect 14952 9760 15016 9764
rect 15032 9820 15096 9824
rect 15032 9764 15036 9820
rect 15036 9764 15092 9820
rect 15092 9764 15096 9820
rect 15032 9760 15096 9764
rect 15112 9820 15176 9824
rect 15112 9764 15116 9820
rect 15116 9764 15172 9820
rect 15172 9764 15176 9820
rect 15112 9760 15176 9764
rect 15192 9820 15256 9824
rect 15192 9764 15196 9820
rect 15196 9764 15252 9820
rect 15252 9764 15256 9820
rect 15192 9760 15256 9764
rect 24285 9820 24349 9824
rect 24285 9764 24289 9820
rect 24289 9764 24345 9820
rect 24345 9764 24349 9820
rect 24285 9760 24349 9764
rect 24365 9820 24429 9824
rect 24365 9764 24369 9820
rect 24369 9764 24425 9820
rect 24425 9764 24429 9820
rect 24365 9760 24429 9764
rect 24445 9820 24509 9824
rect 24445 9764 24449 9820
rect 24449 9764 24505 9820
rect 24505 9764 24509 9820
rect 24445 9760 24509 9764
rect 24525 9820 24589 9824
rect 24525 9764 24529 9820
rect 24529 9764 24585 9820
rect 24585 9764 24589 9820
rect 24525 9760 24589 9764
rect 6684 9696 6698 9752
rect 6698 9696 6748 9752
rect 6684 9692 6748 9696
rect 9260 9556 9324 9620
rect 19380 9616 19444 9620
rect 19380 9560 19430 9616
rect 19430 9560 19444 9616
rect 19380 9556 19444 9560
rect 22876 9556 22940 9620
rect 25452 9556 25516 9620
rect 26372 9616 26436 9620
rect 26372 9560 26386 9616
rect 26386 9560 26436 9616
rect 26372 9556 26436 9560
rect 13860 9284 13924 9348
rect 20668 9284 20732 9348
rect 10285 9276 10349 9280
rect 10285 9220 10289 9276
rect 10289 9220 10345 9276
rect 10345 9220 10349 9276
rect 10285 9216 10349 9220
rect 10365 9276 10429 9280
rect 10365 9220 10369 9276
rect 10369 9220 10425 9276
rect 10425 9220 10429 9276
rect 10365 9216 10429 9220
rect 10445 9276 10509 9280
rect 10445 9220 10449 9276
rect 10449 9220 10505 9276
rect 10505 9220 10509 9276
rect 10445 9216 10509 9220
rect 10525 9276 10589 9280
rect 10525 9220 10529 9276
rect 10529 9220 10585 9276
rect 10585 9220 10589 9276
rect 10525 9216 10589 9220
rect 19618 9276 19682 9280
rect 19618 9220 19622 9276
rect 19622 9220 19678 9276
rect 19678 9220 19682 9276
rect 19618 9216 19682 9220
rect 19698 9276 19762 9280
rect 19698 9220 19702 9276
rect 19702 9220 19758 9276
rect 19758 9220 19762 9276
rect 19698 9216 19762 9220
rect 19778 9276 19842 9280
rect 19778 9220 19782 9276
rect 19782 9220 19838 9276
rect 19838 9220 19842 9276
rect 19778 9216 19842 9220
rect 19858 9276 19922 9280
rect 19858 9220 19862 9276
rect 19862 9220 19918 9276
rect 19918 9220 19922 9276
rect 19858 9216 19922 9220
rect 21220 9148 21284 9212
rect 21956 9148 22020 9212
rect 23980 9012 24044 9076
rect 2452 8876 2516 8940
rect 5396 8740 5460 8804
rect 21772 8800 21836 8804
rect 21772 8744 21822 8800
rect 21822 8744 21836 8800
rect 21772 8740 21836 8744
rect 5618 8732 5682 8736
rect 5618 8676 5622 8732
rect 5622 8676 5678 8732
rect 5678 8676 5682 8732
rect 5618 8672 5682 8676
rect 5698 8732 5762 8736
rect 5698 8676 5702 8732
rect 5702 8676 5758 8732
rect 5758 8676 5762 8732
rect 5698 8672 5762 8676
rect 5778 8732 5842 8736
rect 5778 8676 5782 8732
rect 5782 8676 5838 8732
rect 5838 8676 5842 8732
rect 5778 8672 5842 8676
rect 5858 8732 5922 8736
rect 5858 8676 5862 8732
rect 5862 8676 5918 8732
rect 5918 8676 5922 8732
rect 5858 8672 5922 8676
rect 14952 8732 15016 8736
rect 14952 8676 14956 8732
rect 14956 8676 15012 8732
rect 15012 8676 15016 8732
rect 14952 8672 15016 8676
rect 15032 8732 15096 8736
rect 15032 8676 15036 8732
rect 15036 8676 15092 8732
rect 15092 8676 15096 8732
rect 15032 8672 15096 8676
rect 15112 8732 15176 8736
rect 15112 8676 15116 8732
rect 15116 8676 15172 8732
rect 15172 8676 15176 8732
rect 15112 8672 15176 8676
rect 15192 8732 15256 8736
rect 15192 8676 15196 8732
rect 15196 8676 15252 8732
rect 15252 8676 15256 8732
rect 15192 8672 15256 8676
rect 24285 8732 24349 8736
rect 24285 8676 24289 8732
rect 24289 8676 24345 8732
rect 24345 8676 24349 8732
rect 24285 8672 24349 8676
rect 24365 8732 24429 8736
rect 24365 8676 24369 8732
rect 24369 8676 24425 8732
rect 24425 8676 24429 8732
rect 24365 8672 24429 8676
rect 24445 8732 24509 8736
rect 24445 8676 24449 8732
rect 24449 8676 24505 8732
rect 24505 8676 24509 8732
rect 24445 8672 24509 8676
rect 24525 8732 24589 8736
rect 24525 8676 24529 8732
rect 24529 8676 24585 8732
rect 24585 8676 24589 8732
rect 24525 8672 24589 8676
rect 20668 8528 20732 8532
rect 20668 8472 20682 8528
rect 20682 8472 20732 8528
rect 8156 8196 8220 8260
rect 20668 8468 20732 8472
rect 27292 8604 27356 8668
rect 15516 8392 15580 8396
rect 15516 8336 15566 8392
rect 15566 8336 15580 8392
rect 15516 8332 15580 8336
rect 21956 8332 22020 8396
rect 24900 8196 24964 8260
rect 10285 8188 10349 8192
rect 10285 8132 10289 8188
rect 10289 8132 10345 8188
rect 10345 8132 10349 8188
rect 10285 8128 10349 8132
rect 10365 8188 10429 8192
rect 10365 8132 10369 8188
rect 10369 8132 10425 8188
rect 10425 8132 10429 8188
rect 10365 8128 10429 8132
rect 10445 8188 10509 8192
rect 10445 8132 10449 8188
rect 10449 8132 10505 8188
rect 10505 8132 10509 8188
rect 10445 8128 10509 8132
rect 10525 8188 10589 8192
rect 10525 8132 10529 8188
rect 10529 8132 10585 8188
rect 10585 8132 10589 8188
rect 10525 8128 10589 8132
rect 19618 8188 19682 8192
rect 19618 8132 19622 8188
rect 19622 8132 19678 8188
rect 19678 8132 19682 8188
rect 19618 8128 19682 8132
rect 19698 8188 19762 8192
rect 19698 8132 19702 8188
rect 19702 8132 19758 8188
rect 19758 8132 19762 8188
rect 19698 8128 19762 8132
rect 19778 8188 19842 8192
rect 19778 8132 19782 8188
rect 19782 8132 19838 8188
rect 19838 8132 19842 8188
rect 19778 8128 19842 8132
rect 19858 8188 19922 8192
rect 19858 8132 19862 8188
rect 19862 8132 19918 8188
rect 19918 8132 19922 8188
rect 19858 8128 19922 8132
rect 9996 8060 10060 8124
rect 22876 8060 22940 8124
rect 5618 7644 5682 7648
rect 5618 7588 5622 7644
rect 5622 7588 5678 7644
rect 5678 7588 5682 7644
rect 5618 7584 5682 7588
rect 5698 7644 5762 7648
rect 5698 7588 5702 7644
rect 5702 7588 5758 7644
rect 5758 7588 5762 7644
rect 5698 7584 5762 7588
rect 5778 7644 5842 7648
rect 5778 7588 5782 7644
rect 5782 7588 5838 7644
rect 5838 7588 5842 7644
rect 5778 7584 5842 7588
rect 5858 7644 5922 7648
rect 5858 7588 5862 7644
rect 5862 7588 5918 7644
rect 5918 7588 5922 7644
rect 5858 7584 5922 7588
rect 14952 7644 15016 7648
rect 14952 7588 14956 7644
rect 14956 7588 15012 7644
rect 15012 7588 15016 7644
rect 14952 7584 15016 7588
rect 15032 7644 15096 7648
rect 15032 7588 15036 7644
rect 15036 7588 15092 7644
rect 15092 7588 15096 7644
rect 15032 7584 15096 7588
rect 15112 7644 15176 7648
rect 15112 7588 15116 7644
rect 15116 7588 15172 7644
rect 15172 7588 15176 7644
rect 15112 7584 15176 7588
rect 15192 7644 15256 7648
rect 15192 7588 15196 7644
rect 15196 7588 15252 7644
rect 15252 7588 15256 7644
rect 15192 7584 15256 7588
rect 2820 7516 2884 7580
rect 19380 7788 19444 7852
rect 17724 7652 17788 7716
rect 24285 7644 24349 7648
rect 24285 7588 24289 7644
rect 24289 7588 24345 7644
rect 24345 7588 24349 7644
rect 24285 7584 24349 7588
rect 24365 7644 24429 7648
rect 24365 7588 24369 7644
rect 24369 7588 24425 7644
rect 24425 7588 24429 7644
rect 24365 7584 24429 7588
rect 24445 7644 24509 7648
rect 24445 7588 24449 7644
rect 24449 7588 24505 7644
rect 24505 7588 24509 7644
rect 24445 7584 24509 7588
rect 24525 7644 24589 7648
rect 24525 7588 24529 7644
rect 24529 7588 24585 7644
rect 24585 7588 24589 7644
rect 24525 7584 24589 7588
rect 25820 7576 25884 7580
rect 25820 7520 25834 7576
rect 25834 7520 25884 7576
rect 25820 7516 25884 7520
rect 5396 7108 5460 7172
rect 10285 7100 10349 7104
rect 10285 7044 10289 7100
rect 10289 7044 10345 7100
rect 10345 7044 10349 7100
rect 10285 7040 10349 7044
rect 10365 7100 10429 7104
rect 10365 7044 10369 7100
rect 10369 7044 10425 7100
rect 10425 7044 10429 7100
rect 10365 7040 10429 7044
rect 10445 7100 10509 7104
rect 10445 7044 10449 7100
rect 10449 7044 10505 7100
rect 10505 7044 10509 7100
rect 10445 7040 10509 7044
rect 10525 7100 10589 7104
rect 10525 7044 10529 7100
rect 10529 7044 10585 7100
rect 10585 7044 10589 7100
rect 10525 7040 10589 7044
rect 19618 7100 19682 7104
rect 19618 7044 19622 7100
rect 19622 7044 19678 7100
rect 19678 7044 19682 7100
rect 19618 7040 19682 7044
rect 19698 7100 19762 7104
rect 19698 7044 19702 7100
rect 19702 7044 19758 7100
rect 19758 7044 19762 7100
rect 19698 7040 19762 7044
rect 19778 7100 19842 7104
rect 19778 7044 19782 7100
rect 19782 7044 19838 7100
rect 19838 7044 19842 7100
rect 19778 7040 19842 7044
rect 19858 7100 19922 7104
rect 19858 7044 19862 7100
rect 19862 7044 19918 7100
rect 19918 7044 19922 7100
rect 19858 7040 19922 7044
rect 10732 6564 10796 6628
rect 5618 6556 5682 6560
rect 5618 6500 5622 6556
rect 5622 6500 5678 6556
rect 5678 6500 5682 6556
rect 5618 6496 5682 6500
rect 5698 6556 5762 6560
rect 5698 6500 5702 6556
rect 5702 6500 5758 6556
rect 5758 6500 5762 6556
rect 5698 6496 5762 6500
rect 5778 6556 5842 6560
rect 5778 6500 5782 6556
rect 5782 6500 5838 6556
rect 5838 6500 5842 6556
rect 5778 6496 5842 6500
rect 5858 6556 5922 6560
rect 5858 6500 5862 6556
rect 5862 6500 5918 6556
rect 5918 6500 5922 6556
rect 5858 6496 5922 6500
rect 25268 7108 25332 7172
rect 24900 7032 24964 7036
rect 24900 6976 24950 7032
rect 24950 6976 24964 7032
rect 24900 6972 24964 6976
rect 20300 6760 20364 6764
rect 20300 6704 20350 6760
rect 20350 6704 20364 6760
rect 20300 6700 20364 6704
rect 20668 6760 20732 6764
rect 20668 6704 20682 6760
rect 20682 6704 20732 6760
rect 20668 6700 20732 6704
rect 21956 6564 22020 6628
rect 14952 6556 15016 6560
rect 14952 6500 14956 6556
rect 14956 6500 15012 6556
rect 15012 6500 15016 6556
rect 14952 6496 15016 6500
rect 15032 6556 15096 6560
rect 15032 6500 15036 6556
rect 15036 6500 15092 6556
rect 15092 6500 15096 6556
rect 15032 6496 15096 6500
rect 15112 6556 15176 6560
rect 15112 6500 15116 6556
rect 15116 6500 15172 6556
rect 15172 6500 15176 6556
rect 15112 6496 15176 6500
rect 15192 6556 15256 6560
rect 15192 6500 15196 6556
rect 15196 6500 15252 6556
rect 15252 6500 15256 6556
rect 15192 6496 15256 6500
rect 24285 6556 24349 6560
rect 24285 6500 24289 6556
rect 24289 6500 24345 6556
rect 24345 6500 24349 6556
rect 24285 6496 24349 6500
rect 24365 6556 24429 6560
rect 24365 6500 24369 6556
rect 24369 6500 24425 6556
rect 24425 6500 24429 6556
rect 24365 6496 24429 6500
rect 24445 6556 24509 6560
rect 24445 6500 24449 6556
rect 24449 6500 24505 6556
rect 24505 6500 24509 6556
rect 24445 6496 24509 6500
rect 24525 6556 24589 6560
rect 24525 6500 24529 6556
rect 24529 6500 24585 6556
rect 24585 6500 24589 6556
rect 24525 6496 24589 6500
rect 9996 6156 10060 6220
rect 20668 6428 20732 6492
rect 21588 6488 21652 6492
rect 21588 6432 21602 6488
rect 21602 6432 21652 6488
rect 21588 6428 21652 6432
rect 22876 6020 22940 6084
rect 10285 6012 10349 6016
rect 10285 5956 10289 6012
rect 10289 5956 10345 6012
rect 10345 5956 10349 6012
rect 10285 5952 10349 5956
rect 10365 6012 10429 6016
rect 10365 5956 10369 6012
rect 10369 5956 10425 6012
rect 10425 5956 10429 6012
rect 10365 5952 10429 5956
rect 10445 6012 10509 6016
rect 10445 5956 10449 6012
rect 10449 5956 10505 6012
rect 10505 5956 10509 6012
rect 10445 5952 10509 5956
rect 10525 6012 10589 6016
rect 10525 5956 10529 6012
rect 10529 5956 10585 6012
rect 10585 5956 10589 6012
rect 10525 5952 10589 5956
rect 19618 6012 19682 6016
rect 19618 5956 19622 6012
rect 19622 5956 19678 6012
rect 19678 5956 19682 6012
rect 19618 5952 19682 5956
rect 19698 6012 19762 6016
rect 19698 5956 19702 6012
rect 19702 5956 19758 6012
rect 19758 5956 19762 6012
rect 19698 5952 19762 5956
rect 19778 6012 19842 6016
rect 19778 5956 19782 6012
rect 19782 5956 19838 6012
rect 19838 5956 19842 6012
rect 19778 5952 19842 5956
rect 19858 6012 19922 6016
rect 19858 5956 19862 6012
rect 19862 5956 19918 6012
rect 19918 5956 19922 6012
rect 19858 5952 19922 5956
rect 4108 5672 4172 5676
rect 4108 5616 4122 5672
rect 4122 5616 4172 5672
rect 4108 5612 4172 5616
rect 5618 5468 5682 5472
rect 5618 5412 5622 5468
rect 5622 5412 5678 5468
rect 5678 5412 5682 5468
rect 5618 5408 5682 5412
rect 5698 5468 5762 5472
rect 5698 5412 5702 5468
rect 5702 5412 5758 5468
rect 5758 5412 5762 5468
rect 5698 5408 5762 5412
rect 5778 5468 5842 5472
rect 5778 5412 5782 5468
rect 5782 5412 5838 5468
rect 5838 5412 5842 5468
rect 5778 5408 5842 5412
rect 5858 5468 5922 5472
rect 5858 5412 5862 5468
rect 5862 5412 5918 5468
rect 5918 5412 5922 5468
rect 5858 5408 5922 5412
rect 12388 5340 12452 5404
rect 14952 5468 15016 5472
rect 14952 5412 14956 5468
rect 14956 5412 15012 5468
rect 15012 5412 15016 5468
rect 14952 5408 15016 5412
rect 15032 5468 15096 5472
rect 15032 5412 15036 5468
rect 15036 5412 15092 5468
rect 15092 5412 15096 5468
rect 15032 5408 15096 5412
rect 15112 5468 15176 5472
rect 15112 5412 15116 5468
rect 15116 5412 15172 5468
rect 15172 5412 15176 5468
rect 15112 5408 15176 5412
rect 15192 5468 15256 5472
rect 15192 5412 15196 5468
rect 15196 5412 15252 5468
rect 15252 5412 15256 5468
rect 15192 5408 15256 5412
rect 23612 5476 23676 5540
rect 24285 5468 24349 5472
rect 24285 5412 24289 5468
rect 24289 5412 24345 5468
rect 24345 5412 24349 5468
rect 24285 5408 24349 5412
rect 24365 5468 24429 5472
rect 24365 5412 24369 5468
rect 24369 5412 24425 5468
rect 24425 5412 24429 5468
rect 24365 5408 24429 5412
rect 24445 5468 24509 5472
rect 24445 5412 24449 5468
rect 24449 5412 24505 5468
rect 24505 5412 24509 5468
rect 24445 5408 24509 5412
rect 24525 5468 24589 5472
rect 24525 5412 24529 5468
rect 24529 5412 24585 5468
rect 24585 5412 24589 5468
rect 24525 5408 24589 5412
rect 2084 5068 2148 5132
rect 8156 5128 8220 5132
rect 8156 5072 8170 5128
rect 8170 5072 8220 5128
rect 8156 5068 8220 5072
rect 10285 4924 10349 4928
rect 10285 4868 10289 4924
rect 10289 4868 10345 4924
rect 10345 4868 10349 4924
rect 10285 4864 10349 4868
rect 10365 4924 10429 4928
rect 10365 4868 10369 4924
rect 10369 4868 10425 4924
rect 10425 4868 10429 4924
rect 10365 4864 10429 4868
rect 10445 4924 10509 4928
rect 10445 4868 10449 4924
rect 10449 4868 10505 4924
rect 10505 4868 10509 4924
rect 10445 4864 10509 4868
rect 10525 4924 10589 4928
rect 10525 4868 10529 4924
rect 10529 4868 10585 4924
rect 10585 4868 10589 4924
rect 10525 4864 10589 4868
rect 19618 4924 19682 4928
rect 19618 4868 19622 4924
rect 19622 4868 19678 4924
rect 19678 4868 19682 4924
rect 19618 4864 19682 4868
rect 19698 4924 19762 4928
rect 19698 4868 19702 4924
rect 19702 4868 19758 4924
rect 19758 4868 19762 4924
rect 19698 4864 19762 4868
rect 19778 4924 19842 4928
rect 19778 4868 19782 4924
rect 19782 4868 19838 4924
rect 19838 4868 19842 4924
rect 19778 4864 19842 4868
rect 19858 4924 19922 4928
rect 19858 4868 19862 4924
rect 19862 4868 19918 4924
rect 19918 4868 19922 4924
rect 19858 4864 19922 4868
rect 9628 4796 9692 4860
rect 12388 4796 12452 4860
rect 6684 4720 6748 4724
rect 6684 4664 6698 4720
rect 6698 4664 6748 4720
rect 6684 4660 6748 4664
rect 9260 4660 9324 4724
rect 23796 4660 23860 4724
rect 5618 4380 5682 4384
rect 5618 4324 5622 4380
rect 5622 4324 5678 4380
rect 5678 4324 5682 4380
rect 5618 4320 5682 4324
rect 5698 4380 5762 4384
rect 5698 4324 5702 4380
rect 5702 4324 5758 4380
rect 5758 4324 5762 4380
rect 5698 4320 5762 4324
rect 5778 4380 5842 4384
rect 5778 4324 5782 4380
rect 5782 4324 5838 4380
rect 5838 4324 5842 4380
rect 5778 4320 5842 4324
rect 5858 4380 5922 4384
rect 5858 4324 5862 4380
rect 5862 4324 5918 4380
rect 5918 4324 5922 4380
rect 5858 4320 5922 4324
rect 14952 4380 15016 4384
rect 14952 4324 14956 4380
rect 14956 4324 15012 4380
rect 15012 4324 15016 4380
rect 14952 4320 15016 4324
rect 15032 4380 15096 4384
rect 15032 4324 15036 4380
rect 15036 4324 15092 4380
rect 15092 4324 15096 4380
rect 15032 4320 15096 4324
rect 15112 4380 15176 4384
rect 15112 4324 15116 4380
rect 15116 4324 15172 4380
rect 15172 4324 15176 4380
rect 15112 4320 15176 4324
rect 15192 4380 15256 4384
rect 15192 4324 15196 4380
rect 15196 4324 15252 4380
rect 15252 4324 15256 4380
rect 15192 4320 15256 4324
rect 24285 4380 24349 4384
rect 24285 4324 24289 4380
rect 24289 4324 24345 4380
rect 24345 4324 24349 4380
rect 24285 4320 24349 4324
rect 24365 4380 24429 4384
rect 24365 4324 24369 4380
rect 24369 4324 24425 4380
rect 24425 4324 24429 4380
rect 24365 4320 24429 4324
rect 24445 4380 24509 4384
rect 24445 4324 24449 4380
rect 24449 4324 24505 4380
rect 24505 4324 24509 4380
rect 24445 4320 24509 4324
rect 24525 4380 24589 4384
rect 24525 4324 24529 4380
rect 24529 4324 24585 4380
rect 24585 4324 24589 4380
rect 24525 4320 24589 4324
rect 20668 4252 20732 4316
rect 24716 3980 24780 4044
rect 16436 3844 16500 3908
rect 10285 3836 10349 3840
rect 10285 3780 10289 3836
rect 10289 3780 10345 3836
rect 10345 3780 10349 3836
rect 10285 3776 10349 3780
rect 10365 3836 10429 3840
rect 10365 3780 10369 3836
rect 10369 3780 10425 3836
rect 10425 3780 10429 3836
rect 10365 3776 10429 3780
rect 10445 3836 10509 3840
rect 10445 3780 10449 3836
rect 10449 3780 10505 3836
rect 10505 3780 10509 3836
rect 10445 3776 10509 3780
rect 10525 3836 10589 3840
rect 10525 3780 10529 3836
rect 10529 3780 10585 3836
rect 10585 3780 10589 3836
rect 10525 3776 10589 3780
rect 19618 3836 19682 3840
rect 19618 3780 19622 3836
rect 19622 3780 19678 3836
rect 19678 3780 19682 3836
rect 19618 3776 19682 3780
rect 19698 3836 19762 3840
rect 19698 3780 19702 3836
rect 19702 3780 19758 3836
rect 19758 3780 19762 3836
rect 19698 3776 19762 3780
rect 19778 3836 19842 3840
rect 19778 3780 19782 3836
rect 19782 3780 19838 3836
rect 19838 3780 19842 3836
rect 19778 3776 19842 3780
rect 19858 3836 19922 3840
rect 19858 3780 19862 3836
rect 19862 3780 19918 3836
rect 19918 3780 19922 3836
rect 19858 3776 19922 3780
rect 4660 3572 4724 3636
rect 21036 3768 21100 3772
rect 21036 3712 21050 3768
rect 21050 3712 21100 3768
rect 6684 3436 6748 3500
rect 6316 3300 6380 3364
rect 11836 3572 11900 3636
rect 21036 3708 21100 3712
rect 23612 3360 23676 3364
rect 23612 3304 23662 3360
rect 23662 3304 23676 3360
rect 23612 3300 23676 3304
rect 5618 3292 5682 3296
rect 5618 3236 5622 3292
rect 5622 3236 5678 3292
rect 5678 3236 5682 3292
rect 5618 3232 5682 3236
rect 5698 3292 5762 3296
rect 5698 3236 5702 3292
rect 5702 3236 5758 3292
rect 5758 3236 5762 3292
rect 5698 3232 5762 3236
rect 5778 3292 5842 3296
rect 5778 3236 5782 3292
rect 5782 3236 5838 3292
rect 5838 3236 5842 3292
rect 5778 3232 5842 3236
rect 5858 3292 5922 3296
rect 5858 3236 5862 3292
rect 5862 3236 5918 3292
rect 5918 3236 5922 3292
rect 5858 3232 5922 3236
rect 14952 3292 15016 3296
rect 14952 3236 14956 3292
rect 14956 3236 15012 3292
rect 15012 3236 15016 3292
rect 14952 3232 15016 3236
rect 15032 3292 15096 3296
rect 15032 3236 15036 3292
rect 15036 3236 15092 3292
rect 15092 3236 15096 3292
rect 15032 3232 15096 3236
rect 15112 3292 15176 3296
rect 15112 3236 15116 3292
rect 15116 3236 15172 3292
rect 15172 3236 15176 3292
rect 15112 3232 15176 3236
rect 15192 3292 15256 3296
rect 15192 3236 15196 3292
rect 15196 3236 15252 3292
rect 15252 3236 15256 3292
rect 15192 3232 15256 3236
rect 24285 3292 24349 3296
rect 24285 3236 24289 3292
rect 24289 3236 24345 3292
rect 24345 3236 24349 3292
rect 24285 3232 24349 3236
rect 24365 3292 24429 3296
rect 24365 3236 24369 3292
rect 24369 3236 24425 3292
rect 24425 3236 24429 3292
rect 24365 3232 24429 3236
rect 24445 3292 24509 3296
rect 24445 3236 24449 3292
rect 24449 3236 24505 3292
rect 24505 3236 24509 3292
rect 24445 3232 24509 3236
rect 24525 3292 24589 3296
rect 24525 3236 24529 3292
rect 24529 3236 24585 3292
rect 24585 3236 24589 3292
rect 24525 3232 24589 3236
rect 23428 3224 23492 3228
rect 23428 3168 23478 3224
rect 23478 3168 23492 3224
rect 23428 3164 23492 3168
rect 10285 2748 10349 2752
rect 10285 2692 10289 2748
rect 10289 2692 10345 2748
rect 10345 2692 10349 2748
rect 10285 2688 10349 2692
rect 10365 2748 10429 2752
rect 10365 2692 10369 2748
rect 10369 2692 10425 2748
rect 10425 2692 10429 2748
rect 10365 2688 10429 2692
rect 10445 2748 10509 2752
rect 10445 2692 10449 2748
rect 10449 2692 10505 2748
rect 10505 2692 10509 2748
rect 10445 2688 10509 2692
rect 10525 2748 10589 2752
rect 10525 2692 10529 2748
rect 10529 2692 10585 2748
rect 10585 2692 10589 2748
rect 10525 2688 10589 2692
rect 19618 2748 19682 2752
rect 19618 2692 19622 2748
rect 19622 2692 19678 2748
rect 19678 2692 19682 2748
rect 19618 2688 19682 2692
rect 19698 2748 19762 2752
rect 19698 2692 19702 2748
rect 19702 2692 19758 2748
rect 19758 2692 19762 2748
rect 19698 2688 19762 2692
rect 19778 2748 19842 2752
rect 19778 2692 19782 2748
rect 19782 2692 19838 2748
rect 19838 2692 19842 2748
rect 19778 2688 19842 2692
rect 19858 2748 19922 2752
rect 19858 2692 19862 2748
rect 19862 2692 19918 2748
rect 19918 2692 19922 2748
rect 19858 2688 19922 2692
rect 12388 2620 12452 2684
rect 16804 2484 16868 2548
rect 5618 2204 5682 2208
rect 5618 2148 5622 2204
rect 5622 2148 5678 2204
rect 5678 2148 5682 2204
rect 5618 2144 5682 2148
rect 5698 2204 5762 2208
rect 5698 2148 5702 2204
rect 5702 2148 5758 2204
rect 5758 2148 5762 2204
rect 5698 2144 5762 2148
rect 5778 2204 5842 2208
rect 5778 2148 5782 2204
rect 5782 2148 5838 2204
rect 5838 2148 5842 2204
rect 5778 2144 5842 2148
rect 5858 2204 5922 2208
rect 5858 2148 5862 2204
rect 5862 2148 5918 2204
rect 5918 2148 5922 2204
rect 5858 2144 5922 2148
rect 14952 2204 15016 2208
rect 14952 2148 14956 2204
rect 14956 2148 15012 2204
rect 15012 2148 15016 2204
rect 14952 2144 15016 2148
rect 15032 2204 15096 2208
rect 15032 2148 15036 2204
rect 15036 2148 15092 2204
rect 15092 2148 15096 2204
rect 15032 2144 15096 2148
rect 15112 2204 15176 2208
rect 15112 2148 15116 2204
rect 15116 2148 15172 2204
rect 15172 2148 15176 2204
rect 15112 2144 15176 2148
rect 15192 2204 15256 2208
rect 15192 2148 15196 2204
rect 15196 2148 15252 2204
rect 15252 2148 15256 2204
rect 15192 2144 15256 2148
rect 24285 2204 24349 2208
rect 24285 2148 24289 2204
rect 24289 2148 24345 2204
rect 24345 2148 24349 2204
rect 24285 2144 24349 2148
rect 24365 2204 24429 2208
rect 24365 2148 24369 2204
rect 24369 2148 24425 2204
rect 24425 2148 24429 2204
rect 24365 2144 24429 2148
rect 24445 2204 24509 2208
rect 24445 2148 24449 2204
rect 24449 2148 24505 2204
rect 24505 2148 24509 2204
rect 24445 2144 24509 2148
rect 24525 2204 24589 2208
rect 24525 2148 24529 2204
rect 24529 2148 24585 2204
rect 24585 2148 24589 2204
rect 24525 2144 24589 2148
rect 12388 1804 12452 1868
rect 15516 1804 15580 1868
rect 2084 1668 2148 1732
<< metal4 >>
rect 2819 26076 2885 26077
rect 2819 26012 2820 26076
rect 2884 26012 2885 26076
rect 2819 26011 2885 26012
rect 2635 24716 2701 24717
rect 2635 24652 2636 24716
rect 2700 24652 2701 24716
rect 2635 24651 2701 24652
rect 2083 20908 2149 20909
rect 2083 20844 2084 20908
rect 2148 20844 2149 20908
rect 2083 20843 2149 20844
rect 1718 10301 1778 17902
rect 2086 13021 2146 20843
rect 2270 19277 2330 21982
rect 2638 21589 2698 24651
rect 2635 21588 2701 21589
rect 2635 21524 2636 21588
rect 2700 21524 2701 21588
rect 2635 21523 2701 21524
rect 2267 19276 2333 19277
rect 2267 19212 2268 19276
rect 2332 19212 2333 19276
rect 2267 19211 2333 19212
rect 2083 13020 2149 13021
rect 2083 12956 2084 13020
rect 2148 12956 2149 13020
rect 2083 12955 2149 12956
rect 1715 10300 1781 10301
rect 1715 10236 1716 10300
rect 1780 10236 1781 10300
rect 1715 10235 1781 10236
rect 2454 8941 2514 9742
rect 2451 8940 2517 8941
rect 2451 8876 2452 8940
rect 2516 8876 2517 8940
rect 2451 8875 2517 8876
rect 2822 7581 2882 26011
rect 25819 25668 25885 25669
rect 5610 25056 5931 25616
rect 5610 24992 5618 25056
rect 5682 24992 5698 25056
rect 5762 24992 5778 25056
rect 5842 24992 5858 25056
rect 5922 24992 5931 25056
rect 3187 24852 3253 24853
rect 3187 24788 3188 24852
rect 3252 24788 3253 24852
rect 3187 24787 3253 24788
rect 3739 24852 3805 24853
rect 3739 24788 3740 24852
rect 3804 24788 3805 24852
rect 3739 24787 3805 24788
rect 3190 12205 3250 24787
rect 3187 12204 3253 12205
rect 3187 12140 3188 12204
rect 3252 12140 3253 12204
rect 3187 12139 3253 12140
rect 3742 12069 3802 24787
rect 5610 23968 5931 24992
rect 5610 23904 5618 23968
rect 5682 23904 5698 23968
rect 5762 23904 5778 23968
rect 5842 23904 5858 23968
rect 5922 23904 5931 23968
rect 5610 22880 5931 23904
rect 10277 25600 10597 25616
rect 10277 25536 10285 25600
rect 10349 25536 10365 25600
rect 10429 25536 10445 25600
rect 10509 25536 10525 25600
rect 10589 25536 10597 25600
rect 10277 24512 10597 25536
rect 10915 25260 10981 25261
rect 10915 25196 10916 25260
rect 10980 25196 10981 25260
rect 10915 25195 10981 25196
rect 10277 24448 10285 24512
rect 10349 24448 10365 24512
rect 10429 24448 10445 24512
rect 10509 24448 10525 24512
rect 10589 24448 10597 24512
rect 10277 23424 10597 24448
rect 10277 23360 10285 23424
rect 10349 23360 10365 23424
rect 10429 23360 10445 23424
rect 10509 23360 10525 23424
rect 10589 23360 10597 23424
rect 5610 22816 5618 22880
rect 5682 22816 5698 22880
rect 5762 22816 5778 22880
rect 5842 22816 5858 22880
rect 5922 22816 5931 22880
rect 5610 21792 5931 22816
rect 5610 21728 5618 21792
rect 5682 21728 5698 21792
rect 5762 21728 5778 21792
rect 5842 21728 5858 21792
rect 5922 21728 5931 21792
rect 5610 20704 5931 21728
rect 5610 20640 5618 20704
rect 5682 20640 5698 20704
rect 5762 20640 5778 20704
rect 5842 20640 5858 20704
rect 5922 20640 5931 20704
rect 5610 19616 5931 20640
rect 5610 19552 5618 19616
rect 5682 19552 5698 19616
rect 5762 19552 5778 19616
rect 5842 19552 5858 19616
rect 5922 19552 5931 19616
rect 5610 18528 5931 19552
rect 5610 18464 5618 18528
rect 5682 18464 5698 18528
rect 5762 18464 5778 18528
rect 5842 18464 5858 18528
rect 5922 18464 5931 18528
rect 5610 17440 5931 18464
rect 5610 17376 5618 17440
rect 5682 17376 5698 17440
rect 5762 17376 5778 17440
rect 5842 17376 5858 17440
rect 5922 17376 5931 17440
rect 5610 16352 5931 17376
rect 6131 17172 6132 17222
rect 6196 17172 6197 17222
rect 6131 17171 6197 17172
rect 5610 16288 5618 16352
rect 5682 16288 5698 16352
rect 5762 16288 5778 16352
rect 5842 16288 5858 16352
rect 5922 16288 5931 16352
rect 5610 15264 5931 16288
rect 6131 15740 6197 15741
rect 6131 15676 6132 15740
rect 6196 15676 6197 15740
rect 6131 15675 6197 15676
rect 6134 15418 6194 15675
rect 5610 15200 5618 15264
rect 5682 15200 5698 15264
rect 5762 15200 5778 15264
rect 5842 15200 5858 15264
rect 5922 15200 5931 15264
rect 5610 14176 5931 15200
rect 6315 14788 6381 14789
rect 6315 14724 6316 14788
rect 6380 14724 6381 14788
rect 6315 14723 6381 14724
rect 5610 14112 5618 14176
rect 5682 14112 5698 14176
rect 5762 14112 5778 14176
rect 5842 14112 5858 14176
rect 5922 14112 5931 14176
rect 5211 13700 5277 13701
rect 5211 13636 5212 13700
rect 5276 13636 5277 13700
rect 5211 13635 5277 13636
rect 4843 13020 4909 13021
rect 4843 12956 4844 13020
rect 4908 12956 4909 13020
rect 4843 12955 4909 12956
rect 3739 12068 3805 12069
rect 3739 12004 3740 12068
rect 3804 12004 3805 12068
rect 3739 12003 3805 12004
rect 4846 10573 4906 12955
rect 5214 12018 5274 13635
rect 5610 13088 5931 14112
rect 5610 13024 5618 13088
rect 5682 13024 5698 13088
rect 5762 13024 5778 13088
rect 5842 13024 5858 13088
rect 5922 13024 5931 13088
rect 5610 12000 5931 13024
rect 6131 12884 6197 12885
rect 6131 12820 6132 12884
rect 6196 12820 6197 12884
rect 6131 12819 6197 12820
rect 5610 11936 5618 12000
rect 5682 11936 5698 12000
rect 5762 11936 5778 12000
rect 5842 11936 5858 12000
rect 5922 11936 5931 12000
rect 5214 11253 5274 11782
rect 5211 11252 5277 11253
rect 5211 11188 5212 11252
rect 5276 11188 5277 11252
rect 5211 11187 5277 11188
rect 5610 10912 5931 11936
rect 5610 10848 5618 10912
rect 5682 10848 5698 10912
rect 5762 10848 5778 10912
rect 5842 10848 5858 10912
rect 5922 10848 5931 10912
rect 4843 10572 4909 10573
rect 4843 10508 4844 10572
rect 4908 10508 4909 10572
rect 4843 10507 4909 10508
rect 3003 10028 3069 10029
rect 3003 9964 3004 10028
rect 3068 9964 3069 10028
rect 3003 9963 3069 9964
rect 2819 7580 2885 7581
rect 2819 7516 2820 7580
rect 2884 7516 2885 7580
rect 2819 7515 2885 7516
rect 2086 5133 2146 5662
rect 2083 5132 2149 5133
rect 2083 5068 2084 5132
rect 2148 5068 2149 5132
rect 2083 5067 2149 5068
rect 3006 2498 3066 9963
rect 5610 9824 5931 10848
rect 6134 10165 6194 12819
rect 6131 10164 6197 10165
rect 6131 10100 6132 10164
rect 6196 10100 6197 10164
rect 6131 10099 6197 10100
rect 5610 9760 5618 9824
rect 5682 9760 5698 9824
rect 5762 9760 5778 9824
rect 5842 9760 5858 9824
rect 5922 9760 5931 9824
rect 5398 8805 5458 9062
rect 5395 8804 5461 8805
rect 5395 8740 5396 8804
rect 5460 8740 5461 8804
rect 5395 8739 5461 8740
rect 5610 8736 5931 9760
rect 5610 8672 5618 8736
rect 5682 8672 5698 8736
rect 5762 8672 5778 8736
rect 5842 8672 5858 8736
rect 5922 8672 5931 8736
rect 5610 7648 5931 8672
rect 5610 7584 5618 7648
rect 5682 7584 5698 7648
rect 5762 7584 5778 7648
rect 5842 7584 5858 7648
rect 5922 7584 5931 7648
rect 5610 6560 5931 7584
rect 5610 6496 5618 6560
rect 5682 6496 5698 6560
rect 5762 6496 5778 6560
rect 5842 6496 5858 6560
rect 5922 6496 5931 6560
rect 4107 5676 4173 5677
rect 4107 5612 4108 5676
rect 4172 5612 4173 5676
rect 4107 5611 4173 5612
rect 4110 1138 4170 5611
rect 5610 5472 5931 6496
rect 5610 5408 5618 5472
rect 5682 5408 5698 5472
rect 5762 5408 5778 5472
rect 5842 5408 5858 5472
rect 5922 5408 5931 5472
rect 5610 4384 5931 5408
rect 5610 4320 5618 4384
rect 5682 4320 5698 4384
rect 5762 4320 5778 4384
rect 5842 4320 5858 4384
rect 5922 4320 5931 4384
rect 4659 3572 4660 3622
rect 4724 3572 4725 3622
rect 4659 3571 4725 3572
rect 5610 3296 5931 4320
rect 6318 3365 6378 14723
rect 6502 10709 6562 23342
rect 10277 22336 10597 23360
rect 10277 22272 10285 22336
rect 10349 22272 10365 22336
rect 10429 22272 10445 22336
rect 10509 22272 10525 22336
rect 10589 22272 10597 22336
rect 10277 21248 10597 22272
rect 10277 21184 10285 21248
rect 10349 21184 10365 21248
rect 10429 21184 10445 21248
rect 10509 21184 10525 21248
rect 10589 21184 10597 21248
rect 10277 20160 10597 21184
rect 10918 20229 10978 25195
rect 14944 25056 15264 25616
rect 14944 24992 14952 25056
rect 15016 24992 15032 25056
rect 15096 24992 15112 25056
rect 15176 24992 15192 25056
rect 15256 24992 15264 25056
rect 14227 24852 14293 24853
rect 14227 24788 14228 24852
rect 14292 24788 14293 24852
rect 14227 24787 14293 24788
rect 10915 20228 10981 20229
rect 10915 20164 10916 20228
rect 10980 20164 10981 20228
rect 10915 20163 10981 20164
rect 10277 20096 10285 20160
rect 10349 20096 10365 20160
rect 10429 20096 10445 20160
rect 10509 20096 10525 20160
rect 10589 20096 10597 20160
rect 9075 19548 9141 19549
rect 9075 19498 9076 19548
rect 9140 19498 9141 19548
rect 10277 19072 10597 20096
rect 10731 19684 10797 19685
rect 10731 19620 10732 19684
rect 10796 19620 10797 19684
rect 10731 19619 10797 19620
rect 10277 19008 10285 19072
rect 10349 19008 10365 19072
rect 10429 19008 10445 19072
rect 10509 19008 10525 19072
rect 10589 19008 10597 19072
rect 10277 17984 10597 19008
rect 10277 17920 10285 17984
rect 10349 17920 10365 17984
rect 10429 17920 10445 17984
rect 10509 17920 10525 17984
rect 10589 17920 10597 17984
rect 10277 16896 10597 17920
rect 10277 16832 10285 16896
rect 10349 16832 10365 16896
rect 10429 16832 10445 16896
rect 10509 16832 10525 16896
rect 10589 16832 10597 16896
rect 6683 16420 6749 16421
rect 6683 16356 6684 16420
rect 6748 16356 6749 16420
rect 6683 16355 6749 16356
rect 6499 10708 6565 10709
rect 6499 10644 6500 10708
rect 6564 10644 6565 10708
rect 6499 10643 6565 10644
rect 6499 10436 6565 10437
rect 6499 10372 6500 10436
rect 6564 10372 6565 10436
rect 6499 10371 6565 10372
rect 6502 10029 6562 10371
rect 6499 10028 6565 10029
rect 6499 9964 6500 10028
rect 6564 9964 6565 10028
rect 6499 9963 6565 9964
rect 6686 9757 6746 16355
rect 9630 14653 9690 16542
rect 9995 16284 10061 16285
rect 9995 16220 9996 16284
rect 10060 16220 10061 16284
rect 9995 16219 10061 16220
rect 9627 14652 9693 14653
rect 9627 14588 9628 14652
rect 9692 14588 9693 14652
rect 9627 14587 9693 14588
rect 9630 13565 9690 13822
rect 9811 13700 9877 13701
rect 9811 13636 9812 13700
rect 9876 13636 9877 13700
rect 9811 13635 9877 13636
rect 9627 13564 9693 13565
rect 9627 13500 9628 13564
rect 9692 13500 9693 13564
rect 9627 13499 9693 13500
rect 7603 12340 7669 12341
rect 7603 12276 7604 12340
rect 7668 12276 7669 12340
rect 7603 12275 7669 12276
rect 7606 11933 7666 12275
rect 7235 11932 7301 11933
rect 7235 11868 7236 11932
rect 7300 11868 7301 11932
rect 7235 11867 7301 11868
rect 7603 11932 7669 11933
rect 7603 11868 7604 11932
rect 7668 11868 7669 11932
rect 7603 11867 7669 11868
rect 7238 11338 7298 11867
rect 7235 11052 7236 11102
rect 7300 11052 7301 11102
rect 7235 11051 7301 11052
rect 6683 9756 6749 9757
rect 6683 9692 6684 9756
rect 6748 9692 6749 9756
rect 6683 9691 6749 9692
rect 8158 8261 8218 13142
rect 9259 9620 9325 9621
rect 9259 9556 9260 9620
rect 9324 9556 9325 9620
rect 9259 9555 9325 9556
rect 8155 8260 8221 8261
rect 8155 8196 8156 8260
rect 8220 8196 8221 8260
rect 8155 8195 8221 8196
rect 6686 4725 6746 7702
rect 9262 4725 9322 9555
rect 9814 7170 9874 13635
rect 9998 8125 10058 16219
rect 10277 15808 10597 16832
rect 10277 15744 10285 15808
rect 10349 15744 10365 15808
rect 10429 15744 10445 15808
rect 10509 15744 10525 15808
rect 10589 15744 10597 15808
rect 10277 14720 10597 15744
rect 10277 14656 10285 14720
rect 10349 14656 10365 14720
rect 10429 14656 10445 14720
rect 10509 14656 10525 14720
rect 10589 14656 10597 14720
rect 10277 13632 10597 14656
rect 10277 13568 10285 13632
rect 10349 13568 10365 13632
rect 10429 13568 10445 13632
rect 10509 13568 10525 13632
rect 10589 13568 10597 13632
rect 10277 12544 10597 13568
rect 10277 12480 10285 12544
rect 10349 12480 10365 12544
rect 10429 12480 10445 12544
rect 10509 12480 10525 12544
rect 10589 12480 10597 12544
rect 10277 11456 10597 12480
rect 10277 11392 10285 11456
rect 10349 11392 10365 11456
rect 10429 11392 10445 11456
rect 10509 11392 10525 11456
rect 10589 11392 10597 11456
rect 10277 10368 10597 11392
rect 10277 10304 10285 10368
rect 10349 10304 10365 10368
rect 10429 10304 10445 10368
rect 10509 10304 10525 10368
rect 10589 10304 10597 10368
rect 10277 9280 10597 10304
rect 10277 9216 10285 9280
rect 10349 9216 10365 9280
rect 10429 9216 10445 9280
rect 10509 9216 10525 9280
rect 10589 9216 10597 9280
rect 10277 8192 10597 9216
rect 10277 8128 10285 8192
rect 10349 8128 10365 8192
rect 10429 8128 10445 8192
rect 10509 8128 10525 8192
rect 10589 8128 10597 8192
rect 9995 8124 10061 8125
rect 9995 8060 9996 8124
rect 10060 8060 10061 8124
rect 9995 8059 10061 8060
rect 9814 7110 10058 7170
rect 9630 4861 9690 6342
rect 9998 6221 10058 7110
rect 10277 7104 10597 8128
rect 10277 7040 10285 7104
rect 10349 7040 10365 7104
rect 10429 7040 10445 7104
rect 10509 7040 10525 7104
rect 10589 7040 10597 7104
rect 9995 6220 10061 6221
rect 9995 6156 9996 6220
rect 10060 6156 10061 6220
rect 9995 6155 10061 6156
rect 10277 6016 10597 7040
rect 10734 6629 10794 19619
rect 12939 19140 13005 19141
rect 12939 19076 12940 19140
rect 13004 19076 13005 19140
rect 12939 19075 13005 19076
rect 10915 17916 10981 17917
rect 10915 17852 10916 17916
rect 10980 17852 10981 17916
rect 10915 17851 10981 17852
rect 10918 17373 10978 17851
rect 10915 17372 10981 17373
rect 10915 17308 10916 17372
rect 10980 17308 10981 17372
rect 10915 17307 10981 17308
rect 11099 14108 11165 14109
rect 11099 14058 11100 14108
rect 11164 14058 11165 14108
rect 10915 10572 10981 10573
rect 10915 10508 10916 10572
rect 10980 10570 10981 10572
rect 10980 10510 11198 10570
rect 10980 10508 10981 10510
rect 10915 10507 10981 10508
rect 10915 10300 10981 10301
rect 10915 10236 10916 10300
rect 10980 10236 10981 10300
rect 10915 10235 10981 10236
rect 10731 6628 10797 6629
rect 10731 6564 10732 6628
rect 10796 6564 10797 6628
rect 10731 6563 10797 6564
rect 10277 5952 10285 6016
rect 10349 5952 10365 6016
rect 10429 5952 10445 6016
rect 10509 5952 10525 6016
rect 10589 5952 10597 6016
rect 10277 4928 10597 5952
rect 10918 5898 10978 10235
rect 10277 4864 10285 4928
rect 10349 4864 10365 4928
rect 10429 4864 10445 4928
rect 10509 4864 10525 4928
rect 10589 4864 10597 4928
rect 9627 4860 9693 4861
rect 9627 4796 9628 4860
rect 9692 4796 9693 4860
rect 9627 4795 9693 4796
rect 6683 4724 6749 4725
rect 6683 4660 6684 4724
rect 6748 4660 6749 4724
rect 6683 4659 6749 4660
rect 9259 4724 9325 4725
rect 9259 4660 9260 4724
rect 9324 4660 9325 4724
rect 9259 4659 9325 4660
rect 6686 3501 6746 4302
rect 10277 3840 10597 4864
rect 10277 3776 10285 3840
rect 10349 3776 10365 3840
rect 10429 3776 10445 3840
rect 10509 3776 10525 3840
rect 10589 3776 10597 3840
rect 6683 3500 6749 3501
rect 6683 3436 6684 3500
rect 6748 3436 6749 3500
rect 6683 3435 6749 3436
rect 6315 3364 6381 3365
rect 6315 3300 6316 3364
rect 6380 3300 6381 3364
rect 6315 3299 6381 3300
rect 5610 3232 5618 3296
rect 5682 3232 5698 3296
rect 5762 3232 5778 3296
rect 5842 3232 5858 3296
rect 5922 3232 5931 3296
rect 5610 2208 5931 3232
rect 5610 2144 5618 2208
rect 5682 2144 5698 2208
rect 5762 2144 5778 2208
rect 5842 2144 5858 2208
rect 5922 2144 5931 2208
rect 5610 2128 5931 2144
rect 10277 2752 10597 3776
rect 11838 3637 11898 17222
rect 12942 12613 13002 19075
rect 14230 18818 14290 24787
rect 14944 23968 15264 24992
rect 14944 23904 14952 23968
rect 15016 23904 15032 23968
rect 15096 23904 15112 23968
rect 15176 23904 15192 23968
rect 15256 23904 15264 23968
rect 14944 22880 15264 23904
rect 19610 25600 19930 25616
rect 19610 25536 19618 25600
rect 19682 25536 19698 25600
rect 19762 25536 19778 25600
rect 19842 25536 19858 25600
rect 19922 25536 19930 25600
rect 19610 24512 19930 25536
rect 23979 25396 24045 25397
rect 23979 25332 23980 25396
rect 24044 25332 24045 25396
rect 23979 25331 24045 25332
rect 21219 25260 21285 25261
rect 21219 25196 21220 25260
rect 21284 25196 21285 25260
rect 21219 25195 21285 25196
rect 19610 24448 19618 24512
rect 19682 24448 19698 24512
rect 19762 24448 19778 24512
rect 19842 24448 19858 24512
rect 19922 24448 19930 24512
rect 19610 23424 19930 24448
rect 20115 24444 20181 24445
rect 20115 24380 20116 24444
rect 20180 24380 20181 24444
rect 20115 24379 20181 24380
rect 19610 23360 19618 23424
rect 19682 23360 19698 23424
rect 19762 23360 19778 23424
rect 19842 23360 19858 23424
rect 19922 23360 19930 23424
rect 14944 22816 14952 22880
rect 15016 22816 15032 22880
rect 15096 22816 15112 22880
rect 15176 22816 15192 22880
rect 15256 22816 15264 22880
rect 14944 21792 15264 22816
rect 17723 22540 17789 22541
rect 17723 22476 17724 22540
rect 17788 22476 17789 22540
rect 17723 22475 17789 22476
rect 14944 21728 14952 21792
rect 15016 21728 15032 21792
rect 15096 21728 15112 21792
rect 15176 21728 15192 21792
rect 15256 21728 15264 21792
rect 14944 20704 15264 21728
rect 14944 20640 14952 20704
rect 15016 20640 15032 20704
rect 15096 20640 15112 20704
rect 15176 20640 15192 20704
rect 15256 20640 15264 20704
rect 14779 20364 14845 20365
rect 14779 20300 14780 20364
rect 14844 20300 14845 20364
rect 14779 20299 14845 20300
rect 14782 19549 14842 20299
rect 14944 19616 15264 20640
rect 17726 20093 17786 22475
rect 19610 22336 19930 23360
rect 19610 22272 19618 22336
rect 19682 22272 19698 22336
rect 19762 22272 19778 22336
rect 19842 22272 19858 22336
rect 19922 22272 19930 22336
rect 19610 21248 19930 22272
rect 19610 21184 19618 21248
rect 19682 21184 19698 21248
rect 19762 21184 19778 21248
rect 19842 21184 19858 21248
rect 19922 21184 19930 21248
rect 19610 20160 19930 21184
rect 19610 20096 19618 20160
rect 19682 20096 19698 20160
rect 19762 20096 19778 20160
rect 19842 20096 19858 20160
rect 19922 20096 19930 20160
rect 17723 20092 17789 20093
rect 17723 20028 17724 20092
rect 17788 20028 17789 20092
rect 17723 20027 17789 20028
rect 14944 19552 14952 19616
rect 15016 19552 15032 19616
rect 15096 19552 15112 19616
rect 15176 19552 15192 19616
rect 15256 19552 15264 19616
rect 14779 19548 14845 19549
rect 14779 19484 14780 19548
rect 14844 19484 14845 19548
rect 14779 19483 14845 19484
rect 13859 15132 13860 15182
rect 13924 15132 13925 15182
rect 13859 15131 13925 15132
rect 14230 14245 14290 18582
rect 14944 18528 15264 19552
rect 19379 19140 19445 19141
rect 19379 19076 19380 19140
rect 19444 19076 19445 19140
rect 19379 19075 19445 19076
rect 14944 18464 14952 18528
rect 15016 18464 15032 18528
rect 15096 18464 15112 18528
rect 15176 18464 15192 18528
rect 15256 18464 15264 18528
rect 14944 17440 15264 18464
rect 14944 17376 14952 17440
rect 15016 17376 15032 17440
rect 15096 17376 15112 17440
rect 15176 17376 15192 17440
rect 15256 17376 15264 17440
rect 14944 16352 15264 17376
rect 14944 16288 14952 16352
rect 15016 16288 15032 16352
rect 15096 16288 15112 16352
rect 15176 16288 15192 16352
rect 15256 16288 15264 16352
rect 14595 16284 14661 16285
rect 14595 16220 14596 16284
rect 14660 16220 14661 16284
rect 14595 16219 14661 16220
rect 14598 15418 14658 16219
rect 14944 15264 15264 16288
rect 14944 15200 14952 15264
rect 15016 15200 15032 15264
rect 15096 15200 15112 15264
rect 15176 15200 15192 15264
rect 15256 15200 15264 15264
rect 14227 14244 14293 14245
rect 14227 14180 14228 14244
rect 14292 14180 14293 14244
rect 14227 14179 14293 14180
rect 14944 14176 15264 15200
rect 14944 14112 14952 14176
rect 15016 14112 15032 14176
rect 15096 14112 15112 14176
rect 15176 14112 15192 14176
rect 15256 14112 15264 14176
rect 14944 13088 15264 14112
rect 14944 13024 14952 13088
rect 15016 13024 15032 13088
rect 15096 13024 15112 13088
rect 15176 13024 15192 13088
rect 15256 13024 15264 13088
rect 12939 12612 13005 12613
rect 12939 12548 12940 12612
rect 13004 12548 13005 12612
rect 12939 12547 13005 12548
rect 14944 12000 15264 13024
rect 19382 13021 19442 19075
rect 19610 19072 19930 20096
rect 20118 19821 20178 24379
rect 20667 23492 20733 23493
rect 20667 23428 20668 23492
rect 20732 23428 20733 23492
rect 20667 23427 20733 23428
rect 20115 19820 20181 19821
rect 20115 19756 20116 19820
rect 20180 19756 20181 19820
rect 20115 19755 20181 19756
rect 20299 19140 20365 19141
rect 20299 19076 20300 19140
rect 20364 19076 20365 19140
rect 20299 19075 20365 19076
rect 19610 19008 19618 19072
rect 19682 19008 19698 19072
rect 19762 19008 19778 19072
rect 19842 19008 19858 19072
rect 19922 19008 19930 19072
rect 19610 17984 19930 19008
rect 20302 18818 20362 19075
rect 20299 18052 20365 18053
rect 20299 17988 20300 18052
rect 20364 17988 20365 18052
rect 20299 17987 20365 17988
rect 19610 17920 19618 17984
rect 19682 17920 19698 17984
rect 19762 17920 19778 17984
rect 19842 17920 19858 17984
rect 19922 17920 19930 17984
rect 19610 16896 19930 17920
rect 20115 17780 20181 17781
rect 20115 17716 20116 17780
rect 20180 17716 20181 17780
rect 20115 17715 20181 17716
rect 20118 17101 20178 17715
rect 20115 17100 20181 17101
rect 20115 17036 20116 17100
rect 20180 17036 20181 17100
rect 20115 17035 20181 17036
rect 19610 16832 19618 16896
rect 19682 16832 19698 16896
rect 19762 16832 19778 16896
rect 19842 16832 19858 16896
rect 19922 16832 19930 16896
rect 19610 15808 19930 16832
rect 19610 15744 19618 15808
rect 19682 15744 19698 15808
rect 19762 15744 19778 15808
rect 19842 15744 19858 15808
rect 19922 15744 19930 15808
rect 19610 14720 19930 15744
rect 20302 15061 20362 17987
rect 20670 17458 20730 23427
rect 21035 21860 21101 21861
rect 21035 21796 21036 21860
rect 21100 21796 21101 21860
rect 21035 21795 21101 21796
rect 21038 18053 21098 21795
rect 21035 18052 21101 18053
rect 21035 17988 21036 18052
rect 21100 17988 21101 18052
rect 21035 17987 21101 17988
rect 20483 17100 20549 17101
rect 20483 17036 20484 17100
rect 20548 17036 20549 17100
rect 20483 17035 20549 17036
rect 20299 15060 20365 15061
rect 20299 14996 20300 15060
rect 20364 14996 20365 15060
rect 20299 14995 20365 14996
rect 20486 14925 20546 17035
rect 20670 16965 20730 17222
rect 20667 16964 20733 16965
rect 20667 16900 20668 16964
rect 20732 16900 20733 16964
rect 20667 16899 20733 16900
rect 20854 15877 20914 16542
rect 21035 16012 21101 16013
rect 21035 15948 21036 16012
rect 21100 15948 21101 16012
rect 21035 15947 21101 15948
rect 20851 15876 20917 15877
rect 20851 15812 20852 15876
rect 20916 15812 20917 15876
rect 20851 15811 20917 15812
rect 20483 14924 20549 14925
rect 20483 14860 20484 14924
rect 20548 14860 20549 14924
rect 20483 14859 20549 14860
rect 19610 14656 19618 14720
rect 19682 14656 19698 14720
rect 19762 14656 19778 14720
rect 19842 14656 19858 14720
rect 19922 14656 19930 14720
rect 19610 13632 19930 14656
rect 20854 13837 20914 15811
rect 21038 13837 21098 15947
rect 20851 13836 20917 13837
rect 19610 13568 19618 13632
rect 19682 13568 19698 13632
rect 19762 13568 19778 13632
rect 19842 13568 19858 13632
rect 19922 13568 19930 13632
rect 15883 13020 15949 13021
rect 15883 12956 15884 13020
rect 15948 12956 15949 13020
rect 15883 12955 15949 12956
rect 17723 13020 17789 13021
rect 17723 12956 17724 13020
rect 17788 12956 17789 13020
rect 17723 12955 17789 12956
rect 19379 13020 19445 13021
rect 19379 12956 19380 13020
rect 19444 12956 19445 13020
rect 19379 12955 19445 12956
rect 15518 12205 15578 12462
rect 15515 12204 15581 12205
rect 15515 12140 15516 12204
rect 15580 12140 15581 12204
rect 15515 12139 15581 12140
rect 14944 11936 14952 12000
rect 15016 11936 15032 12000
rect 15096 11936 15112 12000
rect 15176 11936 15192 12000
rect 15256 11936 15264 12000
rect 14043 11732 14044 11782
rect 14108 11732 14109 11782
rect 14043 11731 14109 11732
rect 14595 11660 14661 11661
rect 14595 11596 14596 11660
rect 14660 11596 14661 11660
rect 14595 11595 14661 11596
rect 14598 11338 14658 11595
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 13862 9349 13922 11051
rect 14944 10912 15264 11936
rect 15886 11253 15946 12955
rect 17726 12018 17786 12955
rect 19610 12544 19930 13568
rect 20115 13156 20181 13157
rect 20115 13092 20116 13156
rect 20180 13092 20181 13156
rect 20115 13091 20181 13092
rect 19610 12480 19618 12544
rect 19682 12480 19698 12544
rect 19762 12480 19778 12544
rect 19842 12480 19858 12544
rect 19922 12480 19930 12544
rect 15883 11252 15949 11253
rect 15883 11188 15884 11252
rect 15948 11188 15949 11252
rect 15883 11187 15949 11188
rect 14944 10848 14952 10912
rect 15016 10848 15032 10912
rect 15096 10848 15112 10912
rect 15176 10848 15192 10912
rect 15256 10848 15264 10912
rect 14944 9824 15264 10848
rect 14944 9760 14952 9824
rect 15016 9760 15032 9824
rect 15096 9760 15112 9824
rect 15176 9760 15192 9824
rect 15256 9760 15264 9824
rect 13859 9348 13925 9349
rect 13859 9284 13860 9348
rect 13924 9284 13925 9348
rect 13859 9283 13925 9284
rect 14944 8736 15264 9760
rect 14944 8672 14952 8736
rect 15016 8672 15032 8736
rect 15096 8672 15112 8736
rect 15176 8672 15192 8736
rect 15256 8672 15264 8736
rect 14944 7648 15264 8672
rect 15515 8396 15581 8397
rect 15515 8332 15516 8396
rect 15580 8332 15581 8396
rect 15515 8331 15581 8332
rect 14944 7584 14952 7648
rect 15016 7584 15032 7648
rect 15096 7584 15112 7648
rect 15176 7584 15192 7648
rect 15256 7584 15264 7648
rect 14944 6560 15264 7584
rect 14944 6496 14952 6560
rect 15016 6496 15032 6560
rect 15096 6496 15112 6560
rect 15176 6496 15192 6560
rect 15256 6496 15264 6560
rect 14944 5472 15264 6496
rect 14944 5408 14952 5472
rect 15016 5408 15032 5472
rect 15096 5408 15112 5472
rect 15176 5408 15192 5472
rect 15256 5408 15264 5472
rect 12387 5404 12453 5405
rect 12387 5340 12388 5404
rect 12452 5340 12453 5404
rect 12387 5339 12453 5340
rect 12390 4861 12450 5339
rect 12387 4860 12453 4861
rect 12387 4796 12388 4860
rect 12452 4796 12453 4860
rect 12387 4795 12453 4796
rect 14944 4384 15264 5408
rect 14944 4320 14952 4384
rect 15016 4320 15032 4384
rect 15096 4320 15112 4384
rect 15176 4320 15192 4384
rect 15256 4320 15264 4384
rect 11835 3636 11901 3637
rect 11835 3572 11836 3636
rect 11900 3572 11901 3636
rect 11835 3571 11901 3572
rect 10277 2688 10285 2752
rect 10349 2688 10365 2752
rect 10429 2688 10445 2752
rect 10509 2688 10525 2752
rect 10589 2688 10597 2752
rect 10277 2128 10597 2688
rect 14944 3296 15264 4320
rect 14944 3232 14952 3296
rect 15016 3232 15032 3296
rect 15096 3232 15112 3296
rect 15176 3232 15192 3296
rect 15256 3232 15264 3296
rect 12387 2684 12453 2685
rect 12387 2620 12388 2684
rect 12452 2620 12453 2684
rect 12387 2619 12453 2620
rect 12390 1869 12450 2619
rect 14944 2208 15264 3232
rect 14944 2144 14952 2208
rect 15016 2144 15032 2208
rect 15096 2144 15112 2208
rect 15176 2144 15192 2208
rect 15256 2144 15264 2208
rect 14944 2128 15264 2144
rect 15518 1869 15578 8331
rect 17726 7717 17786 9742
rect 19382 9621 19442 12462
rect 19610 11456 19930 12480
rect 19610 11392 19618 11456
rect 19682 11392 19698 11456
rect 19762 11392 19778 11456
rect 19842 11392 19858 11456
rect 19922 11392 19930 11456
rect 19610 10368 19930 11392
rect 20118 10437 20178 13091
rect 20115 10436 20181 10437
rect 20115 10372 20116 10436
rect 20180 10372 20181 10436
rect 20115 10371 20181 10372
rect 19610 10304 19618 10368
rect 19682 10304 19698 10368
rect 19762 10304 19778 10368
rect 19842 10304 19858 10368
rect 19922 10304 19930 10368
rect 19379 9620 19445 9621
rect 19379 9556 19380 9620
rect 19444 9556 19445 9620
rect 19379 9555 19445 9556
rect 19610 9280 19930 10304
rect 19610 9216 19618 9280
rect 19682 9216 19698 9280
rect 19762 9216 19778 9280
rect 19842 9216 19858 9280
rect 19922 9216 19930 9280
rect 19610 8192 19930 9216
rect 19610 8128 19618 8192
rect 19682 8128 19698 8192
rect 19762 8128 19778 8192
rect 19842 8128 19858 8192
rect 19922 8128 19930 8192
rect 17723 7716 17789 7717
rect 17723 7652 17724 7716
rect 17788 7652 17789 7716
rect 17723 7651 17789 7652
rect 19610 7104 19930 8128
rect 19610 7040 19618 7104
rect 19682 7040 19698 7104
rect 19762 7040 19778 7104
rect 19842 7040 19858 7104
rect 19922 7040 19930 7104
rect 19610 6016 19930 7040
rect 20302 6765 20362 13822
rect 20851 13772 20852 13836
rect 20916 13772 20917 13836
rect 20851 13771 20917 13772
rect 21035 13836 21101 13837
rect 21035 13772 21036 13836
rect 21100 13772 21101 13836
rect 21035 13771 21101 13772
rect 20667 13700 20733 13701
rect 20667 13636 20668 13700
rect 20732 13636 20733 13700
rect 20667 13635 20733 13636
rect 20670 10658 20730 13635
rect 21035 12884 21101 12885
rect 21035 12820 21036 12884
rect 21100 12820 21101 12884
rect 21035 12819 21101 12820
rect 21038 11389 21098 12819
rect 21035 11388 21101 11389
rect 21035 11324 21036 11388
rect 21100 11324 21101 11388
rect 21035 11323 21101 11324
rect 20670 9349 20730 10422
rect 21222 10298 21282 25195
rect 23611 24988 23677 24989
rect 23611 24924 23612 24988
rect 23676 24924 23677 24988
rect 23611 24923 23677 24924
rect 20854 10238 21282 10298
rect 20667 9348 20733 9349
rect 20667 9284 20668 9348
rect 20732 9284 20733 9348
rect 20667 9283 20733 9284
rect 20667 8532 20733 8533
rect 20667 8468 20668 8532
rect 20732 8468 20733 8532
rect 20667 8467 20733 8468
rect 20670 6765 20730 8467
rect 20854 7170 20914 10238
rect 20854 7110 21098 7170
rect 20299 6764 20365 6765
rect 20299 6700 20300 6764
rect 20364 6700 20365 6764
rect 20299 6699 20365 6700
rect 20667 6764 20733 6765
rect 20667 6700 20668 6764
rect 20732 6700 20733 6764
rect 20667 6699 20733 6700
rect 19610 5952 19618 6016
rect 19682 5952 19698 6016
rect 19762 5952 19778 6016
rect 19842 5952 19858 6016
rect 19922 5952 19930 6016
rect 19610 4928 19930 5952
rect 19610 4864 19618 4928
rect 19682 4864 19698 4928
rect 19762 4864 19778 4928
rect 19842 4864 19858 4928
rect 19922 4864 19930 4928
rect 16435 3908 16501 3909
rect 16435 3858 16436 3908
rect 16500 3858 16501 3908
rect 16806 2549 16866 4302
rect 19610 3840 19930 4864
rect 20670 4317 20730 4982
rect 20667 4316 20733 4317
rect 20667 4252 20668 4316
rect 20732 4252 20733 4316
rect 20667 4251 20733 4252
rect 19610 3776 19618 3840
rect 19682 3776 19698 3840
rect 19762 3776 19778 3840
rect 19842 3776 19858 3840
rect 19922 3776 19930 3840
rect 19610 2752 19930 3776
rect 21038 3773 21098 7110
rect 21590 6493 21650 21982
rect 21771 21588 21837 21589
rect 21771 21524 21772 21588
rect 21836 21524 21837 21588
rect 21771 21523 21837 21524
rect 21774 8805 21834 21523
rect 22507 17916 22573 17917
rect 22507 17852 22508 17916
rect 22572 17852 22573 17916
rect 22507 17851 22573 17852
rect 21955 12748 22021 12749
rect 21955 12684 21956 12748
rect 22020 12684 22021 12748
rect 21955 12683 22021 12684
rect 21958 9213 22018 12683
rect 22142 12069 22202 15862
rect 22323 14244 22389 14245
rect 22323 14180 22324 14244
rect 22388 14180 22389 14244
rect 22323 14179 22389 14180
rect 22139 12068 22205 12069
rect 22139 12004 22140 12068
rect 22204 12004 22205 12068
rect 22139 12003 22205 12004
rect 22326 11525 22386 14179
rect 22510 12613 22570 17851
rect 22875 17236 22941 17237
rect 22875 17172 22876 17236
rect 22940 17172 22941 17236
rect 22875 17171 22941 17172
rect 22507 12612 22573 12613
rect 22507 12548 22508 12612
rect 22572 12548 22573 12612
rect 22507 12547 22573 12548
rect 22323 11524 22389 11525
rect 22323 11460 22324 11524
rect 22388 11460 22389 11524
rect 22323 11459 22389 11460
rect 22878 9621 22938 17171
rect 23246 15061 23306 15182
rect 23243 15060 23309 15061
rect 23243 14996 23244 15060
rect 23308 14996 23309 15060
rect 23243 14995 23309 14996
rect 23614 13154 23674 24923
rect 23795 19140 23861 19141
rect 23795 19076 23796 19140
rect 23860 19076 23861 19140
rect 23795 19075 23861 19076
rect 23430 13094 23674 13154
rect 23430 11525 23490 13094
rect 23611 12204 23677 12205
rect 23611 12140 23612 12204
rect 23676 12140 23677 12204
rect 23798 12202 23858 19075
rect 23982 12205 24042 25331
rect 24277 25056 24597 25616
rect 25819 25604 25820 25668
rect 25884 25604 25885 25668
rect 25819 25603 25885 25604
rect 24277 24992 24285 25056
rect 24349 24992 24365 25056
rect 24429 24992 24445 25056
rect 24509 24992 24525 25056
rect 24589 24992 24597 25056
rect 24277 23968 24597 24992
rect 24277 23904 24285 23968
rect 24349 23904 24365 23968
rect 24429 23904 24445 23968
rect 24509 23904 24525 23968
rect 24589 23904 24597 23968
rect 24277 22880 24597 23904
rect 24715 23492 24781 23493
rect 24715 23428 24716 23492
rect 24780 23428 24781 23492
rect 24715 23427 24781 23428
rect 24277 22816 24285 22880
rect 24349 22816 24365 22880
rect 24429 22816 24445 22880
rect 24509 22816 24525 22880
rect 24589 22816 24597 22880
rect 24277 21792 24597 22816
rect 24277 21728 24285 21792
rect 24349 21728 24365 21792
rect 24429 21728 24445 21792
rect 24509 21728 24525 21792
rect 24589 21728 24597 21792
rect 24277 20704 24597 21728
rect 24277 20640 24285 20704
rect 24349 20640 24365 20704
rect 24429 20640 24445 20704
rect 24509 20640 24525 20704
rect 24589 20640 24597 20704
rect 24277 19616 24597 20640
rect 24277 19552 24285 19616
rect 24349 19552 24365 19616
rect 24429 19552 24445 19616
rect 24509 19552 24525 19616
rect 24589 19552 24597 19616
rect 24277 18528 24597 19552
rect 24277 18464 24285 18528
rect 24349 18464 24365 18528
rect 24429 18464 24445 18528
rect 24509 18464 24525 18528
rect 24589 18464 24597 18528
rect 24277 17440 24597 18464
rect 24277 17376 24285 17440
rect 24349 17376 24365 17440
rect 24429 17376 24445 17440
rect 24509 17376 24525 17440
rect 24589 17376 24597 17440
rect 24277 16352 24597 17376
rect 24277 16288 24285 16352
rect 24349 16288 24365 16352
rect 24429 16288 24445 16352
rect 24509 16288 24525 16352
rect 24589 16288 24597 16352
rect 24277 15264 24597 16288
rect 24277 15200 24285 15264
rect 24349 15200 24365 15264
rect 24429 15200 24445 15264
rect 24509 15200 24525 15264
rect 24589 15200 24597 15264
rect 24277 14176 24597 15200
rect 24718 14789 24778 23427
rect 24899 15060 24965 15061
rect 24899 14996 24900 15060
rect 24964 14996 24965 15060
rect 24899 14995 24965 14996
rect 24715 14788 24781 14789
rect 24715 14724 24716 14788
rect 24780 14724 24781 14788
rect 24715 14723 24781 14724
rect 24277 14112 24285 14176
rect 24349 14112 24365 14176
rect 24429 14112 24445 14176
rect 24509 14112 24525 14176
rect 24589 14112 24597 14176
rect 24277 13088 24597 14112
rect 24715 13428 24781 13429
rect 24715 13364 24716 13428
rect 24780 13364 24781 13428
rect 24715 13363 24781 13364
rect 24277 13024 24285 13088
rect 24349 13024 24365 13088
rect 24429 13024 24445 13088
rect 24509 13024 24525 13088
rect 24589 13024 24597 13088
rect 23611 12139 23677 12140
rect 23752 12142 23858 12202
rect 23979 12204 24045 12205
rect 23427 11524 23493 11525
rect 23427 11460 23428 11524
rect 23492 11460 23493 11524
rect 23427 11459 23493 11460
rect 22875 9620 22941 9621
rect 22875 9556 22876 9620
rect 22940 9556 22941 9620
rect 22875 9555 22941 9556
rect 21955 9212 22021 9213
rect 21955 9148 21956 9212
rect 22020 9148 22021 9212
rect 21955 9147 22021 9148
rect 21771 8804 21837 8805
rect 21771 8740 21772 8804
rect 21836 8740 21837 8804
rect 21771 8739 21837 8740
rect 21955 8396 22021 8397
rect 21955 8332 21956 8396
rect 22020 8332 22021 8396
rect 21955 8331 22021 8332
rect 21958 6629 22018 8331
rect 22875 8124 22941 8125
rect 22875 8060 22876 8124
rect 22940 8060 22941 8124
rect 22875 8059 22941 8060
rect 21955 6628 22021 6629
rect 21955 6564 21956 6628
rect 22020 6564 22021 6628
rect 21955 6563 22021 6564
rect 21587 6492 21653 6493
rect 21587 6428 21588 6492
rect 21652 6428 21653 6492
rect 21587 6427 21653 6428
rect 22878 6085 22938 8059
rect 22875 6084 22941 6085
rect 22875 6020 22876 6084
rect 22940 6020 22941 6084
rect 22875 6019 22941 6020
rect 21035 3772 21101 3773
rect 21035 3708 21036 3772
rect 21100 3708 21101 3772
rect 21035 3707 21101 3708
rect 23430 3229 23490 11459
rect 23614 5541 23674 12139
rect 23752 11658 23812 12142
rect 23979 12140 23980 12204
rect 24044 12140 24045 12204
rect 23979 12139 24045 12140
rect 24277 12000 24597 13024
rect 24277 11936 24285 12000
rect 24349 11936 24365 12000
rect 24429 11936 24445 12000
rect 24509 11936 24525 12000
rect 24589 11936 24597 12000
rect 23982 11661 24042 11782
rect 23979 11660 24045 11661
rect 23752 11598 23858 11658
rect 23611 5540 23677 5541
rect 23611 5476 23612 5540
rect 23676 5476 23677 5540
rect 23611 5475 23677 5476
rect 23798 4725 23858 11598
rect 23979 11596 23980 11660
rect 24044 11596 24045 11660
rect 23979 11595 24045 11596
rect 24277 10912 24597 11936
rect 24277 10848 24285 10912
rect 24349 10848 24365 10912
rect 24429 10848 24445 10912
rect 24509 10848 24525 10912
rect 24589 10848 24597 10912
rect 24277 9824 24597 10848
rect 24277 9760 24285 9824
rect 24349 9760 24365 9824
rect 24429 9760 24445 9824
rect 24509 9760 24525 9824
rect 24589 9760 24597 9824
rect 23979 9076 24045 9077
rect 23979 9012 23980 9076
rect 24044 9012 24045 9076
rect 23979 9011 24045 9012
rect 23795 4724 23861 4725
rect 23795 4660 23796 4724
rect 23860 4660 23861 4724
rect 23795 4659 23861 4660
rect 23611 3364 23677 3365
rect 23611 3300 23612 3364
rect 23676 3300 23677 3364
rect 23611 3299 23677 3300
rect 23427 3228 23493 3229
rect 23427 3164 23428 3228
rect 23492 3164 23493 3228
rect 23427 3163 23493 3164
rect 19610 2688 19618 2752
rect 19682 2688 19698 2752
rect 19762 2688 19778 2752
rect 19842 2688 19858 2752
rect 19922 2688 19930 2752
rect 16803 2548 16869 2549
rect 16803 2484 16804 2548
rect 16868 2484 16869 2548
rect 16803 2483 16869 2484
rect 19610 2128 19930 2688
rect 12387 1868 12453 1869
rect 12387 1804 12388 1868
rect 12452 1804 12453 1868
rect 12387 1803 12453 1804
rect 15515 1868 15581 1869
rect 15515 1804 15516 1868
rect 15580 1804 15581 1868
rect 23614 1818 23674 3299
rect 23982 2498 24042 9011
rect 24277 8736 24597 9760
rect 24277 8672 24285 8736
rect 24349 8672 24365 8736
rect 24429 8672 24445 8736
rect 24509 8672 24525 8736
rect 24589 8672 24597 8736
rect 24277 7648 24597 8672
rect 24277 7584 24285 7648
rect 24349 7584 24365 7648
rect 24429 7584 24445 7648
rect 24509 7584 24525 7648
rect 24589 7584 24597 7648
rect 24277 6560 24597 7584
rect 24277 6496 24285 6560
rect 24349 6496 24365 6560
rect 24429 6496 24445 6560
rect 24509 6496 24525 6560
rect 24589 6496 24597 6560
rect 24277 5472 24597 6496
rect 24277 5408 24285 5472
rect 24349 5408 24365 5472
rect 24429 5408 24445 5472
rect 24509 5408 24525 5472
rect 24589 5408 24597 5472
rect 24277 4384 24597 5408
rect 24277 4320 24285 4384
rect 24349 4320 24365 4384
rect 24429 4320 24445 4384
rect 24509 4320 24525 4384
rect 24589 4320 24597 4384
rect 24277 3296 24597 4320
rect 24718 4045 24778 13363
rect 24902 8261 24962 14995
rect 25086 10981 25146 20622
rect 25267 17916 25333 17917
rect 25267 17852 25268 17916
rect 25332 17852 25333 17916
rect 25267 17851 25333 17852
rect 25270 12477 25330 17851
rect 25267 12476 25333 12477
rect 25267 12412 25268 12476
rect 25332 12412 25333 12476
rect 25267 12411 25333 12412
rect 25083 10980 25149 10981
rect 25083 10916 25084 10980
rect 25148 10916 25149 10980
rect 25083 10915 25149 10916
rect 25454 9621 25514 23342
rect 25451 9620 25517 9621
rect 25451 9556 25452 9620
rect 25516 9556 25517 9620
rect 25451 9555 25517 9556
rect 24899 8260 24965 8261
rect 24899 8196 24900 8260
rect 24964 8196 24965 8260
rect 24899 8195 24965 8196
rect 25822 7581 25882 25603
rect 26374 9621 26434 21302
rect 26742 10301 26802 19262
rect 26739 10300 26805 10301
rect 26739 10236 26740 10300
rect 26804 10236 26805 10300
rect 26739 10235 26805 10236
rect 26371 9620 26437 9621
rect 26371 9556 26372 9620
rect 26436 9556 26437 9620
rect 26371 9555 26437 9556
rect 27294 8669 27354 17902
rect 27291 8668 27357 8669
rect 27291 8604 27292 8668
rect 27356 8604 27357 8668
rect 27291 8603 27357 8604
rect 25819 7580 25885 7581
rect 25819 7516 25820 7580
rect 25884 7516 25885 7580
rect 25819 7515 25885 7516
rect 24899 7036 24965 7037
rect 24899 6972 24900 7036
rect 24964 6972 24965 7036
rect 24899 6971 24965 6972
rect 24715 4044 24781 4045
rect 24715 3980 24716 4044
rect 24780 3980 24781 4044
rect 24715 3979 24781 3980
rect 24277 3232 24285 3296
rect 24349 3232 24365 3296
rect 24429 3232 24445 3296
rect 24509 3232 24525 3296
rect 24589 3232 24597 3296
rect 24277 2208 24597 3232
rect 24277 2144 24285 2208
rect 24349 2144 24365 2208
rect 24429 2144 24445 2208
rect 24509 2144 24525 2208
rect 24589 2144 24597 2208
rect 24277 2128 24597 2144
rect 15515 1803 15581 1804
rect 24902 1138 24962 6971
<< via4 >>
rect 2182 21982 2418 22218
rect 1630 17902 1866 18138
rect 2366 13972 2602 14058
rect 2366 13908 2452 13972
rect 2452 13908 2516 13972
rect 2516 13908 2602 13972
rect 2366 13822 2602 13908
rect 2366 9742 2602 9978
rect 4942 22812 5178 22898
rect 4942 22748 5028 22812
rect 5028 22748 5092 22812
rect 5092 22748 5178 22812
rect 4942 22662 5178 22748
rect 6414 23342 6650 23578
rect 5310 20772 5546 20858
rect 5310 20708 5396 20772
rect 5396 20708 5460 20772
rect 5460 20708 5546 20772
rect 5310 20622 5546 20708
rect 6046 17236 6282 17458
rect 6046 17222 6132 17236
rect 6132 17222 6196 17236
rect 6196 17222 6282 17236
rect 6046 15182 6282 15418
rect 5126 11782 5362 12018
rect 1998 5662 2234 5898
rect 5310 9062 5546 9298
rect 5310 7172 5546 7258
rect 5310 7108 5396 7172
rect 5396 7108 5460 7172
rect 5460 7108 5546 7172
rect 5310 7022 5546 7108
rect 2918 2262 3154 2498
rect 1998 1732 2234 1818
rect 1998 1668 2084 1732
rect 2084 1668 2148 1732
rect 2148 1668 2234 1732
rect 1998 1582 2234 1668
rect 4574 3636 4810 3858
rect 4574 3622 4660 3636
rect 4660 3622 4724 3636
rect 4724 3622 4810 3636
rect 9174 21452 9410 21538
rect 9174 21388 9260 21452
rect 9260 21388 9324 21452
rect 9324 21388 9410 21452
rect 9174 21302 9410 21388
rect 8990 19484 9076 19498
rect 9076 19484 9140 19498
rect 9140 19484 9226 19498
rect 8990 19262 9226 19484
rect 9542 16542 9778 16778
rect 9542 13822 9778 14058
rect 8070 13142 8306 13378
rect 7150 11116 7386 11338
rect 7150 11102 7236 11116
rect 7236 11102 7300 11116
rect 7300 11102 7386 11116
rect 6598 7702 6834 7938
rect 8070 5132 8306 5218
rect 8070 5068 8156 5132
rect 8156 5068 8220 5132
rect 8220 5068 8306 5132
rect 8070 4982 8306 5068
rect 9542 6342 9778 6578
rect 11750 17222 11986 17458
rect 11014 14044 11100 14058
rect 11100 14044 11164 14058
rect 11164 14044 11250 14058
rect 11014 13822 11250 14044
rect 11198 10422 11434 10658
rect 10830 5662 11066 5898
rect 6598 4302 6834 4538
rect 15430 22812 15666 22898
rect 15430 22748 15516 22812
rect 15516 22748 15580 22812
rect 15580 22748 15666 22812
rect 15430 22662 15666 22748
rect 14142 18582 14378 18818
rect 13222 16012 13458 16098
rect 13222 15948 13308 16012
rect 13308 15948 13372 16012
rect 13372 15948 13458 16012
rect 13222 15862 13458 15948
rect 13774 15196 14010 15418
rect 13774 15182 13860 15196
rect 13860 15182 13924 15196
rect 13924 15182 14010 15196
rect 14510 15182 14746 15418
rect 13590 13292 13826 13378
rect 13590 13228 13676 13292
rect 13676 13228 13740 13292
rect 13740 13228 13826 13292
rect 13590 13142 13826 13228
rect 13958 11796 14194 12018
rect 13958 11782 14044 11796
rect 14044 11782 14108 11796
rect 14108 11782 14194 11796
rect 20214 18582 20450 18818
rect 20582 17222 20818 17458
rect 20766 16542 21002 16778
rect 20214 13822 20450 14058
rect 15430 12462 15666 12698
rect 14510 11102 14746 11338
rect 19294 12462 19530 12698
rect 17638 11782 17874 12018
rect 17638 9742 17874 9978
rect 19294 7852 19530 7938
rect 19294 7788 19380 7852
rect 19380 7788 19444 7852
rect 19444 7788 19530 7852
rect 19294 7702 19530 7788
rect 20582 10422 20818 10658
rect 21502 21982 21738 22218
rect 21134 9212 21370 9298
rect 21134 9148 21220 9212
rect 21220 9148 21284 9212
rect 21284 9148 21370 9212
rect 21134 9062 21370 9148
rect 20582 6492 20818 6578
rect 20582 6428 20668 6492
rect 20668 6428 20732 6492
rect 20732 6428 20818 6492
rect 20582 6342 20818 6428
rect 20582 4982 20818 5218
rect 16718 4302 16954 4538
rect 16350 3844 16436 3858
rect 16436 3844 16500 3858
rect 16500 3844 16586 3858
rect 16350 3622 16586 3844
rect 22054 15862 22290 16098
rect 23158 15182 23394 15418
rect 25366 23342 25602 23578
rect 24998 20622 25234 20858
rect 23894 11782 24130 12018
rect 26286 21302 26522 21538
rect 26654 19262 26890 19498
rect 27206 17902 27442 18138
rect 25182 7172 25418 7258
rect 25182 7108 25268 7172
rect 25268 7108 25332 7172
rect 25332 7108 25418 7172
rect 25182 7022 25418 7108
rect 23894 2262 24130 2498
rect 23526 1582 23762 1818
rect 4022 902 4258 1138
rect 24814 902 25050 1138
<< metal5 >>
rect 6372 23578 25644 23620
rect 6372 23342 6414 23578
rect 6650 23342 25366 23578
rect 25602 23342 25644 23578
rect 6372 23300 25644 23342
rect 4900 22898 15708 22940
rect 4900 22662 4942 22898
rect 5178 22662 15430 22898
rect 15666 22662 15708 22898
rect 4900 22620 15708 22662
rect 2140 22218 21780 22260
rect 2140 21982 2182 22218
rect 2418 21982 21502 22218
rect 21738 21982 21780 22218
rect 2140 21940 21780 21982
rect 9132 21538 26564 21580
rect 9132 21302 9174 21538
rect 9410 21302 26286 21538
rect 26522 21302 26564 21538
rect 9132 21260 26564 21302
rect 5268 20858 25276 20900
rect 5268 20622 5310 20858
rect 5546 20622 24998 20858
rect 25234 20622 25276 20858
rect 5268 20580 25276 20622
rect 8948 19498 26932 19540
rect 8948 19262 8990 19498
rect 9226 19262 26654 19498
rect 26890 19262 26932 19498
rect 8948 19220 26932 19262
rect 14100 18818 20492 18860
rect 14100 18582 14142 18818
rect 14378 18582 20214 18818
rect 20450 18582 20492 18818
rect 14100 18540 20492 18582
rect 1588 18138 27484 18180
rect 1588 17902 1630 18138
rect 1866 17902 27206 18138
rect 27442 17902 27484 18138
rect 1588 17860 27484 17902
rect 6004 17458 20860 17500
rect 6004 17222 6046 17458
rect 6282 17222 11750 17458
rect 11986 17222 20582 17458
rect 20818 17222 20860 17458
rect 6004 17180 20860 17222
rect 9500 16778 21044 16820
rect 9500 16542 9542 16778
rect 9778 16542 20766 16778
rect 21002 16542 21044 16778
rect 9500 16500 21044 16542
rect 13180 16098 22332 16140
rect 13180 15862 13222 16098
rect 13458 15862 22054 16098
rect 22290 15862 22332 16098
rect 13180 15820 22332 15862
rect 6004 15418 14052 15460
rect 6004 15182 6046 15418
rect 6282 15182 13774 15418
rect 14010 15182 14052 15418
rect 6004 15140 14052 15182
rect 14468 15418 23436 15460
rect 14468 15182 14510 15418
rect 14746 15182 23158 15418
rect 23394 15182 23436 15418
rect 14468 15140 23436 15182
rect 2324 14058 9820 14100
rect 2324 13822 2366 14058
rect 2602 13822 9542 14058
rect 9778 13822 9820 14058
rect 2324 13780 9820 13822
rect 10972 14058 20492 14100
rect 10972 13822 11014 14058
rect 11250 13822 20214 14058
rect 20450 13822 20492 14058
rect 10972 13780 20492 13822
rect 8028 13378 13868 13420
rect 8028 13142 8070 13378
rect 8306 13142 13590 13378
rect 13826 13142 13868 13378
rect 8028 13100 13868 13142
rect 15388 12698 19572 12740
rect 15388 12462 15430 12698
rect 15666 12462 19294 12698
rect 19530 12462 19572 12698
rect 15388 12420 19572 12462
rect 5084 12018 14236 12060
rect 5084 11782 5126 12018
rect 5362 11782 13958 12018
rect 14194 11782 14236 12018
rect 5084 11740 14236 11782
rect 17596 12018 24172 12060
rect 17596 11782 17638 12018
rect 17874 11782 23894 12018
rect 24130 11782 24172 12018
rect 17596 11740 24172 11782
rect 7108 11338 14788 11380
rect 7108 11102 7150 11338
rect 7386 11102 14510 11338
rect 14746 11102 14788 11338
rect 7108 11060 14788 11102
rect 11156 10658 20860 10700
rect 11156 10422 11198 10658
rect 11434 10422 20582 10658
rect 20818 10422 20860 10658
rect 11156 10380 20860 10422
rect 2324 9978 17916 10020
rect 2324 9742 2366 9978
rect 2602 9742 17638 9978
rect 17874 9742 17916 9978
rect 2324 9700 17916 9742
rect 5268 9298 21412 9340
rect 5268 9062 5310 9298
rect 5546 9062 21134 9298
rect 21370 9062 21412 9298
rect 5268 9020 21412 9062
rect 6556 7938 19572 7980
rect 6556 7702 6598 7938
rect 6834 7702 19294 7938
rect 19530 7702 19572 7938
rect 6556 7660 19572 7702
rect 5268 7258 25460 7300
rect 5268 7022 5310 7258
rect 5546 7022 25182 7258
rect 25418 7022 25460 7258
rect 5268 6980 25460 7022
rect 9500 6578 20860 6620
rect 9500 6342 9542 6578
rect 9778 6342 20582 6578
rect 20818 6342 20860 6578
rect 9500 6300 20860 6342
rect 1956 5898 11108 5940
rect 1956 5662 1998 5898
rect 2234 5662 10830 5898
rect 11066 5662 11108 5898
rect 1956 5620 11108 5662
rect 8028 5218 20860 5260
rect 8028 4982 8070 5218
rect 8306 4982 20582 5218
rect 20818 4982 20860 5218
rect 8028 4940 20860 4982
rect 6556 4538 16996 4580
rect 6556 4302 6598 4538
rect 6834 4302 16718 4538
rect 16954 4302 16996 4538
rect 6556 4260 16996 4302
rect 4532 3858 16628 3900
rect 4532 3622 4574 3858
rect 4810 3622 16350 3858
rect 16586 3622 16628 3858
rect 4532 3580 16628 3622
rect 2876 2498 24172 2540
rect 2876 2262 2918 2498
rect 3154 2262 23894 2498
rect 24130 2262 24172 2498
rect 2876 2220 24172 2262
rect 1956 1818 23804 1860
rect 1956 1582 1998 1818
rect 2234 1582 23526 1818
rect 23762 1582 23804 1818
rect 1956 1540 23804 1582
rect 3980 1138 25092 1180
rect 3980 902 4022 1138
rect 4258 902 24814 1138
rect 25050 902 25092 1138
rect 3980 860 25092 902
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__S
timestamp 1604666999
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1932 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1604666999
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10
timestamp 1604666999
transform 1 0 2024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 2208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_22
timestamp 1604666999
transform 1 0 3128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28
timestamp 1604666999
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 1604666999
transform 1 0 3220 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3496 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 3312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 3496 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1604666999
transform 1 0 4692 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1604666999
transform 1 0 4324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1604666999
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 4324 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5060 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A0
timestamp 1604666999
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6072 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1604666999
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604666999
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_52
timestamp 1604666999
transform 1 0 5888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_56
timestamp 1604666999
transform 1 0 6256 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1604666999
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1604666999
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8372 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8832 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1604666999
transform 1 0 8648 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_86
timestamp 1604666999
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604666999
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604666999
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1604666999
transform 1 0 11500 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _113_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1604666999
transform 1 0 11868 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12880 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1604666999
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 1604666999
transform 1 0 14720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_142
timestamp 1604666999
transform 1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1604666999
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 14536 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1604666999
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 14904 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15088 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1604666999
transform 1 0 17204 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_175
timestamp 1604666999
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1604666999
transform 1 0 17572 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604666999
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604666999
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_197
timestamp 1604666999
transform 1 0 19228 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_193
timestamp 1604666999
transform 1 0 18860 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_196
timestamp 1604666999
transform 1 0 19136 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19044 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_208
timestamp 1604666999
transform 1 0 20240 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_203
timestamp 1604666999
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_200
timestamp 1604666999
transform 1 0 19504 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19412 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1604666999
transform 1 0 19872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20608 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1604666999
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_210
timestamp 1604666999
transform 1 0 20424 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 20976 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_214
timestamp 1604666999
transform 1 0 20792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21160 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_227
timestamp 1604666999
transform 1 0 21988 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_227
timestamp 1604666999
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1604666999
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604666999
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1604666999
transform 1 0 22172 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 22172 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_235
timestamp 1604666999
transform 1 0 22724 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 22908 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 22540 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1604666999
transform 1 0 22724 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_239
timestamp 1604666999
transform 1 0 23092 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604666999
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_243
timestamp 1604666999
transform 1 0 23460 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_239
timestamp 1604666999
transform 1 0 23092 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 23644 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1604666999
transform 1 0 23276 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 23368 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_254
timestamp 1604666999
transform 1 0 24472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 24656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_258
timestamp 1604666999
transform 1 0 24840 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_262
timestamp 1604666999
transform 1 0 25208 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_258
timestamp 1604666999
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 25024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 25024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1604666999
transform 1 0 25208 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_266
timestamp 1604666999
transform 1 0 25576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 25392 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25576 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_270
timestamp 1604666999
transform 1 0 25944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_269
timestamp 1604666999
transform 1 0 25852 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 26128 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A
timestamp 1604666999
transform 1 0 25760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_274
timestamp 1604666999
transform 1 0 26312 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 26864 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 26864 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1604666999
transform 1 0 2392 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__S
timestamp 1604666999
transform 1 0 1840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1604666999
transform 1 0 1656 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1604666999
transform 1 0 2024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__S
timestamp 1604666999
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__S
timestamp 1604666999
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604666999
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5796 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A0
timestamp 1604666999
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1604666999
transform 1 0 4876 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1604666999
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7728 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 1604666999
transform 1 0 7544 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1604666999
transform 1 0 7912 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_78
timestamp 1604666999
transform 1 0 8280 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604666999
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1604666999
transform 1 0 11224 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10672 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__S
timestamp 1604666999
transform 1 0 11040 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1604666999
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1604666999
transform 1 0 10856 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp 1604666999
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 12696 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_123
timestamp 1604666999
transform 1 0 12420 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1604666999
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_132
timestamp 1604666999
transform 1 0 13248 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 15640 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15456 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1604666999
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_149
timestamp 1604666999
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 17204 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 16836 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1604666999
transform 1 0 16468 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1604666999
transform 1 0 17020 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18768 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1604666999
transform 1 0 18032 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19780 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 20148 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1604666999
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1604666999
transform 1 0 19964 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 1604666999
transform 1 0 20332 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 22448 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 21896 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 22264 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_224
timestamp 1604666999
transform 1 0 21712 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_228
timestamp 1604666999
transform 1 0 22080 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 24012 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 23828 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 23460 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_241
timestamp 1604666999
transform 1 0 23276 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_245
timestamp 1604666999
transform 1 0 23644 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_258
timestamp 1604666999
transform 1 0 24840 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_262
timestamp 1604666999
transform 1 0 25208 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_266
timestamp 1604666999
transform 1 0 25576 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 25760 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_270
timestamp 1604666999
transform 1 0 25944 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 26128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_274
timestamp 1604666999
transform 1 0 26312 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 26864 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1604666999
transform 1 0 1748 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1604666999
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__S
timestamp 1604666999
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_16
timestamp 1604666999
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1604666999
transform 1 0 3312 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A1
timestamp 1604666999
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1604666999
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1604666999
transform 1 0 4140 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1604666999
transform 1 0 4508 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1604666999
transform 1 0 4876 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_50
timestamp 1604666999
transform 1 0 5704 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_54
timestamp 1604666999
transform 1 0 6072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1604666999
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9292 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9108 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8740 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1604666999
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_85
timestamp 1604666999
transform 1 0 8924 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1604666999
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10304 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10672 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 1604666999
transform 1 0 10488 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_106
timestamp 1604666999
transform 1 0 10856 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604666999
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604666999
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1604666999
transform 1 0 12696 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14260 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_139
timestamp 1604666999
transform 1 0 13892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_152
timestamp 1604666999
transform 1 0 15088 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1604666999
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_170
timestamp 1604666999
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_174
timestamp 1604666999
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp 1604666999
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19044 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1604666999
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1604666999
transform 1 0 19228 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1604666999
transform 1 0 21160 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 20976 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 19412 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_210
timestamp 1604666999
transform 1 0 20424 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1604666999
transform 1 0 20792 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 22172 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 22540 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 22908 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_227
timestamp 1604666999
transform 1 0 21988 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 1604666999
transform 1 0 22356 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_235
timestamp 1604666999
transform 1 0 22724 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1604666999
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_239
timestamp 1604666999
transform 1 0 23092 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_254
timestamp 1604666999
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1604666999
transform 1 0 25208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 26864 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1604666999
transform 1 0 25760 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_258
timestamp 1604666999
transform 1 0 24840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1604666999
transform 1 0 25576 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_270
timestamp 1604666999
transform 1 0 25944 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_274
timestamp 1604666999
transform 1 0 26312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__S
timestamp 1604666999
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1604666999
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1604666999
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604666999
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6532 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__S
timestamp 1604666999
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1604666999
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_55
timestamp 1604666999
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_78
timestamp 1604666999
transform 1 0 8280 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1604666999
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_82
timestamp 1604666999
transform 1 0 8648 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9292 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1604666999
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1604666999
transform 1 0 9476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10212 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 11776 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1604666999
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_108
timestamp 1604666999
transform 1 0 11040 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_112
timestamp 1604666999
transform 1 0 11408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13616 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 12788 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1604666999
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_125
timestamp 1604666999
transform 1 0 12604 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_133
timestamp 1604666999
transform 1 0 13340 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1604666999
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1604666999
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1604666999
transform 1 0 16836 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16284 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 16652 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_163
timestamp 1604666999
transform 1 0 16100 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1604666999
transform 1 0 16468 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18400 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 18032 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_180
timestamp 1604666999
transform 1 0 17664 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1604666999
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_197
timestamp 1604666999
transform 1 0 19228 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 19964 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20332 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_203
timestamp 1604666999
transform 1 0 19780 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_207
timestamp 1604666999
transform 1 0 20148 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1604666999
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 22448 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22264 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604666999
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_228
timestamp 1604666999
transform 1 0 22080 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1604666999
transform 1 0 24472 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 24012 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_241
timestamp 1604666999
transform 1 0 23276 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_247
timestamp 1604666999
transform 1 0 23828 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_258
timestamp 1604666999
transform 1 0 24840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604666999
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_266
timestamp 1604666999
transform 1 0 25576 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25760 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_270
timestamp 1604666999
transform 1 0 25944 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604666999
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 26864 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2576 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1604666999
transform 1 0 2392 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1604666999
transform 1 0 2024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_8
timestamp 1604666999
transform 1 0 1840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_12
timestamp 1604666999
transform 1 0 2208 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4600 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp 1604666999
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604666999
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604666999
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7728 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7544 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1604666999
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1604666999
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8740 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1604666999
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604666999
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_92
timestamp 1604666999
transform 1 0 9568 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1604666999
transform 1 0 10028 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10396 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604666999
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604666999
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1604666999
transform 1 0 12788 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_131
timestamp 1604666999
transform 1 0 13156 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15456 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13892 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 14904 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1604666999
transform 1 0 14720 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1604666999
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1604666999
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 19044 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_179
timestamp 1604666999
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1604666999
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_197
timestamp 1604666999
transform 1 0 19228 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 21160 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 20976 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1604666999
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_214
timestamp 1604666999
transform 1 0 20792 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_227
timestamp 1604666999
transform 1 0 21988 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_231
timestamp 1604666999
transform 1 0 22356 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_234
timestamp 1604666999
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_238
timestamp 1604666999
transform 1 0 23000 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_254
timestamp 1604666999
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1604666999
transform 1 0 25208 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 26864 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1604666999
transform 1 0 25760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1604666999
transform 1 0 26128 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604666999
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_266
timestamp 1604666999
transform 1 0 25576 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_270
timestamp 1604666999
transform 1 0 25944 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_274
timestamp 1604666999
transform 1 0 26312 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_8
timestamp 1604666999
transform 1 0 1840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1604666999
transform 1 0 1748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_3
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__S
timestamp 1604666999
transform 1 0 1656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1604666999
transform 1 0 2024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2208 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1604666999
transform 1 0 2392 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_25
timestamp 1604666999
transform 1 0 3404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1604666999
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604666999
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A1
timestamp 1604666999
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__S
timestamp 1604666999
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1604666999
transform 1 0 4508 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 4692 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1604666999
transform 1 0 4232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 3772 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_48
timestamp 1604666999
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_41
timestamp 1604666999
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5060 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5244 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_56
timestamp 1604666999
transform 1 0 6256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_52
timestamp 1604666999
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_58
timestamp 1604666999
transform 1 0 6440 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1604666999
transform 1 0 6072 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6072 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6808 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7728 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1604666999
transform 1 0 6624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_68
timestamp 1604666999
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_89
timestamp 1604666999
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp 1604666999
transform 1 0 8924 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_81
timestamp 1604666999
transform 1 0 8556 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1604666999
transform 1 0 9844 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_91
timestamp 1604666999
transform 1 0 9476 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10488 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1604666999
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_111
timestamp 1604666999
transform 1 0 11316 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_116
timestamp 1604666999
transform 1 0 11776 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1604666999
transform 1 0 11408 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l5_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1604666999
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12696 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12972 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_122
timestamp 1604666999
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_148
timestamp 1604666999
transform 1 0 14720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1604666999
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_156
timestamp 1604666999
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_152
timestamp 1604666999
transform 1 0 15088 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1604666999
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14904 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_160
timestamp 1604666999
transform 1 0 15824 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_167
timestamp 1604666999
transform 1 0 16468 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_163
timestamp 1604666999
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604666999
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_171
timestamp 1604666999
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16652 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16928 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604666999
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604666999
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604666999
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1604666999
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_191
timestamp 1604666999
transform 1 0 18676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19228 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 18860 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_207
timestamp 1604666999
transform 1 0 20148 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 1604666999
transform 1 0 19780 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 19596 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1604666999
transform 1 0 19412 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_217
timestamp 1604666999
transform 1 0 21068 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_214
timestamp 1604666999
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_210
timestamp 1604666999
transform 1 0 20424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_211
timestamp 1604666999
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20884 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21160 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_227
timestamp 1604666999
transform 1 0 21988 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_228
timestamp 1604666999
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_224
timestamp 1604666999
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 21896 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_235
timestamp 1604666999
transform 1 0 22724 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_231
timestamp 1604666999
transform 1 0 22356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22264 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 22908 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22540 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 22172 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 22448 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_239
timestamp 1604666999
transform 1 0 23092 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 1604666999
transform 1 0 23828 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_241
timestamp 1604666999
transform 1 0 23276 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23644 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_254
timestamp 1604666999
transform 1 0 24472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1604666999
transform 1 0 24656 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24012 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_258
timestamp 1604666999
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_262
timestamp 1604666999
transform 1 0 25208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1604666999
transform 1 0 24840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1604666999
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1604666999
transform 1 0 25208 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_266
timestamp 1604666999
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_266
timestamp 1604666999
transform 1 0 25576 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_270
timestamp 1604666999
transform 1 0 25944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_270
timestamp 1604666999
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 26128 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 26128 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1604666999
transform 1 0 25760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_274
timestamp 1604666999
transform 1 0 26312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_274
timestamp 1604666999
transform 1 0 26312 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 26864 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 26864 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__S
timestamp 1604666999
transform 1 0 1564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 2208 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_7
timestamp 1604666999
transform 1 0 1748 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_11
timestamp 1604666999
transform 1 0 2116 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_1__A0
timestamp 1604666999
transform 1 0 3404 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_23
timestamp 1604666999
transform 1 0 3220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604666999
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6072 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A1
timestamp 1604666999
transform 1 0 5428 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_2__A0
timestamp 1604666999
transform 1 0 5796 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1604666999
transform 1 0 4876 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_45
timestamp 1604666999
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_49
timestamp 1604666999
transform 1 0 5612 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_53
timestamp 1604666999
transform 1 0 5980 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7636 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_63
timestamp 1604666999
transform 1 0 6900 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1604666999
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 1604666999
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_84
timestamp 1604666999
transform 1 0 8832 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1604666999
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1604666999
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10304 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 1604666999
transform 1 0 12052 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_123
timestamp 1604666999
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_136
timestamp 1604666999
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1604666999
transform 1 0 15548 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_140
timestamp 1604666999
transform 1 0 13984 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_145
timestamp 1604666999
transform 1 0 14444 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1604666999
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_154
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16652 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 16100 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 16468 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_161
timestamp 1604666999
transform 1 0 15916 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_165
timestamp 1604666999
transform 1 0 16284 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19136 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1604666999
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_192
timestamp 1604666999
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20148 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1604666999
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 1604666999
transform 1 0 20332 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1604666999
transform 1 0 22448 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21896 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 1604666999
transform 1 0 21712 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_228
timestamp 1604666999
transform 1 0 22080 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1604666999
transform 1 0 24012 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 23644 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1604666999
transform 1 0 24748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_241
timestamp 1604666999
transform 1 0 23276 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_247
timestamp 1604666999
transform 1 0 23828 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_253
timestamp 1604666999
transform 1 0 24380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_259
timestamp 1604666999
transform 1 0 24932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1604666999
transform 1 0 25116 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_265
timestamp 1604666999
transform 1 0 25484 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 25668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_269
timestamp 1604666999
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 26036 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_276
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_273
timestamp 1604666999
transform 1 0 26220 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 26864 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1604666999
transform 1 0 1564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_14
timestamp 1604666999
transform 1 0 2392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1604666999
transform 1 0 2760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1604666999
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1604666999
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1604666999
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__S
timestamp 1604666999
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604666999
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1604666999
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5704 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1604666999
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_52
timestamp 1604666999
transform 1 0 5888 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_56
timestamp 1604666999
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 7636 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_67
timestamp 1604666999
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9200 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_80
timestamp 1604666999
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_84
timestamp 1604666999
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 1604666999
transform 1 0 10028 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1604666999
transform 1 0 10764 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11868 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1604666999
transform 1 0 10396 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_114
timestamp 1604666999
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1604666999
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13340 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13156 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12788 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1604666999
transform 1 0 12972 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1604666999
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1604666999
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1604666999
transform 1 0 15824 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_169
timestamp 1604666999
transform 1 0 16652 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604666999
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18124 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1604666999
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604666999
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_194
timestamp 1604666999
transform 1 0 18952 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1604666999
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_211
timestamp 1604666999
transform 1 0 20516 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1604666999
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21252 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22448 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 22816 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_228
timestamp 1604666999
transform 1 0 22080 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_234
timestamp 1604666999
transform 1 0 22632 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_238
timestamp 1604666999
transform 1 0 23000 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1604666999
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1604666999
transform 1 0 24564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23184 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_242
timestamp 1604666999
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_249
timestamp 1604666999
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_253
timestamp 1604666999
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 26864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1604666999
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A0
timestamp 1604666999
transform 1 0 25668 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A1
timestamp 1604666999
transform 1 0 26036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A1
timestamp 1604666999
transform 1 0 26404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_261
timestamp 1604666999
transform 1 0 25116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_265
timestamp 1604666999
transform 1 0 25484 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_269
timestamp 1604666999
transform 1 0 25852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_273
timestamp 1604666999
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__S
timestamp 1604666999
transform 1 0 2208 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_6
timestamp 1604666999
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1604666999
transform 1 0 2024 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1604666999
transform 1 0 4600 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A0
timestamp 1604666999
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604666999
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1604666999
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5244 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__S
timestamp 1604666999
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1604666999
transform 1 0 4784 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_44
timestamp 1604666999
transform 1 0 5152 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_64
timestamp 1604666999
transform 1 0 6992 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1604666999
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_73
timestamp 1604666999
transform 1 0 7820 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9752 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9016 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1604666999
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1604666999
transform 1 0 9200 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_103
timestamp 1604666999
transform 1 0 10580 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_107
timestamp 1604666999
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_111
timestamp 1604666999
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1604666999
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13800 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1604666999
transform 1 0 13616 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1604666999
transform 1 0 14628 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14168 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_140
timestamp 1604666999
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_144
timestamp 1604666999
transform 1 0 14352 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1604666999
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17204 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1604666999
transform 1 0 17020 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_177
timestamp 1604666999
transform 1 0 17388 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1604666999
transform 1 0 19320 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 17756 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18768 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17572 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19136 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_190
timestamp 1604666999
transform 1 0 18584 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1604666999
transform 1 0 18952 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 19872 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_202
timestamp 1604666999
transform 1 0 19688 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_206
timestamp 1604666999
transform 1 0 20056 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_210
timestamp 1604666999
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 22448 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1604666999
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_228
timestamp 1604666999
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1604666999
transform 1 0 24012 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 24564 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_241
timestamp 1604666999
transform 1 0 23276 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_245
timestamp 1604666999
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1604666999
transform 1 0 24380 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_257
timestamp 1604666999
transform 1 0 24748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_1__A1
timestamp 1604666999
transform 1 0 24932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1604666999
transform 1 0 25116 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_265
timestamp 1604666999
transform 1 0 25484 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l5_in_0__A0
timestamp 1604666999
transform 1 0 25668 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_269
timestamp 1604666999
transform 1 0 25852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_2__A0
timestamp 1604666999
transform 1 0 26036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_273
timestamp 1604666999
transform 1 0 26220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 26864 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1604666999
transform 1 0 2852 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1604666999
transform 1 0 2392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__A1
timestamp 1604666999
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_7
timestamp 1604666999
transform 1 0 1748 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_12
timestamp 1604666999
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_16
timestamp 1604666999
transform 1 0 2576 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1604666999
transform 1 0 4416 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1604666999
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1604666999
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_28
timestamp 1604666999
transform 1 0 3680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_32
timestamp 1604666999
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__S
timestamp 1604666999
transform 1 0 5428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_45
timestamp 1604666999
transform 1 0 5244 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_49
timestamp 1604666999
transform 1 0 5612 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_56
timestamp 1604666999
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7636 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604666999
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_67
timestamp 1604666999
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10212 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9568 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1604666999
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_94
timestamp 1604666999
transform 1 0 9752 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1604666999
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1604666999
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_116
timestamp 1604666999
transform 1 0 11776 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13248 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 13064 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12696 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_128
timestamp 1604666999
transform 1 0 12880 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 15180 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_151
timestamp 1604666999
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 1604666999
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 16744 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_168
timestamp 1604666999
transform 1 0 16560 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_172
timestamp 1604666999
transform 1 0 16928 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_176
timestamp 1604666999
transform 1 0 17296 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_179
timestamp 1604666999
transform 1 0 17572 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1604666999
transform 1 0 20516 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1604666999
transform 1 0 19964 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1604666999
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1604666999
transform 1 0 20148 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1604666999
transform 1 0 22080 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1604666999
transform 1 0 22632 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 21528 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 21896 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_220
timestamp 1604666999
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_224
timestamp 1604666999
transform 1 0 21712 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_232
timestamp 1604666999
transform 1 0 22448 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_236
timestamp 1604666999
transform 1 0 22816 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24104 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1604666999
transform 1 0 24472 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604666999
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_248
timestamp 1604666999
transform 1 0 23920 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_252
timestamp 1604666999
transform 1 0 24288 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_259
timestamp 1604666999
transform 1 0 24932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_263
timestamp 1604666999
transform 1 0 25300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A1
timestamp 1604666999
transform 1 0 25484 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_267
timestamp 1604666999
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_3__A0
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_271
timestamp 1604666999
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_275
timestamp 1604666999
transform 1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 26864 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1604666999
transform 1 0 2392 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2208 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A1
timestamp 1604666999
transform 1 0 1840 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_6
timestamp 1604666999
transform 1 0 1656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_10
timestamp 1604666999
transform 1 0 2024 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_7__S
timestamp 1604666999
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l3_in_3__A0
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 1604666999
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 1604666999
transform 1 0 4416 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6440 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4876 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5888 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1604666999
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_40
timestamp 1604666999
transform 1 0 4784 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_50
timestamp 1604666999
transform 1 0 5704 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1604666999
transform 1 0 6072 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1604666999
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_81
timestamp 1604666999
transform 1 0 8556 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1604666999
transform 1 0 8924 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1604666999
transform 1 0 9200 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_96
timestamp 1604666999
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10672 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_12_101
timestamp 1604666999
transform 1 0 10396 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1604666999
transform 1 0 12420 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1604666999
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14168 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1604666999
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1604666999
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_148
timestamp 1604666999
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1604666999
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 1604666999
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17756 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17572 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_190
timestamp 1604666999
transform 1 0 18584 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_194
timestamp 1604666999
transform 1 0 18952 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1604666999
transform 1 0 19228 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1604666999
transform 1 0 19688 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20240 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_201
timestamp 1604666999
transform 1 0 19596 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1604666999
transform 1 0 20056 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_210
timestamp 1604666999
transform 1 0 20424 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22448 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 21896 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 22264 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22908 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 1604666999
transform 1 0 21712 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_228
timestamp 1604666999
transform 1 0 22080 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_235
timestamp 1604666999
transform 1 0 22724 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1604666999
transform 1 0 24564 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24012 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 24380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_239
timestamp 1604666999
transform 1 0 23092 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_243
timestamp 1604666999
transform 1 0 23460 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_247
timestamp 1604666999
transform 1 0 23828 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_251
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_259
timestamp 1604666999
transform 1 0 24932 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25116 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_263
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25484 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_267
timestamp 1604666999
transform 1 0 25668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_271
timestamp 1604666999
transform 1 0 26036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_276
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 26864 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1604666999
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 1748 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_10
timestamp 1604666999
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_16
timestamp 1604666999
transform 1 0 2576 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2760 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 3312 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3128 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_20
timestamp 1604666999
transform 1 0 2944 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1604666999
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 1604666999
transform 1 0 4876 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_47
timestamp 1604666999
transform 1 0 5428 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_43
timestamp 1604666999
transform 1 0 5060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 5244 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_54
timestamp 1604666999
transform 1 0 6072 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1604666999
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604666999
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604666999
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1604666999
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5796 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6164 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_69
timestamp 1604666999
transform 1 0 7452 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_64
timestamp 1604666999
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 7268 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7084 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_78
timestamp 1604666999
transform 1 0 8280 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1604666999
transform 1 0 7912 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7728 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_89
timestamp 1604666999
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1604666999
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_81
timestamp 1604666999
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1604666999
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 8464 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 1604666999
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_14_100
timestamp 1604666999
transform 1 0 10304 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_109
timestamp 1604666999
transform 1 0 11132 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1604666999
transform 1 0 10764 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10948 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1604666999
transform 1 0 10856 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1604666999
transform 1 0 11684 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_113
timestamp 1604666999
transform 1 0 11500 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11868 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 11316 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1604666999
transform 1 0 12052 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_136
timestamp 1604666999
transform 1 0 13616 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_132
timestamp 1604666999
transform 1 0 13248 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1604666999
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_140
timestamp 1604666999
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_147
timestamp 1604666999
transform 1 0 14628 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_143
timestamp 1604666999
transform 1 0 14260 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14720 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1604666999
transform 1 0 14168 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1604666999
transform 1 0 13984 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_158
timestamp 1604666999
transform 1 0 15640 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1604666999
transform 1 0 14812 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1604666999
transform 1 0 14904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 15456 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15272 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_167
timestamp 1604666999
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_163
timestamp 1604666999
transform 1 0 16100 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 16284 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1604666999
transform 1 0 15916 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_174
timestamp 1604666999
transform 1 0 17112 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1604666999
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_174
timestamp 1604666999
transform 1 0 17112 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 16928 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1604666999
transform 1 0 17480 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1604666999
transform 1 0 16836 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_187
timestamp 1604666999
transform 1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1604666999
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_197
timestamp 1604666999
transform 1 0 19228 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_193
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 18492 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19044 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1604666999
transform 1 0 19044 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_208
timestamp 1604666999
transform 1 0 20240 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_204
timestamp 1604666999
transform 1 0 19872 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1604666999
transform 1 0 19596 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_217
timestamp 1604666999
transform 1 0 21068 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_214
timestamp 1604666999
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_210
timestamp 1604666999
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21160 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604666999
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_228
timestamp 1604666999
transform 1 0 22080 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_227
timestamp 1604666999
transform 1 0 21988 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 22172 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_232
timestamp 1604666999
transform 1 0 22448 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_231
timestamp 1604666999
transform 1 0 22356 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 22264 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 22540 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 22540 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_236
timestamp 1604666999
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_235
timestamp 1604666999
transform 1 0 22724 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22908 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp 1604666999
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_239
timestamp 1604666999
transform 1 0 23092 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 23276 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_247
timestamp 1604666999
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1604666999
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_251
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_249
timestamp 1604666999
transform 1 0 24012 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1604666999
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1604666999
transform 1 0 24564 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1604666999
transform 1 0 24564 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_259
timestamp 1604666999
transform 1 0 24932 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604666999
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25116 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1604666999
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_263
timestamp 1604666999
transform 1 0 25300 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_263
timestamp 1604666999
transform 1 0 25300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 25484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 25484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_267
timestamp 1604666999
transform 1 0 25668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_267
timestamp 1604666999
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_271
timestamp 1604666999
transform 1 0 26036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_271
timestamp 1604666999
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 26220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604666999
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 26864 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2668 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1604666999
transform 1 0 1932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1604666999
transform 1 0 1748 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_11
timestamp 1604666999
transform 1 0 2116 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604666999
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1604666999
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604666999
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1604666999
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1604666999
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1604666999
transform 1 0 9108 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_80
timestamp 1604666999
transform 1 0 8464 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 1604666999
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604666999
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10672 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 10488 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 13432 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1604666999
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_136
timestamp 1604666999
transform 1 0 13616 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 14260 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14076 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_140
timestamp 1604666999
transform 1 0 13984 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1604666999
transform 1 0 16744 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 16560 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604666999
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1604666999
transform 1 0 16376 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_173
timestamp 1604666999
transform 1 0 17020 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 19596 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1604666999
transform 1 0 21160 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19412 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_210
timestamp 1604666999
transform 1 0 20424 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_214
timestamp 1604666999
transform 1 0 20792 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 22540 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_227
timestamp 1604666999
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 1604666999
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_235
timestamp 1604666999
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1604666999
transform 1 0 24564 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23276 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24012 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 24380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_239
timestamp 1604666999
transform 1 0 23092 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_243
timestamp 1604666999
transform 1 0 23460 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_245
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_251
timestamp 1604666999
transform 1 0 24196 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_259
timestamp 1604666999
transform 1 0 24932 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1604666999
transform 1 0 25116 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_263
timestamp 1604666999
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_267
timestamp 1604666999
transform 1 0 25668 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_271
timestamp 1604666999
transform 1 0 26036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 26220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_275
timestamp 1604666999
transform 1 0 26404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 26864 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1604666999
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_10
timestamp 1604666999
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4508 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_36
timestamp 1604666999
transform 1 0 4416 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A0
timestamp 1604666999
transform 1 0 6440 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_56
timestamp 1604666999
transform 1 0 6256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1604666999
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_60
timestamp 1604666999
transform 1 0 6624 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_64
timestamp 1604666999
transform 1 0 6992 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_69
timestamp 1604666999
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1604666999
transform 1 0 10212 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_82
timestamp 1604666999
transform 1 0 8648 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_86
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_89
timestamp 1604666999
transform 1 0 9292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_97
timestamp 1604666999
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10488 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11500 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11868 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1604666999
transform 1 0 10396 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_111
timestamp 1604666999
transform 1 0 11316 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_115
timestamp 1604666999
transform 1 0 11684 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1604666999
transform 1 0 12052 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12696 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 12420 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_125
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_149
timestamp 1604666999
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_157
timestamp 1604666999
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16560 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 16192 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_161
timestamp 1604666999
transform 1 0 15916 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1604666999
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19044 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1604666999
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_191
timestamp 1604666999
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_204
timestamp 1604666999
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_208
timestamp 1604666999
transform 1 0 20240 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 22448 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 22264 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604666999
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_228
timestamp 1604666999
transform 1 0 22080 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24012 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23644 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_241
timestamp 1604666999
transform 1 0 23276 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_247
timestamp 1604666999
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_258
timestamp 1604666999
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_262
timestamp 1604666999
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25392 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_266
timestamp 1604666999
transform 1 0 25576 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25760 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_270
timestamp 1604666999
transform 1 0 25944 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_276
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 26864 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1748 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1604666999
transform 1 0 2576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 3312 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 3128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_20
timestamp 1604666999
transform 1 0 2944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5520 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1604666999
transform 1 0 5060 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_47
timestamp 1604666999
transform 1 0 5428 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_50
timestamp 1604666999
transform 1 0 5704 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_54
timestamp 1604666999
transform 1 0 6072 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9752 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 9568 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9200 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_81
timestamp 1604666999
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_85
timestamp 1604666999
transform 1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_90
timestamp 1604666999
transform 1 0 9384 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604666999
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_117
timestamp 1604666999
transform 1 0 11868 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15456 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14720 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1604666999
transform 1 0 14168 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_146
timestamp 1604666999
transform 1 0 14536 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_150
timestamp 1604666999
transform 1 0 14904 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20608 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19964 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1604666999
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1604666999
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_211
timestamp 1604666999
transform 1 0 20516 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_215
timestamp 1604666999
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21620 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 22632 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_219
timestamp 1604666999
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_232
timestamp 1604666999
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_236
timestamp 1604666999
transform 1 0 22816 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604666999
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_254
timestamp 1604666999
transform 1 0 24472 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1604666999
transform 1 0 25208 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 26864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1604666999
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_258
timestamp 1604666999
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_266
timestamp 1604666999
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_270
timestamp 1604666999
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_274
timestamp 1604666999
transform 1 0 26312 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2024 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp 1604666999
transform 1 0 1656 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1604666999
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1604666999
transform 1 0 4600 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A0
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604666999
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_36
timestamp 1604666999
transform 1 0 4416 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5520 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5152 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1604666999
transform 1 0 4784 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_46
timestamp 1604666999
transform 1 0 5336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_57
timestamp 1604666999
transform 1 0 6348 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7084 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6808 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_61
timestamp 1604666999
transform 1 0 6716 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_64
timestamp 1604666999
transform 1 0 6992 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1604666999
transform 1 0 7912 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1604666999
transform 1 0 8280 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9936 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp 1604666999
transform 1 0 8924 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_89
timestamp 1604666999
transform 1 0 9292 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_98
timestamp 1604666999
transform 1 0 10120 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10396 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 12604 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1604666999
transform 1 0 12144 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_124
timestamp 1604666999
transform 1 0 12512 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_127
timestamp 1604666999
transform 1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_140
timestamp 1604666999
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 14168 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1604666999
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 14536 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_148
timestamp 1604666999
transform 1 0 14720 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14904 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1604666999
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_158
timestamp 1604666999
transform 1 0 15640 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1604666999
transform 1 0 16192 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 15916 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 17204 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1604666999
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_173
timestamp 1604666999
transform 1 0 17020 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_177
timestamp 1604666999
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1604666999
transform 1 0 17848 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1604666999
transform 1 0 18860 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18676 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17572 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_181
timestamp 1604666999
transform 1 0 17756 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1604666999
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_189
timestamp 1604666999
transform 1 0 18492 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19872 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1604666999
transform 1 0 19688 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21528 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22908 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 21344 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 22540 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_219
timestamp 1604666999
transform 1 0 21252 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1604666999
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_235
timestamp 1604666999
transform 1 0 22724 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 24656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23092 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 24472 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_248
timestamp 1604666999
transform 1 0 23920 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_252
timestamp 1604666999
transform 1 0 24288 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 26864 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 26036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_265
timestamp 1604666999
transform 1 0 25484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_269
timestamp 1604666999
transform 1 0 25852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_273
timestamp 1604666999
transform 1 0 26220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_276
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_7
timestamp 1604666999
transform 1 0 1748 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__S
timestamp 1604666999
transform 1 0 1564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 1840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1604666999
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_17
timestamp 1604666999
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_19
timestamp 1604666999
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2024 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_25
timestamp 1604666999
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1604666999
transform 1 0 3036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp 1604666999
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_1__A1
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__S
timestamp 1604666999
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_37
timestamp 1604666999
transform 1 0 4508 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_36
timestamp 1604666999
transform 1 0 4416 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4324 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_40
timestamp 1604666999
transform 1 0 4784 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4968 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 4876 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1604666999
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_50
timestamp 1604666999
transform 1 0 5704 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1604666999
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_53
timestamp 1604666999
transform 1 0 5980 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5888 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6440 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6440 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1604666999
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1604666999
transform 1 0 8188 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604666999
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604666999
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8372 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1604666999
transform 1 0 9292 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp 1604666999
transform 1 0 8924 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1604666999
transform 1 0 8556 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_88
timestamp 1604666999
transform 1 0 9200 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8740 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1604666999
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9384 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9936 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604666999
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_102
timestamp 1604666999
transform 1 0 10488 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_109
timestamp 1604666999
transform 1 0 11132 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1604666999
transform 1 0 10764 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604666999
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1604666999
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1604666999
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604666999
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12788 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_136
timestamp 1604666999
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1604666999
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 13800 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1604666999
transform 1 0 12972 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_148
timestamp 1604666999
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1604666999
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_140
timestamp 1604666999
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1604666999
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14168 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 14536 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1604666999
transform 1 0 15640 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604666999
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1604666999
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 15548 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_163
timestamp 1604666999
transform 1 0 16100 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_159
timestamp 1604666999
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 15732 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 15916 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_178
timestamp 1604666999
transform 1 0 17480 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_174
timestamp 1604666999
transform 1 0 17112 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 1604666999
transform 1 0 16744 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604666999
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17296 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16928 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_183
timestamp 1604666999
transform 1 0 17940 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1604666999
transform 1 0 18124 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 18308 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_189
timestamp 1604666999
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 18308 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18676 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604666999
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604666999
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_217
timestamp 1604666999
transform 1 0 21068 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_214
timestamp 1604666999
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_210
timestamp 1604666999
transform 1 0 20424 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20884 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_224
timestamp 1604666999
transform 1 0 21712 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_221
timestamp 1604666999
transform 1 0 21436 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 21528 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 21988 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21712 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1604666999
transform 1 0 22172 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_237
timestamp 1604666999
transform 1 0 22908 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1604666999
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1604666999
transform 1 0 22540 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_247
timestamp 1604666999
transform 1 0 23828 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_242
timestamp 1604666999
transform 1 0 23368 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_241
timestamp 1604666999
transform 1 0 23276 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23644 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_254
timestamp 1604666999
transform 1 0 24472 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 24656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24104 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_259
timestamp 1604666999
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_258
timestamp 1604666999
transform 1 0 24840 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 25024 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 25116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1604666999
transform 1 0 25208 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604666999
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_263
timestamp 1604666999
transform 1 0 25300 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_266
timestamp 1604666999
transform 1 0 25576 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25484 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_271
timestamp 1604666999
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_270
timestamp 1604666999
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 26128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1604666999
transform 1 0 25760 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_276
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_274
timestamp 1604666999
transform 1 0 26312 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 26864 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 26864 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1604666999
transform 1 0 1564 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1604666999
transform 1 0 2392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_18
timestamp 1604666999
transform 1 0 2760 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 3404 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3220 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_22
timestamp 1604666999
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_34
timestamp 1604666999
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_38
timestamp 1604666999
transform 1 0 4600 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4968 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4784 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_51
timestamp 1604666999
transform 1 0 5796 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_55
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7176 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 6992 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604666999
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9844 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 9108 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1604666999
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_89
timestamp 1604666999
transform 1 0 9292 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 13984 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_149
timestamp 1604666999
transform 1 0 14812 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1604666999
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1604666999
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1604666999
transform 1 0 15824 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 16836 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17204 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1604666999
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1604666999
transform 1 0 17020 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_177
timestamp 1604666999
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1604666999
transform 1 0 18308 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19320 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_190
timestamp 1604666999
transform 1 0 18584 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_217
timestamp 1604666999
transform 1 0 21068 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 21804 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1604666999
transform 1 0 21252 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1604666999
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_234
timestamp 1604666999
transform 1 0 22632 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_238
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 24656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_254
timestamp 1604666999
transform 1 0 24472 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1604666999
transform 1 0 25208 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 26864 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1604666999
transform 1 0 25760 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 26128 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604666999
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_266
timestamp 1604666999
transform 1 0 25576 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_270
timestamp 1604666999
transform 1 0 25944 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_274
timestamp 1604666999
transform 1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 2208 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 1604666999
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_10
timestamp 1604666999
transform 1 0 2024 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4324 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_23
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l5_in_0__A1
timestamp 1604666999
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_54
timestamp 1604666999
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1604666999
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1604666999
transform 1 0 6808 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_66
timestamp 1604666999
transform 1 0 7176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_70
timestamp 1604666999
transform 1 0 7544 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9936 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604666999
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 11684 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_105
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1604666999
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_113
timestamp 1604666999
transform 1 0 11500 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1604666999
transform 1 0 11868 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 12144 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_22_139
timestamp 1604666999
transform 1 0 13892 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1604666999
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_157
timestamp 1604666999
transform 1 0 15548 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 16468 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 15824 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_162
timestamp 1604666999
transform 1 0 16008 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_166
timestamp 1604666999
transform 1 0 16376 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 18952 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 18768 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_186
timestamp 1604666999
transform 1 0 18216 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_190
timestamp 1604666999
transform 1 0 18584 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19964 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1604666999
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1604666999
transform 1 0 19780 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_207
timestamp 1604666999
transform 1 0 20148 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_211
timestamp 1604666999
transform 1 0 20516 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21988 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 21804 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_219
timestamp 1604666999
transform 1 0 21252 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_223
timestamp 1604666999
transform 1 0 21620 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1604666999
transform 1 0 24472 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 23920 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 24288 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_246
timestamp 1604666999
transform 1 0 23736 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1604666999
transform 1 0 24104 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 26864 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_263
timestamp 1604666999
transform 1 0 25300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_276
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2576 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1604666999
transform 1 0 1932 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 2392 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_11
timestamp 1604666999
transform 1 0 2116 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4140 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3956 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_25
timestamp 1604666999
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_29
timestamp 1604666999
transform 1 0 3772 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6072 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_52
timestamp 1604666999
transform 1 0 5888 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_56
timestamp 1604666999
transform 1 0 6256 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7084 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8096 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_78
timestamp 1604666999
transform 1 0 8280 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8648 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1604666999
transform 1 0 11132 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10856 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_105
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_108
timestamp 1604666999
transform 1 0 11040 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1604666999
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_116
timestamp 1604666999
transform 1 0 11776 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12512 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1604666999
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1604666999
transform 1 0 13708 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15456 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14076 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1604666999
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_148
timestamp 1604666999
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1604666999
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1604666999
transform 1 0 17204 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1604666999
transform 1 0 18308 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 18860 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1604666999
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_191
timestamp 1604666999
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1604666999
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19412 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 1604666999
transform 1 0 21160 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 21896 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 21712 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 21344 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 22908 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1604666999
transform 1 0 21528 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_235
timestamp 1604666999
transform 1 0 22724 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_239
timestamp 1604666999
transform 1 0 23092 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_254
timestamp 1604666999
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1604666999
transform 1 0 25208 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 26864 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1604666999
transform 1 0 25760 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 25024 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_258
timestamp 1604666999
transform 1 0 24840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_266
timestamp 1604666999
transform 1 0 25576 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_270
timestamp 1604666999
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_274
timestamp 1604666999
transform 1 0 26312 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 2392 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2024 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_6
timestamp 1604666999
transform 1 0 1656 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1604666999
transform 1 0 2208 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1604666999
transform 1 0 3220 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4876 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7084 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 7452 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_60
timestamp 1604666999
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1604666999
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_67
timestamp 1604666999
transform 1 0 7268 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1604666999
transform 1 0 7636 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604666999
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_96
timestamp 1604666999
transform 1 0 9936 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10856 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10488 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_100
timestamp 1604666999
transform 1 0 10304 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1604666999
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1604666999
transform 1 0 13340 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13156 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604666999
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_129
timestamp 1604666999
transform 1 0 12972 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 15456 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14720 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_142
timestamp 1604666999
transform 1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1604666999
transform 1 0 14536 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1604666999
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_158
timestamp 1604666999
transform 1 0 15640 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15732 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1604666999
transform 1 0 17480 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18216 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 17664 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19228 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1604666999
transform 1 0 17848 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_195
timestamp 1604666999
transform 1 0 19044 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 19780 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20240 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1604666999
transform 1 0 19412 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1604666999
transform 1 0 20056 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1604666999
transform 1 0 20424 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 21804 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_219
timestamp 1604666999
transform 1 0 21252 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_223
timestamp 1604666999
transform 1 0 21620 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1604666999
transform 1 0 24472 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 23920 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24288 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_246
timestamp 1604666999
transform 1 0 23736 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1604666999
transform 1 0 24104 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 26864 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25484 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_263
timestamp 1604666999
transform 1 0 25300 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_267
timestamp 1604666999
transform 1 0 25668 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_276
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2024 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1604666999
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1604666999
transform 1 0 2852 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 3036 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1604666999
transform 1 0 3220 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1604666999
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_40
timestamp 1604666999
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 8188 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1604666999
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1604666999
transform 1 0 7176 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_70
timestamp 1604666999
transform 1 0 7544 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 9752 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 9568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 9200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_86
timestamp 1604666999
transform 1 0 9016 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_90
timestamp 1604666999
transform 1 0 9384 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1604666999
transform 1 0 11316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1604666999
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_107
timestamp 1604666999
transform 1 0 10948 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12512 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_133
timestamp 1604666999
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_137
timestamp 1604666999
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 14812 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_141
timestamp 1604666999
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_145
timestamp 1604666999
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_158
timestamp 1604666999
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_162
timestamp 1604666999
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_175
timestamp 1604666999
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 19044 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604666999
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_193
timestamp 1604666999
transform 1 0 18860 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1604666999
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21160 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 19596 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1604666999
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_214
timestamp 1604666999
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 22724 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 22356 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_227
timestamp 1604666999
transform 1 0 21988 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1604666999
transform 1 0 22540 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1604666999
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 24656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1604666999
transform 1 0 23276 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_254
timestamp 1604666999
transform 1 0 24472 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1604666999
transform 1 0 25208 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 26864 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1604666999
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1604666999
transform 1 0 25024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 26128 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_258
timestamp 1604666999
transform 1 0 24840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_266
timestamp 1604666999
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_270
timestamp 1604666999
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_274
timestamp 1604666999
transform 1 0 26312 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_6
timestamp 1604666999
transform 1 0 1656 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_12
timestamp 1604666999
transform 1 0 2208 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 2024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 2116 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1604666999
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_30
timestamp 1604666999
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4232 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_27_40
timestamp 1604666999
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1604666999
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_53
timestamp 1604666999
transform 1 0 5980 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_55
timestamp 1604666999
transform 1 0 6164 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1604666999
transform 1 0 5796 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6440 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6532 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1604666999
transform 1 0 8280 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1604666999
transform 1 0 6624 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_85
timestamp 1604666999
transform 1 0 8924 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_81
timestamp 1604666999
transform 1 0 8556 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_88
timestamp 1604666999
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_82
timestamp 1604666999
transform 1 0 8648 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 8464 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8740 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 9292 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1604666999
transform 1 0 9476 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_97
timestamp 1604666999
transform 1 0 10028 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9660 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9844 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10304 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1604666999
transform 1 0 12052 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604666999
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12420 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_125
timestamp 1604666999
transform 1 0 12604 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1604666999
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1604666999
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_140
timestamp 1604666999
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_146
timestamp 1604666999
transform 1 0 14536 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1604666999
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14536 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_148
timestamp 1604666999
transform 1 0 14720 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1604666999
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_154
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1604666999
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_158
timestamp 1604666999
transform 1 0 15640 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15548 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1604666999
transform 1 0 15364 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_162
timestamp 1604666999
transform 1 0 16008 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1604666999
transform 1 0 16560 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_162
timestamp 1604666999
transform 1 0 16008 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16376 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 16192 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 16376 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1604666999
transform 1 0 15732 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1604666999
transform 1 0 16744 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_179
timestamp 1604666999
transform 1 0 17572 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_183
timestamp 1604666999
transform 1 0 17940 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604666999
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_186
timestamp 1604666999
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_187
timestamp 1604666999
transform 1 0 18308 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1604666999
transform 1 0 18676 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_196
timestamp 1604666999
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 18860 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 18492 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 19044 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_26_204
timestamp 1604666999
transform 1 0 19872 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_200
timestamp 1604666999
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19688 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_218
timestamp 1604666999
transform 1 0 21160 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_214
timestamp 1604666999
transform 1 0 20792 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604666999
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_228
timestamp 1604666999
transform 1 0 22080 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_224
timestamp 1604666999
transform 1 0 21712 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 21896 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 21344 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 21528 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604666999
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_231
timestamp 1604666999
transform 1 0 22356 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_232
timestamp 1604666999
transform 1 0 22448 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 22540 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 22632 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 22724 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 24656 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_254
timestamp 1604666999
transform 1 0 24472 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604666999
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1604666999
transform 1 0 24472 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_266
timestamp 1604666999
transform 1 0 25576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_258
timestamp 1604666999
transform 1 0 24840 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_266
timestamp 1604666999
transform 1 0 25576 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_258
timestamp 1604666999
transform 1 0 24840 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 25024 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1604666999
transform 1 0 25024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1604666999
transform 1 0 25208 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1604666999
transform 1 0 25208 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_270 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25944 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_274
timestamp 1604666999
transform 1 0 26312 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1604666999
transform 1 0 25760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_276
timestamp 1604666999
transform 1 0 26496 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_276
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 26864 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 26864 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1472 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4692 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 4324 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_23
timestamp 1604666999
transform 1 0 3220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604666999
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1604666999
transform 1 0 4508 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6440 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5888 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6256 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_50
timestamp 1604666999
transform 1 0 5704 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_54
timestamp 1604666999
transform 1 0 6072 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1604666999
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1604666999
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9200 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_84
timestamp 1604666999
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_90
timestamp 1604666999
transform 1 0 9384 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 11224 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10764 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_102
timestamp 1604666999
transform 1 0 10488 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_107
timestamp 1604666999
transform 1 0 10948 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_119
timestamp 1604666999
transform 1 0 12052 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 12788 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_123
timestamp 1604666999
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_136
timestamp 1604666999
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14168 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14536 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_140
timestamp 1604666999
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1604666999
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_148
timestamp 1604666999
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1604666999
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1604666999
transform 1 0 17020 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1604666999
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 18308 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A1
timestamp 1604666999
transform 1 0 17572 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__A0
timestamp 1604666999
transform 1 0 17940 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_181
timestamp 1604666999
transform 1 0 17756 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_185
timestamp 1604666999
transform 1 0 18124 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1604666999
transform 1 0 20056 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604666999
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_24.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22724 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 22540 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1604666999
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_228
timestamp 1604666999
transform 1 0 22080 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_232
timestamp 1604666999
transform 1 0 22448 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_254
timestamp 1604666999
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1604666999
transform 1 0 25208 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 26864 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_258
timestamp 1604666999
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_266
timestamp 1604666999
transform 1 0 25576 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604666999
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_276
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2208 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1604666999
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1604666999
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_31
timestamp 1604666999
transform 1 0 3956 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_35
timestamp 1604666999
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_39
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604666999
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604666999
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7544 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7360 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 6992 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_66
timestamp 1604666999
transform 1 0 7176 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1604666999
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1604666999
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 8556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 8924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1604666999
transform 1 0 8740 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_87
timestamp 1604666999
transform 1 0 9108 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_97
timestamp 1604666999
transform 1 0 10028 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604666999
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1604666999
transform 1 0 12512 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 13340 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 12972 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_127
timestamp 1604666999
transform 1 0 12788 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1604666999
transform 1 0 13156 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15088 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14904 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp 1604666999
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_148
timestamp 1604666999
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_171
timestamp 1604666999
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1604666999
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19044 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604666999
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1604666999
transform 1 0 18308 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_191
timestamp 1604666999
transform 1 0 18676 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20976 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_214
timestamp 1604666999
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1604666999
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21528 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_231
timestamp 1604666999
transform 1 0 22356 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_235
timestamp 1604666999
transform 1 0 22724 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 24656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604666999
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_254
timestamp 1604666999
transform 1 0 24472 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1604666999
transform 1 0 25208 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 26864 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1604666999
transform 1 0 25760 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1604666999
transform 1 0 25024 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_258
timestamp 1604666999
transform 1 0 24840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_266
timestamp 1604666999
transform 1 0 25576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_270
timestamp 1604666999
transform 1 0 25944 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_276
timestamp 1604666999
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2208 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 1840 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_6
timestamp 1604666999
transform 1 0 1656 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1604666999
transform 1 0 2024 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__S
timestamp 1604666999
transform 1 0 3404 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_23
timestamp 1604666999
transform 1 0 3220 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604666999
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604666999
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5336 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 5152 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_40
timestamp 1604666999
transform 1 0 4784 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7820 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_65
timestamp 1604666999
transform 1 0 7084 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1604666999
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10212 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604666999
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_88
timestamp 1604666999
transform 1 0 9200 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1604666999
transform 1 0 10028 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10764 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_101
timestamp 1604666999
transform 1 0 10396 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 13340 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_124
timestamp 1604666999
transform 1 0 12512 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_128
timestamp 1604666999
transform 1 0 12880 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1604666999
transform 1 0 14168 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_146
timestamp 1604666999
transform 1 0 14536 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_150
timestamp 1604666999
transform 1 0 14904 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_157
timestamp 1604666999
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16284 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15732 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 16100 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_161
timestamp 1604666999
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18768 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1604666999
transform 1 0 18032 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1604666999
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20976 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_201
timestamp 1604666999
transform 1 0 19596 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1604666999
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_209
timestamp 1604666999
transform 1 0 20332 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 22540 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21988 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_225
timestamp 1604666999
transform 1 0 21804 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_229
timestamp 1604666999
transform 1 0 22172 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 24472 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_252
timestamp 1604666999
transform 1 0 24288 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_256
timestamp 1604666999
transform 1 0 24656 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1604666999
transform 1 0 25024 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 26864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_264
timestamp 1604666999
transform 1 0 25392 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_272
timestamp 1604666999
transform 1 0 26128 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_276
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2668 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1604666999
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_11
timestamp 1604666999
transform 1 0 2116 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4232 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1604666999
transform 1 0 4048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_26
timestamp 1604666999
transform 1 0 3496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_30
timestamp 1604666999
transform 1 0 3864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_53
timestamp 1604666999
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8004 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1604666999
transform 1 0 7360 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 7820 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1604666999
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_70
timestamp 1604666999
transform 1 0 7544 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_94
timestamp 1604666999
transform 1 0 9752 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_98
timestamp 1604666999
transform 1 0 10120 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604666999
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604666999
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 13156 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12696 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_128
timestamp 1604666999
transform 1 0 12880 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 15088 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 14904 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1604666999
transform 1 0 13984 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_144
timestamp 1604666999
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1604666999
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16928 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 16100 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1604666999
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__S
timestamp 1604666999
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_161
timestamp 1604666999
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_165
timestamp 1604666999
transform 1 0 16284 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1604666999
transform 1 0 16652 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1604666999
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 18584 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 18400 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1604666999
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20148 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19964 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21160 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_199
timestamp 1604666999
transform 1 0 19412 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1604666999
transform 1 0 19780 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1604666999
transform 1 0 20976 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1604666999
transform 1 0 21988 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21528 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_220
timestamp 1604666999
transform 1 0 21344 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_224
timestamp 1604666999
transform 1 0 21712 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1604666999
transform 1 0 22816 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 24656 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604666999
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_254
timestamp 1604666999
transform 1 0 24472 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1604666999
transform 1 0 25208 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 26864 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A
timestamp 1604666999
transform 1 0 25760 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25024 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_258
timestamp 1604666999
transform 1 0 24840 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_266
timestamp 1604666999
transform 1 0 25576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_270
timestamp 1604666999
transform 1 0 25944 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_276
timestamp 1604666999
transform 1 0 26496 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A0
timestamp 1604666999
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_6
timestamp 1604666999
transform 1 0 1656 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_11
timestamp 1604666999
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4600 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1604666999
transform 1 0 4416 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5520 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__S
timestamp 1604666999
transform 1 0 5336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1604666999
transform 1 0 4784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7820 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7452 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1604666999
transform 1 0 7268 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1604666999
transform 1 0 7636 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604666999
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1604666999
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_96
timestamp 1604666999
transform 1 0 9936 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10672 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11684 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12052 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp 1604666999
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1604666999
transform 1 0 11500 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1604666999
transform 1 0 11868 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12696 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1604666999
transform 1 0 12236 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_125
timestamp 1604666999
transform 1 0 12604 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1604666999
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1604666999
transform 1 0 14812 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1604666999
transform 1 0 17020 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A0
timestamp 1604666999
transform 1 0 16376 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16836 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_163
timestamp 1604666999
transform 1 0 16100 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_168
timestamp 1604666999
transform 1 0 16560 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18584 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_182
timestamp 1604666999
transform 1 0 17848 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1604666999
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1604666999
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_203
timestamp 1604666999
transform 1 0 19780 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_209
timestamp 1604666999
transform 1 0 20332 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 22816 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_234
timestamp 1604666999
transform 1 0 22632 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_238
timestamp 1604666999
transform 1 0 23000 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23368 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 23184 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 26864 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 25116 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604666999
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_276
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A1
timestamp 1604666999
transform 1 0 1748 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_4__A1
timestamp 1604666999
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1604666999
transform 1 0 1932 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1604666999
transform 1 0 1932 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_18
timestamp 1604666999
transform 1 0 2760 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_18
timestamp 1604666999
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_28
timestamp 1604666999
transform 1 0 3680 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_24
timestamp 1604666999
transform 1 0 3312 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_26
timestamp 1604666999
transform 1 0 3496 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_22
timestamp 1604666999
transform 1 0 3128 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 3128 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3496 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1604666999
transform 1 0 3312 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A1
timestamp 1604666999
transform 1 0 2944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 3772 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_45
timestamp 1604666999
transform 1 0 5244 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1604666999
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1604666999
transform 1 0 5520 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 5428 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1604666999
transform 1 0 5612 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_58
timestamp 1604666999
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_56
timestamp 1604666999
transform 1 0 6256 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_52
timestamp 1604666999
transform 1 0 5888 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 6440 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 6072 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 5704 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6992 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1604666999
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_62
timestamp 1604666999
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7268 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_65
timestamp 1604666999
transform 1 0 7084 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1604666999
transform 1 0 7452 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 7176 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_79
timestamp 1604666999
transform 1 0 8372 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_75
timestamp 1604666999
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7820 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_87
timestamp 1604666999
transform 1 0 9108 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_83
timestamp 1604666999
transform 1 0 8740 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9292 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8556 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604666999
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_96
timestamp 1604666999
transform 1 0 9936 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_92
timestamp 1604666999
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10120 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_33_109
timestamp 1604666999
transform 1 0 11132 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10304 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp 1604666999
transform 1 0 11776 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_112
timestamp 1604666999
transform 1 0 11408 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_118
timestamp 1604666999
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_113
timestamp 1604666999
transform 1 0 11500 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11592 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11960 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 11316 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12144 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_136
timestamp 1604666999
transform 1 0 13616 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_133
timestamp 1604666999
transform 1 0 13340 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_129
timestamp 1604666999
transform 1 0 12972 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1604666999
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604666999
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13800 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_140
timestamp 1604666999
transform 1 0 13984 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14628 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 13984 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _133_
timestamp 1604666999
transform 1 0 14076 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1604666999
transform 1 0 14812 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_156
timestamp 1604666999
transform 1 0 15456 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_153
timestamp 1604666999
transform 1 0 15180 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_149
timestamp 1604666999
transform 1 0 14812 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1604666999
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_163
timestamp 1604666999
transform 1 0 16100 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_160
timestamp 1604666999
transform 1 0 15824 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__S
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1604666999
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1604666999
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604666999
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A1
timestamp 1604666999
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_3__S
timestamp 1604666999
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1604666999
transform 1 0 16928 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_185
timestamp 1604666999
transform 1 0 18124 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_181
timestamp 1604666999
transform 1 0 17756 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_188
timestamp 1604666999
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604666999
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A0
timestamp 1604666999
transform 1 0 17940 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__S
timestamp 1604666999
transform 1 0 18308 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _130_
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_198
timestamp 1604666999
transform 1 0 19320 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_192
timestamp 1604666999
transform 1 0 18768 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 18952 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1604666999
transform 1 0 18584 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18492 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19136 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_202
timestamp 1604666999
transform 1 0 19688 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19504 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1604666999
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 19872 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1604666999
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1604666999
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 21068 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1604666999
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_225
timestamp 1604666999
transform 1 0 21804 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_222
timestamp 1604666999
transform 1 0 21528 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_219
timestamp 1604666999
transform 1 0 21252 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21620 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21436 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21620 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_236
timestamp 1604666999
transform 1 0 22816 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_232
timestamp 1604666999
transform 1 0 22448 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 23000 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_16.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21896 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_34_245
timestamp 1604666999
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_240
timestamp 1604666999
transform 1 0 23184 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 23828 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_249
timestamp 1604666999
transform 1 0 24012 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_254
timestamp 1604666999
transform 1 0 24472 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 24656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1604666999
transform 1 0 24380 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_33_266
timestamp 1604666999
transform 1 0 25576 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_258
timestamp 1604666999
transform 1 0 24840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 25024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1604666999
transform 1 0 25208 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1604666999
transform 1 0 26312 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_274
timestamp 1604666999
transform 1 0 26312 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_270
timestamp 1604666999
transform 1 0 25944 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 26128 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A
timestamp 1604666999
transform 1 0 25760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 26864 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 26864 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1604666999
transform 1 0 25208 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1604666999
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A1
timestamp 1604666999
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1604666999
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1604666999
transform 1 0 3496 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 3312 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__A0
timestamp 1604666999
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_22
timestamp 1604666999
transform 1 0 3128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_35
timestamp 1604666999
transform 1 0 4324 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_39
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6072 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1604666999
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7636 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_60
timestamp 1604666999
transform 1 0 6624 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_66
timestamp 1604666999
transform 1 0 7176 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10120 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__A
timestamp 1604666999
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_90
timestamp 1604666999
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_35_95
timestamp 1604666999
transform 1 0 9844 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11132 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11500 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11868 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_107
timestamp 1604666999
transform 1 0 10948 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_111
timestamp 1604666999
transform 1 0 11316 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_115
timestamp 1604666999
transform 1 0 11684 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_119
timestamp 1604666999
transform 1 0 12052 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 13248 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13064 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 12696 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_123
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_128
timestamp 1604666999
transform 1 0 12880 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 15272 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_151
timestamp 1604666999
transform 1 0 14996 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_156
timestamp 1604666999
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1604666999
transform 1 0 16376 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__S
timestamp 1604666999
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__A1
timestamp 1604666999
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_160
timestamp 1604666999
transform 1 0 15824 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1604666999
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1604666999
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_1__S
timestamp 1604666999
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1604666999
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_184
timestamp 1604666999
transform 1 0 18032 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_196
timestamp 1604666999
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1604666999
transform 1 0 19872 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 19688 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20976 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_200
timestamp 1604666999
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_213
timestamp 1604666999
transform 1 0 20700 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_218
timestamp 1604666999
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21620 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_222
timestamp 1604666999
transform 1 0 21528 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_232
timestamp 1604666999
transform 1 0 22448 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_238
timestamp 1604666999
transform 1 0 23000 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1604666999
transform 1 0 23644 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_242
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_254
timestamp 1604666999
transform 1 0 24472 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1604666999
transform 1 0 25208 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 26864 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1604666999
transform 1 0 25760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 26128 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_258
timestamp 1604666999
transform 1 0 24840 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_266
timestamp 1604666999
transform 1 0 25576 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_270
timestamp 1604666999
transform 1 0 25944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_274
timestamp 1604666999
transform 1 0 26312 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1604666999
transform 1 0 1932 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__A0
timestamp 1604666999
transform 1 0 1748 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_18
timestamp 1604666999
transform 1 0 2760 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4232 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 2944 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 3496 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_22
timestamp 1604666999
transform 1 0 3128 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_28
timestamp 1604666999
transform 1 0 3680 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6440 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 5244 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5612 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 6256 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_43
timestamp 1604666999
transform 1 0 5060 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_47
timestamp 1604666999
transform 1 0 5428 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_51
timestamp 1604666999
transform 1 0 5796 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_55
timestamp 1604666999
transform 1 0 6164 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7636 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_67
timestamp 1604666999
transform 1 0 7268 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_73
timestamp 1604666999
transform 1 0 7820 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_84
timestamp 1604666999
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604666999
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_97
timestamp 1604666999
transform 1 0 10028 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10948 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10580 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_101
timestamp 1604666999
transform 1 0 10396 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_105
timestamp 1604666999
transform 1 0 10764 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13432 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 13248 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12880 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_126
timestamp 1604666999
transform 1 0 12696 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_130
timestamp 1604666999
transform 1 0 13064 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15272 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1604666999
transform 1 0 14260 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_147
timestamp 1604666999
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1604666999
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_173
timestamp 1604666999
transform 1 0 17020 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_177
timestamp 1604666999
transform 1 0 17388 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _128_
timestamp 1604666999
transform 1 0 19320 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1604666999
transform 1 0 17756 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 18952 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A1
timestamp 1604666999
transform 1 0 17572 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_190
timestamp 1604666999
transform 1 0 18584 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_196
timestamp 1604666999
transform 1 0 19136 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21068 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_202
timestamp 1604666999
transform 1 0 19688 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_206
timestamp 1604666999
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_210
timestamp 1604666999
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_215
timestamp 1604666999
transform 1 0 20884 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1604666999
transform 1 0 22816 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1604666999
transform 1 0 21252 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 22632 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 22264 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_228
timestamp 1604666999
transform 1 0 22080 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_232
timestamp 1604666999
transform 1 0 22448 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1604666999
transform 1 0 24380 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 23828 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_245
timestamp 1604666999
transform 1 0 23644 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_249
timestamp 1604666999
transform 1 0 24012 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_256
timestamp 1604666999
transform 1 0 24656 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25392 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 26864 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_267
timestamp 1604666999
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_276
timestamp 1604666999
transform 1 0 26496 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2668 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1604666999
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_7
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1604666999
transform 1 0 2116 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4232 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 3680 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4048 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_26
timestamp 1604666999
transform 1 0 3496 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_30
timestamp 1604666999
transform 1 0 3864 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604666999
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604666999
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8372 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8004 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_71
timestamp 1604666999
transform 1 0 7636 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_77
timestamp 1604666999
transform 1 0 8188 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_17.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8556 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _134_
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_100
timestamp 1604666999
transform 1 0 10304 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_106
timestamp 1604666999
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604666999
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604666999
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_132
timestamp 1604666999
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_136
timestamp 1604666999
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 14352 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14168 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_140
timestamp 1604666999
transform 1 0 13984 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _129_
timestamp 1604666999
transform 1 0 16836 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1604666999
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16468 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1604666999
transform 1 0 16100 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1604666999
transform 1 0 16652 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1604666999
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4_
timestamp 1604666999
transform 1 0 18860 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4__CLK
timestamp 1604666999
transform 1 0 18676 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_4__D
timestamp 1604666999
transform 1 0 18308 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l5_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1604666999
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_184
timestamp 1604666999
transform 1 0 18032 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_189
timestamp 1604666999
transform 1 0 18492 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 21160 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 20792 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_212
timestamp 1604666999
transform 1 0 20608 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_216
timestamp 1604666999
transform 1 0 20976 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21344 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_229
timestamp 1604666999
transform 1 0 22172 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_234
timestamp 1604666999
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_238
timestamp 1604666999
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _120_
timestamp 1604666999
transform 1 0 23644 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24748 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1604666999
transform 1 0 24196 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1604666999
transform 1 0 24564 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 23184 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_242
timestamp 1604666999
transform 1 0 23368 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_249
timestamp 1604666999
transform 1 0 24012 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_253
timestamp 1604666999
transform 1 0 24380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 26864 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25208 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_260
timestamp 1604666999
transform 1 0 25024 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_264
timestamp 1604666999
transform 1 0 25392 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_276
timestamp 1604666999
transform 1 0 26496 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1604666999
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_7__S
timestamp 1604666999
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_6
timestamp 1604666999
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_10
timestamp 1604666999
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A1
timestamp 1604666999
transform 1 0 4508 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3404 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_23
timestamp 1604666999
transform 1 0 3220 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_27
timestamp 1604666999
transform 1 0 3588 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_36
timestamp 1604666999
transform 1 0 4416 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_39
timestamp 1604666999
transform 1 0 4692 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4876 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7176 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_60
timestamp 1604666999
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_64
timestamp 1604666999
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_68
timestamp 1604666999
transform 1 0 7360 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_72
timestamp 1604666999
transform 1 0 7728 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 9016 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_84
timestamp 1604666999
transform 1 0 8832 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_88
timestamp 1604666999
transform 1 0 9200 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1604666999
transform 1 0 11224 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_102
timestamp 1604666999
transform 1 0 10488 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_38_107
timestamp 1604666999
transform 1 0 10948 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_119
timestamp 1604666999
transform 1 0 12052 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12788 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_125
timestamp 1604666999
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_136
timestamp 1604666999
transform 1 0 13616 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _127_
timestamp 1604666999
transform 1 0 15272 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14352 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14720 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_140
timestamp 1604666999
transform 1 0 13984 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_146
timestamp 1604666999
transform 1 0 14536 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1604666999
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_158
timestamp 1604666999
transform 1 0 15640 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16468 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 15824 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 16284 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_162
timestamp 1604666999
transform 1 0 16008 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 18952 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 18768 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_186
timestamp 1604666999
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_190
timestamp 1604666999
transform 1 0 18584 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20516 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 20148 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_203
timestamp 1604666999
transform 1 0 19780 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_209
timestamp 1604666999
transform 1 0 20332 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1604666999
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1604666999
transform 1 0 22448 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_224
timestamp 1604666999
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_228
timestamp 1604666999
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _117_
timestamp 1604666999
transform 1 0 24564 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 23460 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_241
timestamp 1604666999
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_245
timestamp 1604666999
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1604666999
transform 1 0 24380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 26864 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1604666999
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_259
timestamp 1604666999
transform 1 0 24932 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_271
timestamp 1604666999
transform 1 0 26036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_276
timestamp 1604666999
transform 1 0 26496 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1604666999
transform 1 0 1656 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1604666999
transform 1 0 1656 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_19
timestamp 1604666999
transform 1 0 2852 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_15
timestamp 1604666999
transform 1 0 2484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_19
timestamp 1604666999
transform 1 0 2852 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_15
timestamp 1604666999
transform 1 0 2484 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__S
timestamp 1604666999
transform 1 0 2668 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_6__S
timestamp 1604666999
transform 1 0 2668 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_27
timestamp 1604666999
transform 1 0 3588 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_23
timestamp 1604666999
transform 1 0 3220 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_23
timestamp 1604666999
transform 1 0 3220 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3772 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__S
timestamp 1604666999
transform 1 0 3036 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_32
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_36
timestamp 1604666999
transform 1 0 4416 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__S
timestamp 1604666999
transform 1 0 4324 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1604666999
transform 1 0 4508 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_46
timestamp 1604666999
transform 1 0 5336 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_40
timestamp 1604666999
transform 1 0 4784 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5520 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4968 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_54
timestamp 1604666999
transform 1 0 6072 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_50
timestamp 1604666999
transform 1 0 5704 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1604666999
transform 1 0 6348 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_53
timestamp 1604666999
transform 1 0 5980 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A0
timestamp 1604666999
transform 1 0 5888 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6440 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_3__A0
timestamp 1604666999
transform 1 0 6164 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_66
timestamp 1604666999
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__A
timestamp 1604666999
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_79
timestamp 1604666999
transform 1 0 8372 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_74
timestamp 1604666999
transform 1 0 7912 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_70
timestamp 1604666999
transform 1 0 7544 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8004 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_33.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6624 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8188 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_40_83
timestamp 1604666999
transform 1 0 8740 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1604666999
transform 1 0 9292 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1604666999
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_97
timestamp 1604666999
transform 1 0 10028 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_96
timestamp 1604666999
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10120 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10488 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10488 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11776 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10304 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_100
timestamp 1604666999
transform 1 0 10304 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_104
timestamp 1604666999
transform 1 0 10672 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_114
timestamp 1604666999
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1604666999
transform 1 0 11960 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_track_25.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A1
timestamp 1604666999
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_121
timestamp 1604666999
transform 1 0 12236 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_127
timestamp 1604666999
transform 1 0 12788 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_138
timestamp 1604666999
transform 1 0 13800 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_143
timestamp 1604666999
transform 1 0 14260 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_146
timestamp 1604666999
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1604666999
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_2__A0
timestamp 1604666999
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_158
timestamp 1604666999
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1604666999
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_150
timestamp 1604666999
transform 1 0 14904 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1604666999
transform 1 0 15088 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1604666999
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _121_
timestamp 1604666999
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 16560 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 15824 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__S
timestamp 1604666999
transform 1 0 16376 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_173
timestamp 1604666999
transform 1 0 17020 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_162
timestamp 1604666999
transform 1 0 16008 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_177
timestamp 1604666999
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_181
timestamp 1604666999
transform 1 0 17756 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1604666999
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17572 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A0
timestamp 1604666999
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1604666999
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 18124 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_198
timestamp 1604666999
transform 1 0 19320 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1604666999
transform 1 0 18952 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 19136 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_track_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 18032 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_40_206
timestamp 1604666999
transform 1 0 20056 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1604666999
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1604666999
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 19504 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1604666999
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _124_
timestamp 1604666999
transform 1 0 19688 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1604666999
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_210
timestamp 1604666999
transform 1 0 20424 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20516 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1604666999
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 20516 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_228
timestamp 1604666999
transform 1 0 22080 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1604666999
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_224
timestamp 1604666999
transform 1 0 21712 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_220
timestamp 1604666999
transform 1 0 21344 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 21528 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1604666999
transform 1 0 21896 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _126_
timestamp 1604666999
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_236
timestamp 1604666999
transform 1 0 22816 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_232
timestamp 1604666999
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1604666999
transform 1 0 22632 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _122_
timestamp 1604666999
transform 1 0 22448 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_236
timestamp 1604666999
transform 1 0 22816 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _116_
timestamp 1604666999
transform 1 0 24564 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _118_
timestamp 1604666999
transform 1 0 24472 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1604666999
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1604666999
transform 1 0 24380 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1604666999
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_40_248
timestamp 1604666999
transform 1 0 23920 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_259
timestamp 1604666999
transform 1 0 24932 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A
timestamp 1604666999
transform 1 0 25116 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_276
timestamp 1604666999
transform 1 0 26496 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_274
timestamp 1604666999
transform 1 0 26312 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_270
timestamp 1604666999
transform 1 0 25944 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_275
timestamp 1604666999
transform 1 0 26404 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1604666999
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 26864 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 26864 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_258
timestamp 1604666999
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_263
timestamp 1604666999
transform 1 0 25300 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1604666999
transform 1 0 2484 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1604666999
transform 1 0 1932 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1604666999
transform 1 0 2300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1604666999
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_11
timestamp 1604666999
transform 1 0 2116 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_19
timestamp 1604666999
transform 1 0 2852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4600 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 3588 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A
timestamp 1604666999
transform 1 0 3036 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__A
timestamp 1604666999
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A
timestamp 1604666999
transform 1 0 3404 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_23
timestamp 1604666999
transform 1 0 3220 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_30
timestamp 1604666999
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_34
timestamp 1604666999
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 5612 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A1
timestamp 1604666999
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_47
timestamp 1604666999
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_51
timestamp 1604666999
transform 1 0 5796 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_55
timestamp 1604666999
transform 1 0 6164 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _131_
timestamp 1604666999
transform 1 0 7084 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8188 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 8004 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_69
timestamp 1604666999
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_73
timestamp 1604666999
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1604666999
transform 1 0 9752 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 9568 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 9200 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_86
timestamp 1604666999
transform 1 0 9016 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_90
timestamp 1604666999
transform 1 0 9384 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1604666999
transform 1 0 11316 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1604666999
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10948 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_103
timestamp 1604666999
transform 1 0 10580 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1604666999
transform 1 0 11132 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1604666999
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1604666999
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12512 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_133
timestamp 1604666999
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_137
timestamp 1604666999
transform 1 0 13708 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 14076 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1604666999
transform 1 0 15088 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 13892 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_150
timestamp 1604666999
transform 1 0 14904 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_154
timestamp 1604666999
transform 1 0 15272 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1604666999
transform 1 0 15732 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1604666999
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1604666999
transform 1 0 17112 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_168
timestamp 1604666999
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_172
timestamp 1604666999
transform 1 0 16928 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_176
timestamp 1604666999
transform 1 0 17296 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1604666999
transform 1 0 18032 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1604666999
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19044 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_180
timestamp 1604666999
transform 1 0 17664 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_193
timestamp 1604666999
transform 1 0 18860 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_197
timestamp 1604666999
transform 1 0 19228 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 19596 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1604666999
transform 1 0 21160 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 19412 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_210
timestamp 1604666999
transform 1 0 20424 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_214
timestamp 1604666999
transform 1 0 20792 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _123_
timestamp 1604666999
transform 1 0 21620 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1604666999
transform 1 0 22172 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_220
timestamp 1604666999
transform 1 0 21344 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_227
timestamp 1604666999
transform 1 0 21988 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_231
timestamp 1604666999
transform 1 0 22356 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 1604666999
transform 1 0 23920 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1604666999
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1604666999
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1604666999
transform 1 0 23460 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_245
timestamp 1604666999
transform 1 0 23644 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_252
timestamp 1604666999
transform 1 0 24288 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_256
timestamp 1604666999
transform 1 0 24656 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 26864 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_268
timestamp 1604666999
transform 1 0 25760 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_276
timestamp 1604666999
transform 1 0 26496 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1604666999
transform 1 0 2484 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_2__A1
timestamp 1604666999
transform 1 0 1932 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_7
timestamp 1604666999
transform 1 0 1748 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_11
timestamp 1604666999
transform 1 0 2116 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_19
timestamp 1604666999
transform 1 0 2852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3588 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 4600 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1604666999
transform 1 0 3220 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_29
timestamp 1604666999
transform 1 0 3772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_36
timestamp 1604666999
transform 1 0 4416 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1604666999
transform 1 0 5152 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4968 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l3_in_3__A0
timestamp 1604666999
transform 1 0 5612 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_40
timestamp 1604666999
transform 1 0 4784 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_47
timestamp 1604666999
transform 1 0 5428 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_51
timestamp 1604666999
transform 1 0 5796 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_59
timestamp 1604666999
transform 1 0 6532 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1604666999
transform 1 0 7452 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 7268 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1604666999
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_63
timestamp 1604666999
transform 1 0 6900 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_78
timestamp 1604666999
transform 1 0 8280 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1604666999
transform 1 0 8648 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_86
timestamp 1604666999
transform 1 0 9016 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_90
timestamp 1604666999
transform 1 0 9384 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1604666999
transform 1 0 9476 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_94
timestamp 1604666999
transform 1 0 9752 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _135_
timestamp 1604666999
transform 1 0 9844 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_99
timestamp 1604666999
transform 1 0 10212 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10948 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__S
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10396 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_103
timestamp 1604666999
transform 1 0 10580 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_116
timestamp 1604666999
transform 1 0 11776 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1604666999
transform 1 0 12604 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1604666999
transform 1 0 12512 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 12328 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_120
timestamp 1604666999
transform 1 0 12144 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_134
timestamp 1604666999
transform 1 0 13432 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _132_
timestamp 1604666999
transform 1 0 14260 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1604666999
transform 1 0 15364 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 14076 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1604666999
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_140
timestamp 1604666999
transform 1 0 13984 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1604666999
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_151
timestamp 1604666999
transform 1 0 14996 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_156
timestamp 1604666999
transform 1 0 15456 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1604666999
transform 1 0 16468 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 15732 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1604666999
transform 1 0 16100 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_161
timestamp 1604666999
transform 1 0 15916 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1604666999
transform 1 0 16284 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_176
timestamp 1604666999
transform 1 0 17296 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 18584 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1604666999
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__A1
timestamp 1604666999
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_4__S
timestamp 1604666999
transform 1 0 17664 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_182
timestamp 1604666999
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_187
timestamp 1604666999
transform 1 0 18308 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _125_
timestamp 1604666999
transform 1 0 21160 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1604666999
transform 1 0 21068 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19596 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19964 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_199
timestamp 1604666999
transform 1 0 19412 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_203
timestamp 1604666999
transform 1 0 19780 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_207
timestamp 1604666999
transform 1 0 20148 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1604666999
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_222
timestamp 1604666999
transform 1 0 21528 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_234
timestamp 1604666999
transform 1 0 22632 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1604666999
transform 1 0 23920 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_246
timestamp 1604666999
transform 1 0 23736 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_249
timestamp 1604666999
transform 1 0 24012 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 26864 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1604666999
transform 1 0 25116 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_273
timestamp 1604666999
transform 1 0 26220 0 -1 25568
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_34_
port 0 nsew default input
rlabel metal2 s 662 0 718 480 6 bottom_left_grid_pin_35_
port 1 nsew default input
rlabel metal2 s 1214 0 1270 480 6 bottom_left_grid_pin_36_
port 2 nsew default input
rlabel metal2 s 1766 0 1822 480 6 bottom_left_grid_pin_37_
port 3 nsew default input
rlabel metal2 s 2318 0 2374 480 6 bottom_left_grid_pin_38_
port 4 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_39_
port 5 nsew default input
rlabel metal2 s 3422 0 3478 480 6 bottom_left_grid_pin_40_
port 6 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_left_grid_pin_41_
port 7 nsew default input
rlabel metal2 s 5078 0 5134 480 6 ccff_head
port 8 nsew default input
rlabel metal2 s 5630 0 5686 480 6 ccff_tail
port 9 nsew default tristate
rlabel metal3 s 0 280 480 400 6 chanx_left_in[0]
port 10 nsew default input
rlabel metal3 s 0 5992 480 6112 6 chanx_left_in[10]
port 11 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[11]
port 12 nsew default input
rlabel metal3 s 0 7216 480 7336 6 chanx_left_in[12]
port 13 nsew default input
rlabel metal3 s 0 7760 480 7880 6 chanx_left_in[13]
port 14 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[14]
port 15 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[15]
port 16 nsew default input
rlabel metal3 s 0 9528 480 9648 6 chanx_left_in[16]
port 17 nsew default input
rlabel metal3 s 0 10072 480 10192 6 chanx_left_in[17]
port 18 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[18]
port 19 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[19]
port 20 nsew default input
rlabel metal3 s 0 824 480 944 6 chanx_left_in[1]
port 21 nsew default input
rlabel metal3 s 0 1368 480 1488 6 chanx_left_in[2]
port 22 nsew default input
rlabel metal3 s 0 1912 480 2032 6 chanx_left_in[3]
port 23 nsew default input
rlabel metal3 s 0 2592 480 2712 6 chanx_left_in[4]
port 24 nsew default input
rlabel metal3 s 0 3136 480 3256 6 chanx_left_in[5]
port 25 nsew default input
rlabel metal3 s 0 3680 480 3800 6 chanx_left_in[6]
port 26 nsew default input
rlabel metal3 s 0 4360 480 4480 6 chanx_left_in[7]
port 27 nsew default input
rlabel metal3 s 0 4904 480 5024 6 chanx_left_in[8]
port 28 nsew default input
rlabel metal3 s 0 5448 480 5568 6 chanx_left_in[9]
port 29 nsew default input
rlabel metal3 s 0 11840 480 11960 6 chanx_left_out[0]
port 30 nsew default tristate
rlabel metal3 s 0 17688 480 17808 6 chanx_left_out[10]
port 31 nsew default tristate
rlabel metal3 s 0 18368 480 18488 6 chanx_left_out[11]
port 32 nsew default tristate
rlabel metal3 s 0 18912 480 19032 6 chanx_left_out[12]
port 33 nsew default tristate
rlabel metal3 s 0 19456 480 19576 6 chanx_left_out[13]
port 34 nsew default tristate
rlabel metal3 s 0 20000 480 20120 6 chanx_left_out[14]
port 35 nsew default tristate
rlabel metal3 s 0 20680 480 20800 6 chanx_left_out[15]
port 36 nsew default tristate
rlabel metal3 s 0 21224 480 21344 6 chanx_left_out[16]
port 37 nsew default tristate
rlabel metal3 s 0 21768 480 21888 6 chanx_left_out[17]
port 38 nsew default tristate
rlabel metal3 s 0 22448 480 22568 6 chanx_left_out[18]
port 39 nsew default tristate
rlabel metal3 s 0 22992 480 23112 6 chanx_left_out[19]
port 40 nsew default tristate
rlabel metal3 s 0 12520 480 12640 6 chanx_left_out[1]
port 41 nsew default tristate
rlabel metal3 s 0 13064 480 13184 6 chanx_left_out[2]
port 42 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[3]
port 43 nsew default tristate
rlabel metal3 s 0 14288 480 14408 6 chanx_left_out[4]
port 44 nsew default tristate
rlabel metal3 s 0 14832 480 14952 6 chanx_left_out[5]
port 45 nsew default tristate
rlabel metal3 s 0 15376 480 15496 6 chanx_left_out[6]
port 46 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[7]
port 47 nsew default tristate
rlabel metal3 s 0 16600 480 16720 6 chanx_left_out[8]
port 48 nsew default tristate
rlabel metal3 s 0 17144 480 17264 6 chanx_left_out[9]
port 49 nsew default tristate
rlabel metal3 s 27520 280 28000 400 6 chanx_right_in[0]
port 50 nsew default input
rlabel metal3 s 27520 5992 28000 6112 6 chanx_right_in[10]
port 51 nsew default input
rlabel metal3 s 27520 6672 28000 6792 6 chanx_right_in[11]
port 52 nsew default input
rlabel metal3 s 27520 7216 28000 7336 6 chanx_right_in[12]
port 53 nsew default input
rlabel metal3 s 27520 7760 28000 7880 6 chanx_right_in[13]
port 54 nsew default input
rlabel metal3 s 27520 8440 28000 8560 6 chanx_right_in[14]
port 55 nsew default input
rlabel metal3 s 27520 8984 28000 9104 6 chanx_right_in[15]
port 56 nsew default input
rlabel metal3 s 27520 9528 28000 9648 6 chanx_right_in[16]
port 57 nsew default input
rlabel metal3 s 27520 10072 28000 10192 6 chanx_right_in[17]
port 58 nsew default input
rlabel metal3 s 27520 10752 28000 10872 6 chanx_right_in[18]
port 59 nsew default input
rlabel metal3 s 27520 11296 28000 11416 6 chanx_right_in[19]
port 60 nsew default input
rlabel metal3 s 27520 824 28000 944 6 chanx_right_in[1]
port 61 nsew default input
rlabel metal3 s 27520 1368 28000 1488 6 chanx_right_in[2]
port 62 nsew default input
rlabel metal3 s 27520 1912 28000 2032 6 chanx_right_in[3]
port 63 nsew default input
rlabel metal3 s 27520 2592 28000 2712 6 chanx_right_in[4]
port 64 nsew default input
rlabel metal3 s 27520 3136 28000 3256 6 chanx_right_in[5]
port 65 nsew default input
rlabel metal3 s 27520 3680 28000 3800 6 chanx_right_in[6]
port 66 nsew default input
rlabel metal3 s 27520 4360 28000 4480 6 chanx_right_in[7]
port 67 nsew default input
rlabel metal3 s 27520 4904 28000 5024 6 chanx_right_in[8]
port 68 nsew default input
rlabel metal3 s 27520 5448 28000 5568 6 chanx_right_in[9]
port 69 nsew default input
rlabel metal3 s 27520 11840 28000 11960 6 chanx_right_out[0]
port 70 nsew default tristate
rlabel metal3 s 27520 17688 28000 17808 6 chanx_right_out[10]
port 71 nsew default tristate
rlabel metal3 s 27520 18368 28000 18488 6 chanx_right_out[11]
port 72 nsew default tristate
rlabel metal3 s 27520 18912 28000 19032 6 chanx_right_out[12]
port 73 nsew default tristate
rlabel metal3 s 27520 19456 28000 19576 6 chanx_right_out[13]
port 74 nsew default tristate
rlabel metal3 s 27520 20000 28000 20120 6 chanx_right_out[14]
port 75 nsew default tristate
rlabel metal3 s 27520 20680 28000 20800 6 chanx_right_out[15]
port 76 nsew default tristate
rlabel metal3 s 27520 21224 28000 21344 6 chanx_right_out[16]
port 77 nsew default tristate
rlabel metal3 s 27520 21768 28000 21888 6 chanx_right_out[17]
port 78 nsew default tristate
rlabel metal3 s 27520 22448 28000 22568 6 chanx_right_out[18]
port 79 nsew default tristate
rlabel metal3 s 27520 22992 28000 23112 6 chanx_right_out[19]
port 80 nsew default tristate
rlabel metal3 s 27520 12520 28000 12640 6 chanx_right_out[1]
port 81 nsew default tristate
rlabel metal3 s 27520 13064 28000 13184 6 chanx_right_out[2]
port 82 nsew default tristate
rlabel metal3 s 27520 13608 28000 13728 6 chanx_right_out[3]
port 83 nsew default tristate
rlabel metal3 s 27520 14288 28000 14408 6 chanx_right_out[4]
port 84 nsew default tristate
rlabel metal3 s 27520 14832 28000 14952 6 chanx_right_out[5]
port 85 nsew default tristate
rlabel metal3 s 27520 15376 28000 15496 6 chanx_right_out[6]
port 86 nsew default tristate
rlabel metal3 s 27520 15920 28000 16040 6 chanx_right_out[7]
port 87 nsew default tristate
rlabel metal3 s 27520 16600 28000 16720 6 chanx_right_out[8]
port 88 nsew default tristate
rlabel metal3 s 27520 17144 28000 17264 6 chanx_right_out[9]
port 89 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_in[0]
port 90 nsew default input
rlabel metal2 s 11702 0 11758 480 6 chany_bottom_in[10]
port 91 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[11]
port 92 nsew default input
rlabel metal2 s 12806 0 12862 480 6 chany_bottom_in[12]
port 93 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 94 nsew default input
rlabel metal2 s 13910 0 13966 480 6 chany_bottom_in[14]
port 95 nsew default input
rlabel metal2 s 14370 0 14426 480 6 chany_bottom_in[15]
port 96 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[16]
port 97 nsew default input
rlabel metal2 s 15474 0 15530 480 6 chany_bottom_in[17]
port 98 nsew default input
rlabel metal2 s 16026 0 16082 480 6 chany_bottom_in[18]
port 99 nsew default input
rlabel metal2 s 16578 0 16634 480 6 chany_bottom_in[19]
port 100 nsew default input
rlabel metal2 s 6734 0 6790 480 6 chany_bottom_in[1]
port 101 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[2]
port 102 nsew default input
rlabel metal2 s 7838 0 7894 480 6 chany_bottom_in[3]
port 103 nsew default input
rlabel metal2 s 8390 0 8446 480 6 chany_bottom_in[4]
port 104 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[5]
port 105 nsew default input
rlabel metal2 s 9494 0 9550 480 6 chany_bottom_in[6]
port 106 nsew default input
rlabel metal2 s 10046 0 10102 480 6 chany_bottom_in[7]
port 107 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[8]
port 108 nsew default input
rlabel metal2 s 11150 0 11206 480 6 chany_bottom_in[9]
port 109 nsew default input
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[0]
port 110 nsew default tristate
rlabel metal2 s 22650 0 22706 480 6 chany_bottom_out[10]
port 111 nsew default tristate
rlabel metal2 s 23202 0 23258 480 6 chany_bottom_out[11]
port 112 nsew default tristate
rlabel metal2 s 23754 0 23810 480 6 chany_bottom_out[12]
port 113 nsew default tristate
rlabel metal2 s 24306 0 24362 480 6 chany_bottom_out[13]
port 114 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 chany_bottom_out[14]
port 115 nsew default tristate
rlabel metal2 s 25410 0 25466 480 6 chany_bottom_out[15]
port 116 nsew default tristate
rlabel metal2 s 25962 0 26018 480 6 chany_bottom_out[16]
port 117 nsew default tristate
rlabel metal2 s 26514 0 26570 480 6 chany_bottom_out[17]
port 118 nsew default tristate
rlabel metal2 s 27066 0 27122 480 6 chany_bottom_out[18]
port 119 nsew default tristate
rlabel metal2 s 27618 0 27674 480 6 chany_bottom_out[19]
port 120 nsew default tristate
rlabel metal2 s 17682 0 17738 480 6 chany_bottom_out[1]
port 121 nsew default tristate
rlabel metal2 s 18234 0 18290 480 6 chany_bottom_out[2]
port 122 nsew default tristate
rlabel metal2 s 18786 0 18842 480 6 chany_bottom_out[3]
port 123 nsew default tristate
rlabel metal2 s 19338 0 19394 480 6 chany_bottom_out[4]
port 124 nsew default tristate
rlabel metal2 s 19890 0 19946 480 6 chany_bottom_out[5]
port 125 nsew default tristate
rlabel metal2 s 20442 0 20498 480 6 chany_bottom_out[6]
port 126 nsew default tristate
rlabel metal2 s 20994 0 21050 480 6 chany_bottom_out[7]
port 127 nsew default tristate
rlabel metal2 s 21546 0 21602 480 6 chany_bottom_out[8]
port 128 nsew default tristate
rlabel metal2 s 22098 0 22154 480 6 chany_bottom_out[9]
port 129 nsew default tristate
rlabel metal2 s 4894 27520 4950 28000 6 chany_top_in[0]
port 130 nsew default input
rlabel metal2 s 10782 27520 10838 28000 6 chany_top_in[10]
port 131 nsew default input
rlabel metal2 s 11334 27520 11390 28000 6 chany_top_in[11]
port 132 nsew default input
rlabel metal2 s 11886 27520 11942 28000 6 chany_top_in[12]
port 133 nsew default input
rlabel metal2 s 12530 27520 12586 28000 6 chany_top_in[13]
port 134 nsew default input
rlabel metal2 s 13082 27520 13138 28000 6 chany_top_in[14]
port 135 nsew default input
rlabel metal2 s 13634 27520 13690 28000 6 chany_top_in[15]
port 136 nsew default input
rlabel metal2 s 14278 27520 14334 28000 6 chany_top_in[16]
port 137 nsew default input
rlabel metal2 s 14830 27520 14886 28000 6 chany_top_in[17]
port 138 nsew default input
rlabel metal2 s 15382 27520 15438 28000 6 chany_top_in[18]
port 139 nsew default input
rlabel metal2 s 16026 27520 16082 28000 6 chany_top_in[19]
port 140 nsew default input
rlabel metal2 s 5538 27520 5594 28000 6 chany_top_in[1]
port 141 nsew default input
rlabel metal2 s 6090 27520 6146 28000 6 chany_top_in[2]
port 142 nsew default input
rlabel metal2 s 6642 27520 6698 28000 6 chany_top_in[3]
port 143 nsew default input
rlabel metal2 s 7286 27520 7342 28000 6 chany_top_in[4]
port 144 nsew default input
rlabel metal2 s 7838 27520 7894 28000 6 chany_top_in[5]
port 145 nsew default input
rlabel metal2 s 8390 27520 8446 28000 6 chany_top_in[6]
port 146 nsew default input
rlabel metal2 s 9034 27520 9090 28000 6 chany_top_in[7]
port 147 nsew default input
rlabel metal2 s 9586 27520 9642 28000 6 chany_top_in[8]
port 148 nsew default input
rlabel metal2 s 10138 27520 10194 28000 6 chany_top_in[9]
port 149 nsew default input
rlabel metal2 s 16578 27520 16634 28000 6 chany_top_out[0]
port 150 nsew default tristate
rlabel metal2 s 22374 27520 22430 28000 6 chany_top_out[10]
port 151 nsew default tristate
rlabel metal2 s 23018 27520 23074 28000 6 chany_top_out[11]
port 152 nsew default tristate
rlabel metal2 s 23570 27520 23626 28000 6 chany_top_out[12]
port 153 nsew default tristate
rlabel metal2 s 24122 27520 24178 28000 6 chany_top_out[13]
port 154 nsew default tristate
rlabel metal2 s 24766 27520 24822 28000 6 chany_top_out[14]
port 155 nsew default tristate
rlabel metal2 s 25318 27520 25374 28000 6 chany_top_out[15]
port 156 nsew default tristate
rlabel metal2 s 25870 27520 25926 28000 6 chany_top_out[16]
port 157 nsew default tristate
rlabel metal2 s 26514 27520 26570 28000 6 chany_top_out[17]
port 158 nsew default tristate
rlabel metal2 s 27066 27520 27122 28000 6 chany_top_out[18]
port 159 nsew default tristate
rlabel metal2 s 27618 27520 27674 28000 6 chany_top_out[19]
port 160 nsew default tristate
rlabel metal2 s 17130 27520 17186 28000 6 chany_top_out[1]
port 161 nsew default tristate
rlabel metal2 s 17774 27520 17830 28000 6 chany_top_out[2]
port 162 nsew default tristate
rlabel metal2 s 18326 27520 18382 28000 6 chany_top_out[3]
port 163 nsew default tristate
rlabel metal2 s 18878 27520 18934 28000 6 chany_top_out[4]
port 164 nsew default tristate
rlabel metal2 s 19522 27520 19578 28000 6 chany_top_out[5]
port 165 nsew default tristate
rlabel metal2 s 20074 27520 20130 28000 6 chany_top_out[6]
port 166 nsew default tristate
rlabel metal2 s 20626 27520 20682 28000 6 chany_top_out[7]
port 167 nsew default tristate
rlabel metal2 s 21270 27520 21326 28000 6 chany_top_out[8]
port 168 nsew default tristate
rlabel metal2 s 21822 27520 21878 28000 6 chany_top_out[9]
port 169 nsew default tristate
rlabel metal3 s 0 23536 480 23656 6 left_top_grid_pin_42_
port 170 nsew default input
rlabel metal3 s 0 24080 480 24200 6 left_top_grid_pin_43_
port 171 nsew default input
rlabel metal3 s 0 24760 480 24880 6 left_top_grid_pin_44_
port 172 nsew default input
rlabel metal3 s 0 25304 480 25424 6 left_top_grid_pin_45_
port 173 nsew default input
rlabel metal3 s 0 25848 480 25968 6 left_top_grid_pin_46_
port 174 nsew default input
rlabel metal3 s 0 26528 480 26648 6 left_top_grid_pin_47_
port 175 nsew default input
rlabel metal3 s 0 27072 480 27192 6 left_top_grid_pin_48_
port 176 nsew default input
rlabel metal3 s 0 27616 480 27736 6 left_top_grid_pin_49_
port 177 nsew default input
rlabel metal2 s 4526 0 4582 480 6 prog_clk
port 178 nsew default input
rlabel metal3 s 27520 23536 28000 23656 6 right_top_grid_pin_42_
port 179 nsew default input
rlabel metal3 s 27520 24080 28000 24200 6 right_top_grid_pin_43_
port 180 nsew default input
rlabel metal3 s 27520 24760 28000 24880 6 right_top_grid_pin_44_
port 181 nsew default input
rlabel metal3 s 27520 25304 28000 25424 6 right_top_grid_pin_45_
port 182 nsew default input
rlabel metal3 s 27520 25848 28000 25968 6 right_top_grid_pin_46_
port 183 nsew default input
rlabel metal3 s 27520 26528 28000 26648 6 right_top_grid_pin_47_
port 184 nsew default input
rlabel metal3 s 27520 27072 28000 27192 6 right_top_grid_pin_48_
port 185 nsew default input
rlabel metal3 s 27520 27616 28000 27736 6 right_top_grid_pin_49_
port 186 nsew default input
rlabel metal2 s 294 27520 350 28000 6 top_left_grid_pin_34_
port 187 nsew default input
rlabel metal2 s 846 27520 902 28000 6 top_left_grid_pin_35_
port 188 nsew default input
rlabel metal2 s 1398 27520 1454 28000 6 top_left_grid_pin_36_
port 189 nsew default input
rlabel metal2 s 2042 27520 2098 28000 6 top_left_grid_pin_37_
port 190 nsew default input
rlabel metal2 s 2594 27520 2650 28000 6 top_left_grid_pin_38_
port 191 nsew default input
rlabel metal2 s 3146 27520 3202 28000 6 top_left_grid_pin_39_
port 192 nsew default input
rlabel metal2 s 3790 27520 3846 28000 6 top_left_grid_pin_40_
port 193 nsew default input
rlabel metal2 s 4342 27520 4398 28000 6 top_left_grid_pin_41_
port 194 nsew default input
rlabel metal4 s 5611 2128 5931 25616 6 VPWR
port 195 nsew default input
rlabel metal4 s 10277 2128 10597 25616 6 VGND
port 196 nsew default input
<< properties >>
string FIXED_BBOX 0 0 28000 28000
<< end >>
