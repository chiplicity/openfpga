magic
tech sky130A
magscale 1 2
timestamp 1605013774
<< locali >>
rect 6469 20247 6503 20417
rect 2697 13311 2731 13481
rect 2237 5695 2271 5865
<< viali >>
rect 7021 21097 7055 21131
rect 21097 21097 21131 21131
rect 20913 20961 20947 20995
rect 23673 20757 23707 20791
rect 1869 20553 1903 20587
rect 20821 20553 20855 20587
rect 21373 20553 21407 20587
rect 26617 20553 26651 20587
rect 6469 20417 6503 20451
rect 7389 20417 7423 20451
rect 16957 20417 16991 20451
rect 23673 20417 23707 20451
rect 1685 20349 1719 20383
rect 2973 20349 3007 20383
rect 2881 20281 2915 20315
rect 3218 20281 3252 20315
rect 6285 20281 6319 20315
rect 8493 20349 8527 20383
rect 13921 20349 13955 20383
rect 16681 20349 16715 20383
rect 17417 20349 17451 20383
rect 19441 20349 19475 20383
rect 26433 20349 26467 20383
rect 26985 20349 27019 20383
rect 7205 20281 7239 20315
rect 8738 20281 8772 20315
rect 13829 20281 13863 20315
rect 14166 20281 14200 20315
rect 19349 20281 19383 20315
rect 19708 20281 19742 20315
rect 23489 20281 23523 20315
rect 23918 20281 23952 20315
rect 2329 20213 2363 20247
rect 4353 20213 4387 20247
rect 6469 20213 6503 20247
rect 6561 20213 6595 20247
rect 6837 20213 6871 20247
rect 7297 20213 7331 20247
rect 8401 20213 8435 20247
rect 9873 20213 9907 20247
rect 15301 20213 15335 20247
rect 25053 20213 25087 20247
rect 6009 20009 6043 20043
rect 6929 20009 6963 20043
rect 7113 20009 7147 20043
rect 8493 20009 8527 20043
rect 13921 20009 13955 20043
rect 19441 20009 19475 20043
rect 23213 20009 23247 20043
rect 24501 20009 24535 20043
rect 24961 20009 24995 20043
rect 26525 20009 26559 20043
rect 26985 20009 27019 20043
rect 10876 19941 10910 19975
rect 4896 19873 4930 19907
rect 7481 19873 7515 19907
rect 10609 19873 10643 19907
rect 16497 19873 16531 19907
rect 22100 19873 22134 19907
rect 26893 19873 26927 19907
rect 4629 19805 4663 19839
rect 7573 19805 7607 19839
rect 7757 19805 7791 19839
rect 16589 19805 16623 19839
rect 16681 19805 16715 19839
rect 17693 19805 17727 19839
rect 21833 19805 21867 19839
rect 25053 19805 25087 19839
rect 25145 19805 25179 19839
rect 27077 19805 27111 19839
rect 3065 19669 3099 19703
rect 11989 19669 12023 19703
rect 15669 19669 15703 19703
rect 16129 19669 16163 19703
rect 23857 19669 23891 19703
rect 24593 19669 24627 19703
rect 10701 19465 10735 19499
rect 14473 19465 14507 19499
rect 17049 19465 17083 19499
rect 23397 19465 23431 19499
rect 24961 19465 24995 19499
rect 25513 19465 25547 19499
rect 26893 19465 26927 19499
rect 7389 19397 7423 19431
rect 10977 19397 11011 19431
rect 26617 19397 26651 19431
rect 8033 19329 8067 19363
rect 16037 19329 16071 19363
rect 16129 19329 16163 19363
rect 24133 19329 24167 19363
rect 24225 19329 24259 19363
rect 26065 19329 26099 19363
rect 27261 19329 27295 19363
rect 6285 19261 6319 19295
rect 8769 19261 8803 19295
rect 13093 19261 13127 19295
rect 15117 19261 15151 19295
rect 15945 19261 15979 19295
rect 23121 19261 23155 19295
rect 24041 19261 24075 19295
rect 4997 19193 5031 19227
rect 6653 19193 6687 19227
rect 7757 19193 7791 19227
rect 8953 19193 8987 19227
rect 13001 19193 13035 19227
rect 13338 19193 13372 19227
rect 15393 19193 15427 19227
rect 21925 19193 21959 19227
rect 22293 19193 22327 19227
rect 25973 19193 26007 19227
rect 4445 19125 4479 19159
rect 5365 19125 5399 19159
rect 7205 19125 7239 19159
rect 7849 19125 7883 19159
rect 8493 19125 8527 19159
rect 15577 19125 15611 19159
rect 16681 19125 16715 19159
rect 20361 19125 20395 19159
rect 23673 19125 23707 19159
rect 25329 19125 25363 19159
rect 25881 19125 25915 19159
rect 7389 18921 7423 18955
rect 13093 18921 13127 18955
rect 14013 18921 14047 18955
rect 16037 18921 16071 18955
rect 23397 18921 23431 18955
rect 25053 18921 25087 18955
rect 26525 18921 26559 18955
rect 7205 18853 7239 18887
rect 10968 18853 11002 18887
rect 1409 18785 1443 18819
rect 4721 18785 4755 18819
rect 7757 18785 7791 18819
rect 10701 18785 10735 18819
rect 16405 18785 16439 18819
rect 18501 18785 18535 18819
rect 21281 18785 21315 18819
rect 21373 18785 21407 18819
rect 23765 18785 23799 18819
rect 4813 18717 4847 18751
rect 4997 18717 5031 18751
rect 7849 18717 7883 18751
rect 8033 18717 8067 18751
rect 14105 18717 14139 18751
rect 14289 18717 14323 18751
rect 16497 18717 16531 18751
rect 16589 18717 16623 18751
rect 18245 18717 18279 18751
rect 21465 18717 21499 18751
rect 23857 18717 23891 18751
rect 23949 18717 23983 18751
rect 24593 18717 24627 18751
rect 1593 18581 1627 18615
rect 2053 18581 2087 18615
rect 2329 18581 2363 18615
rect 3893 18581 3927 18615
rect 4353 18581 4387 18615
rect 8769 18581 8803 18615
rect 9045 18581 9079 18615
rect 12081 18581 12115 18615
rect 13645 18581 13679 18615
rect 15025 18581 15059 18615
rect 15577 18581 15611 18615
rect 19625 18581 19659 18615
rect 20269 18581 20303 18615
rect 20913 18581 20947 18615
rect 25605 18581 25639 18615
rect 3801 18377 3835 18411
rect 4169 18377 4203 18411
rect 7113 18377 7147 18411
rect 8125 18377 8159 18411
rect 11069 18377 11103 18411
rect 14933 18377 14967 18411
rect 16037 18377 16071 18411
rect 16497 18377 16531 18411
rect 18705 18377 18739 18411
rect 21281 18377 21315 18411
rect 22753 18377 22787 18411
rect 23765 18377 23799 18411
rect 27537 18377 27571 18411
rect 3065 18309 3099 18343
rect 6653 18309 6687 18343
rect 10793 18309 10827 18343
rect 14381 18309 14415 18343
rect 14749 18309 14783 18343
rect 21649 18309 21683 18343
rect 23029 18309 23063 18343
rect 4813 18241 4847 18275
rect 5641 18241 5675 18275
rect 6285 18241 6319 18275
rect 7757 18241 7791 18275
rect 8585 18241 8619 18275
rect 9321 18241 9355 18275
rect 15393 18241 15427 18275
rect 15485 18241 15519 18275
rect 16773 18241 16807 18275
rect 20821 18241 20855 18275
rect 24409 18241 24443 18275
rect 1685 18173 1719 18207
rect 4629 18173 4663 18207
rect 9045 18173 9079 18207
rect 12449 18173 12483 18207
rect 20085 18173 20119 18207
rect 20637 18173 20671 18207
rect 22017 18173 22051 18207
rect 26157 18173 26191 18207
rect 1952 18105 1986 18139
rect 7573 18105 7607 18139
rect 12265 18105 12299 18139
rect 12694 18105 12728 18139
rect 20729 18105 20763 18139
rect 26402 18105 26436 18139
rect 4261 18037 4295 18071
rect 4721 18037 4755 18071
rect 5273 18037 5307 18071
rect 7481 18037 7515 18071
rect 8677 18037 8711 18071
rect 9137 18037 9171 18071
rect 13829 18037 13863 18071
rect 15301 18037 15335 18071
rect 18337 18037 18371 18071
rect 20269 18037 20303 18071
rect 23489 18037 23523 18071
rect 24133 18037 24167 18071
rect 24225 18037 24259 18071
rect 24777 18037 24811 18071
rect 25973 18037 26007 18071
rect 2053 17833 2087 17867
rect 3893 17833 3927 17867
rect 4353 17833 4387 17867
rect 4721 17833 4755 17867
rect 7113 17833 7147 17867
rect 8033 17833 8067 17867
rect 9689 17833 9723 17867
rect 12449 17833 12483 17867
rect 13737 17833 13771 17867
rect 14105 17833 14139 17867
rect 14749 17833 14783 17867
rect 15301 17833 15335 17867
rect 20361 17833 20395 17867
rect 21281 17833 21315 17867
rect 23489 17833 23523 17867
rect 23949 17833 23983 17867
rect 26249 17833 26283 17867
rect 7849 17765 7883 17799
rect 17233 17765 17267 17799
rect 23765 17765 23799 17799
rect 1409 17697 1443 17731
rect 4813 17697 4847 17731
rect 7481 17697 7515 17731
rect 8401 17697 8435 17731
rect 10057 17697 10091 17731
rect 15669 17697 15703 17731
rect 20729 17697 20763 17731
rect 24317 17697 24351 17731
rect 26525 17697 26559 17731
rect 2421 17629 2455 17663
rect 4905 17629 4939 17663
rect 8493 17629 8527 17663
rect 8585 17629 8619 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 15117 17629 15151 17663
rect 15761 17629 15795 17663
rect 15853 17629 15887 17663
rect 17325 17629 17359 17663
rect 17417 17629 17451 17663
rect 21373 17629 21407 17663
rect 21465 17629 21499 17663
rect 24409 17629 24443 17663
rect 24593 17629 24627 17663
rect 9137 17561 9171 17595
rect 1593 17493 1627 17527
rect 2697 17493 2731 17527
rect 5365 17493 5399 17527
rect 16865 17493 16899 17527
rect 18521 17493 18555 17527
rect 20913 17493 20947 17527
rect 25053 17493 25087 17527
rect 26709 17493 26743 17527
rect 1685 17289 1719 17323
rect 4077 17289 4111 17323
rect 7757 17289 7791 17323
rect 9045 17289 9079 17323
rect 10793 17289 10827 17323
rect 14565 17289 14599 17323
rect 14933 17289 14967 17323
rect 15117 17289 15151 17323
rect 16129 17289 16163 17323
rect 18245 17289 18279 17323
rect 20177 17289 20211 17323
rect 22569 17289 22603 17323
rect 26525 17289 26559 17323
rect 1869 17221 1903 17255
rect 23121 17221 23155 17255
rect 24501 17221 24535 17255
rect 2421 17153 2455 17187
rect 4445 17153 4479 17187
rect 5273 17153 5307 17187
rect 5457 17153 5491 17187
rect 5825 17153 5859 17187
rect 8493 17153 8527 17187
rect 9689 17153 9723 17187
rect 15669 17153 15703 17187
rect 17877 17153 17911 17187
rect 19073 17153 19107 17187
rect 20637 17153 20671 17187
rect 25053 17153 25087 17187
rect 2237 17085 2271 17119
rect 5181 17085 5215 17119
rect 6285 17085 6319 17119
rect 14289 17085 14323 17119
rect 15577 17085 15611 17119
rect 18797 17085 18831 17119
rect 18889 17085 18923 17119
rect 24041 17085 24075 17119
rect 9505 17017 9539 17051
rect 16957 17017 16991 17051
rect 20882 17017 20916 17051
rect 23489 17017 23523 17051
rect 24961 17017 24995 17051
rect 2329 16949 2363 16983
rect 2881 16949 2915 16983
rect 4813 16949 4847 16983
rect 8033 16949 8067 16983
rect 8861 16949 8895 16983
rect 9413 16949 9447 16983
rect 10057 16949 10091 16983
rect 10425 16949 10459 16983
rect 15485 16949 15519 16983
rect 16589 16949 16623 16983
rect 17325 16949 17359 16983
rect 18429 16949 18463 16983
rect 20453 16949 20487 16983
rect 22017 16949 22051 16983
rect 24317 16949 24351 16983
rect 24869 16949 24903 16983
rect 1869 16745 1903 16779
rect 2329 16745 2363 16779
rect 6193 16745 6227 16779
rect 9689 16745 9723 16779
rect 13737 16745 13771 16779
rect 15117 16745 15151 16779
rect 18429 16745 18463 16779
rect 20913 16745 20947 16779
rect 21281 16745 21315 16779
rect 24041 16745 24075 16779
rect 24501 16745 24535 16779
rect 1777 16677 1811 16711
rect 5080 16677 5114 16711
rect 10057 16677 10091 16711
rect 15945 16677 15979 16711
rect 20637 16677 20671 16711
rect 24869 16677 24903 16711
rect 2237 16609 2271 16643
rect 2973 16609 3007 16643
rect 4353 16609 4387 16643
rect 9137 16609 9171 16643
rect 12357 16609 12391 16643
rect 12624 16609 12658 16643
rect 15853 16609 15887 16643
rect 18797 16609 18831 16643
rect 21373 16609 21407 16643
rect 24961 16609 24995 16643
rect 2513 16541 2547 16575
rect 4813 16541 4847 16575
rect 10149 16541 10183 16575
rect 10333 16541 10367 16575
rect 16037 16541 16071 16575
rect 18889 16541 18923 16575
rect 18981 16541 19015 16575
rect 21557 16541 21591 16575
rect 25053 16541 25087 16575
rect 15485 16473 15519 16507
rect 24409 16405 24443 16439
rect 1869 16201 1903 16235
rect 3617 16201 3651 16235
rect 4905 16201 4939 16235
rect 6561 16201 6595 16235
rect 9413 16201 9447 16235
rect 12265 16201 12299 16235
rect 13829 16201 13863 16235
rect 15485 16201 15519 16235
rect 16589 16201 16623 16235
rect 17877 16201 17911 16235
rect 18429 16201 18463 16235
rect 19809 16201 19843 16235
rect 20177 16201 20211 16235
rect 21649 16201 21683 16235
rect 24317 16201 24351 16235
rect 25329 16201 25363 16235
rect 27261 16201 27295 16235
rect 9873 16133 9907 16167
rect 21373 16133 21407 16167
rect 2237 16065 2271 16099
rect 11529 16065 11563 16099
rect 12449 16065 12483 16099
rect 16129 16065 16163 16099
rect 16865 16065 16899 16099
rect 17233 16065 17267 16099
rect 19073 16065 19107 16099
rect 21005 16065 21039 16099
rect 23489 16065 23523 16099
rect 24961 16065 24995 16099
rect 25881 16065 25915 16099
rect 5273 15997 5307 16031
rect 6837 15997 6871 16031
rect 7093 15997 7127 16031
rect 10057 15997 10091 16031
rect 10701 15997 10735 16031
rect 14657 15997 14691 16031
rect 15853 15997 15887 16031
rect 2504 15929 2538 15963
rect 11897 15929 11931 15963
rect 12694 15929 12728 15963
rect 15393 15929 15427 15963
rect 15945 15929 15979 15963
rect 24777 15929 24811 15963
rect 26126 15929 26160 15963
rect 8217 15861 8251 15895
rect 9781 15861 9815 15895
rect 10333 15861 10367 15895
rect 14933 15861 14967 15895
rect 18337 15861 18371 15895
rect 18797 15861 18831 15895
rect 18889 15861 18923 15895
rect 19441 15861 19475 15895
rect 24133 15861 24167 15895
rect 24685 15861 24719 15895
rect 25697 15861 25731 15895
rect 1777 15657 1811 15691
rect 11069 15657 11103 15691
rect 12817 15657 12851 15691
rect 18889 15657 18923 15691
rect 24961 15657 24995 15691
rect 25973 15657 26007 15691
rect 2145 15589 2179 15623
rect 15546 15589 15580 15623
rect 19349 15589 19383 15623
rect 22262 15589 22296 15623
rect 1685 15521 1719 15555
rect 7297 15521 7331 15555
rect 9689 15521 9723 15555
rect 9956 15521 9990 15555
rect 19257 15521 19291 15555
rect 22017 15521 22051 15555
rect 26525 15521 26559 15555
rect 2237 15453 2271 15487
rect 2421 15453 2455 15487
rect 15301 15453 15335 15487
rect 19533 15453 19567 15487
rect 2789 15317 2823 15351
rect 6929 15317 6963 15351
rect 7113 15317 7147 15351
rect 12541 15317 12575 15351
rect 16681 15317 16715 15351
rect 18521 15317 18555 15351
rect 23397 15317 23431 15351
rect 24593 15317 24627 15351
rect 26709 15317 26743 15351
rect 3065 15113 3099 15147
rect 7205 15113 7239 15147
rect 10057 15113 10091 15147
rect 12173 15113 12207 15147
rect 15209 15113 15243 15147
rect 18613 15113 18647 15147
rect 18797 15113 18831 15147
rect 19349 15113 19383 15147
rect 20913 15113 20947 15147
rect 22017 15113 22051 15147
rect 26525 15113 26559 15147
rect 2053 15045 2087 15079
rect 3433 15045 3467 15079
rect 14473 15045 14507 15079
rect 2697 14977 2731 15011
rect 13001 14977 13035 15011
rect 14841 14977 14875 15011
rect 16313 14977 16347 15011
rect 7665 14909 7699 14943
rect 7932 14909 7966 14943
rect 9781 14909 9815 14943
rect 12817 14909 12851 14943
rect 16037 14909 16071 14943
rect 18337 14909 18371 14943
rect 18981 14909 19015 14943
rect 19533 14909 19567 14943
rect 2421 14841 2455 14875
rect 7573 14841 7607 14875
rect 15577 14841 15611 14875
rect 19778 14841 19812 14875
rect 1961 14773 1995 14807
rect 2513 14773 2547 14807
rect 9045 14773 9079 14807
rect 11621 14773 11655 14807
rect 12449 14773 12483 14807
rect 12909 14773 12943 14807
rect 15669 14773 15703 14807
rect 16129 14773 16163 14807
rect 22477 14773 22511 14807
rect 2237 14569 2271 14603
rect 2605 14569 2639 14603
rect 6377 14569 6411 14603
rect 8309 14569 8343 14603
rect 8861 14569 8895 14603
rect 11897 14569 11931 14603
rect 17509 14569 17543 14603
rect 19993 14569 20027 14603
rect 20545 14569 20579 14603
rect 1869 14501 1903 14535
rect 5264 14501 5298 14535
rect 2973 14433 3007 14467
rect 4997 14433 5031 14467
rect 9045 14433 9079 14467
rect 13461 14433 13495 14467
rect 16129 14433 16163 14467
rect 16396 14433 16430 14467
rect 20729 14433 20763 14467
rect 21465 14433 21499 14467
rect 21732 14433 21766 14467
rect 24205 14433 24239 14467
rect 11437 14365 11471 14399
rect 11989 14365 12023 14399
rect 12173 14365 12207 14399
rect 13553 14365 13587 14399
rect 13645 14365 13679 14399
rect 23949 14365 23983 14399
rect 4445 14229 4479 14263
rect 7757 14229 7791 14263
rect 10885 14229 10919 14263
rect 11529 14229 11563 14263
rect 12633 14229 12667 14263
rect 13001 14229 13035 14263
rect 13093 14229 13127 14263
rect 15669 14229 15703 14263
rect 18981 14229 19015 14263
rect 19625 14229 19659 14263
rect 22845 14229 22879 14263
rect 25329 14229 25363 14263
rect 5825 14025 5859 14059
rect 10793 14025 10827 14059
rect 12449 14025 12483 14059
rect 18797 14025 18831 14059
rect 20637 14025 20671 14059
rect 21833 14025 21867 14059
rect 3249 13957 3283 13991
rect 8217 13957 8251 13991
rect 10701 13957 10735 13991
rect 12173 13957 12207 13991
rect 21557 13957 21591 13991
rect 27445 13957 27479 13991
rect 4905 13889 4939 13923
rect 8769 13889 8803 13923
rect 11437 13889 11471 13923
rect 11897 13889 11931 13923
rect 12909 13889 12943 13923
rect 13001 13889 13035 13923
rect 14933 13889 14967 13923
rect 16405 13889 16439 13923
rect 19165 13889 19199 13923
rect 24409 13889 24443 13923
rect 26065 13889 26099 13923
rect 1869 13821 1903 13855
rect 3893 13821 3927 13855
rect 5457 13821 5491 13855
rect 7757 13821 7791 13855
rect 8677 13821 8711 13855
rect 11253 13821 11287 13855
rect 12817 13821 12851 13855
rect 13829 13821 13863 13855
rect 15577 13821 15611 13855
rect 16221 13821 16255 13855
rect 19257 13821 19291 13855
rect 19524 13821 19558 13855
rect 23949 13821 23983 13855
rect 26321 13821 26355 13855
rect 2114 13753 2148 13787
rect 4261 13753 4295 13787
rect 4721 13753 4755 13787
rect 9229 13753 9263 13787
rect 11161 13753 11195 13787
rect 15301 13753 15335 13787
rect 16129 13753 16163 13787
rect 1777 13685 1811 13719
rect 4353 13685 4387 13719
rect 4813 13685 4847 13719
rect 8125 13685 8159 13719
rect 8585 13685 8619 13719
rect 13461 13685 13495 13719
rect 15761 13685 15795 13719
rect 16865 13685 16899 13719
rect 25881 13685 25915 13719
rect 1777 13481 1811 13515
rect 2697 13481 2731 13515
rect 2881 13481 2915 13515
rect 4629 13481 4663 13515
rect 7481 13481 7515 13515
rect 10793 13481 10827 13515
rect 11253 13481 11287 13515
rect 12449 13481 12483 13515
rect 12817 13481 12851 13515
rect 15117 13481 15151 13515
rect 15669 13481 15703 13515
rect 16865 13481 16899 13515
rect 19717 13481 19751 13515
rect 20545 13481 20579 13515
rect 26065 13481 26099 13515
rect 2329 13413 2363 13447
rect 2237 13345 2271 13379
rect 15761 13413 15795 13447
rect 16405 13413 16439 13447
rect 19533 13413 19567 13447
rect 7849 13345 7883 13379
rect 7941 13345 7975 13379
rect 11621 13345 11655 13379
rect 17233 13345 17267 13379
rect 19901 13345 19935 13379
rect 22753 13345 22787 13379
rect 2513 13277 2547 13311
rect 2697 13277 2731 13311
rect 4721 13277 4755 13311
rect 4813 13277 4847 13311
rect 8125 13277 8159 13311
rect 11713 13277 11747 13311
rect 11897 13277 11931 13311
rect 13277 13277 13311 13311
rect 15945 13277 15979 13311
rect 17325 13277 17359 13311
rect 17509 13277 17543 13311
rect 22845 13277 22879 13311
rect 23029 13277 23063 13311
rect 1869 13141 1903 13175
rect 3801 13141 3835 13175
rect 4261 13141 4295 13175
rect 15301 13141 15335 13175
rect 22385 13141 22419 13175
rect 24225 13141 24259 13175
rect 25789 13141 25823 13175
rect 2973 12937 3007 12971
rect 4721 12937 4755 12971
rect 5089 12937 5123 12971
rect 7573 12937 7607 12971
rect 7849 12937 7883 12971
rect 12081 12937 12115 12971
rect 16313 12937 16347 12971
rect 17601 12937 17635 12971
rect 22385 12937 22419 12971
rect 23213 12937 23247 12971
rect 7205 12869 7239 12903
rect 22845 12869 22879 12903
rect 24133 12869 24167 12903
rect 1777 12801 1811 12835
rect 2329 12801 2363 12835
rect 2513 12801 2547 12835
rect 4261 12801 4295 12835
rect 14381 12801 14415 12835
rect 15669 12801 15703 12835
rect 15853 12801 15887 12835
rect 18981 12801 19015 12835
rect 19533 12801 19567 12835
rect 24041 12801 24075 12835
rect 24685 12801 24719 12835
rect 25513 12801 25547 12835
rect 26249 12801 26283 12835
rect 2237 12733 2271 12767
rect 4077 12733 4111 12767
rect 5457 12733 5491 12767
rect 8585 12733 8619 12767
rect 11253 12733 11287 12767
rect 11713 12733 11747 12767
rect 19789 12733 19823 12767
rect 24501 12733 24535 12767
rect 26065 12733 26099 12767
rect 8493 12665 8527 12699
rect 8830 12665 8864 12699
rect 15025 12665 15059 12699
rect 15577 12665 15611 12699
rect 16957 12665 16991 12699
rect 1869 12597 1903 12631
rect 3341 12597 3375 12631
rect 3709 12597 3743 12631
rect 4169 12597 4203 12631
rect 9965 12597 9999 12631
rect 14749 12597 14783 12631
rect 15209 12597 15243 12631
rect 17325 12597 17359 12631
rect 19441 12597 19475 12631
rect 20913 12597 20947 12631
rect 24593 12597 24627 12631
rect 25697 12597 25731 12631
rect 26157 12597 26191 12631
rect 27261 12597 27295 12631
rect 2053 12393 2087 12427
rect 3065 12393 3099 12427
rect 4353 12393 4387 12427
rect 7665 12393 7699 12427
rect 8585 12393 8619 12427
rect 15117 12393 15151 12427
rect 23213 12393 23247 12427
rect 24317 12393 24351 12427
rect 24777 12393 24811 12427
rect 26249 12393 26283 12427
rect 14749 12325 14783 12359
rect 15761 12325 15795 12359
rect 26893 12325 26927 12359
rect 2789 12257 2823 12291
rect 6552 12257 6586 12291
rect 11253 12257 11287 12291
rect 15669 12257 15703 12291
rect 16681 12257 16715 12291
rect 18337 12257 18371 12291
rect 18604 12257 18638 12291
rect 20729 12257 20763 12291
rect 21281 12257 21315 12291
rect 23121 12257 23155 12291
rect 24685 12257 24719 12291
rect 26985 12257 27019 12291
rect 2145 12189 2179 12223
rect 2329 12189 2363 12223
rect 4905 12189 4939 12223
rect 4997 12189 5031 12223
rect 6285 12189 6319 12223
rect 11345 12189 11379 12223
rect 11529 12189 11563 12223
rect 15853 12189 15887 12223
rect 21373 12189 21407 12223
rect 21465 12189 21499 12223
rect 23397 12189 23431 12223
rect 24869 12189 24903 12223
rect 27169 12189 27203 12223
rect 1685 12121 1719 12155
rect 19717 12121 19751 12155
rect 22753 12121 22787 12155
rect 24133 12121 24167 12155
rect 25789 12121 25823 12155
rect 26525 12121 26559 12155
rect 3709 12053 3743 12087
rect 8217 12053 8251 12087
rect 10885 12053 10919 12087
rect 15301 12053 15335 12087
rect 16313 12053 16347 12087
rect 18153 12053 18187 12087
rect 20913 12053 20947 12087
rect 22017 12053 22051 12087
rect 7665 11849 7699 11883
rect 9597 11849 9631 11883
rect 13829 11849 13863 11883
rect 15209 11849 15243 11883
rect 19717 11849 19751 11883
rect 21465 11849 21499 11883
rect 22845 11849 22879 11883
rect 24041 11849 24075 11883
rect 25605 11849 25639 11883
rect 26157 11849 26191 11883
rect 9689 11781 9723 11815
rect 25973 11781 26007 11815
rect 27537 11781 27571 11815
rect 5365 11713 5399 11747
rect 8401 11713 8435 11747
rect 10241 11713 10275 11747
rect 11253 11713 11287 11747
rect 11713 11713 11747 11747
rect 16405 11713 16439 11747
rect 17509 11713 17543 11747
rect 18889 11713 18923 11747
rect 20453 11713 20487 11747
rect 21281 11713 21315 11747
rect 22017 11713 22051 11747
rect 24317 11713 24351 11747
rect 25053 11713 25087 11747
rect 26709 11713 26743 11747
rect 1685 11645 1719 11679
rect 5181 11645 5215 11679
rect 6377 11645 6411 11679
rect 8217 11645 8251 11679
rect 10057 11645 10091 11679
rect 13921 11645 13955 11679
rect 16221 11645 16255 11679
rect 17877 11645 17911 11679
rect 20269 11645 20303 11679
rect 21925 11645 21959 11679
rect 24869 11645 24903 11679
rect 26525 11645 26559 11679
rect 1952 11577 1986 11611
rect 3617 11577 3651 11611
rect 4721 11577 4755 11611
rect 5273 11577 5307 11611
rect 8309 11577 8343 11611
rect 9229 11577 9263 11611
rect 10149 11577 10183 11611
rect 16129 11577 16163 11611
rect 18705 11577 18739 11611
rect 21005 11577 21039 11611
rect 21833 11577 21867 11611
rect 24961 11577 24995 11611
rect 26617 11577 26651 11611
rect 3065 11509 3099 11543
rect 4261 11509 4295 11543
rect 4813 11509 4847 11543
rect 5917 11509 5951 11543
rect 7389 11509 7423 11543
rect 7849 11509 7883 11543
rect 10885 11509 10919 11543
rect 12173 11509 12207 11543
rect 15761 11509 15795 11543
rect 16865 11509 16899 11543
rect 18337 11509 18371 11543
rect 18797 11509 18831 11543
rect 19349 11509 19383 11543
rect 19901 11509 19935 11543
rect 20361 11509 20395 11543
rect 23397 11509 23431 11543
rect 24501 11509 24535 11543
rect 27169 11509 27203 11543
rect 2053 11305 2087 11339
rect 2421 11305 2455 11339
rect 2697 11305 2731 11339
rect 4629 11305 4663 11339
rect 7849 11305 7883 11339
rect 9965 11305 9999 11339
rect 10609 11305 10643 11339
rect 18153 11305 18187 11339
rect 19901 11305 19935 11339
rect 20361 11305 20395 11339
rect 20729 11305 20763 11339
rect 21373 11305 21407 11339
rect 22845 11305 22879 11339
rect 23213 11305 23247 11339
rect 24961 11305 24995 11339
rect 25329 11305 25363 11339
rect 26709 11305 26743 11339
rect 3065 11237 3099 11271
rect 16037 11237 16071 11271
rect 18061 11237 18095 11271
rect 21189 11237 21223 11271
rect 24593 11237 24627 11271
rect 1409 11169 1443 11203
rect 2513 11169 2547 11203
rect 6193 11169 6227 11203
rect 7757 11169 7791 11203
rect 8217 11169 8251 11203
rect 10977 11169 11011 11203
rect 13165 11169 13199 11203
rect 15945 11169 15979 11203
rect 18521 11169 18555 11203
rect 21741 11169 21775 11203
rect 26525 11169 26559 11203
rect 4721 11101 4755 11135
rect 4813 11101 4847 11135
rect 6285 11101 6319 11135
rect 6469 11101 6503 11135
rect 8309 11101 8343 11135
rect 8493 11101 8527 11135
rect 11069 11101 11103 11135
rect 11161 11101 11195 11135
rect 12909 11101 12943 11135
rect 16129 11101 16163 11135
rect 16589 11101 16623 11135
rect 18613 11101 18647 11135
rect 18797 11101 18831 11135
rect 21833 11101 21867 11135
rect 22017 11101 22051 11135
rect 1593 11033 1627 11067
rect 5825 11033 5859 11067
rect 15025 11033 15059 11067
rect 26157 11033 26191 11067
rect 4261 10965 4295 10999
rect 5273 10965 5307 10999
rect 8861 10965 8895 10999
rect 14289 10965 14323 10999
rect 15577 10965 15611 10999
rect 19165 10965 19199 10999
rect 23949 10965 23983 10999
rect 1593 10761 1627 10795
rect 6561 10761 6595 10795
rect 8217 10761 8251 10795
rect 13277 10761 13311 10795
rect 15945 10761 15979 10795
rect 16313 10761 16347 10795
rect 18337 10761 18371 10795
rect 21097 10761 21131 10795
rect 22293 10761 22327 10795
rect 27353 10761 27387 10795
rect 3433 10693 3467 10727
rect 5917 10693 5951 10727
rect 9781 10693 9815 10727
rect 13001 10693 13035 10727
rect 14749 10693 14783 10727
rect 19717 10693 19751 10727
rect 21373 10693 21407 10727
rect 4445 10625 4479 10659
rect 5089 10625 5123 10659
rect 8677 10625 8711 10659
rect 8861 10625 8895 10659
rect 10333 10625 10367 10659
rect 15485 10625 15519 10659
rect 16497 10625 16531 10659
rect 17509 10625 17543 10659
rect 18981 10625 19015 10659
rect 21741 10625 21775 10659
rect 23121 10625 23155 10659
rect 24501 10625 24535 10659
rect 2053 10557 2087 10591
rect 4905 10557 4939 10591
rect 7757 10557 7791 10591
rect 8125 10557 8159 10591
rect 14105 10557 14139 10591
rect 15301 10557 15335 10591
rect 18705 10557 18739 10591
rect 23489 10557 23523 10591
rect 26433 10557 26467 10591
rect 26985 10557 27019 10591
rect 27537 10557 27571 10591
rect 28089 10557 28123 10591
rect 2298 10489 2332 10523
rect 3985 10489 4019 10523
rect 4997 10489 5031 10523
rect 7113 10489 7147 10523
rect 8585 10489 8619 10523
rect 9689 10489 9723 10523
rect 14473 10489 14507 10523
rect 15393 10489 15427 10523
rect 24317 10489 24351 10523
rect 4537 10421 4571 10455
rect 6193 10421 6227 10455
rect 7481 10421 7515 10455
rect 7941 10421 7975 10455
rect 9229 10421 9263 10455
rect 10149 10421 10183 10455
rect 10241 10421 10275 10455
rect 10885 10421 10919 10455
rect 11253 10421 11287 10455
rect 14933 10421 14967 10455
rect 17877 10421 17911 10455
rect 18797 10421 18831 10455
rect 19349 10421 19383 10455
rect 23857 10421 23891 10455
rect 24225 10421 24259 10455
rect 26617 10421 26651 10455
rect 27721 10421 27755 10455
rect 2145 10217 2179 10251
rect 2513 10217 2547 10251
rect 4353 10217 4387 10251
rect 4721 10217 4755 10251
rect 4997 10217 5031 10251
rect 7573 10217 7607 10251
rect 7849 10217 7883 10251
rect 8033 10217 8067 10251
rect 12449 10217 12483 10251
rect 15761 10217 15795 10251
rect 18337 10217 18371 10251
rect 22293 10217 22327 10251
rect 25329 10217 25363 10251
rect 8401 10149 8435 10183
rect 18245 10149 18279 10183
rect 24133 10149 24167 10183
rect 1409 10081 1443 10115
rect 8493 10081 8527 10115
rect 11325 10081 11359 10115
rect 15669 10081 15703 10115
rect 18705 10081 18739 10115
rect 21169 10081 21203 10115
rect 26525 10081 26559 10115
rect 8677 10013 8711 10047
rect 10609 10013 10643 10047
rect 11069 10013 11103 10047
rect 15853 10013 15887 10047
rect 18797 10013 18831 10047
rect 18981 10013 19015 10047
rect 20913 10013 20947 10047
rect 24225 10013 24259 10047
rect 24409 10013 24443 10047
rect 1593 9877 1627 9911
rect 2881 9877 2915 9911
rect 9873 9877 9907 9911
rect 14933 9877 14967 9911
rect 15301 9877 15335 9911
rect 19349 9877 19383 9911
rect 23765 9877 23799 9911
rect 24869 9877 24903 9911
rect 26709 9877 26743 9911
rect 2421 9673 2455 9707
rect 3985 9673 4019 9707
rect 8125 9673 8159 9707
rect 15393 9673 15427 9707
rect 15669 9673 15703 9707
rect 16037 9673 16071 9707
rect 18613 9673 18647 9707
rect 23857 9673 23891 9707
rect 26617 9673 26651 9707
rect 7481 9605 7515 9639
rect 14657 9605 14691 9639
rect 19993 9605 20027 9639
rect 26065 9605 26099 9639
rect 27353 9605 27387 9639
rect 8493 9537 8527 9571
rect 9505 9537 9539 9571
rect 11069 9537 11103 9571
rect 13277 9537 13311 9571
rect 19073 9537 19107 9571
rect 19257 9537 19291 9571
rect 21925 9537 21959 9571
rect 22661 9537 22695 9571
rect 23489 9537 23523 9571
rect 1409 9469 1443 9503
rect 3617 9469 3651 9503
rect 4077 9469 4111 9503
rect 4333 9469 4367 9503
rect 7757 9469 7791 9503
rect 9321 9469 9355 9503
rect 17785 9469 17819 9503
rect 20361 9469 20395 9503
rect 22477 9469 22511 9503
rect 24685 9469 24719 9503
rect 27169 9469 27203 9503
rect 27721 9469 27755 9503
rect 9413 9401 9447 9435
rect 13185 9401 13219 9435
rect 13544 9401 13578 9435
rect 17509 9401 17543 9435
rect 19717 9401 19751 9435
rect 21557 9401 21591 9435
rect 22385 9401 22419 9435
rect 24930 9401 24964 9435
rect 1593 9333 1627 9367
rect 2053 9333 2087 9367
rect 5457 9333 5491 9367
rect 7573 9333 7607 9367
rect 8769 9333 8803 9367
rect 8953 9333 8987 9367
rect 11529 9333 11563 9367
rect 18429 9333 18463 9367
rect 18981 9333 19015 9367
rect 20177 9333 20211 9367
rect 20913 9333 20947 9367
rect 22017 9333 22051 9367
rect 24225 9333 24259 9367
rect 4813 9129 4847 9163
rect 7665 9129 7699 9163
rect 8125 9129 8159 9163
rect 9045 9129 9079 9163
rect 9689 9129 9723 9163
rect 13277 9129 13311 9163
rect 18613 9129 18647 9163
rect 18981 9129 19015 9163
rect 22109 9129 22143 9163
rect 26709 9129 26743 9163
rect 15546 9061 15580 9095
rect 1409 8993 1443 9027
rect 5724 8993 5758 9027
rect 9505 8993 9539 9027
rect 10057 8993 10091 9027
rect 19073 8993 19107 9027
rect 23857 8993 23891 9027
rect 26525 8993 26559 9027
rect 5457 8925 5491 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 15301 8925 15335 8959
rect 19257 8925 19291 8959
rect 23949 8925 23983 8959
rect 24133 8925 24167 8959
rect 18337 8857 18371 8891
rect 1593 8789 1627 8823
rect 6837 8789 6871 8823
rect 9321 8789 9355 8823
rect 16681 8789 16715 8823
rect 21189 8789 21223 8823
rect 23489 8789 23523 8823
rect 24685 8789 24719 8823
rect 2421 8585 2455 8619
rect 4629 8585 4663 8619
rect 8585 8585 8619 8619
rect 10517 8585 10551 8619
rect 14473 8585 14507 8619
rect 15209 8585 15243 8619
rect 18705 8585 18739 8619
rect 19073 8585 19107 8619
rect 19441 8585 19475 8619
rect 23857 8585 23891 8619
rect 1593 8517 1627 8551
rect 24041 8517 24075 8551
rect 2053 8449 2087 8483
rect 4261 8449 4295 8483
rect 5273 8449 5307 8483
rect 5733 8449 5767 8483
rect 8953 8449 8987 8483
rect 14841 8449 14875 8483
rect 16221 8449 16255 8483
rect 23489 8449 23523 8483
rect 24593 8449 24627 8483
rect 1409 8381 1443 8415
rect 5181 8381 5215 8415
rect 9137 8381 9171 8415
rect 15577 8381 15611 8415
rect 16129 8381 16163 8415
rect 21097 8381 21131 8415
rect 21373 8381 21407 8415
rect 24409 8381 24443 8415
rect 25421 8381 25455 8415
rect 5089 8313 5123 8347
rect 6193 8313 6227 8347
rect 9382 8313 9416 8347
rect 23121 8313 23155 8347
rect 24501 8313 24535 8347
rect 25053 8313 25087 8347
rect 26617 8313 26651 8347
rect 4721 8245 4755 8279
rect 8309 8245 8343 8279
rect 15669 8245 15703 8279
rect 16037 8245 16071 8279
rect 20913 8245 20947 8279
rect 1593 8041 1627 8075
rect 4537 8041 4571 8075
rect 9229 8041 9263 8075
rect 10333 8041 10367 8075
rect 24317 8041 24351 8075
rect 24685 8041 24719 8075
rect 26157 8041 26191 8075
rect 26709 8041 26743 8075
rect 16282 7973 16316 8007
rect 21272 7973 21306 8007
rect 24133 7973 24167 8007
rect 1409 7905 1443 7939
rect 11980 7905 12014 7939
rect 16037 7905 16071 7939
rect 18705 7905 18739 7939
rect 21005 7905 21039 7939
rect 26525 7905 26559 7939
rect 4629 7837 4663 7871
rect 4813 7837 4847 7871
rect 5273 7837 5307 7871
rect 5825 7837 5859 7871
rect 11713 7837 11747 7871
rect 24777 7837 24811 7871
rect 24961 7837 24995 7871
rect 15669 7769 15703 7803
rect 18521 7769 18555 7803
rect 2053 7701 2087 7735
rect 4169 7701 4203 7735
rect 9965 7701 9999 7735
rect 13093 7701 13127 7735
rect 17417 7701 17451 7735
rect 22385 7701 22419 7735
rect 25421 7701 25455 7735
rect 4261 7497 4295 7531
rect 9689 7497 9723 7531
rect 15209 7497 15243 7531
rect 16681 7497 16715 7531
rect 18613 7497 18647 7531
rect 20913 7497 20947 7531
rect 21465 7497 21499 7531
rect 23489 7497 23523 7531
rect 24593 7497 24627 7531
rect 27537 7497 27571 7531
rect 3893 7361 3927 7395
rect 4721 7361 4755 7395
rect 5825 7361 5859 7395
rect 8309 7361 8343 7395
rect 13277 7361 13311 7395
rect 16129 7361 16163 7395
rect 16221 7361 16255 7395
rect 22569 7361 22603 7395
rect 24409 7361 24443 7395
rect 25237 7361 25271 7395
rect 26157 7361 26191 7395
rect 1593 7293 1627 7327
rect 1860 7293 1894 7327
rect 5549 7293 5583 7327
rect 13093 7293 13127 7327
rect 19533 7293 19567 7327
rect 24961 7293 24995 7327
rect 5089 7225 5123 7259
rect 8217 7225 8251 7259
rect 8554 7225 8588 7259
rect 12173 7225 12207 7259
rect 13001 7225 13035 7259
rect 15577 7225 15611 7259
rect 16037 7225 16071 7259
rect 19441 7225 19475 7259
rect 19778 7225 19812 7259
rect 21833 7225 21867 7259
rect 22385 7225 22419 7259
rect 25053 7225 25087 7259
rect 26402 7225 26436 7259
rect 2973 7157 3007 7191
rect 5181 7157 5215 7191
rect 5641 7157 5675 7191
rect 11437 7157 11471 7191
rect 11805 7157 11839 7191
rect 12633 7157 12667 7191
rect 14197 7157 14231 7191
rect 15669 7157 15703 7191
rect 18061 7157 18095 7191
rect 22017 7157 22051 7191
rect 22477 7157 22511 7191
rect 24133 7157 24167 7191
rect 25697 7157 25731 7191
rect 25973 7157 26007 7191
rect 1961 6953 1995 6987
rect 2421 6953 2455 6987
rect 6193 6953 6227 6987
rect 8309 6953 8343 6987
rect 11713 6953 11747 6987
rect 13001 6953 13035 6987
rect 13829 6953 13863 6987
rect 16037 6953 16071 6987
rect 19533 6953 19567 6987
rect 22109 6953 22143 6987
rect 22661 6953 22695 6987
rect 23029 6953 23063 6987
rect 25237 6953 25271 6987
rect 4629 6885 4663 6919
rect 10057 6885 10091 6919
rect 22385 6885 22419 6919
rect 1409 6817 1443 6851
rect 3893 6817 3927 6851
rect 6285 6817 6319 6851
rect 12265 6817 12299 6851
rect 17877 6817 17911 6851
rect 18521 6817 18555 6851
rect 23121 6817 23155 6851
rect 24685 6817 24719 6851
rect 26525 6817 26559 6851
rect 4721 6749 4755 6783
rect 4813 6749 4847 6783
rect 6469 6749 6503 6783
rect 10149 6749 10183 6783
rect 10241 6749 10275 6783
rect 12357 6749 12391 6783
rect 12541 6749 12575 6783
rect 13921 6749 13955 6783
rect 14105 6749 14139 6783
rect 17969 6749 18003 6783
rect 18061 6749 18095 6783
rect 23213 6749 23247 6783
rect 25329 6749 25363 6783
rect 25513 6749 25547 6783
rect 1593 6681 1627 6715
rect 11897 6681 11931 6715
rect 24869 6681 24903 6715
rect 26709 6681 26743 6715
rect 4261 6613 4295 6647
rect 5825 6613 5859 6647
rect 7665 6613 7699 6647
rect 9689 6613 9723 6647
rect 13461 6613 13495 6647
rect 15669 6613 15703 6647
rect 16497 6613 16531 6647
rect 17509 6613 17543 6647
rect 20085 6613 20119 6647
rect 21189 6613 21223 6647
rect 26249 6613 26283 6647
rect 1685 6409 1719 6443
rect 3801 6409 3835 6443
rect 5825 6409 5859 6443
rect 6285 6409 6319 6443
rect 6653 6409 6687 6443
rect 7389 6409 7423 6443
rect 9045 6409 9079 6443
rect 10057 6409 10091 6443
rect 11621 6409 11655 6443
rect 12633 6409 12667 6443
rect 13921 6409 13955 6443
rect 17785 6409 17819 6443
rect 22661 6409 22695 6443
rect 23121 6409 23155 6443
rect 23489 6409 23523 6443
rect 24869 6409 24903 6443
rect 25329 6409 25363 6443
rect 25697 6409 25731 6443
rect 26985 6409 27019 6443
rect 4077 6341 4111 6375
rect 9689 6341 9723 6375
rect 17417 6341 17451 6375
rect 4721 6273 4755 6307
rect 4813 6273 4847 6307
rect 5273 6273 5307 6307
rect 8125 6273 8159 6307
rect 10609 6273 10643 6307
rect 11897 6273 11931 6307
rect 16957 6273 16991 6307
rect 18613 6273 18647 6307
rect 19073 6273 19107 6307
rect 20453 6273 20487 6307
rect 20545 6273 20579 6307
rect 1777 6205 1811 6239
rect 8033 6205 8067 6239
rect 13461 6205 13495 6239
rect 15945 6205 15979 6239
rect 16773 6205 16807 6239
rect 18429 6205 18463 6239
rect 18521 6205 18555 6239
rect 19901 6205 19935 6239
rect 26433 6205 26467 6239
rect 2044 6137 2078 6171
rect 10425 6137 10459 6171
rect 11069 6137 11103 6171
rect 16313 6137 16347 6171
rect 19533 6137 19567 6171
rect 20361 6137 20395 6171
rect 26249 6137 26283 6171
rect 3157 6069 3191 6103
rect 4261 6069 4295 6103
rect 4629 6069 4663 6103
rect 7113 6069 7147 6103
rect 7573 6069 7607 6103
rect 7941 6069 7975 6103
rect 9413 6069 9447 6103
rect 10517 6069 10551 6103
rect 14289 6069 14323 6103
rect 16405 6069 16439 6103
rect 16865 6069 16899 6103
rect 18061 6069 18095 6103
rect 19993 6069 20027 6103
rect 26617 6069 26651 6103
rect 2053 5865 2087 5899
rect 2237 5865 2271 5899
rect 3525 5865 3559 5899
rect 5089 5865 5123 5899
rect 9505 5865 9539 5899
rect 10057 5865 10091 5899
rect 10701 5865 10735 5899
rect 11253 5865 11287 5899
rect 12357 5865 12391 5899
rect 12725 5865 12759 5899
rect 17601 5865 17635 5899
rect 18245 5865 18279 5899
rect 20913 5865 20947 5899
rect 21281 5865 21315 5899
rect 1409 5729 1443 5763
rect 3893 5797 3927 5831
rect 4997 5797 5031 5831
rect 11161 5797 11195 5831
rect 18153 5797 18187 5831
rect 7941 5729 7975 5763
rect 13737 5729 13771 5763
rect 15301 5729 15335 5763
rect 15557 5729 15591 5763
rect 22733 5729 22767 5763
rect 25329 5729 25363 5763
rect 26525 5729 26559 5763
rect 2237 5661 2271 5695
rect 2329 5661 2363 5695
rect 5273 5661 5307 5695
rect 8033 5661 8067 5695
rect 8125 5661 8159 5695
rect 11345 5661 11379 5695
rect 12817 5661 12851 5695
rect 13001 5661 13035 5695
rect 18337 5661 18371 5695
rect 18797 5661 18831 5695
rect 19809 5661 19843 5695
rect 21373 5661 21407 5695
rect 21465 5661 21499 5695
rect 22477 5661 22511 5695
rect 1593 5593 1627 5627
rect 10793 5593 10827 5627
rect 25513 5593 25547 5627
rect 4353 5525 4387 5559
rect 4629 5525 4663 5559
rect 7297 5525 7331 5559
rect 7573 5525 7607 5559
rect 13461 5525 13495 5559
rect 16681 5525 16715 5559
rect 17785 5525 17819 5559
rect 20545 5525 20579 5559
rect 23857 5525 23891 5559
rect 26709 5525 26743 5559
rect 2421 5321 2455 5355
rect 2973 5321 3007 5355
rect 5089 5321 5123 5355
rect 5457 5321 5491 5355
rect 7113 5321 7147 5355
rect 10793 5321 10827 5355
rect 14473 5321 14507 5355
rect 15393 5321 15427 5355
rect 17877 5321 17911 5355
rect 18245 5321 18279 5355
rect 18613 5321 18647 5355
rect 20361 5321 20395 5355
rect 20545 5321 20579 5355
rect 21649 5321 21683 5355
rect 25145 5321 25179 5355
rect 26617 5321 26651 5355
rect 27169 5321 27203 5355
rect 10701 5253 10735 5287
rect 2053 5185 2087 5219
rect 9689 5185 9723 5219
rect 11345 5185 11379 5219
rect 13093 5185 13127 5219
rect 16681 5185 16715 5219
rect 16773 5185 16807 5219
rect 21097 5185 21131 5219
rect 1409 5117 1443 5151
rect 3065 5117 3099 5151
rect 3321 5117 3355 5151
rect 7205 5117 7239 5151
rect 15761 5117 15795 5151
rect 16589 5117 16623 5151
rect 21005 5117 21039 5151
rect 25237 5117 25271 5151
rect 7450 5049 7484 5083
rect 9137 5049 9171 5083
rect 11161 5049 11195 5083
rect 13360 5049 13394 5083
rect 16129 5049 16163 5083
rect 21925 5049 21959 5083
rect 22477 5049 22511 5083
rect 25482 5049 25516 5083
rect 1593 4981 1627 5015
rect 4445 4981 4479 5015
rect 8585 4981 8619 5015
rect 10333 4981 10367 5015
rect 11253 4981 11287 5015
rect 11897 4981 11931 5015
rect 12173 4981 12207 5015
rect 12725 4981 12759 5015
rect 16221 4981 16255 5015
rect 19993 4981 20027 5015
rect 20913 4981 20947 5015
rect 22937 4981 22971 5015
rect 24777 4981 24811 5015
rect 3065 4777 3099 4811
rect 4537 4777 4571 4811
rect 5181 4777 5215 4811
rect 7849 4777 7883 4811
rect 10793 4777 10827 4811
rect 11253 4777 11287 4811
rect 11345 4777 11379 4811
rect 11805 4777 11839 4811
rect 12909 4777 12943 4811
rect 13369 4777 13403 4811
rect 16221 4777 16255 4811
rect 16589 4777 16623 4811
rect 19257 4777 19291 4811
rect 21373 4777 21407 4811
rect 21925 4777 21959 4811
rect 25421 4777 25455 4811
rect 4445 4709 4479 4743
rect 7757 4709 7791 4743
rect 11713 4709 11747 4743
rect 15577 4709 15611 4743
rect 20545 4709 20579 4743
rect 21281 4709 21315 4743
rect 23734 4709 23768 4743
rect 1409 4641 1443 4675
rect 2513 4641 2547 4675
rect 13277 4641 13311 4675
rect 19625 4641 19659 4675
rect 19717 4641 19751 4675
rect 23489 4641 23523 4675
rect 26525 4641 26559 4675
rect 4629 4573 4663 4607
rect 7941 4573 7975 4607
rect 8401 4573 8435 4607
rect 11989 4573 12023 4607
rect 12449 4573 12483 4607
rect 13553 4573 13587 4607
rect 19809 4573 19843 4607
rect 21557 4573 21591 4607
rect 24869 4505 24903 4539
rect 1593 4437 1627 4471
rect 2697 4437 2731 4471
rect 4077 4437 4111 4471
rect 6929 4437 6963 4471
rect 7205 4437 7239 4471
rect 7389 4437 7423 4471
rect 20913 4437 20947 4471
rect 26709 4437 26743 4471
rect 4077 4233 4111 4267
rect 4445 4233 4479 4267
rect 7941 4233 7975 4267
rect 11437 4233 11471 4267
rect 13645 4233 13679 4267
rect 15945 4233 15979 4267
rect 19073 4233 19107 4267
rect 23857 4233 23891 4267
rect 24317 4233 24351 4267
rect 26985 4233 27019 4267
rect 13001 4165 13035 4199
rect 2329 4097 2363 4131
rect 4813 4097 4847 4131
rect 6653 4097 6687 4131
rect 16865 4097 16899 4131
rect 16957 4097 16991 4131
rect 18705 4097 18739 4131
rect 19717 4097 19751 4131
rect 20453 4097 20487 4131
rect 21005 4097 21039 4131
rect 21925 4097 21959 4131
rect 22017 4097 22051 4131
rect 1409 4029 1443 4063
rect 2513 4029 2547 4063
rect 3157 4029 3191 4063
rect 6837 4029 6871 4063
rect 8677 4029 8711 4063
rect 9413 4029 9447 4063
rect 16773 4029 16807 4063
rect 19441 4029 19475 4063
rect 21281 4029 21315 4063
rect 21833 4029 21867 4063
rect 22477 4029 22511 4063
rect 26433 4029 26467 4063
rect 27537 4029 27571 4063
rect 28089 4029 28123 4063
rect 2053 3961 2087 3995
rect 7113 3961 7147 3995
rect 8953 3961 8987 3995
rect 16313 3961 16347 3995
rect 20269 3961 20303 3995
rect 1593 3893 1627 3927
rect 2697 3893 2731 3927
rect 7573 3893 7607 3927
rect 11713 3893 11747 3927
rect 12173 3893 12207 3927
rect 13277 3893 13311 3927
rect 16405 3893 16439 3927
rect 19901 3893 19935 3927
rect 20361 3893 20395 3927
rect 21465 3893 21499 3927
rect 26341 3893 26375 3927
rect 26617 3893 26651 3927
rect 27721 3893 27755 3927
rect 1961 3689 1995 3723
rect 3157 3689 3191 3723
rect 4261 3689 4295 3723
rect 7757 3689 7791 3723
rect 12541 3689 12575 3723
rect 17693 3689 17727 3723
rect 19349 3689 19383 3723
rect 20729 3689 20763 3723
rect 21649 3689 21683 3723
rect 4690 3621 4724 3655
rect 1409 3553 1443 3587
rect 2513 3553 2547 3587
rect 4445 3553 4479 3587
rect 9873 3553 9907 3587
rect 10609 3553 10643 3587
rect 11161 3553 11195 3587
rect 11428 3553 11462 3587
rect 16313 3553 16347 3587
rect 16580 3553 16614 3587
rect 19533 3553 19567 3587
rect 20913 3553 20947 3587
rect 23489 3553 23523 3587
rect 26525 3553 26559 3587
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 10149 3485 10183 3519
rect 19809 3485 19843 3519
rect 21189 3485 21223 3519
rect 1593 3349 1627 3383
rect 2697 3349 2731 3383
rect 5825 3349 5859 3383
rect 7113 3349 7147 3383
rect 7389 3349 7423 3383
rect 20269 3349 20303 3383
rect 23673 3349 23707 3383
rect 26709 3349 26743 3383
rect 2421 3145 2455 3179
rect 2789 3145 2823 3179
rect 3801 3145 3835 3179
rect 7021 3145 7055 3179
rect 10793 3145 10827 3179
rect 11345 3145 11379 3179
rect 11713 3145 11747 3179
rect 15485 3145 15519 3179
rect 16405 3145 16439 3179
rect 19073 3145 19107 3179
rect 19349 3145 19383 3179
rect 19533 3145 19567 3179
rect 22477 3145 22511 3179
rect 24777 3145 24811 3179
rect 27353 3145 27387 3179
rect 4353 3077 4387 3111
rect 5733 3077 5767 3111
rect 8033 3077 8067 3111
rect 8401 3077 8435 3111
rect 16681 3077 16715 3111
rect 2053 3009 2087 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 6561 3009 6595 3043
rect 7573 3009 7607 3043
rect 20085 3009 20119 3043
rect 20545 3009 20579 3043
rect 20913 3009 20947 3043
rect 1409 2941 1443 2975
rect 3065 2941 3099 2975
rect 4721 2941 4755 2975
rect 7389 2941 7423 2975
rect 8769 2941 8803 2975
rect 9413 2941 9447 2975
rect 14749 2941 14783 2975
rect 17877 2941 17911 2975
rect 18245 2941 18279 2975
rect 19901 2941 19935 2975
rect 21097 2941 21131 2975
rect 21353 2941 21387 2975
rect 24041 2941 24075 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 3341 2873 3375 2907
rect 6285 2873 6319 2907
rect 7481 2873 7515 2907
rect 9229 2873 9263 2907
rect 9658 2873 9692 2907
rect 15025 2873 15059 2907
rect 18521 2873 18555 2907
rect 19993 2873 20027 2907
rect 24317 2873 24351 2907
rect 1593 2805 1627 2839
rect 4261 2805 4295 2839
rect 4813 2805 4847 2839
rect 23949 2805 23983 2839
rect 26617 2805 26651 2839
rect 27721 2805 27755 2839
rect 3525 2601 3559 2635
rect 4629 2601 4663 2635
rect 5641 2601 5675 2635
rect 6285 2601 6319 2635
rect 7021 2601 7055 2635
rect 7389 2601 7423 2635
rect 8401 2601 8435 2635
rect 9505 2601 9539 2635
rect 17693 2601 17727 2635
rect 18061 2601 18095 2635
rect 19717 2601 19751 2635
rect 20269 2601 20303 2635
rect 20913 2601 20947 2635
rect 21465 2601 21499 2635
rect 24869 2601 24903 2635
rect 25605 2601 25639 2635
rect 2973 2533 3007 2567
rect 11989 2533 12023 2567
rect 18582 2533 18616 2567
rect 1409 2465 1443 2499
rect 2697 2465 2731 2499
rect 5089 2465 5123 2499
rect 5549 2465 5583 2499
rect 6745 2465 6779 2499
rect 7481 2465 7515 2499
rect 8033 2465 8067 2499
rect 9781 2465 9815 2499
rect 10517 2465 10551 2499
rect 11253 2465 11287 2499
rect 13829 2465 13863 2499
rect 14565 2465 14599 2499
rect 16405 2465 16439 2499
rect 17141 2465 17175 2499
rect 18337 2465 18371 2499
rect 21833 2465 21867 2499
rect 22569 2465 22603 2499
rect 24133 2465 24167 2499
rect 25421 2465 25455 2499
rect 25973 2465 26007 2499
rect 26893 2465 26927 2499
rect 27445 2465 27479 2499
rect 2053 2397 2087 2431
rect 5825 2397 5859 2431
rect 7573 2397 7607 2431
rect 9965 2397 9999 2431
rect 11529 2397 11563 2431
rect 14105 2397 14139 2431
rect 16681 2397 16715 2431
rect 22109 2397 22143 2431
rect 24409 2397 24443 2431
rect 5181 2329 5215 2363
rect 1593 2261 1627 2295
rect 4261 2261 4295 2295
rect 27077 2261 27111 2295
<< metal1 >>
rect 3418 22244 3424 22296
rect 3476 22284 3482 22296
rect 12158 22284 12164 22296
rect 3476 22256 12164 22284
rect 3476 22244 3482 22256
rect 12158 22244 12164 22256
rect 12216 22244 12222 22296
rect 2958 22108 2964 22160
rect 3016 22148 3022 22160
rect 5810 22148 5816 22160
rect 3016 22120 5816 22148
rect 3016 22108 3022 22120
rect 5810 22108 5816 22120
rect 5868 22108 5874 22160
rect 20530 22108 20536 22160
rect 20588 22148 20594 22160
rect 25406 22148 25412 22160
rect 20588 22120 25412 22148
rect 20588 22108 20594 22120
rect 25406 22108 25412 22120
rect 25464 22108 25470 22160
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 7009 21131 7067 21137
rect 7009 21097 7021 21131
rect 7055 21128 7067 21131
rect 8294 21128 8300 21140
rect 7055 21100 8300 21128
rect 7055 21097 7067 21100
rect 7009 21091 7067 21097
rect 8294 21088 8300 21100
rect 8352 21088 8358 21140
rect 21085 21131 21143 21137
rect 21085 21097 21097 21131
rect 21131 21128 21143 21131
rect 21634 21128 21640 21140
rect 21131 21100 21640 21128
rect 21131 21097 21143 21100
rect 21085 21091 21143 21097
rect 21634 21088 21640 21100
rect 21692 21088 21698 21140
rect 3694 20952 3700 21004
rect 3752 20992 3758 21004
rect 10502 20992 10508 21004
rect 3752 20964 10508 20992
rect 3752 20952 3758 20964
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 20901 20995 20959 21001
rect 20901 20992 20913 20995
rect 20864 20964 20913 20992
rect 20864 20952 20870 20964
rect 20901 20961 20913 20964
rect 20947 20961 20959 20995
rect 20901 20955 20959 20961
rect 4062 20748 4068 20800
rect 4120 20788 4126 20800
rect 7650 20788 7656 20800
rect 4120 20760 7656 20788
rect 4120 20748 4126 20760
rect 7650 20748 7656 20760
rect 7708 20748 7714 20800
rect 23658 20788 23664 20800
rect 23619 20760 23664 20788
rect 23658 20748 23664 20760
rect 23716 20748 23722 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 1854 20584 1860 20596
rect 1815 20556 1860 20584
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 20806 20584 20812 20596
rect 20767 20556 20812 20584
rect 20806 20544 20812 20556
rect 20864 20584 20870 20596
rect 21361 20587 21419 20593
rect 21361 20584 21373 20587
rect 20864 20556 21373 20584
rect 20864 20544 20870 20556
rect 21361 20553 21373 20556
rect 21407 20553 21419 20587
rect 21361 20547 21419 20553
rect 26605 20587 26663 20593
rect 26605 20553 26617 20587
rect 26651 20584 26663 20587
rect 28258 20584 28264 20596
rect 26651 20556 28264 20584
rect 26651 20553 26663 20556
rect 26605 20547 26663 20553
rect 28258 20544 28264 20556
rect 28316 20544 28322 20596
rect 6457 20451 6515 20457
rect 6457 20417 6469 20451
rect 6503 20448 6515 20451
rect 7377 20451 7435 20457
rect 7377 20448 7389 20451
rect 6503 20420 7389 20448
rect 6503 20417 6515 20420
rect 6457 20411 6515 20417
rect 7377 20417 7389 20420
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 18322 20448 18328 20460
rect 16991 20420 18328 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 18322 20408 18328 20420
rect 18380 20408 18386 20460
rect 23382 20408 23388 20460
rect 23440 20448 23446 20460
rect 23658 20448 23664 20460
rect 23440 20420 23664 20448
rect 23440 20408 23446 20420
rect 23658 20408 23664 20420
rect 23716 20408 23722 20460
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20380 1731 20383
rect 2958 20380 2964 20392
rect 1719 20352 2360 20380
rect 2919 20352 2964 20380
rect 1719 20349 1731 20352
rect 1673 20343 1731 20349
rect 2332 20253 2360 20352
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 8478 20380 8484 20392
rect 8439 20352 8484 20380
rect 8478 20340 8484 20352
rect 8536 20340 8542 20392
rect 13906 20380 13912 20392
rect 13867 20352 13912 20380
rect 13906 20340 13912 20352
rect 13964 20340 13970 20392
rect 16666 20380 16672 20392
rect 16627 20352 16672 20380
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 17405 20383 17463 20389
rect 17405 20380 17417 20383
rect 16724 20352 17417 20380
rect 16724 20340 16730 20352
rect 17405 20349 17417 20352
rect 17451 20349 17463 20383
rect 19426 20380 19432 20392
rect 19387 20352 19432 20380
rect 17405 20343 17463 20349
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 26418 20380 26424 20392
rect 26379 20352 26424 20380
rect 26418 20340 26424 20352
rect 26476 20380 26482 20392
rect 26973 20383 27031 20389
rect 26973 20380 26985 20383
rect 26476 20352 26985 20380
rect 26476 20340 26482 20352
rect 26973 20349 26985 20352
rect 27019 20349 27031 20383
rect 26973 20343 27031 20349
rect 2869 20315 2927 20321
rect 2869 20281 2881 20315
rect 2915 20312 2927 20315
rect 3206 20315 3264 20321
rect 3206 20312 3218 20315
rect 2915 20284 3218 20312
rect 2915 20281 2927 20284
rect 2869 20275 2927 20281
rect 3206 20281 3218 20284
rect 3252 20312 3264 20315
rect 4062 20312 4068 20324
rect 3252 20284 4068 20312
rect 3252 20281 3264 20284
rect 3206 20275 3264 20281
rect 4062 20272 4068 20284
rect 4120 20272 4126 20324
rect 6273 20315 6331 20321
rect 6273 20281 6285 20315
rect 6319 20312 6331 20315
rect 7098 20312 7104 20324
rect 6319 20284 7104 20312
rect 6319 20281 6331 20284
rect 6273 20275 6331 20281
rect 7098 20272 7104 20284
rect 7156 20312 7162 20324
rect 7193 20315 7251 20321
rect 7193 20312 7205 20315
rect 7156 20284 7205 20312
rect 7156 20272 7162 20284
rect 7193 20281 7205 20284
rect 7239 20281 7251 20315
rect 8726 20315 8784 20321
rect 8726 20312 8738 20315
rect 7193 20275 7251 20281
rect 8404 20284 8738 20312
rect 8404 20256 8432 20284
rect 8726 20281 8738 20284
rect 8772 20281 8784 20315
rect 8726 20275 8784 20281
rect 13817 20315 13875 20321
rect 13817 20281 13829 20315
rect 13863 20312 13875 20315
rect 14154 20315 14212 20321
rect 14154 20312 14166 20315
rect 13863 20284 14166 20312
rect 13863 20281 13875 20284
rect 13817 20275 13875 20281
rect 14154 20281 14166 20284
rect 14200 20312 14212 20315
rect 14458 20312 14464 20324
rect 14200 20284 14464 20312
rect 14200 20281 14212 20284
rect 14154 20275 14212 20281
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 19702 20321 19708 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 19696 20312 19708 20321
rect 19383 20284 19708 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 19696 20275 19708 20284
rect 19702 20272 19708 20275
rect 19760 20272 19766 20324
rect 23477 20315 23535 20321
rect 23477 20281 23489 20315
rect 23523 20312 23535 20315
rect 23906 20315 23964 20321
rect 23906 20312 23918 20315
rect 23523 20284 23918 20312
rect 23523 20281 23535 20284
rect 23477 20275 23535 20281
rect 23906 20281 23918 20284
rect 23952 20312 23964 20315
rect 24670 20312 24676 20324
rect 23952 20284 24676 20312
rect 23952 20281 23964 20284
rect 23906 20275 23964 20281
rect 24670 20272 24676 20284
rect 24728 20272 24734 20324
rect 2317 20247 2375 20253
rect 2317 20213 2329 20247
rect 2363 20244 2375 20247
rect 2590 20244 2596 20256
rect 2363 20216 2596 20244
rect 2363 20213 2375 20216
rect 2317 20207 2375 20213
rect 2590 20204 2596 20216
rect 2648 20204 2654 20256
rect 4338 20244 4344 20256
rect 4299 20216 4344 20244
rect 4338 20204 4344 20216
rect 4396 20204 4402 20256
rect 5994 20204 6000 20256
rect 6052 20244 6058 20256
rect 6457 20247 6515 20253
rect 6457 20244 6469 20247
rect 6052 20216 6469 20244
rect 6052 20204 6058 20216
rect 6457 20213 6469 20216
rect 6503 20244 6515 20247
rect 6549 20247 6607 20253
rect 6549 20244 6561 20247
rect 6503 20216 6561 20244
rect 6503 20213 6515 20216
rect 6457 20207 6515 20213
rect 6549 20213 6561 20216
rect 6595 20213 6607 20247
rect 6822 20244 6828 20256
rect 6783 20216 6828 20244
rect 6549 20207 6607 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 6914 20204 6920 20256
rect 6972 20244 6978 20256
rect 7285 20247 7343 20253
rect 7285 20244 7297 20247
rect 6972 20216 7297 20244
rect 6972 20204 6978 20216
rect 7285 20213 7297 20216
rect 7331 20213 7343 20247
rect 8386 20244 8392 20256
rect 8347 20216 8392 20244
rect 7285 20207 7343 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 9858 20244 9864 20256
rect 9819 20216 9864 20244
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 15194 20204 15200 20256
rect 15252 20244 15258 20256
rect 15289 20247 15347 20253
rect 15289 20244 15301 20247
rect 15252 20216 15301 20244
rect 15252 20204 15258 20216
rect 15289 20213 15301 20216
rect 15335 20213 15347 20247
rect 15289 20207 15347 20213
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25041 20247 25099 20253
rect 25041 20244 25053 20247
rect 24912 20216 25053 20244
rect 24912 20204 24918 20216
rect 25041 20213 25053 20216
rect 25087 20213 25099 20247
rect 25041 20207 25099 20213
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 1670 20000 1676 20052
rect 1728 20040 1734 20052
rect 2406 20040 2412 20052
rect 1728 20012 2412 20040
rect 1728 20000 1734 20012
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 5994 20040 6000 20052
rect 5955 20012 6000 20040
rect 5994 20000 6000 20012
rect 6052 20000 6058 20052
rect 6914 20040 6920 20052
rect 6875 20012 6920 20040
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7098 20040 7104 20052
rect 7059 20012 7104 20040
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 8478 20040 8484 20052
rect 8439 20012 8484 20040
rect 8478 20000 8484 20012
rect 8536 20000 8542 20052
rect 13906 20040 13912 20052
rect 13867 20012 13912 20040
rect 13906 20000 13912 20012
rect 13964 20000 13970 20052
rect 19426 20040 19432 20052
rect 19387 20012 19432 20040
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 23198 20040 23204 20052
rect 23159 20012 23204 20040
rect 23198 20000 23204 20012
rect 23256 20000 23262 20052
rect 24489 20043 24547 20049
rect 24489 20009 24501 20043
rect 24535 20040 24547 20043
rect 24949 20043 25007 20049
rect 24949 20040 24961 20043
rect 24535 20012 24961 20040
rect 24535 20009 24547 20012
rect 24489 20003 24547 20009
rect 24949 20009 24961 20012
rect 24995 20040 25007 20043
rect 26513 20043 26571 20049
rect 26513 20040 26525 20043
rect 24995 20012 26525 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 26513 20009 26525 20012
rect 26559 20009 26571 20043
rect 26970 20040 26976 20052
rect 26931 20012 26976 20040
rect 26513 20003 26571 20009
rect 26970 20000 26976 20012
rect 27028 20000 27034 20052
rect 4890 19913 4896 19916
rect 4884 19904 4896 19913
rect 4851 19876 4896 19904
rect 4884 19867 4896 19876
rect 4890 19864 4896 19867
rect 4948 19864 4954 19916
rect 7466 19904 7472 19916
rect 7427 19876 7472 19904
rect 7466 19864 7472 19876
rect 7524 19864 7530 19916
rect 8496 19904 8524 20000
rect 10686 19932 10692 19984
rect 10744 19972 10750 19984
rect 10864 19975 10922 19981
rect 10864 19972 10876 19975
rect 10744 19944 10876 19972
rect 10744 19932 10750 19944
rect 10864 19941 10876 19944
rect 10910 19972 10922 19975
rect 11606 19972 11612 19984
rect 10910 19944 11612 19972
rect 10910 19941 10922 19944
rect 10864 19935 10922 19941
rect 11606 19932 11612 19944
rect 11664 19932 11670 19984
rect 10594 19904 10600 19916
rect 8496 19876 10600 19904
rect 10594 19864 10600 19876
rect 10652 19864 10658 19916
rect 22094 19913 22100 19916
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 16531 19876 17080 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 17052 19848 17080 19876
rect 22088 19867 22100 19913
rect 22152 19904 22158 19916
rect 26878 19904 26884 19916
rect 22152 19876 22188 19904
rect 26839 19876 26884 19904
rect 22094 19864 22100 19867
rect 22152 19864 22158 19876
rect 26878 19864 26884 19876
rect 26936 19864 26942 19916
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 7558 19836 7564 19848
rect 7519 19808 7564 19836
rect 4617 19799 4675 19805
rect 2958 19660 2964 19712
rect 3016 19700 3022 19712
rect 3053 19703 3111 19709
rect 3053 19700 3065 19703
rect 3016 19672 3065 19700
rect 3016 19660 3022 19672
rect 3053 19669 3065 19672
rect 3099 19700 3111 19703
rect 4632 19700 4660 19799
rect 7558 19796 7564 19808
rect 7616 19796 7622 19848
rect 7742 19836 7748 19848
rect 7703 19808 7748 19836
rect 7742 19796 7748 19808
rect 7800 19796 7806 19848
rect 16390 19796 16396 19848
rect 16448 19836 16454 19848
rect 16577 19839 16635 19845
rect 16577 19836 16589 19839
rect 16448 19808 16589 19836
rect 16448 19796 16454 19808
rect 16577 19805 16589 19808
rect 16623 19805 16635 19839
rect 16577 19799 16635 19805
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19805 16727 19839
rect 16669 19799 16727 19805
rect 16482 19728 16488 19780
rect 16540 19768 16546 19780
rect 16684 19768 16712 19799
rect 17034 19796 17040 19848
rect 17092 19836 17098 19848
rect 17681 19839 17739 19845
rect 17681 19836 17693 19839
rect 17092 19808 17693 19836
rect 17092 19796 17098 19808
rect 17681 19805 17693 19808
rect 17727 19805 17739 19839
rect 21818 19836 21824 19848
rect 21779 19808 21824 19836
rect 17681 19799 17739 19805
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 25038 19836 25044 19848
rect 24999 19808 25044 19836
rect 25038 19796 25044 19808
rect 25096 19796 25102 19848
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19805 25191 19839
rect 27062 19836 27068 19848
rect 27023 19808 27068 19836
rect 25133 19799 25191 19805
rect 16540 19740 16712 19768
rect 16540 19728 16546 19740
rect 24854 19728 24860 19780
rect 24912 19768 24918 19780
rect 25148 19768 25176 19799
rect 27062 19796 27068 19808
rect 27120 19796 27126 19848
rect 24912 19740 25176 19768
rect 24912 19728 24918 19740
rect 5350 19700 5356 19712
rect 3099 19672 5356 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 11330 19660 11336 19712
rect 11388 19700 11394 19712
rect 11977 19703 12035 19709
rect 11977 19700 11989 19703
rect 11388 19672 11989 19700
rect 11388 19660 11394 19672
rect 11977 19669 11989 19672
rect 12023 19669 12035 19703
rect 15654 19700 15660 19712
rect 15615 19672 15660 19700
rect 11977 19663 12035 19669
rect 15654 19660 15660 19672
rect 15712 19660 15718 19712
rect 15838 19660 15844 19712
rect 15896 19700 15902 19712
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15896 19672 16129 19700
rect 15896 19660 15902 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 23842 19700 23848 19712
rect 23803 19672 23848 19700
rect 16117 19663 16175 19669
rect 23842 19660 23848 19672
rect 23900 19660 23906 19712
rect 24026 19660 24032 19712
rect 24084 19700 24090 19712
rect 24581 19703 24639 19709
rect 24581 19700 24593 19703
rect 24084 19672 24593 19700
rect 24084 19660 24090 19672
rect 24581 19669 24593 19672
rect 24627 19669 24639 19703
rect 24581 19663 24639 19669
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 10686 19496 10692 19508
rect 10647 19468 10692 19496
rect 10686 19456 10692 19468
rect 10744 19456 10750 19508
rect 14458 19496 14464 19508
rect 14419 19468 14464 19496
rect 14458 19456 14464 19468
rect 14516 19456 14522 19508
rect 17034 19496 17040 19508
rect 16995 19468 17040 19496
rect 17034 19456 17040 19468
rect 17092 19456 17098 19508
rect 23198 19456 23204 19508
rect 23256 19496 23262 19508
rect 23385 19499 23443 19505
rect 23385 19496 23397 19499
rect 23256 19468 23397 19496
rect 23256 19456 23262 19468
rect 23385 19465 23397 19468
rect 23431 19465 23443 19499
rect 23385 19459 23443 19465
rect 7377 19431 7435 19437
rect 7377 19397 7389 19431
rect 7423 19428 7435 19431
rect 7466 19428 7472 19440
rect 7423 19400 7472 19428
rect 7423 19397 7435 19400
rect 7377 19391 7435 19397
rect 7466 19388 7472 19400
rect 7524 19428 7530 19440
rect 7524 19400 7880 19428
rect 7524 19388 7530 19400
rect 6273 19295 6331 19301
rect 6273 19261 6285 19295
rect 6319 19292 6331 19295
rect 7558 19292 7564 19304
rect 6319 19264 7564 19292
rect 6319 19261 6331 19264
rect 6273 19255 6331 19261
rect 7558 19252 7564 19264
rect 7616 19252 7622 19304
rect 7852 19292 7880 19400
rect 10594 19388 10600 19440
rect 10652 19428 10658 19440
rect 10965 19431 11023 19437
rect 10965 19428 10977 19431
rect 10652 19400 10977 19428
rect 10652 19388 10658 19400
rect 10965 19397 10977 19400
rect 11011 19397 11023 19431
rect 14476 19428 14504 19456
rect 23400 19428 23428 19459
rect 24670 19456 24676 19508
rect 24728 19496 24734 19508
rect 24949 19499 25007 19505
rect 24949 19496 24961 19499
rect 24728 19468 24961 19496
rect 24728 19456 24734 19468
rect 24949 19465 24961 19468
rect 24995 19465 25007 19499
rect 24949 19459 25007 19465
rect 14476 19400 16160 19428
rect 23400 19400 24256 19428
rect 10965 19391 11023 19397
rect 8021 19363 8079 19369
rect 8021 19329 8033 19363
rect 8067 19360 8079 19363
rect 8478 19360 8484 19372
rect 8067 19332 8484 19360
rect 8067 19329 8079 19332
rect 8021 19323 8079 19329
rect 8478 19320 8484 19332
rect 8536 19320 8542 19372
rect 15654 19320 15660 19372
rect 15712 19360 15718 19372
rect 16022 19360 16028 19372
rect 15712 19332 16028 19360
rect 15712 19320 15718 19332
rect 16022 19320 16028 19332
rect 16080 19320 16086 19372
rect 16132 19369 16160 19400
rect 16117 19363 16175 19369
rect 16117 19329 16129 19363
rect 16163 19329 16175 19363
rect 16117 19323 16175 19329
rect 21818 19320 21824 19372
rect 21876 19360 21882 19372
rect 21876 19332 22140 19360
rect 21876 19320 21882 19332
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 7852 19264 8769 19292
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 13078 19292 13084 19304
rect 12991 19264 13084 19292
rect 8757 19255 8815 19261
rect 13078 19252 13084 19264
rect 13136 19292 13142 19304
rect 13722 19292 13728 19304
rect 13136 19264 13728 19292
rect 13136 19252 13142 19264
rect 13722 19252 13728 19264
rect 13780 19252 13786 19304
rect 15105 19295 15163 19301
rect 15105 19261 15117 19295
rect 15151 19292 15163 19295
rect 15838 19292 15844 19304
rect 15151 19264 15844 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15838 19252 15844 19264
rect 15896 19292 15902 19304
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15896 19264 15945 19292
rect 15896 19252 15902 19264
rect 15933 19261 15945 19264
rect 15979 19261 15991 19295
rect 15933 19255 15991 19261
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 4985 19227 5043 19233
rect 4985 19224 4997 19227
rect 4948 19196 4997 19224
rect 4948 19184 4954 19196
rect 4985 19193 4997 19196
rect 5031 19224 5043 19227
rect 5718 19224 5724 19236
rect 5031 19196 5724 19224
rect 5031 19193 5043 19196
rect 4985 19187 5043 19193
rect 5718 19184 5724 19196
rect 5776 19184 5782 19236
rect 6641 19227 6699 19233
rect 6641 19193 6653 19227
rect 6687 19224 6699 19227
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 6687 19196 7757 19224
rect 6687 19193 6699 19196
rect 6641 19187 6699 19193
rect 7745 19193 7757 19196
rect 7791 19224 7803 19227
rect 8941 19227 8999 19233
rect 8941 19224 8953 19227
rect 7791 19196 8953 19224
rect 7791 19193 7803 19196
rect 7745 19187 7803 19193
rect 8941 19193 8953 19196
rect 8987 19193 8999 19227
rect 8941 19187 8999 19193
rect 12989 19227 13047 19233
rect 12989 19193 13001 19227
rect 13035 19224 13047 19227
rect 13326 19227 13384 19233
rect 13326 19224 13338 19227
rect 13035 19196 13338 19224
rect 13035 19193 13047 19196
rect 12989 19187 13047 19193
rect 13326 19193 13338 19196
rect 13372 19224 13384 19227
rect 13538 19224 13544 19236
rect 13372 19196 13544 19224
rect 13372 19193 13384 19196
rect 13326 19187 13384 19193
rect 13538 19184 13544 19196
rect 13596 19224 13602 19236
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 13596 19196 15393 19224
rect 13596 19184 13602 19196
rect 15381 19193 15393 19196
rect 15427 19193 15439 19227
rect 15381 19187 15439 19193
rect 21913 19227 21971 19233
rect 21913 19193 21925 19227
rect 21959 19224 21971 19227
rect 22002 19224 22008 19236
rect 21959 19196 22008 19224
rect 21959 19193 21971 19196
rect 21913 19187 21971 19193
rect 22002 19184 22008 19196
rect 22060 19184 22066 19236
rect 22112 19224 22140 19332
rect 23842 19320 23848 19372
rect 23900 19360 23906 19372
rect 24228 19369 24256 19400
rect 24121 19363 24179 19369
rect 24121 19360 24133 19363
rect 23900 19332 24133 19360
rect 23900 19320 23906 19332
rect 24121 19329 24133 19332
rect 24167 19329 24179 19363
rect 24121 19323 24179 19329
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19329 24271 19363
rect 24964 19360 24992 19459
rect 25038 19456 25044 19508
rect 25096 19496 25102 19508
rect 25501 19499 25559 19505
rect 25501 19496 25513 19499
rect 25096 19468 25513 19496
rect 25096 19456 25102 19468
rect 25501 19465 25513 19468
rect 25547 19465 25559 19499
rect 26878 19496 26884 19508
rect 26839 19468 26884 19496
rect 25501 19459 25559 19465
rect 26878 19456 26884 19468
rect 26936 19456 26942 19508
rect 26605 19431 26663 19437
rect 26605 19397 26617 19431
rect 26651 19428 26663 19431
rect 26970 19428 26976 19440
rect 26651 19400 26976 19428
rect 26651 19397 26663 19400
rect 26605 19391 26663 19397
rect 26970 19388 26976 19400
rect 27028 19388 27034 19440
rect 26053 19363 26111 19369
rect 26053 19360 26065 19363
rect 24964 19332 26065 19360
rect 24213 19323 24271 19329
rect 26053 19329 26065 19332
rect 26099 19360 26111 19363
rect 27062 19360 27068 19372
rect 26099 19332 27068 19360
rect 26099 19329 26111 19332
rect 26053 19323 26111 19329
rect 27062 19320 27068 19332
rect 27120 19360 27126 19372
rect 27249 19363 27307 19369
rect 27249 19360 27261 19363
rect 27120 19332 27261 19360
rect 27120 19320 27126 19332
rect 27249 19329 27261 19332
rect 27295 19329 27307 19363
rect 27249 19323 27307 19329
rect 23109 19295 23167 19301
rect 23109 19261 23121 19295
rect 23155 19292 23167 19295
rect 24026 19292 24032 19304
rect 23155 19264 24032 19292
rect 23155 19261 23167 19264
rect 23109 19255 23167 19261
rect 24026 19252 24032 19264
rect 24084 19252 24090 19304
rect 22281 19227 22339 19233
rect 22281 19224 22293 19227
rect 22112 19196 22293 19224
rect 22281 19193 22293 19196
rect 22327 19224 22339 19227
rect 23382 19224 23388 19236
rect 22327 19196 23388 19224
rect 22327 19193 22339 19196
rect 22281 19187 22339 19193
rect 23382 19184 23388 19196
rect 23440 19184 23446 19236
rect 25590 19184 25596 19236
rect 25648 19224 25654 19236
rect 25961 19227 26019 19233
rect 25961 19224 25973 19227
rect 25648 19196 25973 19224
rect 25648 19184 25654 19196
rect 25961 19193 25973 19196
rect 26007 19193 26019 19227
rect 25961 19187 26019 19193
rect 4430 19156 4436 19168
rect 4391 19128 4436 19156
rect 4430 19116 4436 19128
rect 4488 19116 4494 19168
rect 5353 19159 5411 19165
rect 5353 19125 5365 19159
rect 5399 19156 5411 19159
rect 5442 19156 5448 19168
rect 5399 19128 5448 19156
rect 5399 19125 5411 19128
rect 5353 19119 5411 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 7190 19156 7196 19168
rect 7151 19128 7196 19156
rect 7190 19116 7196 19128
rect 7248 19156 7254 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7248 19128 7849 19156
rect 7248 19116 7254 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 8478 19156 8484 19168
rect 8439 19128 8484 19156
rect 7837 19119 7895 19125
rect 8478 19116 8484 19128
rect 8536 19116 8542 19168
rect 15562 19156 15568 19168
rect 15523 19128 15568 19156
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16390 19116 16396 19168
rect 16448 19156 16454 19168
rect 16666 19156 16672 19168
rect 16448 19128 16672 19156
rect 16448 19116 16454 19128
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 20346 19156 20352 19168
rect 20307 19128 20352 19156
rect 20346 19116 20352 19128
rect 20404 19116 20410 19168
rect 23661 19159 23719 19165
rect 23661 19125 23673 19159
rect 23707 19156 23719 19159
rect 24486 19156 24492 19168
rect 23707 19128 24492 19156
rect 23707 19125 23719 19128
rect 23661 19119 23719 19125
rect 24486 19116 24492 19128
rect 24544 19116 24550 19168
rect 25314 19156 25320 19168
rect 25275 19128 25320 19156
rect 25314 19116 25320 19128
rect 25372 19156 25378 19168
rect 25869 19159 25927 19165
rect 25869 19156 25881 19159
rect 25372 19128 25881 19156
rect 25372 19116 25378 19128
rect 25869 19125 25881 19128
rect 25915 19125 25927 19159
rect 25869 19119 25927 19125
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18952 7435 18955
rect 7558 18952 7564 18964
rect 7423 18924 7564 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 7558 18912 7564 18924
rect 7616 18912 7622 18964
rect 7742 18912 7748 18964
rect 7800 18912 7806 18964
rect 13078 18952 13084 18964
rect 13039 18924 13084 18952
rect 13078 18912 13084 18924
rect 13136 18912 13142 18964
rect 14001 18955 14059 18961
rect 14001 18921 14013 18955
rect 14047 18952 14059 18955
rect 14090 18952 14096 18964
rect 14047 18924 14096 18952
rect 14047 18921 14059 18924
rect 14001 18915 14059 18921
rect 14090 18912 14096 18924
rect 14148 18952 14154 18964
rect 15562 18952 15568 18964
rect 14148 18924 15568 18952
rect 14148 18912 14154 18924
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16022 18952 16028 18964
rect 15983 18924 16028 18952
rect 16022 18912 16028 18924
rect 16080 18912 16086 18964
rect 23385 18955 23443 18961
rect 23385 18921 23397 18955
rect 23431 18952 23443 18955
rect 23842 18952 23848 18964
rect 23431 18924 23848 18952
rect 23431 18921 23443 18924
rect 23385 18915 23443 18921
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 25038 18952 25044 18964
rect 24999 18924 25044 18952
rect 25038 18912 25044 18924
rect 25096 18912 25102 18964
rect 26513 18955 26571 18961
rect 26513 18921 26525 18955
rect 26559 18952 26571 18955
rect 26878 18952 26884 18964
rect 26559 18924 26884 18952
rect 26559 18921 26571 18924
rect 26513 18915 26571 18921
rect 26878 18912 26884 18924
rect 26936 18912 26942 18964
rect 7193 18887 7251 18893
rect 7193 18853 7205 18887
rect 7239 18884 7251 18887
rect 7760 18884 7788 18912
rect 7239 18856 7788 18884
rect 7239 18853 7251 18856
rect 7193 18847 7251 18853
rect 10778 18844 10784 18896
rect 10836 18884 10842 18896
rect 10956 18887 11014 18893
rect 10956 18884 10968 18887
rect 10836 18856 10968 18884
rect 10836 18844 10842 18856
rect 10956 18853 10968 18856
rect 11002 18884 11014 18887
rect 11330 18884 11336 18896
rect 11002 18856 11336 18884
rect 11002 18853 11014 18856
rect 10956 18847 11014 18853
rect 11330 18844 11336 18856
rect 11388 18844 11394 18896
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2130 18816 2136 18828
rect 1443 18788 2136 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2130 18776 2136 18788
rect 2188 18776 2194 18828
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 4430 18816 4436 18828
rect 3844 18788 4436 18816
rect 3844 18776 3850 18788
rect 4430 18776 4436 18788
rect 4488 18816 4494 18828
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4488 18788 4721 18816
rect 4488 18776 4494 18788
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 7650 18776 7656 18828
rect 7708 18816 7714 18828
rect 7745 18819 7803 18825
rect 7745 18816 7757 18819
rect 7708 18788 7757 18816
rect 7708 18776 7714 18788
rect 7745 18785 7757 18788
rect 7791 18785 7803 18819
rect 7745 18779 7803 18785
rect 10594 18776 10600 18828
rect 10652 18816 10658 18828
rect 10689 18819 10747 18825
rect 10689 18816 10701 18819
rect 10652 18788 10701 18816
rect 10652 18776 10658 18788
rect 10689 18785 10701 18788
rect 10735 18785 10747 18819
rect 10689 18779 10747 18785
rect 15838 18776 15844 18828
rect 15896 18816 15902 18828
rect 16393 18819 16451 18825
rect 16393 18816 16405 18819
rect 15896 18788 16405 18816
rect 15896 18776 15902 18788
rect 16393 18785 16405 18788
rect 16439 18785 16451 18819
rect 16393 18779 16451 18785
rect 18322 18776 18328 18828
rect 18380 18816 18386 18828
rect 18489 18819 18547 18825
rect 18489 18816 18501 18819
rect 18380 18788 18501 18816
rect 18380 18776 18386 18788
rect 18489 18785 18501 18788
rect 18535 18785 18547 18819
rect 21266 18816 21272 18828
rect 21227 18788 21272 18816
rect 18489 18779 18547 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 21361 18819 21419 18825
rect 21361 18785 21373 18819
rect 21407 18816 21419 18819
rect 21634 18816 21640 18828
rect 21407 18788 21640 18816
rect 21407 18785 21419 18788
rect 21361 18779 21419 18785
rect 21634 18776 21640 18788
rect 21692 18776 21698 18828
rect 23750 18816 23756 18828
rect 23711 18788 23756 18816
rect 23750 18776 23756 18788
rect 23808 18776 23814 18828
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 4985 18751 5043 18757
rect 4985 18717 4997 18751
rect 5031 18748 5043 18751
rect 5258 18748 5264 18760
rect 5031 18720 5264 18748
rect 5031 18717 5043 18720
rect 4985 18711 5043 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 7834 18748 7840 18760
rect 7795 18720 7840 18748
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 8021 18751 8079 18757
rect 8021 18717 8033 18751
rect 8067 18748 8079 18751
rect 8478 18748 8484 18760
rect 8067 18720 8484 18748
rect 8067 18717 8079 18720
rect 8021 18711 8079 18717
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 13814 18708 13820 18760
rect 13872 18748 13878 18760
rect 14093 18751 14151 18757
rect 14093 18748 14105 18751
rect 13872 18720 14105 18748
rect 13872 18708 13878 18720
rect 14093 18717 14105 18720
rect 14139 18717 14151 18751
rect 14093 18711 14151 18717
rect 14277 18751 14335 18757
rect 14277 18717 14289 18751
rect 14323 18748 14335 18751
rect 14366 18748 14372 18760
rect 14323 18720 14372 18748
rect 14323 18717 14335 18720
rect 14277 18711 14335 18717
rect 14366 18708 14372 18720
rect 14424 18748 14430 18760
rect 15102 18748 15108 18760
rect 14424 18720 15108 18748
rect 14424 18708 14430 18720
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 16574 18708 16580 18760
rect 16632 18748 16638 18760
rect 18230 18748 18236 18760
rect 16632 18720 16677 18748
rect 18191 18720 18236 18748
rect 16632 18708 16638 18720
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 21453 18751 21511 18757
rect 21453 18748 21465 18751
rect 20272 18720 21465 18748
rect 20272 18624 20300 18720
rect 21453 18717 21465 18720
rect 21499 18717 21511 18751
rect 23842 18748 23848 18760
rect 23803 18720 23848 18748
rect 21453 18711 21511 18717
rect 23842 18708 23848 18720
rect 23900 18708 23906 18760
rect 23934 18708 23940 18760
rect 23992 18748 23998 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 23992 18720 24593 18748
rect 23992 18708 23998 18720
rect 24581 18717 24593 18720
rect 24627 18748 24639 18751
rect 24762 18748 24768 18760
rect 24627 18720 24768 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 24762 18708 24768 18720
rect 24820 18708 24826 18760
rect 1394 18572 1400 18624
rect 1452 18612 1458 18624
rect 1581 18615 1639 18621
rect 1581 18612 1593 18615
rect 1452 18584 1593 18612
rect 1452 18572 1458 18584
rect 1581 18581 1593 18584
rect 1627 18581 1639 18615
rect 2038 18612 2044 18624
rect 1999 18584 2044 18612
rect 1581 18575 1639 18581
rect 2038 18572 2044 18584
rect 2096 18572 2102 18624
rect 2314 18612 2320 18624
rect 2275 18584 2320 18612
rect 2314 18572 2320 18584
rect 2372 18572 2378 18624
rect 3881 18615 3939 18621
rect 3881 18581 3893 18615
rect 3927 18612 3939 18615
rect 4341 18615 4399 18621
rect 4341 18612 4353 18615
rect 3927 18584 4353 18612
rect 3927 18581 3939 18584
rect 3881 18575 3939 18581
rect 4341 18581 4353 18584
rect 4387 18612 4399 18615
rect 4614 18612 4620 18624
rect 4387 18584 4620 18612
rect 4387 18581 4399 18584
rect 4341 18575 4399 18581
rect 4614 18572 4620 18584
rect 4672 18572 4678 18624
rect 8754 18612 8760 18624
rect 8715 18584 8760 18612
rect 8754 18572 8760 18584
rect 8812 18572 8818 18624
rect 9030 18612 9036 18624
rect 8991 18584 9036 18612
rect 9030 18572 9036 18584
rect 9088 18572 9094 18624
rect 12066 18612 12072 18624
rect 12027 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 13354 18572 13360 18624
rect 13412 18612 13418 18624
rect 13633 18615 13691 18621
rect 13633 18612 13645 18615
rect 13412 18584 13645 18612
rect 13412 18572 13418 18584
rect 13633 18581 13645 18584
rect 13679 18581 13691 18615
rect 15010 18612 15016 18624
rect 14971 18584 15016 18612
rect 13633 18575 13691 18581
rect 15010 18572 15016 18584
rect 15068 18572 15074 18624
rect 15562 18612 15568 18624
rect 15523 18584 15568 18612
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 19334 18572 19340 18624
rect 19392 18612 19398 18624
rect 19613 18615 19671 18621
rect 19613 18612 19625 18615
rect 19392 18584 19625 18612
rect 19392 18572 19398 18584
rect 19613 18581 19625 18584
rect 19659 18581 19671 18615
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 19613 18575 19671 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20806 18572 20812 18624
rect 20864 18612 20870 18624
rect 20901 18615 20959 18621
rect 20901 18612 20913 18615
rect 20864 18584 20913 18612
rect 20864 18572 20870 18584
rect 20901 18581 20913 18584
rect 20947 18581 20959 18615
rect 25590 18612 25596 18624
rect 25551 18584 25596 18612
rect 20901 18575 20959 18581
rect 25590 18572 25596 18584
rect 25648 18572 25654 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 3786 18408 3792 18420
rect 3747 18380 3792 18408
rect 3786 18368 3792 18380
rect 3844 18368 3850 18420
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 4798 18408 4804 18420
rect 4203 18380 4804 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 4798 18368 4804 18380
rect 4856 18368 4862 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 7101 18411 7159 18417
rect 7101 18408 7113 18411
rect 6972 18380 7113 18408
rect 6972 18368 6978 18380
rect 7101 18377 7113 18380
rect 7147 18377 7159 18411
rect 7101 18371 7159 18377
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 8113 18411 8171 18417
rect 8113 18408 8125 18411
rect 7708 18380 8125 18408
rect 7708 18368 7714 18380
rect 8113 18377 8125 18380
rect 8159 18377 8171 18411
rect 8113 18371 8171 18377
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10652 18380 11069 18408
rect 10652 18368 10658 18380
rect 11057 18377 11069 18380
rect 11103 18408 11115 18411
rect 13078 18408 13084 18420
rect 11103 18380 13084 18408
rect 11103 18377 11115 18380
rect 11057 18371 11115 18377
rect 3053 18343 3111 18349
rect 3053 18309 3065 18343
rect 3099 18309 3111 18343
rect 3053 18303 3111 18309
rect 6641 18343 6699 18349
rect 6641 18309 6653 18343
rect 6687 18340 6699 18343
rect 10778 18340 10784 18352
rect 6687 18312 8524 18340
rect 10739 18312 10784 18340
rect 6687 18309 6699 18312
rect 6641 18303 6699 18309
rect 2682 18232 2688 18284
rect 2740 18272 2746 18284
rect 3068 18272 3096 18303
rect 8496 18284 8524 18312
rect 10778 18300 10784 18312
rect 10836 18300 10842 18352
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 2740 18244 4813 18272
rect 2740 18232 2746 18244
rect 4801 18241 4813 18244
rect 4847 18272 4859 18275
rect 5074 18272 5080 18284
rect 4847 18244 5080 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5074 18232 5080 18244
rect 5132 18272 5138 18284
rect 5629 18275 5687 18281
rect 5629 18272 5641 18275
rect 5132 18244 5641 18272
rect 5132 18232 5138 18244
rect 5629 18241 5641 18244
rect 5675 18241 5687 18275
rect 5629 18235 5687 18241
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 6273 18275 6331 18281
rect 6273 18272 6285 18275
rect 5776 18244 6285 18272
rect 5776 18232 5782 18244
rect 6273 18241 6285 18244
rect 6319 18272 6331 18275
rect 7742 18272 7748 18284
rect 6319 18244 7748 18272
rect 6319 18241 6331 18244
rect 6273 18235 6331 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 8478 18232 8484 18284
rect 8536 18272 8542 18284
rect 8573 18275 8631 18281
rect 8573 18272 8585 18275
rect 8536 18244 8585 18272
rect 8536 18232 8542 18244
rect 8573 18241 8585 18244
rect 8619 18272 8631 18275
rect 9306 18272 9312 18284
rect 8619 18244 9312 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 9306 18232 9312 18244
rect 9364 18232 9370 18284
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 1762 18204 1768 18216
rect 1719 18176 1768 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 1762 18164 1768 18176
rect 1820 18204 1826 18216
rect 2314 18204 2320 18216
rect 1820 18176 2320 18204
rect 1820 18164 1826 18176
rect 2314 18164 2320 18176
rect 2372 18164 2378 18216
rect 4614 18204 4620 18216
rect 4575 18176 4620 18204
rect 4614 18164 4620 18176
rect 4672 18164 4678 18216
rect 9030 18204 9036 18216
rect 8991 18176 9036 18204
rect 9030 18164 9036 18176
rect 9088 18204 9094 18216
rect 9674 18204 9680 18216
rect 9088 18176 9680 18204
rect 9088 18164 9094 18176
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 12360 18204 12388 18380
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13814 18368 13820 18420
rect 13872 18408 13878 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 13872 18380 14933 18408
rect 13872 18368 13878 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 16025 18411 16083 18417
rect 16025 18408 16037 18411
rect 15896 18380 16037 18408
rect 15896 18368 15902 18380
rect 16025 18377 16037 18380
rect 16071 18377 16083 18411
rect 16482 18408 16488 18420
rect 16443 18380 16488 18408
rect 16025 18371 16083 18377
rect 16482 18368 16488 18380
rect 16540 18368 16546 18420
rect 18230 18368 18236 18420
rect 18288 18408 18294 18420
rect 18690 18408 18696 18420
rect 18288 18380 18696 18408
rect 18288 18368 18294 18380
rect 18690 18368 18696 18380
rect 18748 18408 18754 18420
rect 19242 18408 19248 18420
rect 18748 18380 19248 18408
rect 18748 18368 18754 18380
rect 19242 18368 19248 18380
rect 19300 18368 19306 18420
rect 21266 18408 21272 18420
rect 21227 18380 21272 18408
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 22741 18411 22799 18417
rect 22741 18377 22753 18411
rect 22787 18408 22799 18411
rect 23750 18408 23756 18420
rect 22787 18380 23756 18408
rect 22787 18377 22799 18380
rect 22741 18371 22799 18377
rect 23750 18368 23756 18380
rect 23808 18368 23814 18420
rect 27062 18368 27068 18420
rect 27120 18408 27126 18420
rect 27525 18411 27583 18417
rect 27525 18408 27537 18411
rect 27120 18380 27537 18408
rect 27120 18368 27126 18380
rect 27525 18377 27537 18380
rect 27571 18377 27583 18411
rect 27525 18371 27583 18377
rect 14366 18340 14372 18352
rect 14327 18312 14372 18340
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 14737 18343 14795 18349
rect 14737 18340 14749 18343
rect 14516 18312 14749 18340
rect 14516 18300 14522 18312
rect 14737 18309 14749 18312
rect 14783 18340 14795 18343
rect 15562 18340 15568 18352
rect 14783 18312 15568 18340
rect 14783 18309 14795 18312
rect 14737 18303 14795 18309
rect 15010 18232 15016 18284
rect 15068 18272 15074 18284
rect 15488 18281 15516 18312
rect 15562 18300 15568 18312
rect 15620 18300 15626 18352
rect 21634 18340 21640 18352
rect 21595 18312 21640 18340
rect 21634 18300 21640 18312
rect 21692 18300 21698 18352
rect 22002 18300 22008 18352
rect 22060 18340 22066 18352
rect 23017 18343 23075 18349
rect 23017 18340 23029 18343
rect 22060 18312 23029 18340
rect 22060 18300 22066 18312
rect 23017 18309 23029 18312
rect 23063 18340 23075 18343
rect 23934 18340 23940 18352
rect 23063 18312 23940 18340
rect 23063 18309 23075 18312
rect 23017 18303 23075 18309
rect 23934 18300 23940 18312
rect 23992 18300 23998 18352
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15068 18244 15393 18272
rect 15068 18232 15074 18244
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15838 18232 15844 18284
rect 15896 18272 15902 18284
rect 16574 18272 16580 18284
rect 15896 18244 16580 18272
rect 15896 18232 15902 18244
rect 16574 18232 16580 18244
rect 16632 18272 16638 18284
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 16632 18244 16773 18272
rect 16632 18232 16638 18244
rect 16761 18241 16773 18244
rect 16807 18241 16819 18275
rect 16761 18235 16819 18241
rect 18322 18232 18328 18284
rect 18380 18272 18386 18284
rect 20254 18272 20260 18284
rect 18380 18244 20260 18272
rect 18380 18232 18386 18244
rect 20254 18232 20260 18244
rect 20312 18272 20318 18284
rect 20809 18275 20867 18281
rect 20809 18272 20821 18275
rect 20312 18244 20821 18272
rect 20312 18232 20318 18244
rect 20809 18241 20821 18244
rect 20855 18272 20867 18275
rect 24397 18275 24455 18281
rect 20855 18244 22048 18272
rect 20855 18241 20867 18244
rect 20809 18235 20867 18241
rect 12434 18204 12440 18216
rect 12360 18176 12440 18204
rect 12434 18164 12440 18176
rect 12492 18204 12498 18216
rect 20070 18204 20076 18216
rect 12492 18176 12585 18204
rect 20031 18176 20076 18204
rect 12492 18164 12498 18176
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 22020 18213 22048 18244
rect 24397 18241 24409 18275
rect 24443 18272 24455 18275
rect 24670 18272 24676 18284
rect 24443 18244 24676 18272
rect 24443 18241 24455 18244
rect 24397 18235 24455 18241
rect 24670 18232 24676 18244
rect 24728 18232 24734 18284
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20404 18176 20637 18204
rect 20404 18164 20410 18176
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 22005 18207 22063 18213
rect 22005 18173 22017 18207
rect 22051 18173 22063 18207
rect 22005 18167 22063 18173
rect 25774 18164 25780 18216
rect 25832 18204 25838 18216
rect 26142 18204 26148 18216
rect 25832 18176 26148 18204
rect 25832 18164 25838 18176
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 1940 18139 1998 18145
rect 1940 18105 1952 18139
rect 1986 18136 1998 18139
rect 2038 18136 2044 18148
rect 1986 18108 2044 18136
rect 1986 18105 1998 18108
rect 1940 18099 1998 18105
rect 2038 18096 2044 18108
rect 2096 18136 2102 18148
rect 2498 18136 2504 18148
rect 2096 18108 2504 18136
rect 2096 18096 2102 18108
rect 2498 18096 2504 18108
rect 2556 18096 2562 18148
rect 7561 18139 7619 18145
rect 7561 18105 7573 18139
rect 7607 18136 7619 18139
rect 7834 18136 7840 18148
rect 7607 18108 7840 18136
rect 7607 18105 7619 18108
rect 7561 18099 7619 18105
rect 7834 18096 7840 18108
rect 7892 18136 7898 18148
rect 12253 18139 12311 18145
rect 7892 18108 8708 18136
rect 7892 18096 7898 18108
rect 4246 18068 4252 18080
rect 4207 18040 4252 18068
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 4338 18028 4344 18080
rect 4396 18068 4402 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4396 18040 4721 18068
rect 4396 18028 4402 18040
rect 4709 18037 4721 18040
rect 4755 18037 4767 18071
rect 5258 18068 5264 18080
rect 5219 18040 5264 18068
rect 4709 18031 4767 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 7466 18068 7472 18080
rect 7427 18040 7472 18068
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 8680 18077 8708 18108
rect 12253 18105 12265 18139
rect 12299 18136 12311 18139
rect 12682 18139 12740 18145
rect 12682 18136 12694 18139
rect 12299 18108 12694 18136
rect 12299 18105 12311 18108
rect 12253 18099 12311 18105
rect 12682 18105 12694 18108
rect 12728 18136 12740 18139
rect 13446 18136 13452 18148
rect 12728 18108 13452 18136
rect 12728 18105 12740 18108
rect 12682 18099 12740 18105
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 20088 18136 20116 18164
rect 20530 18136 20536 18148
rect 20088 18108 20536 18136
rect 20530 18096 20536 18108
rect 20588 18136 20594 18148
rect 20717 18139 20775 18145
rect 20717 18136 20729 18139
rect 20588 18108 20729 18136
rect 20588 18096 20594 18108
rect 20717 18105 20729 18108
rect 20763 18105 20775 18139
rect 26390 18139 26448 18145
rect 26390 18136 26402 18139
rect 20717 18099 20775 18105
rect 25976 18108 26402 18136
rect 8665 18071 8723 18077
rect 8665 18037 8677 18071
rect 8711 18037 8723 18071
rect 8665 18031 8723 18037
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9125 18071 9183 18077
rect 9125 18068 9137 18071
rect 8812 18040 9137 18068
rect 8812 18028 8818 18040
rect 9125 18037 9137 18040
rect 9171 18068 9183 18071
rect 9582 18068 9588 18080
rect 9171 18040 9588 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 13817 18071 13875 18077
rect 13817 18068 13829 18071
rect 13596 18040 13829 18068
rect 13596 18028 13602 18040
rect 13817 18037 13829 18040
rect 13863 18068 13875 18071
rect 14550 18068 14556 18080
rect 13863 18040 14556 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 14550 18028 14556 18040
rect 14608 18028 14614 18080
rect 15286 18068 15292 18080
rect 15247 18040 15292 18068
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 18322 18068 18328 18080
rect 18283 18040 18328 18068
rect 18322 18028 18328 18040
rect 18380 18028 18386 18080
rect 20257 18071 20315 18077
rect 20257 18037 20269 18071
rect 20303 18068 20315 18071
rect 20622 18068 20628 18080
rect 20303 18040 20628 18068
rect 20303 18037 20315 18040
rect 20257 18031 20315 18037
rect 20622 18028 20628 18040
rect 20680 18028 20686 18080
rect 23477 18071 23535 18077
rect 23477 18037 23489 18071
rect 23523 18068 23535 18071
rect 24118 18068 24124 18080
rect 23523 18040 24124 18068
rect 23523 18037 23535 18040
rect 23477 18031 23535 18037
rect 24118 18028 24124 18040
rect 24176 18028 24182 18080
rect 24210 18028 24216 18080
rect 24268 18068 24274 18080
rect 24765 18071 24823 18077
rect 24765 18068 24777 18071
rect 24268 18040 24777 18068
rect 24268 18028 24274 18040
rect 24765 18037 24777 18040
rect 24811 18037 24823 18071
rect 24765 18031 24823 18037
rect 25038 18028 25044 18080
rect 25096 18068 25102 18080
rect 25976 18077 26004 18108
rect 26390 18105 26402 18108
rect 26436 18105 26448 18139
rect 26390 18099 26448 18105
rect 25961 18071 26019 18077
rect 25961 18068 25973 18071
rect 25096 18040 25973 18068
rect 25096 18028 25102 18040
rect 25961 18037 25973 18040
rect 26007 18037 26019 18071
rect 25961 18031 26019 18037
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 2041 17867 2099 17873
rect 2041 17833 2053 17867
rect 2087 17864 2099 17867
rect 2130 17864 2136 17876
rect 2087 17836 2136 17864
rect 2087 17833 2099 17836
rect 2041 17827 2099 17833
rect 2130 17824 2136 17836
rect 2188 17824 2194 17876
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 4338 17864 4344 17876
rect 3927 17836 4344 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4706 17864 4712 17876
rect 4667 17836 4712 17864
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 7101 17867 7159 17873
rect 7101 17833 7113 17867
rect 7147 17864 7159 17867
rect 7466 17864 7472 17876
rect 7147 17836 7472 17864
rect 7147 17833 7159 17836
rect 7101 17827 7159 17833
rect 7466 17824 7472 17836
rect 7524 17864 7530 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7524 17836 8033 17864
rect 7524 17824 7530 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 9674 17864 9680 17876
rect 9635 17836 9680 17864
rect 8021 17827 8079 17833
rect 9674 17824 9680 17836
rect 9732 17824 9738 17876
rect 12434 17824 12440 17876
rect 12492 17864 12498 17876
rect 13722 17864 13728 17876
rect 12492 17836 12537 17864
rect 13683 17836 13728 17864
rect 12492 17824 12498 17836
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14090 17864 14096 17876
rect 14051 17836 14096 17864
rect 14090 17824 14096 17836
rect 14148 17824 14154 17876
rect 14737 17867 14795 17873
rect 14737 17833 14749 17867
rect 14783 17864 14795 17867
rect 15286 17864 15292 17876
rect 14783 17836 15292 17864
rect 14783 17833 14795 17836
rect 14737 17827 14795 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20714 17824 20720 17876
rect 20772 17864 20778 17876
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 20772 17836 21281 17864
rect 20772 17824 20778 17836
rect 21269 17833 21281 17836
rect 21315 17864 21327 17867
rect 22554 17864 22560 17876
rect 21315 17836 22560 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 23477 17867 23535 17873
rect 23477 17833 23489 17867
rect 23523 17864 23535 17867
rect 23842 17864 23848 17876
rect 23523 17836 23848 17864
rect 23523 17833 23535 17836
rect 23477 17827 23535 17833
rect 23842 17824 23848 17836
rect 23900 17864 23906 17876
rect 23937 17867 23995 17873
rect 23937 17864 23949 17867
rect 23900 17836 23949 17864
rect 23900 17824 23906 17836
rect 23937 17833 23949 17836
rect 23983 17833 23995 17867
rect 26234 17864 26240 17876
rect 26195 17836 26240 17864
rect 23937 17827 23995 17833
rect 26234 17824 26240 17836
rect 26292 17824 26298 17876
rect 7834 17796 7840 17808
rect 7795 17768 7840 17796
rect 7834 17756 7840 17768
rect 7892 17756 7898 17808
rect 17221 17799 17279 17805
rect 17221 17765 17233 17799
rect 17267 17796 17279 17799
rect 17310 17796 17316 17808
rect 17267 17768 17316 17796
rect 17267 17765 17279 17768
rect 17221 17759 17279 17765
rect 17310 17756 17316 17768
rect 17368 17756 17374 17808
rect 23753 17799 23811 17805
rect 23753 17765 23765 17799
rect 23799 17796 23811 17799
rect 24026 17796 24032 17808
rect 23799 17768 24032 17796
rect 23799 17765 23811 17768
rect 23753 17759 23811 17765
rect 24026 17756 24032 17768
rect 24084 17796 24090 17808
rect 24670 17796 24676 17808
rect 24084 17768 24676 17796
rect 24084 17756 24090 17768
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1670 17728 1676 17740
rect 1443 17700 1676 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 4062 17688 4068 17740
rect 4120 17728 4126 17740
rect 4801 17731 4859 17737
rect 4801 17728 4813 17731
rect 4120 17700 4813 17728
rect 4120 17688 4126 17700
rect 4801 17697 4813 17700
rect 4847 17728 4859 17731
rect 7469 17731 7527 17737
rect 7469 17728 7481 17731
rect 4847 17700 7481 17728
rect 4847 17697 4859 17700
rect 4801 17691 4859 17697
rect 7469 17697 7481 17700
rect 7515 17728 7527 17731
rect 7926 17728 7932 17740
rect 7515 17700 7932 17728
rect 7515 17697 7527 17700
rect 7469 17691 7527 17697
rect 7926 17688 7932 17700
rect 7984 17688 7990 17740
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8076 17700 8401 17728
rect 8076 17688 8082 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10410 17728 10416 17740
rect 10091 17700 10416 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10410 17688 10416 17700
rect 10468 17688 10474 17740
rect 15654 17728 15660 17740
rect 15615 17700 15660 17728
rect 15654 17688 15660 17700
rect 15712 17688 15718 17740
rect 20622 17688 20628 17740
rect 20680 17728 20686 17740
rect 20717 17731 20775 17737
rect 20717 17728 20729 17731
rect 20680 17700 20729 17728
rect 20680 17688 20686 17700
rect 20717 17697 20729 17700
rect 20763 17728 20775 17731
rect 21818 17728 21824 17740
rect 20763 17700 21824 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 21818 17688 21824 17700
rect 21876 17688 21882 17740
rect 24302 17728 24308 17740
rect 24263 17700 24308 17728
rect 24302 17688 24308 17700
rect 24360 17688 24366 17740
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2409 17663 2467 17669
rect 2409 17660 2421 17663
rect 2372 17632 2421 17660
rect 2372 17620 2378 17632
rect 2409 17629 2421 17632
rect 2455 17660 2467 17663
rect 2682 17660 2688 17672
rect 2455 17632 2688 17660
rect 2455 17629 2467 17632
rect 2409 17623 2467 17629
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 4893 17663 4951 17669
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 5258 17660 5264 17672
rect 4939 17632 5264 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 4154 17552 4160 17604
rect 4212 17592 4218 17604
rect 4908 17592 4936 17623
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8570 17620 8576 17672
rect 8628 17660 8634 17672
rect 10134 17660 10140 17672
rect 8628 17632 8673 17660
rect 10095 17632 10140 17660
rect 8628 17620 8634 17632
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 10778 17660 10784 17672
rect 10367 17632 10784 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 4212 17564 4936 17592
rect 9125 17595 9183 17601
rect 4212 17552 4218 17564
rect 9125 17561 9137 17595
rect 9171 17592 9183 17595
rect 10336 17592 10364 17623
rect 10778 17620 10784 17632
rect 10836 17620 10842 17672
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15562 17660 15568 17672
rect 15151 17632 15568 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15562 17620 15568 17632
rect 15620 17660 15626 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15620 17632 15761 17660
rect 15620 17620 15626 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 15749 17623 15807 17629
rect 15838 17620 15844 17672
rect 15896 17660 15902 17672
rect 15896 17632 15941 17660
rect 15896 17620 15902 17632
rect 17218 17620 17224 17672
rect 17276 17660 17282 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 17276 17632 17325 17660
rect 17276 17620 17282 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 9171 17564 10364 17592
rect 9171 17561 9183 17564
rect 9125 17555 9183 17561
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 17420 17592 17448 17623
rect 20162 17620 20168 17672
rect 20220 17660 20226 17672
rect 20806 17660 20812 17672
rect 20220 17632 20812 17660
rect 20220 17620 20226 17632
rect 20806 17620 20812 17632
rect 20864 17660 20870 17672
rect 21361 17663 21419 17669
rect 21361 17660 21373 17663
rect 20864 17632 21373 17660
rect 20864 17620 20870 17632
rect 21361 17629 21373 17632
rect 21407 17629 21419 17663
rect 21361 17623 21419 17629
rect 21450 17620 21456 17672
rect 21508 17660 21514 17672
rect 24394 17660 24400 17672
rect 21508 17632 21553 17660
rect 24355 17632 24400 17660
rect 21508 17620 21514 17632
rect 24394 17620 24400 17632
rect 24452 17620 24458 17672
rect 24596 17669 24624 17768
rect 24670 17756 24676 17768
rect 24728 17756 24734 17808
rect 26510 17728 26516 17740
rect 26471 17700 26516 17728
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17629 24639 17663
rect 24581 17623 24639 17629
rect 16632 17564 17448 17592
rect 16632 17552 16638 17564
rect 1486 17484 1492 17536
rect 1544 17524 1550 17536
rect 1581 17527 1639 17533
rect 1581 17524 1593 17527
rect 1544 17496 1593 17524
rect 1544 17484 1550 17496
rect 1581 17493 1593 17496
rect 1627 17493 1639 17527
rect 2682 17524 2688 17536
rect 2643 17496 2688 17524
rect 1581 17487 1639 17493
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 5350 17524 5356 17536
rect 5311 17496 5356 17524
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 16850 17524 16856 17536
rect 16811 17496 16856 17524
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18874 17524 18880 17536
rect 18555 17496 18880 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18874 17484 18880 17496
rect 18932 17484 18938 17536
rect 20901 17527 20959 17533
rect 20901 17493 20913 17527
rect 20947 17524 20959 17527
rect 21266 17524 21272 17536
rect 20947 17496 21272 17524
rect 20947 17493 20959 17496
rect 20901 17487 20959 17493
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 25038 17524 25044 17536
rect 24999 17496 25044 17524
rect 25038 17484 25044 17496
rect 25096 17484 25102 17536
rect 26697 17527 26755 17533
rect 26697 17493 26709 17527
rect 26743 17524 26755 17527
rect 26878 17524 26884 17536
rect 26743 17496 26884 17524
rect 26743 17493 26755 17496
rect 26697 17487 26755 17493
rect 26878 17484 26884 17496
rect 26936 17484 26942 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 1670 17320 1676 17332
rect 1583 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17320 1734 17332
rect 4062 17320 4068 17332
rect 1728 17292 4068 17320
rect 1728 17280 1734 17292
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 7745 17323 7803 17329
rect 7745 17289 7757 17323
rect 7791 17320 7803 17323
rect 8478 17320 8484 17332
rect 7791 17292 8484 17320
rect 7791 17289 7803 17292
rect 7745 17283 7803 17289
rect 8478 17280 8484 17292
rect 8536 17320 8542 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8536 17292 9045 17320
rect 8536 17280 8542 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 10778 17320 10784 17332
rect 10739 17292 10784 17320
rect 9033 17283 9091 17289
rect 10778 17280 10784 17292
rect 10836 17280 10842 17332
rect 14550 17320 14556 17332
rect 14511 17292 14556 17320
rect 14550 17280 14556 17292
rect 14608 17320 14614 17332
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14608 17292 14933 17320
rect 14608 17280 14614 17292
rect 14921 17289 14933 17292
rect 14967 17289 14979 17323
rect 14921 17283 14979 17289
rect 1857 17255 1915 17261
rect 1857 17221 1869 17255
rect 1903 17252 1915 17255
rect 5350 17252 5356 17264
rect 1903 17224 5356 17252
rect 1903 17221 1915 17224
rect 1857 17215 1915 17221
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2372 17156 2421 17184
rect 2372 17144 2378 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4706 17184 4712 17196
rect 4479 17156 4712 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 5276 17193 5304 17224
rect 5350 17212 5356 17224
rect 5408 17212 5414 17264
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5813 17187 5871 17193
rect 5813 17184 5825 17187
rect 5491 17156 5825 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 5813 17153 5825 17156
rect 5859 17184 5871 17187
rect 6178 17184 6184 17196
rect 5859 17156 6184 17184
rect 5859 17153 5871 17156
rect 5813 17147 5871 17153
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 8570 17184 8576 17196
rect 8527 17156 8576 17184
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 9398 17144 9404 17196
rect 9456 17184 9462 17196
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 9456 17156 9689 17184
rect 9456 17144 9462 17156
rect 9677 17153 9689 17156
rect 9723 17184 9735 17187
rect 10778 17184 10784 17196
rect 9723 17156 10784 17184
rect 9723 17153 9735 17156
rect 9677 17147 9735 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 14936 17184 14964 17283
rect 15010 17280 15016 17332
rect 15068 17320 15074 17332
rect 15105 17323 15163 17329
rect 15105 17320 15117 17323
rect 15068 17292 15117 17320
rect 15068 17280 15074 17292
rect 15105 17289 15117 17292
rect 15151 17289 15163 17323
rect 15105 17283 15163 17289
rect 15654 17280 15660 17332
rect 15712 17320 15718 17332
rect 16117 17323 16175 17329
rect 16117 17320 16129 17323
rect 15712 17292 16129 17320
rect 15712 17280 15718 17292
rect 16117 17289 16129 17292
rect 16163 17289 16175 17323
rect 18230 17320 18236 17332
rect 18191 17292 18236 17320
rect 16117 17283 16175 17289
rect 18230 17280 18236 17292
rect 18288 17280 18294 17332
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 22554 17320 22560 17332
rect 22515 17292 22560 17320
rect 22554 17280 22560 17292
rect 22612 17280 22618 17332
rect 26510 17320 26516 17332
rect 26471 17292 26516 17320
rect 26510 17280 26516 17292
rect 26568 17280 26574 17332
rect 23109 17255 23167 17261
rect 23109 17221 23121 17255
rect 23155 17252 23167 17255
rect 24302 17252 24308 17264
rect 23155 17224 24308 17252
rect 23155 17221 23167 17224
rect 23109 17215 23167 17221
rect 24302 17212 24308 17224
rect 24360 17252 24366 17264
rect 24489 17255 24547 17261
rect 24489 17252 24501 17255
rect 24360 17224 24501 17252
rect 24360 17212 24366 17224
rect 24489 17221 24501 17224
rect 24535 17221 24547 17255
rect 24489 17215 24547 17221
rect 24946 17212 24952 17264
rect 25004 17252 25010 17264
rect 25314 17252 25320 17264
rect 25004 17224 25320 17252
rect 25004 17212 25010 17224
rect 25314 17212 25320 17224
rect 25372 17212 25378 17264
rect 15657 17187 15715 17193
rect 15657 17184 15669 17187
rect 14936 17156 15669 17184
rect 15657 17153 15669 17156
rect 15703 17184 15715 17187
rect 15838 17184 15844 17196
rect 15703 17156 15844 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 15838 17144 15844 17156
rect 15896 17144 15902 17196
rect 17865 17187 17923 17193
rect 17865 17153 17877 17187
rect 17911 17184 17923 17187
rect 18322 17184 18328 17196
rect 17911 17156 18328 17184
rect 17911 17153 17923 17156
rect 17865 17147 17923 17153
rect 18322 17144 18328 17156
rect 18380 17184 18386 17196
rect 19058 17184 19064 17196
rect 18380 17156 19064 17184
rect 18380 17144 18386 17156
rect 19058 17144 19064 17156
rect 19116 17144 19122 17196
rect 20622 17184 20628 17196
rect 20583 17156 20628 17184
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 25038 17184 25044 17196
rect 24999 17156 25044 17184
rect 25038 17144 25044 17156
rect 25096 17144 25102 17196
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2225 17119 2283 17125
rect 2225 17116 2237 17119
rect 1912 17088 2237 17116
rect 1912 17076 1918 17088
rect 2225 17085 2237 17088
rect 2271 17116 2283 17119
rect 2682 17116 2688 17128
rect 2271 17088 2688 17116
rect 2271 17085 2283 17088
rect 2225 17079 2283 17085
rect 2682 17076 2688 17088
rect 2740 17076 2746 17128
rect 4246 17076 4252 17128
rect 4304 17116 4310 17128
rect 5169 17119 5227 17125
rect 5169 17116 5181 17119
rect 4304 17088 5181 17116
rect 4304 17076 4310 17088
rect 5169 17085 5181 17088
rect 5215 17116 5227 17119
rect 6273 17119 6331 17125
rect 6273 17116 6285 17119
rect 5215 17088 6285 17116
rect 5215 17085 5227 17088
rect 5169 17079 5227 17085
rect 6273 17085 6285 17088
rect 6319 17085 6331 17119
rect 6273 17079 6331 17085
rect 14277 17119 14335 17125
rect 14277 17085 14289 17119
rect 14323 17116 14335 17119
rect 15565 17119 15623 17125
rect 15565 17116 15577 17119
rect 14323 17088 15577 17116
rect 14323 17085 14335 17088
rect 14277 17079 14335 17085
rect 15565 17085 15577 17088
rect 15611 17116 15623 17119
rect 16850 17116 16856 17128
rect 15611 17088 16856 17116
rect 15611 17085 15623 17088
rect 15565 17079 15623 17085
rect 16850 17076 16856 17088
rect 16908 17076 16914 17128
rect 18230 17076 18236 17128
rect 18288 17116 18294 17128
rect 18782 17116 18788 17128
rect 18288 17088 18788 17116
rect 18288 17076 18294 17088
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 18874 17076 18880 17128
rect 18932 17116 18938 17128
rect 18932 17088 18977 17116
rect 18932 17076 18938 17088
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24029 17119 24087 17125
rect 24029 17116 24041 17119
rect 23992 17088 24041 17116
rect 23992 17076 23998 17088
rect 24029 17085 24041 17088
rect 24075 17116 24087 17119
rect 24854 17116 24860 17128
rect 24075 17088 24860 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 24854 17076 24860 17088
rect 24912 17076 24918 17128
rect 9493 17051 9551 17057
rect 9493 17048 9505 17051
rect 8864 17020 9505 17048
rect 8864 16992 8892 17020
rect 9493 17017 9505 17020
rect 9539 17017 9551 17051
rect 9493 17011 9551 17017
rect 9858 17008 9864 17060
rect 9916 17048 9922 17060
rect 16945 17051 17003 17057
rect 16945 17048 16957 17051
rect 9916 17020 16957 17048
rect 9916 17008 9922 17020
rect 16945 17017 16957 17020
rect 16991 17048 17003 17051
rect 17218 17048 17224 17060
rect 16991 17020 17224 17048
rect 16991 17017 17003 17020
rect 16945 17011 17003 17017
rect 17218 17008 17224 17020
rect 17276 17048 17282 17060
rect 17862 17048 17868 17060
rect 17276 17020 17868 17048
rect 17276 17008 17282 17020
rect 17862 17008 17868 17020
rect 17920 17008 17926 17060
rect 20870 17051 20928 17057
rect 20870 17048 20882 17051
rect 20456 17020 20882 17048
rect 20456 16992 20484 17020
rect 20870 17017 20882 17020
rect 20916 17048 20928 17051
rect 21450 17048 21456 17060
rect 20916 17020 21456 17048
rect 20916 17017 20928 17020
rect 20870 17011 20928 17017
rect 21450 17008 21456 17020
rect 21508 17008 21514 17060
rect 23477 17051 23535 17057
rect 23477 17017 23489 17051
rect 23523 17048 23535 17051
rect 24394 17048 24400 17060
rect 23523 17020 24400 17048
rect 23523 17017 23535 17020
rect 23477 17011 23535 17017
rect 24394 17008 24400 17020
rect 24452 17008 24458 17060
rect 24949 17051 25007 17057
rect 24949 17048 24961 17051
rect 24504 17020 24961 17048
rect 2222 16940 2228 16992
rect 2280 16980 2286 16992
rect 2317 16983 2375 16989
rect 2317 16980 2329 16983
rect 2280 16952 2329 16980
rect 2280 16940 2286 16952
rect 2317 16949 2329 16952
rect 2363 16980 2375 16983
rect 2869 16983 2927 16989
rect 2869 16980 2881 16983
rect 2363 16952 2881 16980
rect 2363 16949 2375 16952
rect 2317 16943 2375 16949
rect 2869 16949 2881 16952
rect 2915 16949 2927 16983
rect 2869 16943 2927 16949
rect 4706 16940 4712 16992
rect 4764 16980 4770 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 4764 16952 4813 16980
rect 4764 16940 4770 16952
rect 4801 16949 4813 16952
rect 4847 16949 4859 16983
rect 8018 16980 8024 16992
rect 7979 16952 8024 16980
rect 4801 16943 4859 16949
rect 8018 16940 8024 16952
rect 8076 16940 8082 16992
rect 8846 16980 8852 16992
rect 8807 16952 8852 16980
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9401 16983 9459 16989
rect 9401 16980 9413 16983
rect 9180 16952 9413 16980
rect 9180 16940 9186 16952
rect 9401 16949 9413 16952
rect 9447 16949 9459 16983
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 9401 16943 9459 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10410 16980 10416 16992
rect 10371 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16940 10474 16992
rect 15470 16980 15476 16992
rect 15431 16952 15476 16980
rect 15470 16940 15476 16952
rect 15528 16940 15534 16992
rect 16574 16980 16580 16992
rect 16535 16952 16580 16980
rect 16574 16940 16580 16952
rect 16632 16940 16638 16992
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 18414 16980 18420 16992
rect 18375 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 20438 16980 20444 16992
rect 20399 16952 20444 16980
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 21634 16940 21640 16992
rect 21692 16980 21698 16992
rect 22005 16983 22063 16989
rect 22005 16980 22017 16983
rect 21692 16952 22017 16980
rect 21692 16940 21698 16952
rect 22005 16949 22017 16952
rect 22051 16949 22063 16983
rect 24302 16980 24308 16992
rect 24263 16952 24308 16980
rect 22005 16943 22063 16949
rect 24302 16940 24308 16952
rect 24360 16980 24366 16992
rect 24504 16980 24532 17020
rect 24949 17017 24961 17020
rect 24995 17017 25007 17051
rect 24949 17011 25007 17017
rect 24854 16980 24860 16992
rect 24360 16952 24532 16980
rect 24815 16952 24860 16980
rect 24360 16940 24366 16952
rect 24854 16940 24860 16952
rect 24912 16940 24918 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2314 16776 2320 16788
rect 2275 16748 2320 16776
rect 2314 16736 2320 16748
rect 2372 16736 2378 16788
rect 6178 16776 6184 16788
rect 6139 16748 6184 16776
rect 6178 16736 6184 16748
rect 6236 16736 6242 16788
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 13446 16736 13452 16788
rect 13504 16776 13510 16788
rect 13725 16779 13783 16785
rect 13725 16776 13737 16779
rect 13504 16748 13737 16776
rect 13504 16736 13510 16748
rect 13725 16745 13737 16748
rect 13771 16745 13783 16779
rect 13725 16739 13783 16745
rect 15105 16779 15163 16785
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15470 16776 15476 16788
rect 15151 16748 15476 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 18417 16779 18475 16785
rect 18417 16745 18429 16779
rect 18463 16776 18475 16779
rect 20901 16779 20959 16785
rect 18463 16748 20852 16776
rect 18463 16745 18475 16748
rect 18417 16739 18475 16745
rect 1765 16711 1823 16717
rect 1765 16677 1777 16711
rect 1811 16708 1823 16711
rect 2332 16708 2360 16736
rect 5074 16717 5080 16720
rect 5068 16708 5080 16717
rect 1811 16680 2360 16708
rect 5035 16680 5080 16708
rect 1811 16677 1823 16680
rect 1765 16671 1823 16677
rect 5068 16671 5080 16680
rect 5074 16668 5080 16671
rect 5132 16668 5138 16720
rect 10045 16711 10103 16717
rect 10045 16677 10057 16711
rect 10091 16708 10103 16711
rect 10318 16708 10324 16720
rect 10091 16680 10324 16708
rect 10091 16677 10103 16680
rect 10045 16671 10103 16677
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15933 16711 15991 16717
rect 15933 16708 15945 16711
rect 15344 16680 15945 16708
rect 15344 16668 15350 16680
rect 15933 16677 15945 16680
rect 15979 16677 15991 16711
rect 15933 16671 15991 16677
rect 19334 16668 19340 16720
rect 19392 16708 19398 16720
rect 20438 16708 20444 16720
rect 19392 16680 20444 16708
rect 19392 16668 19398 16680
rect 20438 16668 20444 16680
rect 20496 16708 20502 16720
rect 20625 16711 20683 16717
rect 20625 16708 20637 16711
rect 20496 16680 20637 16708
rect 20496 16668 20502 16680
rect 20625 16677 20637 16680
rect 20671 16677 20683 16711
rect 20625 16671 20683 16677
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 2225 16643 2283 16649
rect 2225 16640 2237 16643
rect 1636 16612 2237 16640
rect 1636 16600 1642 16612
rect 2225 16609 2237 16612
rect 2271 16640 2283 16643
rect 2682 16640 2688 16652
rect 2271 16612 2688 16640
rect 2271 16609 2283 16612
rect 2225 16603 2283 16609
rect 2682 16600 2688 16612
rect 2740 16600 2746 16652
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2792 16612 2973 16640
rect 2498 16572 2504 16584
rect 2459 16544 2504 16572
rect 2498 16532 2504 16544
rect 2556 16532 2562 16584
rect 2792 16572 2820 16612
rect 2961 16609 2973 16612
rect 3007 16640 3019 16643
rect 3007 16612 4108 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 2700 16544 2820 16572
rect 4080 16572 4108 16612
rect 4154 16600 4160 16652
rect 4212 16640 4218 16652
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 4212 16612 4353 16640
rect 4212 16600 4218 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 9122 16640 9128 16652
rect 9083 16612 9128 16640
rect 4341 16603 4399 16609
rect 9122 16600 9128 16612
rect 9180 16600 9186 16652
rect 12342 16640 12348 16652
rect 12303 16612 12348 16640
rect 12342 16600 12348 16612
rect 12400 16600 12406 16652
rect 12434 16600 12440 16652
rect 12492 16640 12498 16652
rect 12612 16643 12670 16649
rect 12612 16640 12624 16643
rect 12492 16612 12624 16640
rect 12492 16600 12498 16612
rect 12612 16609 12624 16612
rect 12658 16640 12670 16643
rect 13722 16640 13728 16652
rect 12658 16612 13728 16640
rect 12658 16609 12670 16612
rect 12612 16603 12670 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 15562 16640 15568 16652
rect 15488 16612 15568 16640
rect 4798 16572 4804 16584
rect 4080 16544 4804 16572
rect 1762 16464 1768 16516
rect 1820 16504 1826 16516
rect 2130 16504 2136 16516
rect 1820 16476 2136 16504
rect 1820 16464 1826 16476
rect 2130 16464 2136 16476
rect 2188 16504 2194 16516
rect 2700 16504 2728 16544
rect 4798 16532 4804 16544
rect 4856 16532 4862 16584
rect 9858 16532 9864 16584
rect 9916 16572 9922 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 9916 16544 10149 16572
rect 9916 16532 9922 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10778 16572 10784 16584
rect 10367 16544 10784 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10778 16532 10784 16544
rect 10836 16532 10842 16584
rect 15488 16513 15516 16612
rect 15562 16600 15568 16612
rect 15620 16600 15626 16652
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16640 15899 16643
rect 15887 16612 16712 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16684 16584 16712 16612
rect 18414 16600 18420 16652
rect 18472 16640 18478 16652
rect 18785 16643 18843 16649
rect 18785 16640 18797 16643
rect 18472 16612 18797 16640
rect 18472 16600 18478 16612
rect 18785 16609 18797 16612
rect 18831 16640 18843 16643
rect 20824 16640 20852 16748
rect 20901 16745 20913 16779
rect 20947 16745 20959 16779
rect 21266 16776 21272 16788
rect 21227 16748 21272 16776
rect 20901 16739 20959 16745
rect 20916 16708 20944 16739
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 24026 16776 24032 16788
rect 23987 16748 24032 16776
rect 24026 16736 24032 16748
rect 24084 16736 24090 16788
rect 24394 16736 24400 16788
rect 24452 16776 24458 16788
rect 24489 16779 24547 16785
rect 24489 16776 24501 16779
rect 24452 16748 24501 16776
rect 24452 16736 24458 16748
rect 24489 16745 24501 16748
rect 24535 16745 24547 16779
rect 24489 16739 24547 16745
rect 21542 16708 21548 16720
rect 20916 16680 21548 16708
rect 21542 16668 21548 16680
rect 21600 16668 21606 16720
rect 24857 16711 24915 16717
rect 24857 16677 24869 16711
rect 24903 16708 24915 16711
rect 25406 16708 25412 16720
rect 24903 16680 25412 16708
rect 24903 16677 24915 16680
rect 24857 16671 24915 16677
rect 25406 16668 25412 16680
rect 25464 16668 25470 16720
rect 21358 16640 21364 16652
rect 18831 16612 19380 16640
rect 20824 16612 21364 16640
rect 18831 16609 18843 16612
rect 18785 16603 18843 16609
rect 16022 16572 16028 16584
rect 15983 16544 16028 16572
rect 16022 16532 16028 16544
rect 16080 16572 16086 16584
rect 16574 16572 16580 16584
rect 16080 16544 16580 16572
rect 16080 16532 16086 16544
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 18874 16572 18880 16584
rect 18835 16544 18880 16572
rect 18874 16532 18880 16544
rect 18932 16532 18938 16584
rect 18969 16575 19027 16581
rect 18969 16541 18981 16575
rect 19015 16541 19027 16575
rect 19352 16572 19380 16612
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 24762 16600 24768 16652
rect 24820 16640 24826 16652
rect 24949 16643 25007 16649
rect 24949 16640 24961 16643
rect 24820 16612 24961 16640
rect 24820 16600 24826 16612
rect 24949 16609 24961 16612
rect 24995 16609 25007 16643
rect 24949 16603 25007 16609
rect 20162 16572 20168 16584
rect 19352 16544 20168 16572
rect 18969 16535 19027 16541
rect 2188 16476 2728 16504
rect 15473 16507 15531 16513
rect 2188 16464 2194 16476
rect 15473 16473 15485 16507
rect 15519 16473 15531 16507
rect 15473 16467 15531 16473
rect 17862 16464 17868 16516
rect 17920 16504 17926 16516
rect 18984 16504 19012 16535
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 21545 16575 21603 16581
rect 21545 16541 21557 16575
rect 21591 16572 21603 16575
rect 21634 16572 21640 16584
rect 21591 16544 21640 16572
rect 21591 16541 21603 16544
rect 21545 16535 21603 16541
rect 21634 16532 21640 16544
rect 21692 16532 21698 16584
rect 25038 16572 25044 16584
rect 24999 16544 25044 16572
rect 25038 16532 25044 16544
rect 25096 16532 25102 16584
rect 19334 16504 19340 16516
rect 17920 16476 19340 16504
rect 17920 16464 17926 16476
rect 19334 16464 19340 16476
rect 19392 16464 19398 16516
rect 24397 16439 24455 16445
rect 24397 16405 24409 16439
rect 24443 16436 24455 16439
rect 24670 16436 24676 16448
rect 24443 16408 24676 16436
rect 24443 16405 24455 16408
rect 24397 16399 24455 16405
rect 24670 16396 24676 16408
rect 24728 16396 24734 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 1578 16192 1584 16244
rect 1636 16232 1642 16244
rect 1857 16235 1915 16241
rect 1857 16232 1869 16235
rect 1636 16204 1869 16232
rect 1636 16192 1642 16204
rect 1857 16201 1869 16204
rect 1903 16201 1915 16235
rect 1857 16195 1915 16201
rect 2498 16192 2504 16244
rect 2556 16232 2562 16244
rect 3605 16235 3663 16241
rect 3605 16232 3617 16235
rect 2556 16204 3617 16232
rect 2556 16192 2562 16204
rect 3605 16201 3617 16204
rect 3651 16232 3663 16235
rect 4154 16232 4160 16244
rect 3651 16204 4160 16232
rect 3651 16201 3663 16204
rect 3605 16195 3663 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 4893 16235 4951 16241
rect 4893 16201 4905 16235
rect 4939 16232 4951 16235
rect 5074 16232 5080 16244
rect 4939 16204 5080 16232
rect 4939 16201 4951 16204
rect 4893 16195 4951 16201
rect 5074 16192 5080 16204
rect 5132 16192 5138 16244
rect 6270 16192 6276 16244
rect 6328 16232 6334 16244
rect 6549 16235 6607 16241
rect 6549 16232 6561 16235
rect 6328 16204 6561 16232
rect 6328 16192 6334 16204
rect 6549 16201 6561 16204
rect 6595 16201 6607 16235
rect 9398 16232 9404 16244
rect 9359 16204 9404 16232
rect 6549 16195 6607 16201
rect 2130 16056 2136 16108
rect 2188 16096 2194 16108
rect 2225 16099 2283 16105
rect 2225 16096 2237 16099
rect 2188 16068 2237 16096
rect 2188 16056 2194 16068
rect 2225 16065 2237 16068
rect 2271 16065 2283 16099
rect 6564 16096 6592 16195
rect 9398 16192 9404 16204
rect 9456 16192 9462 16244
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 12342 16232 12348 16244
rect 12299 16204 12348 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 12342 16192 12348 16204
rect 12400 16192 12406 16244
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 13817 16235 13875 16241
rect 13817 16232 13829 16235
rect 13780 16204 13829 16232
rect 13780 16192 13786 16204
rect 13817 16201 13829 16204
rect 13863 16201 13875 16235
rect 15470 16232 15476 16244
rect 15431 16204 15476 16232
rect 13817 16195 13875 16201
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 16577 16235 16635 16241
rect 16577 16201 16589 16235
rect 16623 16232 16635 16235
rect 16666 16232 16672 16244
rect 16623 16204 16672 16232
rect 16623 16201 16635 16204
rect 16577 16195 16635 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 17862 16232 17868 16244
rect 17823 16204 17868 16232
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 18417 16235 18475 16241
rect 18417 16201 18429 16235
rect 18463 16232 18475 16235
rect 18874 16232 18880 16244
rect 18463 16204 18880 16232
rect 18463 16201 18475 16204
rect 18417 16195 18475 16201
rect 18874 16192 18880 16204
rect 18932 16232 18938 16244
rect 19797 16235 19855 16241
rect 19797 16232 19809 16235
rect 18932 16204 19809 16232
rect 18932 16192 18938 16204
rect 19797 16201 19809 16204
rect 19843 16201 19855 16235
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 19797 16195 19855 16201
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 21266 16192 21272 16244
rect 21324 16232 21330 16244
rect 21637 16235 21695 16241
rect 21637 16232 21649 16235
rect 21324 16204 21649 16232
rect 21324 16192 21330 16204
rect 21637 16201 21649 16204
rect 21683 16201 21695 16235
rect 21637 16195 21695 16201
rect 24210 16192 24216 16244
rect 24268 16232 24274 16244
rect 24305 16235 24363 16241
rect 24305 16232 24317 16235
rect 24268 16204 24317 16232
rect 24268 16192 24274 16204
rect 24305 16201 24317 16204
rect 24351 16201 24363 16235
rect 24305 16195 24363 16201
rect 24762 16192 24768 16244
rect 24820 16232 24826 16244
rect 25317 16235 25375 16241
rect 25317 16232 25329 16235
rect 24820 16204 25329 16232
rect 24820 16192 24826 16204
rect 25317 16201 25329 16204
rect 25363 16201 25375 16235
rect 27249 16235 27307 16241
rect 27249 16232 27261 16235
rect 25317 16195 25375 16201
rect 25424 16204 27261 16232
rect 9861 16167 9919 16173
rect 9861 16133 9873 16167
rect 9907 16133 9919 16167
rect 21358 16164 21364 16176
rect 21319 16136 21364 16164
rect 9861 16127 9919 16133
rect 6564 16068 6960 16096
rect 2225 16059 2283 16065
rect 4798 15988 4804 16040
rect 4856 16028 4862 16040
rect 5261 16031 5319 16037
rect 5261 16028 5273 16031
rect 4856 16000 5273 16028
rect 4856 15988 4862 16000
rect 5261 15997 5273 16000
rect 5307 16028 5319 16031
rect 5442 16028 5448 16040
rect 5307 16000 5448 16028
rect 5307 15997 5319 16000
rect 5261 15991 5319 15997
rect 5442 15988 5448 16000
rect 5500 16028 5506 16040
rect 6822 16028 6828 16040
rect 5500 16000 6828 16028
rect 5500 15988 5506 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6932 16028 6960 16068
rect 9674 16056 9680 16108
rect 9732 16096 9738 16108
rect 9876 16096 9904 16127
rect 21358 16124 21364 16136
rect 21416 16124 21422 16176
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 9732 16068 11529 16096
rect 9732 16056 9738 16068
rect 11517 16065 11529 16068
rect 11563 16096 11575 16099
rect 12250 16096 12256 16108
rect 11563 16068 12256 16096
rect 11563 16065 11575 16068
rect 11517 16059 11575 16065
rect 12250 16056 12256 16068
rect 12308 16096 12314 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12308 16068 12449 16096
rect 12308 16056 12314 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 12437 16059 12495 16065
rect 16117 16099 16175 16105
rect 16117 16065 16129 16099
rect 16163 16096 16175 16099
rect 16574 16096 16580 16108
rect 16163 16068 16580 16096
rect 16163 16065 16175 16068
rect 16117 16059 16175 16065
rect 16574 16056 16580 16068
rect 16632 16096 16638 16108
rect 16853 16099 16911 16105
rect 16853 16096 16865 16099
rect 16632 16068 16865 16096
rect 16632 16056 16638 16068
rect 16853 16065 16865 16068
rect 16899 16096 16911 16099
rect 17221 16099 17279 16105
rect 17221 16096 17233 16099
rect 16899 16068 17233 16096
rect 16899 16065 16911 16068
rect 16853 16059 16911 16065
rect 17221 16065 17233 16068
rect 17267 16065 17279 16099
rect 19058 16096 19064 16108
rect 19019 16068 19064 16096
rect 17221 16059 17279 16065
rect 19058 16056 19064 16068
rect 19116 16056 19122 16108
rect 20993 16099 21051 16105
rect 20993 16065 21005 16099
rect 21039 16096 21051 16099
rect 21634 16096 21640 16108
rect 21039 16068 21640 16096
rect 21039 16065 21051 16068
rect 20993 16059 21051 16065
rect 21634 16056 21640 16068
rect 21692 16056 21698 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 24946 16096 24952 16108
rect 23523 16068 24952 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 24946 16056 24952 16068
rect 25004 16096 25010 16108
rect 25038 16096 25044 16108
rect 25004 16068 25044 16096
rect 25004 16056 25010 16068
rect 25038 16056 25044 16068
rect 25096 16096 25102 16108
rect 25424 16096 25452 16204
rect 27249 16201 27261 16204
rect 27295 16201 27307 16235
rect 27249 16195 27307 16201
rect 25096 16068 25452 16096
rect 25096 16056 25102 16068
rect 25682 16056 25688 16108
rect 25740 16096 25746 16108
rect 25869 16099 25927 16105
rect 25869 16096 25881 16099
rect 25740 16068 25881 16096
rect 25740 16056 25746 16068
rect 25869 16065 25881 16068
rect 25915 16065 25927 16099
rect 25869 16059 25927 16065
rect 7081 16031 7139 16037
rect 7081 16028 7093 16031
rect 6932 16000 7093 16028
rect 7081 15997 7093 16000
rect 7127 15997 7139 16031
rect 7081 15991 7139 15997
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 10045 16031 10103 16037
rect 10045 16028 10057 16031
rect 9640 16000 10057 16028
rect 9640 15988 9646 16000
rect 10045 15997 10057 16000
rect 10091 16028 10103 16031
rect 10689 16031 10747 16037
rect 10689 16028 10701 16031
rect 10091 16000 10701 16028
rect 10091 15997 10103 16000
rect 10045 15991 10103 15997
rect 10689 15997 10701 16000
rect 10735 15997 10747 16031
rect 14642 16028 14648 16040
rect 14555 16000 14648 16028
rect 10689 15991 10747 15997
rect 14642 15988 14648 16000
rect 14700 16028 14706 16040
rect 15841 16031 15899 16037
rect 15841 16028 15853 16031
rect 14700 16000 15853 16028
rect 14700 15988 14706 16000
rect 15841 15997 15853 16000
rect 15887 16028 15899 16031
rect 16390 16028 16396 16040
rect 15887 16000 16396 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 16390 15988 16396 16000
rect 16448 15988 16454 16040
rect 24394 15988 24400 16040
rect 24452 16028 24458 16040
rect 25498 16028 25504 16040
rect 24452 16000 25504 16028
rect 24452 15988 24458 16000
rect 25498 15988 25504 16000
rect 25556 15988 25562 16040
rect 25884 16028 25912 16059
rect 25958 16028 25964 16040
rect 25884 16000 25964 16028
rect 25958 15988 25964 16000
rect 26016 15988 26022 16040
rect 2492 15963 2550 15969
rect 2492 15929 2504 15963
rect 2538 15960 2550 15963
rect 2682 15960 2688 15972
rect 2538 15932 2688 15960
rect 2538 15929 2550 15932
rect 2492 15923 2550 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 11882 15960 11888 15972
rect 10284 15932 11744 15960
rect 11795 15932 11888 15960
rect 10284 15920 10290 15932
rect 8202 15892 8208 15904
rect 8163 15864 8208 15892
rect 8202 15852 8208 15864
rect 8260 15852 8266 15904
rect 9769 15895 9827 15901
rect 9769 15861 9781 15895
rect 9815 15892 9827 15895
rect 9858 15892 9864 15904
rect 9815 15864 9864 15892
rect 9815 15861 9827 15864
rect 9769 15855 9827 15861
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 11716 15892 11744 15932
rect 11882 15920 11888 15932
rect 11940 15960 11946 15972
rect 12682 15963 12740 15969
rect 12682 15960 12694 15963
rect 11940 15932 12694 15960
rect 11940 15920 11946 15932
rect 12682 15929 12694 15932
rect 12728 15929 12740 15963
rect 15378 15960 15384 15972
rect 15291 15932 15384 15960
rect 12682 15923 12740 15929
rect 15378 15920 15384 15932
rect 15436 15960 15442 15972
rect 15933 15963 15991 15969
rect 15933 15960 15945 15963
rect 15436 15932 15945 15960
rect 15436 15920 15442 15932
rect 15933 15929 15945 15932
rect 15979 15960 15991 15963
rect 24765 15963 24823 15969
rect 24765 15960 24777 15963
rect 15979 15932 18368 15960
rect 15979 15929 15991 15932
rect 15933 15923 15991 15929
rect 14921 15895 14979 15901
rect 14921 15892 14933 15895
rect 11716 15864 14933 15892
rect 14921 15861 14933 15864
rect 14967 15892 14979 15895
rect 15286 15892 15292 15904
rect 14967 15864 15292 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 18340 15901 18368 15932
rect 24136 15932 24777 15960
rect 24136 15904 24164 15932
rect 24765 15929 24777 15932
rect 24811 15929 24823 15963
rect 24765 15923 24823 15929
rect 24854 15920 24860 15972
rect 24912 15960 24918 15972
rect 25038 15960 25044 15972
rect 24912 15932 25044 15960
rect 24912 15920 24918 15932
rect 25038 15920 25044 15932
rect 25096 15920 25102 15972
rect 26114 15963 26172 15969
rect 26114 15960 26126 15963
rect 25700 15932 26126 15960
rect 25700 15904 25728 15932
rect 26114 15929 26126 15932
rect 26160 15929 26172 15963
rect 26114 15923 26172 15929
rect 18325 15895 18383 15901
rect 18325 15861 18337 15895
rect 18371 15892 18383 15895
rect 18782 15892 18788 15904
rect 18371 15864 18788 15892
rect 18371 15861 18383 15864
rect 18325 15855 18383 15861
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 18932 15864 19441 15892
rect 18932 15852 18938 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 24118 15892 24124 15904
rect 24079 15864 24124 15892
rect 19429 15855 19487 15861
rect 24118 15852 24124 15864
rect 24176 15852 24182 15904
rect 24670 15892 24676 15904
rect 24631 15864 24676 15892
rect 24670 15852 24676 15864
rect 24728 15852 24734 15904
rect 25682 15892 25688 15904
rect 25643 15864 25688 15892
rect 25682 15852 25688 15864
rect 25740 15852 25746 15904
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 1765 15691 1823 15697
rect 1765 15657 1777 15691
rect 1811 15688 1823 15691
rect 2222 15688 2228 15700
rect 1811 15660 2228 15688
rect 1811 15657 1823 15660
rect 1765 15651 1823 15657
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 11057 15691 11115 15697
rect 11057 15657 11069 15691
rect 11103 15688 11115 15691
rect 11882 15688 11888 15700
rect 11103 15660 11888 15688
rect 11103 15657 11115 15660
rect 11057 15651 11115 15657
rect 11882 15648 11888 15660
rect 11940 15648 11946 15700
rect 12250 15648 12256 15700
rect 12308 15688 12314 15700
rect 12805 15691 12863 15697
rect 12805 15688 12817 15691
rect 12308 15660 12817 15688
rect 12308 15648 12314 15660
rect 12805 15657 12817 15660
rect 12851 15657 12863 15691
rect 18874 15688 18880 15700
rect 18835 15660 18880 15688
rect 12805 15651 12863 15657
rect 18874 15648 18880 15660
rect 18932 15648 18938 15700
rect 24946 15688 24952 15700
rect 24907 15660 24952 15688
rect 24946 15648 24952 15660
rect 25004 15648 25010 15700
rect 25498 15648 25504 15700
rect 25556 15688 25562 15700
rect 25958 15688 25964 15700
rect 25556 15660 25964 15688
rect 25556 15648 25562 15660
rect 25958 15648 25964 15660
rect 26016 15648 26022 15700
rect 2130 15620 2136 15632
rect 2091 15592 2136 15620
rect 2130 15580 2136 15592
rect 2188 15580 2194 15632
rect 15194 15580 15200 15632
rect 15252 15620 15258 15632
rect 15534 15623 15592 15629
rect 15534 15620 15546 15623
rect 15252 15592 15546 15620
rect 15252 15580 15258 15592
rect 15534 15589 15546 15592
rect 15580 15589 15592 15623
rect 15534 15583 15592 15589
rect 17954 15580 17960 15632
rect 18012 15620 18018 15632
rect 19334 15620 19340 15632
rect 18012 15592 19340 15620
rect 18012 15580 18018 15592
rect 19334 15580 19340 15592
rect 19392 15580 19398 15632
rect 21634 15580 21640 15632
rect 21692 15620 21698 15632
rect 22250 15623 22308 15629
rect 22250 15620 22262 15623
rect 21692 15592 22262 15620
rect 21692 15580 21698 15592
rect 22250 15589 22262 15592
rect 22296 15589 22308 15623
rect 22250 15583 22308 15589
rect 1673 15555 1731 15561
rect 1673 15521 1685 15555
rect 1719 15552 1731 15555
rect 7282 15552 7288 15564
rect 1719 15524 2452 15552
rect 7243 15524 7288 15552
rect 1719 15521 1731 15524
rect 1673 15515 1731 15521
rect 2222 15484 2228 15496
rect 2183 15456 2228 15484
rect 2222 15444 2228 15456
rect 2280 15444 2286 15496
rect 2424 15493 2452 15524
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 9674 15552 9680 15564
rect 9635 15524 9680 15552
rect 9674 15512 9680 15524
rect 9732 15512 9738 15564
rect 9950 15561 9956 15564
rect 9944 15552 9956 15561
rect 9911 15524 9956 15552
rect 9944 15515 9956 15524
rect 9950 15512 9956 15515
rect 10008 15512 10014 15564
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 19242 15552 19248 15564
rect 18656 15524 19248 15552
rect 18656 15512 18662 15524
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 21818 15512 21824 15564
rect 21876 15552 21882 15564
rect 22005 15555 22063 15561
rect 22005 15552 22017 15555
rect 21876 15524 22017 15552
rect 21876 15512 21882 15524
rect 22005 15521 22017 15524
rect 22051 15521 22063 15555
rect 22005 15515 22063 15521
rect 24946 15512 24952 15564
rect 25004 15552 25010 15564
rect 25222 15552 25228 15564
rect 25004 15524 25228 15552
rect 25004 15512 25010 15524
rect 25222 15512 25228 15524
rect 25280 15512 25286 15564
rect 26510 15552 26516 15564
rect 26471 15524 26516 15552
rect 26510 15512 26516 15524
rect 26568 15512 26574 15564
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15484 2467 15487
rect 2498 15484 2504 15496
rect 2455 15456 2504 15484
rect 2455 15453 2467 15456
rect 2409 15447 2467 15453
rect 2498 15444 2504 15456
rect 2556 15484 2562 15496
rect 3050 15484 3056 15496
rect 2556 15456 3056 15484
rect 2556 15444 2562 15456
rect 3050 15444 3056 15456
rect 3108 15444 3114 15496
rect 15286 15484 15292 15496
rect 15247 15456 15292 15484
rect 15286 15444 15292 15456
rect 15344 15444 15350 15496
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15484 19579 15487
rect 19610 15484 19616 15496
rect 19567 15456 19616 15484
rect 19567 15453 19579 15456
rect 19521 15447 19579 15453
rect 19610 15444 19616 15456
rect 19668 15444 19674 15496
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2777 15351 2835 15357
rect 2777 15348 2789 15351
rect 2740 15320 2789 15348
rect 2740 15308 2746 15320
rect 2777 15317 2789 15320
rect 2823 15317 2835 15351
rect 2777 15311 2835 15317
rect 6822 15308 6828 15360
rect 6880 15348 6886 15360
rect 6917 15351 6975 15357
rect 6917 15348 6929 15351
rect 6880 15320 6929 15348
rect 6880 15308 6886 15320
rect 6917 15317 6929 15320
rect 6963 15348 6975 15351
rect 7101 15351 7159 15357
rect 7101 15348 7113 15351
rect 6963 15320 7113 15348
rect 6963 15317 6975 15320
rect 6917 15311 6975 15317
rect 7101 15317 7113 15320
rect 7147 15348 7159 15351
rect 7650 15348 7656 15360
rect 7147 15320 7656 15348
rect 7147 15317 7159 15320
rect 7101 15311 7159 15317
rect 7650 15308 7656 15320
rect 7708 15308 7714 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12802 15348 12808 15360
rect 12575 15320 12808 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 16666 15348 16672 15360
rect 16627 15320 16672 15348
rect 16666 15308 16672 15320
rect 16724 15308 16730 15360
rect 18509 15351 18567 15357
rect 18509 15317 18521 15351
rect 18555 15348 18567 15351
rect 19058 15348 19064 15360
rect 18555 15320 19064 15348
rect 18555 15317 18567 15320
rect 18509 15311 18567 15317
rect 19058 15308 19064 15320
rect 19116 15348 19122 15360
rect 20714 15348 20720 15360
rect 19116 15320 20720 15348
rect 19116 15308 19122 15320
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 23382 15348 23388 15360
rect 23343 15320 23388 15348
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 24578 15348 24584 15360
rect 24491 15320 24584 15348
rect 24578 15308 24584 15320
rect 24636 15348 24642 15360
rect 25406 15348 25412 15360
rect 24636 15320 25412 15348
rect 24636 15308 24642 15320
rect 25406 15308 25412 15320
rect 25464 15308 25470 15360
rect 26697 15351 26755 15357
rect 26697 15317 26709 15351
rect 26743 15348 26755 15351
rect 26786 15348 26792 15360
rect 26743 15320 26792 15348
rect 26743 15317 26755 15320
rect 26697 15311 26755 15317
rect 26786 15308 26792 15320
rect 26844 15308 26850 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 7193 15147 7251 15153
rect 7193 15113 7205 15147
rect 7239 15144 7251 15147
rect 7282 15144 7288 15156
rect 7239 15116 7288 15144
rect 7239 15113 7251 15116
rect 7193 15107 7251 15113
rect 7282 15104 7288 15116
rect 7340 15144 7346 15156
rect 9582 15144 9588 15156
rect 7340 15116 9588 15144
rect 7340 15104 7346 15116
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 9674 15104 9680 15156
rect 9732 15144 9738 15156
rect 10045 15147 10103 15153
rect 10045 15144 10057 15147
rect 9732 15116 10057 15144
rect 9732 15104 9738 15116
rect 10045 15113 10057 15116
rect 10091 15113 10103 15147
rect 12158 15144 12164 15156
rect 12119 15116 12164 15144
rect 10045 15107 10103 15113
rect 12158 15104 12164 15116
rect 12216 15104 12222 15156
rect 15194 15144 15200 15156
rect 15155 15116 15200 15144
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 18598 15144 18604 15156
rect 18559 15116 18604 15144
rect 18598 15104 18604 15116
rect 18656 15104 18662 15156
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18748 15116 18797 15144
rect 18748 15104 18754 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 19334 15144 19340 15156
rect 19295 15116 19340 15144
rect 18785 15107 18843 15113
rect 19334 15104 19340 15116
rect 19392 15144 19398 15156
rect 19702 15144 19708 15156
rect 19392 15116 19708 15144
rect 19392 15104 19398 15116
rect 19702 15104 19708 15116
rect 19760 15104 19766 15156
rect 20714 15104 20720 15156
rect 20772 15144 20778 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 20772 15116 20913 15144
rect 20772 15104 20778 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 21634 15104 21640 15156
rect 21692 15144 21698 15156
rect 22005 15147 22063 15153
rect 22005 15144 22017 15147
rect 21692 15116 22017 15144
rect 21692 15104 21698 15116
rect 22005 15113 22017 15116
rect 22051 15113 22063 15147
rect 26510 15144 26516 15156
rect 26471 15116 26516 15144
rect 22005 15107 22063 15113
rect 26510 15104 26516 15116
rect 26568 15104 26574 15156
rect 2041 15079 2099 15085
rect 2041 15045 2053 15079
rect 2087 15076 2099 15079
rect 2222 15076 2228 15088
rect 2087 15048 2228 15076
rect 2087 15045 2099 15048
rect 2041 15039 2099 15045
rect 2222 15036 2228 15048
rect 2280 15076 2286 15088
rect 3421 15079 3479 15085
rect 3421 15076 3433 15079
rect 2280 15048 3433 15076
rect 2280 15036 2286 15048
rect 3421 15045 3433 15048
rect 3467 15045 3479 15079
rect 3421 15039 3479 15045
rect 14461 15079 14519 15085
rect 14461 15045 14473 15079
rect 14507 15076 14519 15079
rect 15286 15076 15292 15088
rect 14507 15048 15292 15076
rect 14507 15045 14519 15048
rect 14461 15039 14519 15045
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 2682 15008 2688 15020
rect 2643 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12636 14980 13001 15008
rect 12636 14952 12664 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 14875 14980 16313 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 16301 14977 16313 14980
rect 16347 15008 16359 15011
rect 16390 15008 16396 15020
rect 16347 14980 16396 15008
rect 16347 14977 16359 14980
rect 16301 14971 16359 14977
rect 16390 14968 16396 14980
rect 16448 15008 16454 15020
rect 16666 15008 16672 15020
rect 16448 14980 16672 15008
rect 16448 14968 16454 14980
rect 16666 14968 16672 14980
rect 16724 14968 16730 15020
rect 7650 14940 7656 14952
rect 7611 14912 7656 14940
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7920 14943 7978 14949
rect 7920 14940 7932 14943
rect 7760 14912 7932 14940
rect 2222 14832 2228 14884
rect 2280 14872 2286 14884
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 2280 14844 2421 14872
rect 2280 14832 2286 14844
rect 2409 14841 2421 14844
rect 2455 14872 2467 14875
rect 2866 14872 2872 14884
rect 2455 14844 2872 14872
rect 2455 14841 2467 14844
rect 2409 14835 2467 14841
rect 2866 14832 2872 14844
rect 2924 14832 2930 14884
rect 7561 14875 7619 14881
rect 7561 14841 7573 14875
rect 7607 14872 7619 14875
rect 7760 14872 7788 14912
rect 7920 14909 7932 14912
rect 7966 14940 7978 14943
rect 8202 14940 8208 14952
rect 7966 14912 8208 14940
rect 7966 14909 7978 14912
rect 7920 14903 7978 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14940 9827 14943
rect 9950 14940 9956 14952
rect 9815 14912 9956 14940
rect 9815 14909 9827 14912
rect 9769 14903 9827 14909
rect 7607 14844 7788 14872
rect 7607 14841 7619 14844
rect 7561 14835 7619 14841
rect 1946 14804 1952 14816
rect 1859 14776 1952 14804
rect 1946 14764 1952 14776
rect 2004 14804 2010 14816
rect 2501 14807 2559 14813
rect 2501 14804 2513 14807
rect 2004 14776 2513 14804
rect 2004 14764 2010 14776
rect 2501 14773 2513 14776
rect 2547 14773 2559 14807
rect 2501 14767 2559 14773
rect 8294 14764 8300 14816
rect 8352 14804 8358 14816
rect 9033 14807 9091 14813
rect 9033 14804 9045 14807
rect 8352 14776 9045 14804
rect 8352 14764 8358 14776
rect 9033 14773 9045 14776
rect 9079 14804 9091 14807
rect 9784 14804 9812 14903
rect 9950 14900 9956 14912
rect 10008 14940 10014 14952
rect 12618 14940 12624 14952
rect 10008 14912 12624 14940
rect 10008 14900 10014 14912
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 12805 14943 12863 14949
rect 12805 14909 12817 14943
rect 12851 14940 12863 14943
rect 12894 14940 12900 14952
rect 12851 14912 12900 14940
rect 12851 14909 12863 14912
rect 12805 14903 12863 14909
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 12820 14872 12848 14903
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 15654 14900 15660 14952
rect 15712 14940 15718 14952
rect 16025 14943 16083 14949
rect 16025 14940 16037 14943
rect 15712 14912 16037 14940
rect 15712 14900 15718 14912
rect 16025 14909 16037 14912
rect 16071 14909 16083 14943
rect 16025 14903 16083 14909
rect 18325 14943 18383 14949
rect 18325 14909 18337 14943
rect 18371 14940 18383 14943
rect 18969 14943 19027 14949
rect 18969 14940 18981 14943
rect 18371 14912 18981 14940
rect 18371 14909 18383 14912
rect 18325 14903 18383 14909
rect 18969 14909 18981 14912
rect 19015 14940 19027 14943
rect 19334 14940 19340 14952
rect 19015 14912 19340 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 19334 14900 19340 14912
rect 19392 14900 19398 14952
rect 19518 14940 19524 14952
rect 19479 14912 19524 14940
rect 19518 14900 19524 14912
rect 19576 14900 19582 14952
rect 12216 14844 12848 14872
rect 15565 14875 15623 14881
rect 12216 14832 12222 14844
rect 15565 14841 15577 14875
rect 15611 14872 15623 14875
rect 15611 14844 16160 14872
rect 15611 14841 15623 14844
rect 15565 14835 15623 14841
rect 9079 14776 9812 14804
rect 11609 14807 11667 14813
rect 9079 14773 9091 14776
rect 9033 14767 9091 14773
rect 11609 14773 11621 14807
rect 11655 14804 11667 14807
rect 11882 14804 11888 14816
rect 11655 14776 11888 14804
rect 11655 14773 11667 14776
rect 11609 14767 11667 14773
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12492 14776 12537 14804
rect 12492 14764 12498 14776
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12860 14776 12909 14804
rect 12860 14764 12866 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 15657 14807 15715 14813
rect 15657 14773 15669 14807
rect 15703 14804 15715 14807
rect 15746 14804 15752 14816
rect 15703 14776 15752 14804
rect 15703 14773 15715 14776
rect 15657 14767 15715 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 16132 14813 16160 14844
rect 19610 14832 19616 14884
rect 19668 14872 19674 14884
rect 19766 14875 19824 14881
rect 19766 14872 19778 14875
rect 19668 14844 19778 14872
rect 19668 14832 19674 14844
rect 19766 14841 19778 14844
rect 19812 14841 19824 14875
rect 19766 14835 19824 14841
rect 16117 14807 16175 14813
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 16482 14804 16488 14816
rect 16163 14776 16488 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 16482 14764 16488 14776
rect 16540 14764 16546 14816
rect 21818 14764 21824 14816
rect 21876 14804 21882 14816
rect 22465 14807 22523 14813
rect 22465 14804 22477 14807
rect 21876 14776 22477 14804
rect 21876 14764 21882 14776
rect 22465 14773 22477 14776
rect 22511 14804 22523 14807
rect 23934 14804 23940 14816
rect 22511 14776 23940 14804
rect 22511 14773 22523 14776
rect 22465 14767 22523 14773
rect 23934 14764 23940 14776
rect 23992 14764 23998 14816
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 2222 14600 2228 14612
rect 2183 14572 2228 14600
rect 2222 14560 2228 14572
rect 2280 14560 2286 14612
rect 2593 14603 2651 14609
rect 2593 14569 2605 14603
rect 2639 14600 2651 14603
rect 2682 14600 2688 14612
rect 2639 14572 2688 14600
rect 2639 14569 2651 14572
rect 2593 14563 2651 14569
rect 2682 14560 2688 14572
rect 2740 14600 2746 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 2740 14572 6377 14600
rect 2740 14560 2746 14572
rect 6365 14569 6377 14572
rect 6411 14569 6423 14603
rect 8294 14600 8300 14612
rect 8255 14572 8300 14600
rect 6365 14563 6423 14569
rect 8294 14560 8300 14572
rect 8352 14560 8358 14612
rect 8849 14603 8907 14609
rect 8849 14569 8861 14603
rect 8895 14600 8907 14603
rect 9582 14600 9588 14612
rect 8895 14572 9588 14600
rect 8895 14569 8907 14572
rect 8849 14563 8907 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 11882 14600 11888 14612
rect 11843 14572 11888 14600
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 17497 14603 17555 14609
rect 17497 14600 17509 14603
rect 16632 14572 17509 14600
rect 16632 14560 16638 14572
rect 17497 14569 17509 14572
rect 17543 14569 17555 14603
rect 17497 14563 17555 14569
rect 19518 14560 19524 14612
rect 19576 14600 19582 14612
rect 19981 14603 20039 14609
rect 19981 14600 19993 14603
rect 19576 14572 19993 14600
rect 19576 14560 19582 14572
rect 19981 14569 19993 14572
rect 20027 14600 20039 14603
rect 20533 14603 20591 14609
rect 20533 14600 20545 14603
rect 20027 14572 20545 14600
rect 20027 14569 20039 14572
rect 19981 14563 20039 14569
rect 20533 14569 20545 14572
rect 20579 14600 20591 14603
rect 21818 14600 21824 14612
rect 20579 14572 21824 14600
rect 20579 14569 20591 14572
rect 20533 14563 20591 14569
rect 1857 14535 1915 14541
rect 1857 14501 1869 14535
rect 1903 14532 1915 14535
rect 2130 14532 2136 14544
rect 1903 14504 2136 14532
rect 1903 14501 1915 14504
rect 1857 14495 1915 14501
rect 2130 14492 2136 14504
rect 2188 14492 2194 14544
rect 5252 14535 5310 14541
rect 5252 14501 5264 14535
rect 5298 14532 5310 14535
rect 5442 14532 5448 14544
rect 5298 14504 5448 14532
rect 5298 14501 5310 14504
rect 5252 14495 5310 14501
rect 5442 14492 5448 14504
rect 5500 14492 5506 14544
rect 15286 14492 15292 14544
rect 15344 14532 15350 14544
rect 16666 14532 16672 14544
rect 15344 14504 16672 14532
rect 15344 14492 15350 14504
rect 2774 14424 2780 14476
rect 2832 14464 2838 14476
rect 2961 14467 3019 14473
rect 2961 14464 2973 14467
rect 2832 14436 2973 14464
rect 2832 14424 2838 14436
rect 2961 14433 2973 14436
rect 3007 14464 3019 14467
rect 4985 14467 5043 14473
rect 4985 14464 4997 14467
rect 3007 14436 4997 14464
rect 3007 14433 3019 14436
rect 2961 14427 3019 14433
rect 4985 14433 4997 14436
rect 5031 14464 5043 14467
rect 5074 14464 5080 14476
rect 5031 14436 5080 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 5074 14424 5080 14436
rect 5132 14424 5138 14476
rect 9030 14464 9036 14476
rect 8991 14436 9036 14464
rect 9030 14424 9036 14436
rect 9088 14424 9094 14476
rect 13449 14467 13507 14473
rect 13449 14433 13461 14467
rect 13495 14464 13507 14467
rect 13722 14464 13728 14476
rect 13495 14436 13728 14464
rect 13495 14433 13507 14436
rect 13449 14427 13507 14433
rect 13722 14424 13728 14436
rect 13780 14424 13786 14476
rect 16132 14473 16160 14504
rect 16666 14492 16672 14504
rect 16724 14532 16730 14544
rect 18782 14532 18788 14544
rect 16724 14504 18788 14532
rect 16724 14492 16730 14504
rect 18782 14492 18788 14504
rect 18840 14492 18846 14544
rect 16390 14473 16396 14476
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14433 16175 14467
rect 16384 14464 16396 14473
rect 16351 14436 16396 14464
rect 16117 14427 16175 14433
rect 16384 14427 16396 14436
rect 16390 14424 16396 14427
rect 16448 14424 16454 14476
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 21468 14473 21496 14572
rect 21818 14560 21824 14572
rect 21876 14560 21882 14612
rect 23382 14532 23388 14544
rect 21735 14504 23388 14532
rect 21735 14476 21763 14504
rect 23382 14492 23388 14504
rect 23440 14492 23446 14544
rect 21726 14473 21732 14476
rect 20717 14467 20775 14473
rect 20717 14464 20729 14467
rect 19392 14436 20729 14464
rect 19392 14424 19398 14436
rect 20717 14433 20729 14436
rect 20763 14433 20775 14467
rect 20717 14427 20775 14433
rect 21453 14467 21511 14473
rect 21453 14433 21465 14467
rect 21499 14433 21511 14467
rect 21453 14427 21511 14433
rect 21720 14427 21732 14473
rect 21784 14464 21790 14476
rect 21784 14436 21868 14464
rect 21726 14424 21732 14427
rect 21784 14424 21790 14436
rect 23290 14424 23296 14476
rect 23348 14464 23354 14476
rect 24193 14467 24251 14473
rect 24193 14464 24205 14467
rect 23348 14436 24205 14464
rect 23348 14424 23354 14436
rect 24193 14433 24205 14436
rect 24239 14433 24251 14467
rect 24193 14427 24251 14433
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 11425 14399 11483 14405
rect 11425 14396 11437 14399
rect 10836 14368 11437 14396
rect 10836 14356 10842 14368
rect 11425 14365 11437 14368
rect 11471 14396 11483 14399
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11471 14368 11989 14396
rect 11471 14365 11483 14368
rect 11425 14359 11483 14365
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12342 14396 12348 14408
rect 12207 14368 12348 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 13538 14396 13544 14408
rect 13499 14368 13544 14396
rect 13538 14356 13544 14368
rect 13596 14356 13602 14408
rect 13633 14399 13691 14405
rect 13633 14365 13645 14399
rect 13679 14365 13691 14399
rect 23934 14396 23940 14408
rect 23895 14368 23940 14396
rect 13633 14359 13691 14365
rect 13648 14328 13676 14359
rect 23934 14356 23940 14368
rect 23992 14356 23998 14408
rect 25038 14356 25044 14408
rect 25096 14396 25102 14408
rect 25774 14396 25780 14408
rect 25096 14368 25780 14396
rect 25096 14356 25102 14368
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 12636 14300 13676 14328
rect 12636 14272 12664 14300
rect 4433 14263 4491 14269
rect 4433 14229 4445 14263
rect 4479 14260 4491 14263
rect 4982 14260 4988 14272
rect 4479 14232 4988 14260
rect 4479 14229 4491 14232
rect 4433 14223 4491 14229
rect 4982 14220 4988 14232
rect 5040 14220 5046 14272
rect 7650 14220 7656 14272
rect 7708 14260 7714 14272
rect 7745 14263 7803 14269
rect 7745 14260 7757 14263
rect 7708 14232 7757 14260
rect 7708 14220 7714 14232
rect 7745 14229 7757 14232
rect 7791 14260 7803 14263
rect 8570 14260 8576 14272
rect 7791 14232 8576 14260
rect 7791 14229 7803 14232
rect 7745 14223 7803 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11054 14260 11060 14272
rect 10919 14232 11060 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11514 14260 11520 14272
rect 11475 14232 11520 14260
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 12618 14260 12624 14272
rect 12579 14232 12624 14260
rect 12618 14220 12624 14232
rect 12676 14220 12682 14272
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 12989 14263 13047 14269
rect 12989 14260 13001 14263
rect 12860 14232 13001 14260
rect 12860 14220 12866 14232
rect 12989 14229 13001 14232
rect 13035 14260 13047 14263
rect 13081 14263 13139 14269
rect 13081 14260 13093 14263
rect 13035 14232 13093 14260
rect 13035 14229 13047 14232
rect 12989 14223 13047 14229
rect 13081 14229 13093 14232
rect 13127 14229 13139 14263
rect 15654 14260 15660 14272
rect 15615 14232 15660 14260
rect 13081 14223 13139 14229
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 18969 14263 19027 14269
rect 18969 14229 18981 14263
rect 19015 14260 19027 14263
rect 19610 14260 19616 14272
rect 19015 14232 19616 14260
rect 19015 14229 19027 14232
rect 18969 14223 19027 14229
rect 19610 14220 19616 14232
rect 19668 14220 19674 14272
rect 22833 14263 22891 14269
rect 22833 14229 22845 14263
rect 22879 14260 22891 14263
rect 23290 14260 23296 14272
rect 22879 14232 23296 14260
rect 22879 14229 22891 14232
rect 22833 14223 22891 14229
rect 23290 14220 23296 14232
rect 23348 14220 23354 14272
rect 25317 14263 25375 14269
rect 25317 14229 25329 14263
rect 25363 14260 25375 14263
rect 25866 14260 25872 14272
rect 25363 14232 25872 14260
rect 25363 14229 25375 14232
rect 25317 14223 25375 14229
rect 25866 14220 25872 14232
rect 25924 14220 25930 14272
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 5813 14059 5871 14065
rect 5813 14056 5825 14059
rect 5132 14028 5825 14056
rect 5132 14016 5138 14028
rect 5813 14025 5825 14028
rect 5859 14056 5871 14059
rect 7650 14056 7656 14068
rect 5859 14028 7656 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 10778 14056 10784 14068
rect 10739 14028 10784 14056
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 11940 14028 12449 14056
rect 11940 14016 11946 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 18782 14056 18788 14068
rect 18743 14028 18788 14056
rect 12437 14019 12495 14025
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19610 14016 19616 14068
rect 19668 14056 19674 14068
rect 20625 14059 20683 14065
rect 20625 14056 20637 14059
rect 19668 14028 20637 14056
rect 19668 14016 19674 14028
rect 20625 14025 20637 14028
rect 20671 14025 20683 14059
rect 21818 14056 21824 14068
rect 21779 14028 21824 14056
rect 20625 14019 20683 14025
rect 21818 14016 21824 14028
rect 21876 14016 21882 14068
rect 3237 13991 3295 13997
rect 3237 13957 3249 13991
rect 3283 13988 3295 13991
rect 4062 13988 4068 14000
rect 3283 13960 4068 13988
rect 3283 13957 3295 13960
rect 3237 13951 3295 13957
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 8202 13988 8208 14000
rect 8163 13960 8208 13988
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 11974 13988 11980 14000
rect 10735 13960 11980 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13852 1915 13855
rect 1903 13824 2820 13852
rect 1903 13821 1915 13824
rect 1857 13815 1915 13821
rect 2792 13796 2820 13824
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3881 13855 3939 13861
rect 3881 13852 3893 13855
rect 2924 13824 3893 13852
rect 2924 13812 2930 13824
rect 3881 13821 3893 13824
rect 3927 13852 3939 13855
rect 4430 13852 4436 13864
rect 3927 13824 4436 13852
rect 3927 13821 3939 13824
rect 3881 13815 3939 13821
rect 4430 13812 4436 13824
rect 4488 13852 4494 13864
rect 4908 13852 4936 13883
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 11440 13929 11468 13960
rect 11974 13948 11980 13960
rect 12032 13988 12038 14000
rect 12161 13991 12219 13997
rect 12161 13988 12173 13991
rect 12032 13960 12173 13988
rect 12032 13948 12038 13960
rect 12161 13957 12173 13960
rect 12207 13988 12219 13991
rect 21545 13991 21603 13997
rect 12207 13960 13032 13988
rect 12207 13957 12219 13960
rect 12161 13951 12219 13957
rect 8757 13923 8815 13929
rect 8757 13920 8769 13923
rect 8352 13892 8769 13920
rect 8352 13880 8358 13892
rect 8757 13889 8769 13892
rect 8803 13889 8815 13923
rect 8757 13883 8815 13889
rect 11425 13923 11483 13929
rect 11425 13889 11437 13923
rect 11471 13889 11483 13923
rect 11425 13883 11483 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12342 13920 12348 13932
rect 11931 13892 12348 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 12434 13880 12440 13932
rect 12492 13920 12498 13932
rect 13004 13929 13032 13960
rect 21545 13957 21557 13991
rect 21591 13988 21603 13991
rect 21726 13988 21732 14000
rect 21591 13960 21732 13988
rect 21591 13957 21603 13960
rect 21545 13951 21603 13957
rect 21726 13948 21732 13960
rect 21784 13948 21790 14000
rect 23934 13948 23940 14000
rect 23992 13988 23998 14000
rect 27430 13988 27436 14000
rect 23992 13960 24440 13988
rect 27391 13960 27436 13988
rect 23992 13948 23998 13960
rect 12897 13923 12955 13929
rect 12897 13920 12909 13923
rect 12492 13892 12909 13920
rect 12492 13880 12498 13892
rect 12897 13889 12909 13892
rect 12943 13889 12955 13923
rect 12897 13883 12955 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13889 13047 13923
rect 12989 13883 13047 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 16390 13920 16396 13932
rect 14967 13892 16396 13920
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 16390 13880 16396 13892
rect 16448 13920 16454 13932
rect 24412 13929 24440 13960
rect 27430 13948 27436 13960
rect 27488 13948 27494 14000
rect 19153 13923 19211 13929
rect 16448 13892 16896 13920
rect 16448 13880 16454 13892
rect 5442 13852 5448 13864
rect 4488 13824 4936 13852
rect 5403 13824 5448 13852
rect 4488 13812 4494 13824
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 7466 13812 7472 13864
rect 7524 13852 7530 13864
rect 7745 13855 7803 13861
rect 7745 13852 7757 13855
rect 7524 13824 7757 13852
rect 7524 13812 7530 13824
rect 7745 13821 7757 13824
rect 7791 13852 7803 13855
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 7791 13824 8677 13852
rect 7791 13821 7803 13824
rect 7745 13815 7803 13821
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 11241 13855 11299 13861
rect 11241 13852 11253 13855
rect 8665 13815 8723 13821
rect 10980 13824 11253 13852
rect 2102 13787 2160 13793
rect 2102 13784 2114 13787
rect 1780 13756 2114 13784
rect 1780 13728 1808 13756
rect 2102 13753 2114 13756
rect 2148 13753 2160 13787
rect 2102 13747 2160 13753
rect 2774 13744 2780 13796
rect 2832 13744 2838 13796
rect 4246 13784 4252 13796
rect 4159 13756 4252 13784
rect 4246 13744 4252 13756
rect 4304 13784 4310 13796
rect 4709 13787 4767 13793
rect 4304 13756 4660 13784
rect 4304 13744 4310 13756
rect 1762 13716 1768 13728
rect 1723 13688 1768 13716
rect 1762 13676 1768 13688
rect 1820 13676 1826 13728
rect 4338 13716 4344 13728
rect 4299 13688 4344 13716
rect 4338 13676 4344 13688
rect 4396 13676 4402 13728
rect 4632 13716 4660 13756
rect 4709 13753 4721 13787
rect 4755 13784 4767 13787
rect 4982 13784 4988 13796
rect 4755 13756 4988 13784
rect 4755 13753 4767 13756
rect 4709 13747 4767 13753
rect 4982 13744 4988 13756
rect 5040 13744 5046 13796
rect 8386 13744 8392 13796
rect 8444 13784 8450 13796
rect 9030 13784 9036 13796
rect 8444 13756 9036 13784
rect 8444 13744 8450 13756
rect 9030 13744 9036 13756
rect 9088 13784 9094 13796
rect 9217 13787 9275 13793
rect 9217 13784 9229 13787
rect 9088 13756 9229 13784
rect 9088 13744 9094 13756
rect 9217 13753 9229 13756
rect 9263 13753 9275 13787
rect 9217 13747 9275 13753
rect 10778 13744 10784 13796
rect 10836 13784 10842 13796
rect 10980 13784 11008 13824
rect 11241 13821 11253 13824
rect 11287 13821 11299 13855
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 11241 13815 11299 13821
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13722 13812 13728 13864
rect 13780 13852 13786 13864
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 13780 13824 13829 13852
rect 13780 13812 13786 13824
rect 13817 13821 13829 13824
rect 13863 13821 13875 13855
rect 15562 13852 15568 13864
rect 15523 13824 15568 13852
rect 13817 13815 13875 13821
rect 15562 13812 15568 13824
rect 15620 13852 15626 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 15620 13824 16221 13852
rect 15620 13812 15626 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 10836 13756 11008 13784
rect 10836 13744 10842 13756
rect 11054 13744 11060 13796
rect 11112 13784 11118 13796
rect 11149 13787 11207 13793
rect 11149 13784 11161 13787
rect 11112 13756 11161 13784
rect 11112 13744 11118 13756
rect 11149 13753 11161 13756
rect 11195 13784 11207 13787
rect 11330 13784 11336 13796
rect 11195 13756 11336 13784
rect 11195 13753 11207 13756
rect 11149 13747 11207 13753
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 15286 13784 15292 13796
rect 15199 13756 15292 13784
rect 15286 13744 15292 13756
rect 15344 13784 15350 13796
rect 16117 13787 16175 13793
rect 16117 13784 16129 13787
rect 15344 13756 16129 13784
rect 15344 13744 15350 13756
rect 16117 13753 16129 13756
rect 16163 13784 16175 13787
rect 16298 13784 16304 13796
rect 16163 13756 16304 13784
rect 16163 13753 16175 13756
rect 16117 13747 16175 13753
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 4801 13719 4859 13725
rect 4801 13716 4813 13719
rect 4632 13688 4813 13716
rect 4801 13685 4813 13688
rect 4847 13716 4859 13719
rect 5626 13716 5632 13728
rect 4847 13688 5632 13716
rect 4847 13685 4859 13688
rect 4801 13679 4859 13685
rect 5626 13676 5632 13688
rect 5684 13676 5690 13728
rect 8113 13719 8171 13725
rect 8113 13685 8125 13719
rect 8159 13716 8171 13719
rect 8202 13716 8208 13728
rect 8159 13688 8208 13716
rect 8159 13685 8171 13688
rect 8113 13679 8171 13685
rect 8202 13676 8208 13688
rect 8260 13716 8266 13728
rect 8573 13719 8631 13725
rect 8573 13716 8585 13719
rect 8260 13688 8585 13716
rect 8260 13676 8266 13688
rect 8573 13685 8585 13688
rect 8619 13716 8631 13719
rect 9582 13716 9588 13728
rect 8619 13688 9588 13716
rect 8619 13685 8631 13688
rect 8573 13679 8631 13685
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 12250 13676 12256 13728
rect 12308 13716 12314 13728
rect 13449 13719 13507 13725
rect 13449 13716 13461 13719
rect 12308 13688 13461 13716
rect 12308 13676 12314 13688
rect 13449 13685 13461 13688
rect 13495 13716 13507 13719
rect 13538 13716 13544 13728
rect 13495 13688 13544 13716
rect 13495 13685 13507 13688
rect 13449 13679 13507 13685
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 15654 13676 15660 13728
rect 15712 13716 15718 13728
rect 16868 13725 16896 13892
rect 19153 13889 19165 13923
rect 19199 13920 19211 13923
rect 24397 13923 24455 13929
rect 19199 13892 19380 13920
rect 19199 13889 19211 13892
rect 19153 13883 19211 13889
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 18840 13824 19257 13852
rect 18840 13812 18846 13824
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19352 13852 19380 13892
rect 24397 13889 24409 13923
rect 24443 13920 24455 13923
rect 25498 13920 25504 13932
rect 24443 13892 25504 13920
rect 24443 13889 24455 13892
rect 24397 13883 24455 13889
rect 25498 13880 25504 13892
rect 25556 13920 25562 13932
rect 26050 13920 26056 13932
rect 25556 13892 26056 13920
rect 25556 13880 25562 13892
rect 26050 13880 26056 13892
rect 26108 13880 26114 13932
rect 19518 13861 19524 13864
rect 19512 13852 19524 13861
rect 19352 13824 19524 13852
rect 19245 13815 19303 13821
rect 19512 13815 19524 13824
rect 19260 13784 19288 13815
rect 19518 13812 19524 13815
rect 19576 13812 19582 13864
rect 23290 13812 23296 13864
rect 23348 13852 23354 13864
rect 23937 13855 23995 13861
rect 23937 13852 23949 13855
rect 23348 13824 23949 13852
rect 23348 13812 23354 13824
rect 23937 13821 23949 13824
rect 23983 13821 23995 13855
rect 26309 13855 26367 13861
rect 26309 13852 26321 13855
rect 23937 13815 23995 13821
rect 26160 13824 26321 13852
rect 19426 13784 19432 13796
rect 19260 13756 19432 13784
rect 19426 13744 19432 13756
rect 19484 13744 19490 13796
rect 26160 13784 26188 13824
rect 26309 13821 26321 13824
rect 26355 13821 26367 13855
rect 26309 13815 26367 13821
rect 25884 13756 26188 13784
rect 25884 13728 25912 13756
rect 15749 13719 15807 13725
rect 15749 13716 15761 13719
rect 15712 13688 15761 13716
rect 15712 13676 15718 13688
rect 15749 13685 15761 13688
rect 15795 13685 15807 13719
rect 15749 13679 15807 13685
rect 16853 13719 16911 13725
rect 16853 13685 16865 13719
rect 16899 13716 16911 13719
rect 17586 13716 17592 13728
rect 16899 13688 17592 13716
rect 16899 13685 16911 13688
rect 16853 13679 16911 13685
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 25866 13716 25872 13728
rect 25827 13688 25872 13716
rect 25866 13676 25872 13688
rect 25924 13676 25930 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 1762 13512 1768 13524
rect 1675 13484 1768 13512
rect 1762 13472 1768 13484
rect 1820 13512 1826 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 1820 13484 2697 13512
rect 1820 13472 1826 13484
rect 2685 13481 2697 13484
rect 2731 13512 2743 13515
rect 2866 13512 2872 13524
rect 2731 13484 2872 13512
rect 2731 13481 2743 13484
rect 2685 13475 2743 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4580 13484 4629 13512
rect 4580 13472 4586 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 4617 13475 4675 13481
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 10778 13512 10784 13524
rect 10739 13484 10784 13512
rect 10778 13472 10784 13484
rect 10836 13472 10842 13524
rect 11241 13515 11299 13521
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11330 13512 11336 13524
rect 11287 13484 11336 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12805 13515 12863 13521
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 13722 13512 13728 13524
rect 12851 13484 13728 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 15105 13515 15163 13521
rect 15105 13481 15117 13515
rect 15151 13512 15163 13515
rect 15657 13515 15715 13521
rect 15657 13512 15669 13515
rect 15151 13484 15669 13512
rect 15151 13481 15163 13484
rect 15105 13475 15163 13481
rect 15657 13481 15669 13484
rect 15703 13512 15715 13515
rect 16853 13515 16911 13521
rect 16853 13512 16865 13515
rect 15703 13484 16865 13512
rect 15703 13481 15715 13484
rect 15657 13475 15715 13481
rect 16853 13481 16865 13484
rect 16899 13481 16911 13515
rect 16853 13475 16911 13481
rect 19334 13472 19340 13524
rect 19392 13512 19398 13524
rect 19705 13515 19763 13521
rect 19705 13512 19717 13515
rect 19392 13484 19717 13512
rect 19392 13472 19398 13484
rect 19705 13481 19717 13484
rect 19751 13512 19763 13515
rect 20533 13515 20591 13521
rect 20533 13512 20545 13515
rect 19751 13484 20545 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 20533 13481 20545 13484
rect 20579 13481 20591 13515
rect 26050 13512 26056 13524
rect 26011 13484 26056 13512
rect 20533 13475 20591 13481
rect 26050 13472 26056 13484
rect 26108 13472 26114 13524
rect 2317 13447 2375 13453
rect 2317 13413 2329 13447
rect 2363 13444 2375 13447
rect 2958 13444 2964 13456
rect 2363 13416 2964 13444
rect 2363 13413 2375 13416
rect 2317 13407 2375 13413
rect 2958 13404 2964 13416
rect 3016 13404 3022 13456
rect 15194 13404 15200 13456
rect 15252 13444 15258 13456
rect 15746 13444 15752 13456
rect 15252 13416 15752 13444
rect 15252 13404 15258 13416
rect 15746 13404 15752 13416
rect 15804 13404 15810 13456
rect 16393 13447 16451 13453
rect 16393 13413 16405 13447
rect 16439 13444 16451 13447
rect 16666 13444 16672 13456
rect 16439 13416 16672 13444
rect 16439 13413 16451 13416
rect 16393 13407 16451 13413
rect 16666 13404 16672 13416
rect 16724 13404 16730 13456
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 19521 13447 19579 13453
rect 19521 13444 19533 13447
rect 19484 13416 19533 13444
rect 19484 13404 19490 13416
rect 19521 13413 19533 13416
rect 19567 13413 19579 13447
rect 19521 13407 19579 13413
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 3326 13376 3332 13388
rect 2271 13348 3332 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 3326 13336 3332 13348
rect 3384 13336 3390 13388
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 7834 13376 7840 13388
rect 4212 13348 4844 13376
rect 7795 13348 7840 13376
rect 4212 13336 4218 13348
rect 2498 13308 2504 13320
rect 2411 13280 2504 13308
rect 2498 13268 2504 13280
rect 2556 13308 2562 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2556 13280 2697 13308
rect 2556 13268 2562 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 4338 13268 4344 13320
rect 4396 13308 4402 13320
rect 4816 13317 4844 13348
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 7984 13348 8029 13376
rect 7984 13336 7990 13348
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 11296 13348 11621 13376
rect 11296 13336 11302 13348
rect 11609 13345 11621 13348
rect 11655 13345 11667 13379
rect 17218 13376 17224 13388
rect 17179 13348 17224 13376
rect 11609 13339 11667 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 19978 13376 19984 13388
rect 19935 13348 19984 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 19978 13336 19984 13348
rect 20036 13336 20042 13388
rect 22741 13379 22799 13385
rect 22741 13345 22753 13379
rect 22787 13376 22799 13379
rect 22922 13376 22928 13388
rect 22787 13348 22928 13376
rect 22787 13345 22799 13348
rect 22741 13339 22799 13345
rect 22922 13336 22928 13348
rect 22980 13336 22986 13388
rect 4709 13311 4767 13317
rect 4709 13308 4721 13311
rect 4396 13280 4721 13308
rect 4396 13268 4402 13280
rect 4709 13277 4721 13280
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5074 13308 5080 13320
rect 4847 13280 5080 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7742 13308 7748 13320
rect 7616 13280 7748 13308
rect 7616 13268 7622 13280
rect 7742 13268 7748 13280
rect 7800 13308 7806 13320
rect 7944 13308 7972 13336
rect 8110 13308 8116 13320
rect 7800 13280 7972 13308
rect 8071 13280 8116 13308
rect 7800 13268 7806 13280
rect 8110 13268 8116 13280
rect 8168 13268 8174 13320
rect 11698 13308 11704 13320
rect 11659 13280 11704 13308
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11885 13311 11943 13317
rect 11885 13277 11897 13311
rect 11931 13308 11943 13311
rect 12066 13308 12072 13320
rect 11931 13280 12072 13308
rect 11931 13277 11943 13280
rect 11885 13271 11943 13277
rect 12066 13268 12072 13280
rect 12124 13308 12130 13320
rect 12618 13308 12624 13320
rect 12124 13280 12624 13308
rect 12124 13268 12130 13280
rect 12618 13268 12624 13280
rect 12676 13308 12682 13320
rect 13265 13311 13323 13317
rect 13265 13308 13277 13311
rect 12676 13280 13277 13308
rect 12676 13268 12682 13280
rect 13265 13277 13277 13280
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16482 13308 16488 13320
rect 15979 13280 16488 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 17313 13311 17371 13317
rect 17313 13277 17325 13311
rect 17359 13308 17371 13311
rect 17402 13308 17408 13320
rect 17359 13280 17408 13308
rect 17359 13277 17371 13280
rect 17313 13271 17371 13277
rect 17402 13268 17408 13280
rect 17460 13268 17466 13320
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13308 17555 13311
rect 17586 13308 17592 13320
rect 17543 13280 17592 13308
rect 17543 13277 17555 13280
rect 17497 13271 17555 13277
rect 17586 13268 17592 13280
rect 17644 13268 17650 13320
rect 22278 13268 22284 13320
rect 22336 13308 22342 13320
rect 22833 13311 22891 13317
rect 22833 13308 22845 13311
rect 22336 13280 22845 13308
rect 22336 13268 22342 13280
rect 22833 13277 22845 13280
rect 22879 13277 22891 13311
rect 22833 13271 22891 13277
rect 23017 13311 23075 13317
rect 23017 13277 23029 13311
rect 23063 13308 23075 13311
rect 23382 13308 23388 13320
rect 23063 13280 23388 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23382 13268 23388 13280
rect 23440 13268 23446 13320
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 3786 13172 3792 13184
rect 3747 13144 3792 13172
rect 3786 13132 3792 13144
rect 3844 13132 3850 13184
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 4249 13135 4307 13141
rect 15289 13175 15347 13181
rect 15289 13141 15301 13175
rect 15335 13172 15347 13175
rect 15746 13172 15752 13184
rect 15335 13144 15752 13172
rect 15335 13141 15347 13144
rect 15289 13135 15347 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 22370 13172 22376 13184
rect 22331 13144 22376 13172
rect 22370 13132 22376 13144
rect 22428 13132 22434 13184
rect 24210 13172 24216 13184
rect 24171 13144 24216 13172
rect 24210 13132 24216 13144
rect 24268 13132 24274 13184
rect 25774 13172 25780 13184
rect 25735 13144 25780 13172
rect 25774 13132 25780 13144
rect 25832 13132 25838 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 2958 12968 2964 12980
rect 2919 12940 2964 12968
rect 2958 12928 2964 12940
rect 3016 12928 3022 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4580 12940 4721 12968
rect 4580 12928 4586 12940
rect 4709 12937 4721 12940
rect 4755 12937 4767 12971
rect 5074 12968 5080 12980
rect 5035 12940 5080 12968
rect 4709 12931 4767 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 7558 12968 7564 12980
rect 7519 12940 7564 12968
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 7834 12968 7840 12980
rect 7795 12940 7840 12968
rect 7834 12928 7840 12940
rect 7892 12928 7898 12980
rect 12066 12968 12072 12980
rect 12027 12940 12072 12968
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 16482 12968 16488 12980
rect 16347 12940 16488 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 566 12860 572 12912
rect 624 12900 630 12912
rect 7006 12900 7012 12912
rect 624 12872 7012 12900
rect 624 12860 630 12872
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 7193 12903 7251 12909
rect 7193 12869 7205 12903
rect 7239 12900 7251 12903
rect 8110 12900 8116 12912
rect 7239 12872 8116 12900
rect 7239 12869 7251 12872
rect 7193 12863 7251 12869
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12832 1823 12835
rect 2314 12832 2320 12844
rect 1811 12804 2320 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2314 12792 2320 12804
rect 2372 12792 2378 12844
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4249 12835 4307 12841
rect 4249 12832 4261 12835
rect 3936 12804 4261 12832
rect 3936 12792 3942 12804
rect 4249 12801 4261 12804
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 14369 12835 14427 12841
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 15654 12832 15660 12844
rect 14415 12804 15660 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 15841 12835 15899 12841
rect 15841 12801 15853 12835
rect 15887 12832 15899 12835
rect 16316 12832 16344 12931
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 17586 12968 17592 12980
rect 17547 12940 17592 12968
rect 17586 12928 17592 12940
rect 17644 12928 17650 12980
rect 22278 12928 22284 12980
rect 22336 12968 22342 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 22336 12940 22385 12968
rect 22336 12928 22342 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 22373 12931 22431 12937
rect 23201 12971 23259 12977
rect 23201 12937 23213 12971
rect 23247 12968 23259 12971
rect 23382 12968 23388 12980
rect 23247 12940 23388 12968
rect 23247 12937 23259 12940
rect 23201 12931 23259 12937
rect 23382 12928 23388 12940
rect 23440 12928 23446 12980
rect 22002 12860 22008 12912
rect 22060 12900 22066 12912
rect 22833 12903 22891 12909
rect 22833 12900 22845 12903
rect 22060 12872 22845 12900
rect 22060 12860 22066 12872
rect 22833 12869 22845 12872
rect 22879 12900 22891 12903
rect 22922 12900 22928 12912
rect 22879 12872 22928 12900
rect 22879 12869 22891 12872
rect 22833 12863 22891 12869
rect 22922 12860 22928 12872
rect 22980 12860 22986 12912
rect 24121 12903 24179 12909
rect 24121 12869 24133 12903
rect 24167 12900 24179 12903
rect 24946 12900 24952 12912
rect 24167 12872 24952 12900
rect 24167 12869 24179 12872
rect 24121 12863 24179 12869
rect 24946 12860 24952 12872
rect 25004 12860 25010 12912
rect 18966 12832 18972 12844
rect 15887 12804 16344 12832
rect 18927 12804 18972 12832
rect 15887 12801 15899 12804
rect 15841 12795 15899 12801
rect 18966 12792 18972 12804
rect 19024 12792 19030 12844
rect 19058 12792 19064 12844
rect 19116 12832 19122 12844
rect 19426 12832 19432 12844
rect 19116 12804 19432 12832
rect 19116 12792 19122 12804
rect 19426 12792 19432 12804
rect 19484 12832 19490 12844
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 19484 12804 19533 12832
rect 19484 12792 19490 12804
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 24029 12835 24087 12841
rect 24029 12801 24041 12835
rect 24075 12832 24087 12835
rect 24673 12835 24731 12841
rect 24673 12832 24685 12835
rect 24075 12804 24685 12832
rect 24075 12801 24087 12804
rect 24029 12795 24087 12801
rect 24673 12801 24685 12804
rect 24719 12832 24731 12835
rect 25501 12835 25559 12841
rect 25501 12832 25513 12835
rect 24719 12804 25513 12832
rect 24719 12801 24731 12804
rect 24673 12795 24731 12801
rect 25501 12801 25513 12804
rect 25547 12832 25559 12835
rect 25866 12832 25872 12844
rect 25547 12804 25872 12832
rect 25547 12801 25559 12804
rect 25501 12795 25559 12801
rect 25866 12792 25872 12804
rect 25924 12832 25930 12844
rect 26237 12835 26295 12841
rect 26237 12832 26249 12835
rect 25924 12804 26249 12832
rect 25924 12792 25930 12804
rect 26237 12801 26249 12804
rect 26283 12801 26295 12835
rect 26237 12795 26295 12801
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12733 2283 12767
rect 2225 12727 2283 12733
rect 4065 12767 4123 12773
rect 4065 12733 4077 12767
rect 4111 12764 4123 12767
rect 4154 12764 4160 12776
rect 4111 12736 4160 12764
rect 4111 12733 4123 12736
rect 4065 12727 4123 12733
rect 2240 12696 2268 12727
rect 4154 12724 4160 12736
rect 4212 12764 4218 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 4212 12736 5457 12764
rect 4212 12724 4218 12736
rect 5445 12733 5457 12736
rect 5491 12733 5503 12767
rect 8570 12764 8576 12776
rect 8531 12736 8576 12764
rect 5445 12727 5503 12733
rect 8570 12724 8576 12736
rect 8628 12724 8634 12776
rect 11238 12764 11244 12776
rect 11199 12736 11244 12764
rect 11238 12724 11244 12736
rect 11296 12724 11302 12776
rect 11698 12764 11704 12776
rect 11611 12736 11704 12764
rect 11698 12724 11704 12736
rect 11756 12764 11762 12776
rect 17218 12764 17224 12776
rect 11756 12736 17224 12764
rect 11756 12724 11762 12736
rect 17218 12724 17224 12736
rect 17276 12724 17282 12776
rect 19777 12767 19835 12773
rect 19777 12764 19789 12767
rect 19628 12736 19789 12764
rect 2314 12696 2320 12708
rect 2240 12668 2320 12696
rect 2314 12656 2320 12668
rect 2372 12656 2378 12708
rect 2774 12656 2780 12708
rect 2832 12696 2838 12708
rect 3786 12696 3792 12708
rect 2832 12668 3792 12696
rect 2832 12656 2838 12668
rect 3786 12656 3792 12668
rect 3844 12696 3850 12708
rect 8481 12699 8539 12705
rect 3844 12668 4108 12696
rect 3844 12656 3850 12668
rect 1857 12631 1915 12637
rect 1857 12597 1869 12631
rect 1903 12628 1915 12631
rect 2038 12628 2044 12640
rect 1903 12600 2044 12628
rect 1903 12597 1915 12600
rect 1857 12591 1915 12597
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 3326 12628 3332 12640
rect 3287 12600 3332 12628
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 3697 12631 3755 12637
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 3970 12628 3976 12640
rect 3743 12600 3976 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 3970 12588 3976 12600
rect 4028 12588 4034 12640
rect 4080 12628 4108 12668
rect 8481 12665 8493 12699
rect 8527 12696 8539 12699
rect 8818 12699 8876 12705
rect 8818 12696 8830 12699
rect 8527 12668 8830 12696
rect 8527 12665 8539 12668
rect 8481 12659 8539 12665
rect 8818 12665 8830 12668
rect 8864 12696 8876 12699
rect 8938 12696 8944 12708
rect 8864 12668 8944 12696
rect 8864 12665 8876 12668
rect 8818 12659 8876 12665
rect 8938 12656 8944 12668
rect 8996 12656 9002 12708
rect 15010 12696 15016 12708
rect 14971 12668 15016 12696
rect 15010 12656 15016 12668
rect 15068 12696 15074 12708
rect 15565 12699 15623 12705
rect 15565 12696 15577 12699
rect 15068 12668 15577 12696
rect 15068 12656 15074 12668
rect 15565 12665 15577 12668
rect 15611 12696 15623 12699
rect 16574 12696 16580 12708
rect 15611 12668 16580 12696
rect 15611 12665 15623 12668
rect 15565 12659 15623 12665
rect 16574 12656 16580 12668
rect 16632 12656 16638 12708
rect 16945 12699 17003 12705
rect 16945 12665 16957 12699
rect 16991 12696 17003 12699
rect 17402 12696 17408 12708
rect 16991 12668 17408 12696
rect 16991 12665 17003 12668
rect 16945 12659 17003 12665
rect 17402 12656 17408 12668
rect 17460 12696 17466 12708
rect 18874 12696 18880 12708
rect 17460 12668 18880 12696
rect 17460 12656 17466 12668
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 19628 12640 19656 12736
rect 19777 12733 19789 12736
rect 19823 12733 19835 12767
rect 19777 12727 19835 12733
rect 24210 12724 24216 12776
rect 24268 12764 24274 12776
rect 24489 12767 24547 12773
rect 24489 12764 24501 12767
rect 24268 12736 24501 12764
rect 24268 12724 24274 12736
rect 24489 12733 24501 12736
rect 24535 12733 24547 12767
rect 24489 12727 24547 12733
rect 25774 12724 25780 12776
rect 25832 12764 25838 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25832 12736 26065 12764
rect 25832 12724 25838 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 24394 12656 24400 12708
rect 24452 12696 24458 12708
rect 24452 12668 25360 12696
rect 24452 12656 24458 12668
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 4080 12600 4169 12628
rect 4157 12597 4169 12600
rect 4203 12597 4215 12631
rect 9950 12628 9956 12640
rect 9911 12600 9956 12628
rect 4157 12591 4215 12597
rect 9950 12588 9956 12600
rect 10008 12588 10014 12640
rect 14734 12628 14740 12640
rect 14695 12600 14740 12628
rect 14734 12588 14740 12600
rect 14792 12588 14798 12640
rect 15194 12628 15200 12640
rect 15155 12600 15200 12628
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 17218 12588 17224 12640
rect 17276 12628 17282 12640
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 17276 12600 17325 12628
rect 17276 12588 17282 12600
rect 17313 12597 17325 12600
rect 17359 12628 17371 12631
rect 17678 12628 17684 12640
rect 17359 12600 17684 12628
rect 17359 12597 17371 12600
rect 17313 12591 17371 12597
rect 17678 12588 17684 12600
rect 17736 12588 17742 12640
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12628 19487 12631
rect 19610 12628 19616 12640
rect 19475 12600 19616 12628
rect 19475 12597 19487 12600
rect 19429 12591 19487 12597
rect 19610 12588 19616 12600
rect 19668 12588 19674 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 20901 12631 20959 12637
rect 20901 12628 20913 12631
rect 20496 12600 20913 12628
rect 20496 12588 20502 12600
rect 20901 12597 20913 12600
rect 20947 12597 20959 12631
rect 20901 12591 20959 12597
rect 24578 12588 24584 12640
rect 24636 12628 24642 12640
rect 25332 12628 25360 12668
rect 25406 12628 25412 12640
rect 24636 12600 24681 12628
rect 25332 12600 25412 12628
rect 24636 12588 24642 12600
rect 25406 12588 25412 12600
rect 25464 12588 25470 12640
rect 25682 12628 25688 12640
rect 25643 12600 25688 12628
rect 25682 12588 25688 12600
rect 25740 12588 25746 12640
rect 26142 12588 26148 12640
rect 26200 12628 26206 12640
rect 26200 12600 26245 12628
rect 26200 12588 26206 12600
rect 26326 12588 26332 12640
rect 26384 12628 26390 12640
rect 26510 12628 26516 12640
rect 26384 12600 26516 12628
rect 26384 12588 26390 12600
rect 26510 12588 26516 12600
rect 26568 12628 26574 12640
rect 27249 12631 27307 12637
rect 27249 12628 27261 12631
rect 26568 12600 27261 12628
rect 26568 12588 26574 12600
rect 27249 12597 27261 12600
rect 27295 12597 27307 12631
rect 27249 12591 27307 12597
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1912 12396 2053 12424
rect 1912 12384 1918 12396
rect 2041 12393 2053 12396
rect 2087 12424 2099 12427
rect 3053 12427 3111 12433
rect 3053 12424 3065 12427
rect 2087 12396 3065 12424
rect 2087 12393 2099 12396
rect 2041 12387 2099 12393
rect 3053 12393 3065 12396
rect 3099 12393 3111 12427
rect 4338 12424 4344 12436
rect 4299 12396 4344 12424
rect 3053 12387 3111 12393
rect 4338 12384 4344 12396
rect 4396 12384 4402 12436
rect 7650 12424 7656 12436
rect 7611 12396 7656 12424
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8570 12424 8576 12436
rect 8531 12396 8576 12424
rect 8570 12384 8576 12396
rect 8628 12384 8634 12436
rect 15102 12424 15108 12436
rect 15063 12396 15108 12424
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 20438 12424 20444 12436
rect 19576 12396 20444 12424
rect 19576 12384 19582 12396
rect 20438 12384 20444 12396
rect 20496 12384 20502 12436
rect 22370 12384 22376 12436
rect 22428 12424 22434 12436
rect 23198 12424 23204 12436
rect 22428 12396 23204 12424
rect 22428 12384 22434 12396
rect 23198 12384 23204 12396
rect 23256 12384 23262 12436
rect 24210 12384 24216 12436
rect 24268 12424 24274 12436
rect 24305 12427 24363 12433
rect 24305 12424 24317 12427
rect 24268 12396 24317 12424
rect 24268 12384 24274 12396
rect 24305 12393 24317 12396
rect 24351 12393 24363 12427
rect 24762 12424 24768 12436
rect 24723 12396 24768 12424
rect 24305 12387 24363 12393
rect 24762 12384 24768 12396
rect 24820 12384 24826 12436
rect 25498 12384 25504 12436
rect 25556 12424 25562 12436
rect 25866 12424 25872 12436
rect 25556 12396 25872 12424
rect 25556 12384 25562 12396
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 26237 12427 26295 12433
rect 26237 12393 26249 12427
rect 26283 12424 26295 12427
rect 26326 12424 26332 12436
rect 26283 12396 26332 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 26326 12384 26332 12396
rect 26384 12384 26390 12436
rect 14737 12359 14795 12365
rect 14737 12325 14749 12359
rect 14783 12356 14795 12359
rect 15746 12356 15752 12368
rect 14783 12328 15752 12356
rect 14783 12325 14795 12328
rect 14737 12319 14795 12325
rect 15746 12316 15752 12328
rect 15804 12316 15810 12368
rect 15838 12316 15844 12368
rect 15896 12356 15902 12368
rect 16482 12356 16488 12368
rect 15896 12328 16488 12356
rect 15896 12316 15902 12328
rect 16482 12316 16488 12328
rect 16540 12316 16546 12368
rect 19058 12356 19064 12368
rect 18340 12328 19064 12356
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 6546 12297 6552 12300
rect 6540 12288 6552 12297
rect 2832 12260 2877 12288
rect 6507 12260 6552 12288
rect 2832 12248 2838 12260
rect 6540 12251 6552 12260
rect 6546 12248 6552 12251
rect 6604 12248 6610 12300
rect 11238 12288 11244 12300
rect 11199 12260 11244 12288
rect 11238 12248 11244 12260
rect 11296 12248 11302 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15252 12260 15669 12288
rect 15252 12248 15258 12260
rect 15657 12257 15669 12260
rect 15703 12288 15715 12291
rect 16669 12291 16727 12297
rect 16669 12288 16681 12291
rect 15703 12260 16681 12288
rect 15703 12257 15715 12260
rect 15657 12251 15715 12257
rect 16669 12257 16681 12260
rect 16715 12257 16727 12291
rect 16669 12251 16727 12257
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18340 12297 18368 12328
rect 19058 12316 19064 12328
rect 19116 12316 19122 12368
rect 23400 12328 24900 12356
rect 18325 12291 18383 12297
rect 18325 12288 18337 12291
rect 18104 12260 18337 12288
rect 18104 12248 18110 12260
rect 18325 12257 18337 12260
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 18592 12291 18650 12297
rect 18592 12257 18604 12291
rect 18638 12288 18650 12291
rect 18966 12288 18972 12300
rect 18638 12260 18972 12288
rect 18638 12257 18650 12260
rect 18592 12251 18650 12257
rect 18966 12248 18972 12260
rect 19024 12248 19030 12300
rect 20717 12291 20775 12297
rect 20717 12257 20729 12291
rect 20763 12288 20775 12291
rect 21266 12288 21272 12300
rect 20763 12260 21272 12288
rect 20763 12257 20775 12260
rect 20717 12251 20775 12257
rect 21266 12248 21272 12260
rect 21324 12248 21330 12300
rect 22830 12248 22836 12300
rect 22888 12288 22894 12300
rect 23106 12288 23112 12300
rect 22888 12260 23112 12288
rect 22888 12248 22894 12260
rect 23106 12248 23112 12260
rect 23164 12248 23170 12300
rect 23400 12232 23428 12328
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 24673 12291 24731 12297
rect 24673 12288 24685 12291
rect 24360 12260 24685 12288
rect 24360 12248 24366 12260
rect 24673 12257 24685 12260
rect 24719 12257 24731 12291
rect 24673 12251 24731 12257
rect 24872 12232 24900 12328
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 26881 12359 26939 12365
rect 26881 12356 26893 12359
rect 26660 12328 26893 12356
rect 26660 12316 26666 12328
rect 26881 12325 26893 12328
rect 26927 12325 26939 12359
rect 26881 12319 26939 12325
rect 25406 12248 25412 12300
rect 25464 12288 25470 12300
rect 26973 12291 27031 12297
rect 26973 12288 26985 12291
rect 25464 12260 26985 12288
rect 25464 12248 25470 12260
rect 26973 12257 26985 12260
rect 27019 12257 27031 12291
rect 26973 12251 27031 12257
rect 2130 12220 2136 12232
rect 2091 12192 2136 12220
rect 2130 12180 2136 12192
rect 2188 12180 2194 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 2406 12220 2412 12232
rect 2363 12192 2412 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 4985 12223 5043 12229
rect 4985 12220 4997 12223
rect 4939 12192 4997 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 4985 12189 4997 12192
rect 5031 12220 5043 12223
rect 5166 12220 5172 12232
rect 5031 12192 5172 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5592 12192 6285 12220
rect 5592 12180 5598 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 10836 12192 11345 12220
rect 10836 12180 10842 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 12342 12220 12348 12232
rect 11563 12192 12348 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15378 12220 15384 12232
rect 15068 12192 15384 12220
rect 15068 12180 15074 12192
rect 15378 12180 15384 12192
rect 15436 12180 15442 12232
rect 15470 12180 15476 12232
rect 15528 12220 15534 12232
rect 15841 12223 15899 12229
rect 15841 12220 15853 12223
rect 15528 12192 15853 12220
rect 15528 12180 15534 12192
rect 15841 12189 15853 12192
rect 15887 12189 15899 12223
rect 21358 12220 21364 12232
rect 21319 12192 21364 12220
rect 15841 12183 15899 12189
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 23382 12220 23388 12232
rect 21508 12192 21553 12220
rect 23343 12192 23388 12220
rect 21508 12180 21514 12192
rect 23382 12180 23388 12192
rect 23440 12180 23446 12232
rect 24854 12180 24860 12232
rect 24912 12220 24918 12232
rect 27154 12220 27160 12232
rect 24912 12192 25005 12220
rect 27115 12192 27160 12220
rect 24912 12180 24918 12192
rect 27154 12180 27160 12192
rect 27212 12180 27218 12232
rect 1673 12155 1731 12161
rect 1673 12121 1685 12155
rect 1719 12152 1731 12155
rect 2682 12152 2688 12164
rect 1719 12124 2688 12152
rect 1719 12121 1731 12124
rect 1673 12115 1731 12121
rect 2682 12112 2688 12124
rect 2740 12112 2746 12164
rect 19702 12152 19708 12164
rect 19615 12124 19708 12152
rect 19702 12112 19708 12124
rect 19760 12152 19766 12164
rect 21468 12152 21496 12180
rect 19760 12124 21496 12152
rect 22741 12155 22799 12161
rect 19760 12112 19766 12124
rect 22741 12121 22753 12155
rect 22787 12152 22799 12155
rect 24121 12155 24179 12161
rect 24121 12152 24133 12155
rect 22787 12124 24133 12152
rect 22787 12121 22799 12124
rect 22741 12115 22799 12121
rect 24121 12121 24133 12124
rect 24167 12152 24179 12155
rect 24578 12152 24584 12164
rect 24167 12124 24584 12152
rect 24167 12121 24179 12124
rect 24121 12115 24179 12121
rect 24578 12112 24584 12124
rect 24636 12112 24642 12164
rect 25777 12155 25835 12161
rect 25777 12121 25789 12155
rect 25823 12152 25835 12155
rect 26142 12152 26148 12164
rect 25823 12124 26148 12152
rect 25823 12121 25835 12124
rect 25777 12115 25835 12121
rect 26142 12112 26148 12124
rect 26200 12152 26206 12164
rect 26513 12155 26571 12161
rect 26513 12152 26525 12155
rect 26200 12124 26525 12152
rect 26200 12112 26206 12124
rect 26513 12121 26525 12124
rect 26559 12121 26571 12155
rect 26513 12115 26571 12121
rect 3050 12044 3056 12096
rect 3108 12084 3114 12096
rect 3697 12087 3755 12093
rect 3697 12084 3709 12087
rect 3108 12056 3709 12084
rect 3108 12044 3114 12056
rect 3697 12053 3709 12056
rect 3743 12084 3755 12087
rect 3878 12084 3884 12096
rect 3743 12056 3884 12084
rect 3743 12053 3755 12056
rect 3697 12047 3755 12053
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 8202 12084 8208 12096
rect 8163 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12044 8266 12096
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10873 12087 10931 12093
rect 10873 12084 10885 12087
rect 10100 12056 10885 12084
rect 10100 12044 10106 12056
rect 10873 12053 10885 12056
rect 10919 12053 10931 12087
rect 15286 12084 15292 12096
rect 15247 12056 15292 12084
rect 10873 12047 10931 12053
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 16298 12084 16304 12096
rect 16259 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 18138 12084 18144 12096
rect 18099 12056 18144 12084
rect 18138 12044 18144 12056
rect 18196 12044 18202 12096
rect 20898 12084 20904 12096
rect 20859 12056 20904 12084
rect 20898 12044 20904 12056
rect 20956 12044 20962 12096
rect 22002 12084 22008 12096
rect 21963 12056 22008 12084
rect 22002 12044 22008 12056
rect 22060 12044 22066 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 7650 11880 7656 11892
rect 7611 11852 7656 11880
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8478 11840 8484 11892
rect 8536 11880 8542 11892
rect 9585 11883 9643 11889
rect 9585 11880 9597 11883
rect 8536 11852 9597 11880
rect 8536 11840 8542 11852
rect 9585 11849 9597 11852
rect 9631 11880 9643 11883
rect 9950 11880 9956 11892
rect 9631 11852 9956 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14826 11840 14832 11892
rect 14884 11880 14890 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14884 11852 15209 11880
rect 14884 11840 14890 11852
rect 15197 11849 15209 11852
rect 15243 11849 15255 11883
rect 15197 11843 15255 11849
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19705 11883 19763 11889
rect 19705 11880 19717 11883
rect 19576 11852 19717 11880
rect 19576 11840 19582 11852
rect 19705 11849 19717 11852
rect 19751 11849 19763 11883
rect 19705 11843 19763 11849
rect 21266 11840 21272 11892
rect 21324 11880 21330 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 21324 11852 21465 11880
rect 21324 11840 21330 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 22833 11883 22891 11889
rect 22833 11849 22845 11883
rect 22879 11880 22891 11883
rect 23106 11880 23112 11892
rect 22879 11852 23112 11880
rect 22879 11849 22891 11852
rect 22833 11843 22891 11849
rect 23106 11840 23112 11852
rect 23164 11840 23170 11892
rect 24029 11883 24087 11889
rect 24029 11849 24041 11883
rect 24075 11880 24087 11883
rect 24670 11880 24676 11892
rect 24075 11852 24676 11880
rect 24075 11849 24087 11852
rect 24029 11843 24087 11849
rect 4246 11704 4252 11756
rect 4304 11744 4310 11756
rect 5074 11744 5080 11756
rect 4304 11716 5080 11744
rect 4304 11704 4310 11716
rect 5074 11704 5080 11716
rect 5132 11744 5138 11756
rect 5353 11747 5411 11753
rect 5353 11744 5365 11747
rect 5132 11716 5365 11744
rect 5132 11704 5138 11716
rect 5353 11713 5365 11716
rect 5399 11744 5411 11747
rect 6454 11744 6460 11756
rect 5399 11716 6460 11744
rect 5399 11713 5411 11716
rect 5353 11707 5411 11713
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 7668 11744 7696 11840
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 9677 11815 9735 11821
rect 9677 11812 9689 11815
rect 8260 11784 9689 11812
rect 8260 11772 8266 11784
rect 9677 11781 9689 11784
rect 9723 11781 9735 11815
rect 9677 11775 9735 11781
rect 8389 11747 8447 11753
rect 8389 11744 8401 11747
rect 7668 11716 8401 11744
rect 8389 11713 8401 11716
rect 8435 11713 8447 11747
rect 9968 11744 9996 11840
rect 21910 11772 21916 11824
rect 21968 11812 21974 11824
rect 24044 11812 24072 11843
rect 24670 11840 24676 11852
rect 24728 11840 24734 11892
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25593 11883 25651 11889
rect 25593 11880 25605 11883
rect 24912 11852 25605 11880
rect 24912 11840 24918 11852
rect 21968 11784 24072 11812
rect 21968 11772 21974 11784
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 9968 11716 10241 11744
rect 8389 11707 8447 11713
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 11238 11744 11244 11756
rect 11199 11716 11244 11744
rect 10229 11707 10287 11713
rect 11238 11704 11244 11716
rect 11296 11744 11302 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11296 11716 11713 11744
rect 11296 11704 11302 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 16390 11744 16396 11756
rect 16351 11716 16396 11744
rect 11701 11707 11759 11713
rect 16390 11704 16396 11716
rect 16448 11704 16454 11756
rect 17497 11747 17555 11753
rect 17497 11713 17509 11747
rect 17543 11744 17555 11747
rect 18877 11747 18935 11753
rect 18877 11744 18889 11747
rect 17543 11716 18889 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 18877 11713 18889 11716
rect 18923 11744 18935 11747
rect 19702 11744 19708 11756
rect 18923 11716 19708 11744
rect 18923 11713 18935 11716
rect 18877 11707 18935 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 20438 11744 20444 11756
rect 20399 11716 20444 11744
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 20714 11704 20720 11756
rect 20772 11744 20778 11756
rect 21269 11747 21327 11753
rect 21269 11744 21281 11747
rect 20772 11716 21281 11744
rect 20772 11704 20778 11716
rect 21269 11713 21281 11716
rect 21315 11713 21327 11747
rect 22002 11744 22008 11756
rect 21963 11716 22008 11744
rect 21269 11707 21327 11713
rect 1673 11679 1731 11685
rect 1673 11645 1685 11679
rect 1719 11676 1731 11679
rect 5166 11676 5172 11688
rect 1719 11648 2728 11676
rect 5127 11648 5172 11676
rect 1719 11645 1731 11648
rect 1673 11639 1731 11645
rect 1940 11611 1998 11617
rect 1940 11577 1952 11611
rect 1986 11608 1998 11611
rect 2038 11608 2044 11620
rect 1986 11580 2044 11608
rect 1986 11577 1998 11580
rect 1940 11571 1998 11577
rect 2038 11568 2044 11580
rect 2096 11568 2102 11620
rect 2700 11608 2728 11648
rect 5166 11636 5172 11648
rect 5224 11636 5230 11688
rect 6365 11679 6423 11685
rect 6365 11645 6377 11679
rect 6411 11676 6423 11679
rect 6546 11676 6552 11688
rect 6411 11648 6552 11676
rect 6411 11645 6423 11648
rect 6365 11639 6423 11645
rect 6546 11636 6552 11648
rect 6604 11676 6610 11688
rect 7742 11676 7748 11688
rect 6604 11648 7748 11676
rect 6604 11636 6610 11648
rect 7742 11636 7748 11648
rect 7800 11636 7806 11688
rect 8202 11676 8208 11688
rect 8163 11648 8208 11676
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 10042 11676 10048 11688
rect 10003 11648 10048 11676
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 13814 11636 13820 11688
rect 13872 11676 13878 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13872 11648 13921 11676
rect 13872 11636 13878 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 15654 11636 15660 11688
rect 15712 11676 15718 11688
rect 16209 11679 16267 11685
rect 16209 11676 16221 11679
rect 15712 11648 16221 11676
rect 15712 11636 15718 11648
rect 16209 11645 16221 11648
rect 16255 11676 16267 11679
rect 16298 11676 16304 11688
rect 16255 11648 16304 11676
rect 16255 11645 16267 11648
rect 16209 11639 16267 11645
rect 16298 11636 16304 11648
rect 16356 11636 16362 11688
rect 17865 11679 17923 11685
rect 17865 11645 17877 11679
rect 17911 11676 17923 11679
rect 18966 11676 18972 11688
rect 17911 11648 18972 11676
rect 17911 11645 17923 11648
rect 17865 11639 17923 11645
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11676 20315 11679
rect 20346 11676 20352 11688
rect 20303 11648 20352 11676
rect 20303 11645 20315 11648
rect 20257 11639 20315 11645
rect 20346 11636 20352 11648
rect 20404 11676 20410 11688
rect 20898 11676 20904 11688
rect 20404 11648 20904 11676
rect 20404 11636 20410 11648
rect 20898 11636 20904 11648
rect 20956 11636 20962 11688
rect 21284 11676 21312 11707
rect 22002 11704 22008 11716
rect 22060 11704 22066 11756
rect 24302 11744 24308 11756
rect 24263 11716 24308 11744
rect 24302 11704 24308 11716
rect 24360 11704 24366 11756
rect 25038 11744 25044 11756
rect 24999 11716 25044 11744
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25332 11744 25360 11852
rect 25593 11849 25605 11852
rect 25639 11849 25651 11883
rect 25593 11843 25651 11849
rect 25774 11840 25780 11892
rect 25832 11880 25838 11892
rect 26145 11883 26203 11889
rect 26145 11880 26157 11883
rect 25832 11852 26157 11880
rect 25832 11840 25838 11852
rect 26145 11849 26157 11852
rect 26191 11849 26203 11883
rect 26145 11843 26203 11849
rect 25406 11772 25412 11824
rect 25464 11812 25470 11824
rect 25961 11815 26019 11821
rect 25961 11812 25973 11815
rect 25464 11784 25973 11812
rect 25464 11772 25470 11784
rect 25961 11781 25973 11784
rect 26007 11781 26019 11815
rect 27154 11812 27160 11824
rect 25961 11775 26019 11781
rect 26160 11784 27160 11812
rect 26160 11744 26188 11784
rect 26712 11753 26740 11784
rect 27154 11772 27160 11784
rect 27212 11812 27218 11824
rect 27525 11815 27583 11821
rect 27525 11812 27537 11815
rect 27212 11784 27537 11812
rect 27212 11772 27218 11784
rect 27525 11781 27537 11784
rect 27571 11781 27583 11815
rect 27525 11775 27583 11781
rect 25332 11716 26188 11744
rect 26697 11747 26755 11753
rect 26697 11713 26709 11747
rect 26743 11713 26755 11747
rect 26697 11707 26755 11713
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 21284 11648 21925 11676
rect 21913 11645 21925 11648
rect 21959 11645 21971 11679
rect 21913 11639 21971 11645
rect 24857 11679 24915 11685
rect 24857 11645 24869 11679
rect 24903 11676 24915 11679
rect 25682 11676 25688 11688
rect 24903 11648 25688 11676
rect 24903 11645 24915 11648
rect 24857 11639 24915 11645
rect 25682 11636 25688 11648
rect 25740 11636 25746 11688
rect 26510 11676 26516 11688
rect 26471 11648 26516 11676
rect 26510 11636 26516 11648
rect 26568 11636 26574 11688
rect 2774 11608 2780 11620
rect 2700 11580 2780 11608
rect 2774 11568 2780 11580
rect 2832 11608 2838 11620
rect 3605 11611 3663 11617
rect 3605 11608 3617 11611
rect 2832 11580 3617 11608
rect 2832 11568 2838 11580
rect 3605 11577 3617 11580
rect 3651 11577 3663 11611
rect 3605 11571 3663 11577
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11608 4767 11611
rect 5258 11608 5264 11620
rect 4755 11580 5264 11608
rect 4755 11577 4767 11580
rect 4709 11571 4767 11577
rect 5258 11568 5264 11580
rect 5316 11568 5322 11620
rect 8297 11611 8355 11617
rect 8297 11608 8309 11611
rect 7392 11580 8309 11608
rect 7392 11552 7420 11580
rect 8297 11577 8309 11580
rect 8343 11577 8355 11611
rect 8297 11571 8355 11577
rect 9217 11611 9275 11617
rect 9217 11577 9229 11611
rect 9263 11608 9275 11611
rect 10137 11611 10195 11617
rect 10137 11608 10149 11611
rect 9263 11580 10149 11608
rect 9263 11577 9275 11580
rect 9217 11571 9275 11577
rect 10137 11577 10149 11580
rect 10183 11608 10195 11611
rect 10594 11608 10600 11620
rect 10183 11580 10600 11608
rect 10183 11577 10195 11580
rect 10137 11571 10195 11577
rect 10594 11568 10600 11580
rect 10652 11568 10658 11620
rect 15194 11568 15200 11620
rect 15252 11608 15258 11620
rect 16117 11611 16175 11617
rect 16117 11608 16129 11611
rect 15252 11580 16129 11608
rect 15252 11568 15258 11580
rect 16117 11577 16129 11580
rect 16163 11608 16175 11611
rect 16163 11580 16896 11608
rect 16163 11577 16175 11580
rect 16117 11571 16175 11577
rect 16868 11552 16896 11580
rect 18138 11568 18144 11620
rect 18196 11608 18202 11620
rect 18693 11611 18751 11617
rect 18693 11608 18705 11611
rect 18196 11580 18705 11608
rect 18196 11568 18202 11580
rect 18693 11577 18705 11580
rect 18739 11577 18751 11611
rect 18693 11571 18751 11577
rect 20993 11611 21051 11617
rect 20993 11577 21005 11611
rect 21039 11608 21051 11611
rect 21726 11608 21732 11620
rect 21039 11580 21732 11608
rect 21039 11577 21051 11580
rect 20993 11571 21051 11577
rect 21726 11568 21732 11580
rect 21784 11608 21790 11620
rect 21821 11611 21879 11617
rect 21821 11608 21833 11611
rect 21784 11580 21833 11608
rect 21784 11568 21790 11580
rect 21821 11577 21833 11580
rect 21867 11577 21879 11611
rect 24946 11608 24952 11620
rect 24907 11580 24952 11608
rect 21821 11571 21879 11577
rect 24946 11568 24952 11580
rect 25004 11568 25010 11620
rect 26142 11568 26148 11620
rect 26200 11608 26206 11620
rect 26605 11611 26663 11617
rect 26605 11608 26617 11611
rect 26200 11580 26617 11608
rect 26200 11568 26206 11580
rect 26605 11577 26617 11580
rect 26651 11577 26663 11611
rect 26605 11571 26663 11577
rect 3050 11540 3056 11552
rect 3011 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 4246 11540 4252 11552
rect 4207 11512 4252 11540
rect 4246 11500 4252 11512
rect 4304 11500 4310 11552
rect 4798 11540 4804 11552
rect 4759 11512 4804 11540
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 5905 11543 5963 11549
rect 5905 11540 5917 11543
rect 5592 11512 5917 11540
rect 5592 11500 5598 11512
rect 5905 11509 5917 11512
rect 5951 11509 5963 11543
rect 7374 11540 7380 11552
rect 7335 11512 7380 11540
rect 5905 11503 5963 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 7834 11540 7840 11552
rect 7795 11512 7840 11540
rect 7834 11500 7840 11512
rect 7892 11500 7898 11552
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 10873 11543 10931 11549
rect 10873 11540 10885 11543
rect 10836 11512 10885 11540
rect 10836 11500 10842 11512
rect 10873 11509 10885 11512
rect 10919 11509 10931 11543
rect 10873 11503 10931 11509
rect 12161 11543 12219 11549
rect 12161 11509 12173 11543
rect 12207 11540 12219 11543
rect 12342 11540 12348 11552
rect 12207 11512 12348 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15749 11543 15807 11549
rect 15749 11540 15761 11543
rect 15436 11512 15761 11540
rect 15436 11500 15442 11512
rect 15749 11509 15761 11512
rect 15795 11509 15807 11543
rect 16850 11540 16856 11552
rect 16811 11512 16856 11540
rect 15749 11503 15807 11509
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 18322 11540 18328 11552
rect 18283 11512 18328 11540
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 18782 11540 18788 11552
rect 18695 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11540 18846 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 18840 11512 19349 11540
rect 18840 11500 18846 11512
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19337 11503 19395 11509
rect 19889 11543 19947 11549
rect 19889 11509 19901 11543
rect 19935 11540 19947 11543
rect 20070 11540 20076 11552
rect 19935 11512 20076 11540
rect 19935 11509 19947 11512
rect 19889 11503 19947 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20162 11500 20168 11552
rect 20220 11540 20226 11552
rect 20349 11543 20407 11549
rect 20349 11540 20361 11543
rect 20220 11512 20361 11540
rect 20220 11500 20226 11512
rect 20349 11509 20361 11512
rect 20395 11509 20407 11543
rect 20349 11503 20407 11509
rect 22830 11500 22836 11552
rect 22888 11540 22894 11552
rect 23382 11540 23388 11552
rect 22888 11512 23388 11540
rect 22888 11500 22894 11512
rect 23382 11500 23388 11512
rect 23440 11500 23446 11552
rect 24489 11543 24547 11549
rect 24489 11509 24501 11543
rect 24535 11540 24547 11543
rect 24762 11540 24768 11552
rect 24535 11512 24768 11540
rect 24535 11509 24547 11512
rect 24489 11503 24547 11509
rect 24762 11500 24768 11512
rect 24820 11500 24826 11552
rect 26510 11500 26516 11552
rect 26568 11540 26574 11552
rect 27157 11543 27215 11549
rect 27157 11540 27169 11543
rect 26568 11512 27169 11540
rect 26568 11500 26574 11512
rect 27157 11509 27169 11512
rect 27203 11509 27215 11543
rect 27157 11503 27215 11509
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2038 11336 2044 11348
rect 1951 11308 2044 11336
rect 2038 11296 2044 11308
rect 2096 11336 2102 11348
rect 2406 11336 2412 11348
rect 2096 11308 2412 11336
rect 2096 11296 2102 11308
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 4798 11336 4804 11348
rect 4663 11308 4804 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 4798 11296 4804 11308
rect 4856 11296 4862 11348
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 7432 11308 7849 11336
rect 7432 11296 7438 11308
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 10042 11336 10048 11348
rect 9999 11308 10048 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10594 11336 10600 11348
rect 10555 11308 10600 11336
rect 10594 11296 10600 11308
rect 10652 11296 10658 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 19889 11339 19947 11345
rect 19889 11336 19901 11339
rect 18380 11308 19901 11336
rect 18380 11296 18386 11308
rect 19889 11305 19901 11308
rect 19935 11336 19947 11339
rect 20162 11336 20168 11348
rect 19935 11308 20168 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 20717 11339 20775 11345
rect 20717 11305 20729 11339
rect 20763 11336 20775 11339
rect 21358 11336 21364 11348
rect 20763 11308 21364 11336
rect 20763 11305 20775 11308
rect 20717 11299 20775 11305
rect 21358 11296 21364 11308
rect 21416 11296 21422 11348
rect 22830 11336 22836 11348
rect 22791 11308 22836 11336
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 23198 11336 23204 11348
rect 23159 11308 23204 11336
rect 23198 11296 23204 11308
rect 23256 11296 23262 11348
rect 24946 11336 24952 11348
rect 24907 11308 24952 11336
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25317 11339 25375 11345
rect 25317 11305 25329 11339
rect 25363 11336 25375 11339
rect 25682 11336 25688 11348
rect 25363 11308 25688 11336
rect 25363 11305 25375 11308
rect 25317 11299 25375 11305
rect 25682 11296 25688 11308
rect 25740 11296 25746 11348
rect 26694 11336 26700 11348
rect 26655 11308 26700 11336
rect 26694 11296 26700 11308
rect 26752 11296 26758 11348
rect 2130 11228 2136 11280
rect 2188 11268 2194 11280
rect 3053 11271 3111 11277
rect 3053 11268 3065 11271
rect 2188 11240 3065 11268
rect 2188 11228 2194 11240
rect 3053 11237 3065 11240
rect 3099 11237 3111 11271
rect 9582 11268 9588 11280
rect 3053 11231 3111 11237
rect 3804 11240 9588 11268
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 1486 11200 1492 11212
rect 1443 11172 1492 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 1486 11160 1492 11172
rect 1544 11160 1550 11212
rect 2498 11200 2504 11212
rect 2411 11172 2504 11200
rect 2498 11160 2504 11172
rect 2556 11200 2562 11212
rect 3804 11200 3832 11240
rect 9582 11228 9588 11240
rect 9640 11228 9646 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 16022 11268 16028 11280
rect 12308 11240 16028 11268
rect 12308 11228 12314 11240
rect 15856 11212 15884 11240
rect 16022 11228 16028 11240
rect 16080 11228 16086 11280
rect 18046 11268 18052 11280
rect 18007 11240 18052 11268
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 21177 11271 21235 11277
rect 21177 11237 21189 11271
rect 21223 11268 21235 11271
rect 21450 11268 21456 11280
rect 21223 11240 21456 11268
rect 21223 11237 21235 11240
rect 21177 11231 21235 11237
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 24581 11271 24639 11277
rect 24581 11237 24593 11271
rect 24627 11268 24639 11271
rect 25038 11268 25044 11280
rect 24627 11240 25044 11268
rect 24627 11237 24639 11240
rect 24581 11231 24639 11237
rect 25038 11228 25044 11240
rect 25096 11228 25102 11280
rect 2556 11172 3832 11200
rect 2556 11160 2562 11172
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 3936 11172 4844 11200
rect 3936 11160 3942 11172
rect 4816 11141 4844 11172
rect 5810 11160 5816 11212
rect 5868 11200 5874 11212
rect 6181 11203 6239 11209
rect 6181 11200 6193 11203
rect 5868 11172 6193 11200
rect 5868 11160 5874 11172
rect 6181 11169 6193 11172
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 8202 11200 8208 11212
rect 7791 11172 8208 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 10502 11160 10508 11212
rect 10560 11200 10566 11212
rect 10870 11200 10876 11212
rect 10560 11172 10876 11200
rect 10560 11160 10566 11172
rect 10870 11160 10876 11172
rect 10928 11200 10934 11212
rect 10965 11203 11023 11209
rect 10965 11200 10977 11203
rect 10928 11172 10977 11200
rect 10928 11160 10934 11172
rect 10965 11169 10977 11172
rect 11011 11169 11023 11203
rect 10965 11163 11023 11169
rect 12986 11160 12992 11212
rect 13044 11200 13050 11212
rect 13153 11203 13211 11209
rect 13153 11200 13165 11203
rect 13044 11172 13165 11200
rect 13044 11160 13050 11172
rect 13153 11169 13165 11172
rect 13199 11169 13211 11203
rect 13153 11163 13211 11169
rect 15838 11160 15844 11212
rect 15896 11160 15902 11212
rect 15933 11203 15991 11209
rect 15933 11169 15945 11203
rect 15979 11200 15991 11203
rect 16298 11200 16304 11212
rect 15979 11172 16304 11200
rect 15979 11169 15991 11172
rect 15933 11163 15991 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 17954 11160 17960 11212
rect 18012 11200 18018 11212
rect 18509 11203 18567 11209
rect 18509 11200 18521 11203
rect 18012 11172 18521 11200
rect 18012 11160 18018 11172
rect 18509 11169 18521 11172
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 21358 11160 21364 11212
rect 21416 11200 21422 11212
rect 21729 11203 21787 11209
rect 21729 11200 21741 11203
rect 21416 11172 21741 11200
rect 21416 11160 21422 11172
rect 21729 11169 21741 11172
rect 21775 11169 21787 11203
rect 26510 11200 26516 11212
rect 26471 11172 26516 11200
rect 21729 11163 21787 11169
rect 26510 11160 26516 11172
rect 26568 11160 26574 11212
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 4801 11135 4859 11141
rect 4801 11101 4813 11135
rect 4847 11101 4859 11135
rect 6270 11132 6276 11144
rect 6231 11104 6276 11132
rect 4801 11095 4859 11101
rect 1578 11064 1584 11076
rect 1539 11036 1584 11064
rect 1578 11024 1584 11036
rect 1636 11024 1642 11076
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 4724 11064 4752 11095
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6454 11132 6460 11144
rect 6415 11104 6460 11132
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8297 11135 8355 11141
rect 8297 11132 8309 11135
rect 8076 11104 8309 11132
rect 8076 11092 8082 11104
rect 8297 11101 8309 11104
rect 8343 11101 8355 11135
rect 8478 11132 8484 11144
rect 8439 11104 8484 11132
rect 8297 11095 8355 11101
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 11054 11132 11060 11144
rect 11015 11104 11060 11132
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11101 11207 11135
rect 12894 11132 12900 11144
rect 12855 11104 12900 11132
rect 11149 11095 11207 11101
rect 5813 11067 5871 11073
rect 5813 11064 5825 11067
rect 4396 11036 5825 11064
rect 4396 11024 4402 11036
rect 5813 11033 5825 11036
rect 5859 11033 5871 11067
rect 5813 11027 5871 11033
rect 7742 11024 7748 11076
rect 7800 11064 7806 11076
rect 8496 11064 8524 11092
rect 7800 11036 8524 11064
rect 7800 11024 7806 11036
rect 10594 11024 10600 11076
rect 10652 11064 10658 11076
rect 11164 11064 11192 11095
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11132 16175 11135
rect 16390 11132 16396 11144
rect 16163 11104 16396 11132
rect 16163 11101 16175 11104
rect 16117 11095 16175 11101
rect 12342 11064 12348 11076
rect 10652 11036 12348 11064
rect 10652 11024 10658 11036
rect 12342 11024 12348 11036
rect 12400 11024 12406 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14292 11036 15025 11064
rect 14292 11008 14320 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 16132 11064 16160 11095
rect 16390 11092 16396 11104
rect 16448 11132 16454 11144
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16448 11104 16589 11132
rect 16448 11092 16454 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 18598 11132 18604 11144
rect 18559 11104 18604 11132
rect 16577 11095 16635 11101
rect 18598 11092 18604 11104
rect 18656 11092 18662 11144
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11132 18843 11135
rect 18966 11132 18972 11144
rect 18831 11104 18972 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 18966 11092 18972 11104
rect 19024 11092 19030 11144
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21818 11132 21824 11144
rect 20864 11104 21824 11132
rect 20864 11092 20870 11104
rect 21818 11092 21824 11104
rect 21876 11092 21882 11144
rect 22002 11132 22008 11144
rect 21963 11104 22008 11132
rect 22002 11092 22008 11104
rect 22060 11092 22066 11144
rect 15013 11027 15071 11033
rect 15120 11036 16160 11064
rect 4249 10999 4307 11005
rect 4249 10965 4261 10999
rect 4295 10996 4307 10999
rect 4890 10996 4896 11008
rect 4295 10968 4896 10996
rect 4295 10965 4307 10968
rect 4249 10959 4307 10965
rect 4890 10956 4896 10968
rect 4948 10996 4954 11008
rect 5261 10999 5319 11005
rect 5261 10996 5273 10999
rect 4948 10968 5273 10996
rect 4948 10956 4954 10968
rect 5261 10965 5273 10968
rect 5307 10965 5319 10999
rect 5261 10959 5319 10965
rect 8662 10956 8668 11008
rect 8720 10996 8726 11008
rect 8849 10999 8907 11005
rect 8849 10996 8861 10999
rect 8720 10968 8861 10996
rect 8720 10956 8726 10968
rect 8849 10965 8861 10968
rect 8895 10965 8907 10999
rect 14274 10996 14280 11008
rect 14235 10968 14280 10996
rect 8849 10959 8907 10965
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 14734 10956 14740 11008
rect 14792 10996 14798 11008
rect 15120 10996 15148 11036
rect 20714 11024 20720 11076
rect 20772 11064 20778 11076
rect 25130 11064 25136 11076
rect 20772 11036 25136 11064
rect 20772 11024 20778 11036
rect 25130 11024 25136 11036
rect 25188 11064 25194 11076
rect 26142 11064 26148 11076
rect 25188 11036 26148 11064
rect 25188 11024 25194 11036
rect 26142 11024 26148 11036
rect 26200 11024 26206 11076
rect 15562 10996 15568 11008
rect 14792 10968 15148 10996
rect 15523 10968 15568 10996
rect 14792 10956 14798 10968
rect 15562 10956 15568 10968
rect 15620 10956 15626 11008
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 17862 10996 17868 11008
rect 16632 10968 17868 10996
rect 16632 10956 16638 10968
rect 17862 10956 17868 10968
rect 17920 10956 17926 11008
rect 19150 10996 19156 11008
rect 19111 10968 19156 10996
rect 19150 10956 19156 10968
rect 19208 10956 19214 11008
rect 23937 10999 23995 11005
rect 23937 10965 23949 10999
rect 23983 10996 23995 10999
rect 24210 10996 24216 11008
rect 23983 10968 24216 10996
rect 23983 10965 23995 10968
rect 23937 10959 23995 10965
rect 24210 10956 24216 10968
rect 24268 10956 24274 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 1544 10764 1593 10792
rect 1544 10752 1550 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 5074 10752 5080 10804
rect 5132 10792 5138 10804
rect 5718 10792 5724 10804
rect 5132 10764 5724 10792
rect 5132 10752 5138 10764
rect 5718 10752 5724 10764
rect 5776 10752 5782 10804
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 6549 10795 6607 10801
rect 6549 10792 6561 10795
rect 6512 10764 6561 10792
rect 6512 10752 6518 10764
rect 6549 10761 6561 10764
rect 6595 10761 6607 10795
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 6549 10755 6607 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13262 10792 13268 10804
rect 12952 10764 13268 10792
rect 12952 10752 12958 10764
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 15933 10795 15991 10801
rect 15933 10792 15945 10795
rect 15896 10764 15945 10792
rect 15896 10752 15902 10764
rect 15933 10761 15945 10764
rect 15979 10761 15991 10795
rect 16298 10792 16304 10804
rect 16259 10764 16304 10792
rect 15933 10755 15991 10761
rect 16298 10752 16304 10764
rect 16356 10792 16362 10804
rect 18325 10795 18383 10801
rect 16356 10764 16528 10792
rect 16356 10752 16362 10764
rect 3421 10727 3479 10733
rect 3421 10693 3433 10727
rect 3467 10693 3479 10727
rect 5902 10724 5908 10736
rect 5863 10696 5908 10724
rect 3421 10687 3479 10693
rect 3436 10656 3464 10687
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8294 10724 8300 10736
rect 7984 10696 8300 10724
rect 7984 10684 7990 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 8680 10696 9781 10724
rect 8680 10668 8708 10696
rect 9769 10693 9781 10696
rect 9815 10693 9827 10727
rect 12986 10724 12992 10736
rect 12947 10696 12992 10724
rect 9769 10687 9827 10693
rect 12986 10684 12992 10696
rect 13044 10724 13050 10736
rect 14734 10724 14740 10736
rect 13044 10696 14740 10724
rect 13044 10684 13050 10696
rect 14734 10684 14740 10696
rect 14792 10684 14798 10736
rect 3970 10656 3976 10668
rect 3436 10628 3976 10656
rect 3970 10616 3976 10628
rect 4028 10656 4034 10668
rect 4433 10659 4491 10665
rect 4433 10656 4445 10659
rect 4028 10628 4445 10656
rect 4028 10616 4034 10628
rect 4433 10625 4445 10628
rect 4479 10656 4491 10659
rect 5077 10659 5135 10665
rect 5077 10656 5089 10659
rect 4479 10628 5089 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 5077 10625 5089 10628
rect 5123 10625 5135 10659
rect 5077 10619 5135 10625
rect 7558 10616 7564 10668
rect 7616 10656 7622 10668
rect 8386 10656 8392 10668
rect 7616 10628 8392 10656
rect 7616 10616 7622 10628
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2682 10588 2688 10600
rect 2087 10560 2688 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 4890 10588 4896 10600
rect 4851 10560 4896 10588
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 8128 10597 8156 10628
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 8662 10656 8668 10668
rect 8623 10628 8668 10656
rect 8662 10616 8668 10628
rect 8720 10616 8726 10668
rect 8849 10659 8907 10665
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 8938 10656 8944 10668
rect 8895 10628 8944 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 9916 10628 10333 10656
rect 9916 10616 9922 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 14274 10616 14280 10668
rect 14332 10656 14338 10668
rect 15470 10656 15476 10668
rect 14332 10628 15476 10656
rect 14332 10616 14338 10628
rect 15470 10616 15476 10628
rect 15528 10616 15534 10668
rect 16500 10665 16528 10764
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18782 10792 18788 10804
rect 18371 10764 18788 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18782 10752 18788 10764
rect 18840 10752 18846 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 22002 10792 22008 10804
rect 21131 10764 22008 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 18598 10684 18604 10736
rect 18656 10724 18662 10736
rect 19705 10727 19763 10733
rect 19705 10724 19717 10727
rect 18656 10696 19717 10724
rect 18656 10684 18662 10696
rect 19705 10693 19717 10696
rect 19751 10693 19763 10727
rect 19705 10687 19763 10693
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10625 16543 10659
rect 16485 10619 16543 10625
rect 17497 10659 17555 10665
rect 17497 10625 17509 10659
rect 17543 10656 17555 10659
rect 18966 10656 18972 10668
rect 17543 10628 18972 10656
rect 17543 10625 17555 10628
rect 17497 10619 17555 10625
rect 18966 10616 18972 10628
rect 19024 10656 19030 10668
rect 21100 10656 21128 10755
rect 22002 10752 22008 10764
rect 22060 10752 22066 10804
rect 22278 10792 22284 10804
rect 22239 10764 22284 10792
rect 22278 10752 22284 10764
rect 22336 10752 22342 10804
rect 26510 10752 26516 10804
rect 26568 10792 26574 10804
rect 27341 10795 27399 10801
rect 27341 10792 27353 10795
rect 26568 10764 27353 10792
rect 26568 10752 26574 10764
rect 27341 10761 27353 10764
rect 27387 10761 27399 10795
rect 27341 10755 27399 10761
rect 21358 10724 21364 10736
rect 21319 10696 21364 10724
rect 21358 10684 21364 10696
rect 21416 10684 21422 10736
rect 21726 10656 21732 10668
rect 19024 10628 21128 10656
rect 21687 10628 21732 10656
rect 19024 10616 19030 10628
rect 21726 10616 21732 10628
rect 21784 10616 21790 10668
rect 23109 10659 23167 10665
rect 23109 10625 23121 10659
rect 23155 10656 23167 10659
rect 24489 10659 24547 10665
rect 24489 10656 24501 10659
rect 23155 10628 24501 10656
rect 23155 10625 23167 10628
rect 23109 10619 23167 10625
rect 24489 10625 24501 10628
rect 24535 10656 24547 10659
rect 24578 10656 24584 10668
rect 24535 10628 24584 10656
rect 24535 10625 24547 10628
rect 24489 10619 24547 10625
rect 24578 10616 24584 10628
rect 24636 10616 24642 10668
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7708 10560 7757 10588
rect 7708 10548 7714 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 14093 10591 14151 10597
rect 14093 10557 14105 10591
rect 14139 10588 14151 10591
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14139 10560 15301 10588
rect 14139 10557 14151 10560
rect 14093 10551 14151 10557
rect 15289 10557 15301 10560
rect 15335 10588 15347 10591
rect 15562 10588 15568 10600
rect 15335 10560 15568 10588
rect 15335 10557 15347 10560
rect 15289 10551 15347 10557
rect 15562 10548 15568 10560
rect 15620 10548 15626 10600
rect 18598 10548 18604 10600
rect 18656 10588 18662 10600
rect 18693 10591 18751 10597
rect 18693 10588 18705 10591
rect 18656 10560 18705 10588
rect 18656 10548 18662 10560
rect 18693 10557 18705 10560
rect 18739 10588 18751 10591
rect 19150 10588 19156 10600
rect 18739 10560 19156 10588
rect 18739 10557 18751 10560
rect 18693 10551 18751 10557
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 23477 10591 23535 10597
rect 23477 10557 23489 10591
rect 23523 10557 23535 10591
rect 26418 10588 26424 10600
rect 26379 10560 26424 10588
rect 23477 10551 23535 10557
rect 2130 10480 2136 10532
rect 2188 10520 2194 10532
rect 2286 10523 2344 10529
rect 2286 10520 2298 10523
rect 2188 10492 2298 10520
rect 2188 10480 2194 10492
rect 2286 10489 2298 10492
rect 2332 10520 2344 10523
rect 3050 10520 3056 10532
rect 2332 10492 3056 10520
rect 2332 10489 2344 10492
rect 2286 10483 2344 10489
rect 3050 10480 3056 10492
rect 3108 10520 3114 10532
rect 3973 10523 4031 10529
rect 3973 10520 3985 10523
rect 3108 10492 3985 10520
rect 3108 10480 3114 10492
rect 3973 10489 3985 10492
rect 4019 10489 4031 10523
rect 3973 10483 4031 10489
rect 4154 10480 4160 10532
rect 4212 10520 4218 10532
rect 4982 10520 4988 10532
rect 4212 10492 4988 10520
rect 4212 10480 4218 10492
rect 4982 10480 4988 10492
rect 5040 10480 5046 10532
rect 7101 10523 7159 10529
rect 7101 10489 7113 10523
rect 7147 10520 7159 10523
rect 8018 10520 8024 10532
rect 7147 10492 8024 10520
rect 7147 10489 7159 10492
rect 7101 10483 7159 10489
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 8570 10520 8576 10532
rect 8531 10492 8576 10520
rect 8570 10480 8576 10492
rect 8628 10480 8634 10532
rect 9677 10523 9735 10529
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 9723 10492 10272 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 10244 10464 10272 10492
rect 11054 10480 11060 10532
rect 11112 10480 11118 10532
rect 14461 10523 14519 10529
rect 14461 10489 14473 10523
rect 14507 10520 14519 10523
rect 15378 10520 15384 10532
rect 14507 10492 15384 10520
rect 14507 10489 14519 10492
rect 14461 10483 14519 10489
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 23492 10520 23520 10551
rect 26418 10548 26424 10560
rect 26476 10588 26482 10600
rect 26973 10591 27031 10597
rect 26973 10588 26985 10591
rect 26476 10560 26985 10588
rect 26476 10548 26482 10560
rect 26973 10557 26985 10560
rect 27019 10557 27031 10591
rect 27522 10588 27528 10600
rect 27483 10560 27528 10588
rect 26973 10551 27031 10557
rect 27522 10548 27528 10560
rect 27580 10588 27586 10600
rect 28077 10591 28135 10597
rect 28077 10588 28089 10591
rect 27580 10560 28089 10588
rect 27580 10548 27586 10560
rect 28077 10557 28089 10560
rect 28123 10557 28135 10591
rect 28077 10551 28135 10557
rect 24302 10520 24308 10532
rect 23492 10492 24308 10520
rect 24302 10480 24308 10492
rect 24360 10480 24366 10532
rect 4522 10452 4528 10464
rect 4483 10424 4528 10452
rect 4522 10412 4528 10424
rect 4580 10412 4586 10464
rect 6178 10452 6184 10464
rect 6139 10424 6184 10452
rect 6178 10412 6184 10424
rect 6236 10412 6242 10464
rect 7466 10452 7472 10464
rect 7427 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 7926 10452 7932 10464
rect 7887 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 9214 10452 9220 10464
rect 9175 10424 9220 10452
rect 9214 10412 9220 10424
rect 9272 10452 9278 10464
rect 10134 10452 10140 10464
rect 9272 10424 10140 10452
rect 9272 10412 9278 10424
rect 10134 10412 10140 10424
rect 10192 10412 10198 10464
rect 10226 10412 10232 10464
rect 10284 10452 10290 10464
rect 10870 10452 10876 10464
rect 10284 10424 10329 10452
rect 10831 10424 10876 10452
rect 10284 10412 10290 10424
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11072 10452 11100 10480
rect 11241 10455 11299 10461
rect 11241 10452 11253 10455
rect 11072 10424 11253 10452
rect 11241 10421 11253 10424
rect 11287 10452 11299 10455
rect 11606 10452 11612 10464
rect 11287 10424 11612 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11606 10412 11612 10424
rect 11664 10412 11670 10464
rect 14918 10452 14924 10464
rect 14879 10424 14924 10452
rect 14918 10412 14924 10424
rect 14976 10412 14982 10464
rect 17862 10452 17868 10464
rect 17823 10424 17868 10452
rect 17862 10412 17868 10424
rect 17920 10412 17926 10464
rect 18782 10452 18788 10464
rect 18695 10424 18788 10452
rect 18782 10412 18788 10424
rect 18840 10452 18846 10464
rect 19337 10455 19395 10461
rect 19337 10452 19349 10455
rect 18840 10424 19349 10452
rect 18840 10412 18846 10424
rect 19337 10421 19349 10424
rect 19383 10421 19395 10455
rect 19337 10415 19395 10421
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23845 10455 23903 10461
rect 23845 10452 23857 10455
rect 23532 10424 23857 10452
rect 23532 10412 23538 10424
rect 23845 10421 23857 10424
rect 23891 10421 23903 10455
rect 24210 10452 24216 10464
rect 24171 10424 24216 10452
rect 23845 10415 23903 10421
rect 24210 10412 24216 10424
rect 24268 10412 24274 10464
rect 26602 10452 26608 10464
rect 26563 10424 26608 10452
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27706 10452 27712 10464
rect 27667 10424 27712 10452
rect 27706 10412 27712 10424
rect 27764 10412 27770 10464
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 2130 10248 2136 10260
rect 2091 10220 2136 10248
rect 2130 10208 2136 10220
rect 2188 10208 2194 10260
rect 2498 10248 2504 10260
rect 2459 10220 2504 10248
rect 2498 10208 2504 10220
rect 2556 10208 2562 10260
rect 4338 10248 4344 10260
rect 4299 10220 4344 10248
rect 4338 10208 4344 10220
rect 4396 10208 4402 10260
rect 4709 10251 4767 10257
rect 4709 10217 4721 10251
rect 4755 10248 4767 10251
rect 4798 10248 4804 10260
rect 4755 10220 4804 10248
rect 4755 10217 4767 10220
rect 4709 10211 4767 10217
rect 4798 10208 4804 10220
rect 4856 10208 4862 10260
rect 4982 10248 4988 10260
rect 4943 10220 4988 10248
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 7558 10248 7564 10260
rect 7519 10220 7564 10248
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 7837 10251 7895 10257
rect 7837 10248 7849 10251
rect 7800 10220 7849 10248
rect 7800 10208 7806 10220
rect 7837 10217 7849 10220
rect 7883 10217 7895 10251
rect 8018 10248 8024 10260
rect 7979 10220 8024 10248
rect 7837 10211 7895 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 12342 10208 12348 10260
rect 12400 10248 12406 10260
rect 12437 10251 12495 10257
rect 12437 10248 12449 10251
rect 12400 10220 12449 10248
rect 12400 10208 12406 10220
rect 12437 10217 12449 10220
rect 12483 10217 12495 10251
rect 12437 10211 12495 10217
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15654 10248 15660 10260
rect 15344 10220 15660 10248
rect 15344 10208 15350 10220
rect 15654 10208 15660 10220
rect 15712 10248 15718 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15712 10220 15761 10248
rect 15712 10208 15718 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10248 18383 10251
rect 18506 10248 18512 10260
rect 18371 10220 18512 10248
rect 18371 10217 18383 10220
rect 18325 10211 18383 10217
rect 18506 10208 18512 10220
rect 18564 10208 18570 10260
rect 22002 10208 22008 10260
rect 22060 10248 22066 10260
rect 22281 10251 22339 10257
rect 22281 10248 22293 10251
rect 22060 10220 22293 10248
rect 22060 10208 22066 10220
rect 22281 10217 22293 10220
rect 22327 10217 22339 10251
rect 22281 10211 22339 10217
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 25317 10251 25375 10257
rect 25317 10248 25329 10251
rect 24268 10220 25329 10248
rect 24268 10208 24274 10220
rect 25317 10217 25329 10220
rect 25363 10217 25375 10251
rect 25317 10211 25375 10217
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8389 10183 8447 10189
rect 8389 10180 8401 10183
rect 8352 10152 8401 10180
rect 8352 10140 8358 10152
rect 8389 10149 8401 10152
rect 8435 10180 8447 10183
rect 9582 10180 9588 10192
rect 8435 10152 9588 10180
rect 8435 10149 8447 10152
rect 8389 10143 8447 10149
rect 9582 10140 9588 10152
rect 9640 10140 9646 10192
rect 18233 10183 18291 10189
rect 18233 10149 18245 10183
rect 18279 10180 18291 10183
rect 18966 10180 18972 10192
rect 18279 10152 18972 10180
rect 18279 10149 18291 10152
rect 18233 10143 18291 10149
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 23658 10140 23664 10192
rect 23716 10180 23722 10192
rect 24121 10183 24179 10189
rect 24121 10180 24133 10183
rect 23716 10152 24133 10180
rect 23716 10140 23722 10152
rect 24121 10149 24133 10152
rect 24167 10149 24179 10183
rect 24121 10143 24179 10149
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 8481 10115 8539 10121
rect 1443 10084 2452 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 2424 9988 2452 10084
rect 8481 10081 8493 10115
rect 8527 10112 8539 10115
rect 8938 10112 8944 10124
rect 8527 10084 8944 10112
rect 8527 10081 8539 10084
rect 8481 10075 8539 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 11146 10072 11152 10124
rect 11204 10112 11210 10124
rect 11313 10115 11371 10121
rect 11313 10112 11325 10115
rect 11204 10084 11325 10112
rect 11204 10072 11210 10084
rect 11313 10081 11325 10084
rect 11359 10081 11371 10115
rect 11313 10075 11371 10081
rect 14918 10072 14924 10124
rect 14976 10112 14982 10124
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 14976 10084 15669 10112
rect 14976 10072 14982 10084
rect 15657 10081 15669 10084
rect 15703 10112 15715 10115
rect 15746 10112 15752 10124
rect 15703 10084 15752 10112
rect 15703 10081 15715 10084
rect 15657 10075 15715 10081
rect 15746 10072 15752 10084
rect 15804 10072 15810 10124
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18690 10112 18696 10124
rect 18104 10084 18696 10112
rect 18104 10072 18110 10084
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 21157 10115 21215 10121
rect 21157 10112 21169 10115
rect 20864 10084 21169 10112
rect 20864 10072 20870 10084
rect 21157 10081 21169 10084
rect 21203 10081 21215 10115
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 21157 10075 21215 10081
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 7466 10004 7472 10056
rect 7524 10044 7530 10056
rect 8110 10044 8116 10056
rect 7524 10016 8116 10044
rect 7524 10004 7530 10016
rect 8110 10004 8116 10016
rect 8168 10044 8174 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 8168 10016 8677 10044
rect 8168 10004 8174 10016
rect 8665 10013 8677 10016
rect 8711 10044 8723 10047
rect 8846 10044 8852 10056
rect 8711 10016 8852 10044
rect 8711 10013 8723 10016
rect 8665 10007 8723 10013
rect 8846 10004 8852 10016
rect 8904 10044 8910 10056
rect 10594 10044 10600 10056
rect 8904 10016 10600 10044
rect 8904 10004 8910 10016
rect 10594 10004 10600 10016
rect 10652 10004 10658 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10013 11115 10047
rect 11057 10007 11115 10013
rect 2406 9936 2412 9988
rect 2464 9976 2470 9988
rect 7282 9976 7288 9988
rect 2464 9948 7288 9976
rect 2464 9936 2470 9948
rect 7282 9936 7288 9948
rect 7340 9936 7346 9988
rect 1578 9908 1584 9920
rect 1539 9880 1584 9908
rect 1578 9868 1584 9880
rect 1636 9868 1642 9920
rect 2682 9868 2688 9920
rect 2740 9908 2746 9920
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2740 9880 2881 9908
rect 2740 9868 2746 9880
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 9858 9908 9864 9920
rect 9819 9880 9864 9908
rect 2869 9871 2927 9877
rect 9858 9868 9864 9880
rect 9916 9868 9922 9920
rect 11072 9908 11100 10007
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15436 10016 15853 10044
rect 15436 10004 15442 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18785 10047 18843 10053
rect 18785 10044 18797 10047
rect 18380 10016 18797 10044
rect 18380 10004 18386 10016
rect 18785 10013 18797 10016
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10044 19027 10047
rect 20901 10047 20959 10053
rect 19015 10016 19288 10044
rect 19015 10013 19027 10016
rect 18969 10007 19027 10013
rect 19260 9920 19288 10016
rect 20901 10013 20913 10047
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 11698 9908 11704 9920
rect 11072 9880 11704 9908
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 13722 9868 13728 9920
rect 13780 9908 13786 9920
rect 14274 9908 14280 9920
rect 13780 9880 14280 9908
rect 13780 9868 13786 9880
rect 14274 9868 14280 9880
rect 14332 9908 14338 9920
rect 14921 9911 14979 9917
rect 14921 9908 14933 9911
rect 14332 9880 14933 9908
rect 14332 9868 14338 9880
rect 14921 9877 14933 9880
rect 14967 9877 14979 9911
rect 15286 9908 15292 9920
rect 15247 9880 15292 9908
rect 14921 9871 14979 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 19242 9868 19248 9920
rect 19300 9908 19306 9920
rect 19337 9911 19395 9917
rect 19337 9908 19349 9911
rect 19300 9880 19349 9908
rect 19300 9868 19306 9880
rect 19337 9877 19349 9880
rect 19383 9877 19395 9911
rect 20916 9908 20944 10007
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 24210 10044 24216 10056
rect 23624 10016 24216 10044
rect 23624 10004 23630 10016
rect 24210 10004 24216 10016
rect 24268 10004 24274 10056
rect 24397 10047 24455 10053
rect 24397 10013 24409 10047
rect 24443 10044 24455 10047
rect 24578 10044 24584 10056
rect 24443 10016 24584 10044
rect 24443 10013 24455 10016
rect 24397 10007 24455 10013
rect 24578 10004 24584 10016
rect 24636 10004 24642 10056
rect 21634 9908 21640 9920
rect 20916 9880 21640 9908
rect 19337 9871 19395 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 23382 9868 23388 9920
rect 23440 9908 23446 9920
rect 23753 9911 23811 9917
rect 23753 9908 23765 9911
rect 23440 9880 23765 9908
rect 23440 9868 23446 9880
rect 23753 9877 23765 9880
rect 23799 9877 23811 9911
rect 24854 9908 24860 9920
rect 24815 9880 24860 9908
rect 23753 9871 23811 9877
rect 24854 9868 24860 9880
rect 24912 9868 24918 9920
rect 26697 9911 26755 9917
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 26786 9908 26792 9920
rect 26743 9880 26792 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 26786 9868 26792 9880
rect 26844 9868 26850 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2682 9664 2688 9716
rect 2740 9704 2746 9716
rect 3970 9704 3976 9716
rect 2740 9676 3648 9704
rect 3931 9676 3976 9704
rect 2740 9664 2746 9676
rect 3620 9509 3648 9676
rect 3970 9664 3976 9676
rect 4028 9664 4034 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 15654 9704 15660 9716
rect 15615 9676 15660 9704
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 16025 9707 16083 9713
rect 16025 9704 16037 9707
rect 15804 9676 16037 9704
rect 15804 9664 15810 9676
rect 16025 9673 16037 9676
rect 16071 9673 16083 9707
rect 18598 9704 18604 9716
rect 18559 9676 18604 9704
rect 16025 9667 16083 9673
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 23658 9664 23664 9716
rect 23716 9704 23722 9716
rect 23845 9707 23903 9713
rect 23845 9704 23857 9707
rect 23716 9676 23857 9704
rect 23716 9664 23722 9676
rect 23845 9673 23857 9676
rect 23891 9673 23903 9707
rect 23845 9667 23903 9673
rect 3988 9568 4016 9664
rect 7469 9639 7527 9645
rect 7469 9605 7481 9639
rect 7515 9636 7527 9639
rect 8312 9636 8340 9664
rect 7515 9608 8340 9636
rect 14645 9639 14703 9645
rect 7515 9605 7527 9608
rect 7469 9599 7527 9605
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 15396 9636 15424 9664
rect 19702 9636 19708 9648
rect 14691 9608 15424 9636
rect 19076 9608 19708 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 8481 9571 8539 9577
rect 3988 9540 4200 9568
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 3605 9503 3663 9509
rect 1443 9472 2084 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 2056 9373 2084 9472
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4062 9500 4068 9512
rect 3651 9472 4068 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 4172 9500 4200 9540
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 9493 9571 9551 9577
rect 9493 9568 9505 9571
rect 8527 9540 9505 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 9493 9537 9505 9540
rect 9539 9568 9551 9571
rect 9858 9568 9864 9580
rect 9539 9540 9864 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 9858 9528 9864 9540
rect 9916 9568 9922 9580
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 9916 9540 11069 9568
rect 9916 9528 9922 9540
rect 11057 9537 11069 9540
rect 11103 9568 11115 9571
rect 11146 9568 11152 9580
rect 11103 9540 11152 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 11146 9528 11152 9540
rect 11204 9528 11210 9580
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 18874 9568 18880 9580
rect 18472 9540 18880 9568
rect 18472 9528 18478 9540
rect 18874 9528 18880 9540
rect 18932 9568 18938 9580
rect 19076 9577 19104 9608
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 19978 9636 19984 9648
rect 19939 9608 19984 9636
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 23860 9636 23888 9667
rect 26510 9664 26516 9716
rect 26568 9704 26574 9716
rect 26605 9707 26663 9713
rect 26605 9704 26617 9707
rect 26568 9676 26617 9704
rect 26568 9664 26574 9676
rect 26605 9673 26617 9676
rect 26651 9673 26663 9707
rect 26605 9667 26663 9673
rect 26050 9636 26056 9648
rect 23860 9608 24716 9636
rect 26011 9608 26056 9636
rect 19061 9571 19119 9577
rect 19061 9568 19073 9571
rect 18932 9540 19073 9568
rect 18932 9528 18938 9540
rect 19061 9537 19073 9540
rect 19107 9537 19119 9571
rect 19061 9531 19119 9537
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 19245 9531 19303 9537
rect 4321 9503 4379 9509
rect 4321 9500 4333 9503
rect 4172 9472 4333 9500
rect 4321 9469 4333 9472
rect 4367 9469 4379 9503
rect 4321 9463 4379 9469
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 7926 9500 7932 9512
rect 7791 9472 7932 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 9306 9500 9312 9512
rect 9267 9472 9312 9500
rect 9306 9460 9312 9472
rect 9364 9460 9370 9512
rect 10042 9460 10048 9512
rect 10100 9500 10106 9512
rect 17770 9500 17776 9512
rect 10100 9472 17776 9500
rect 10100 9460 10106 9472
rect 17770 9460 17776 9472
rect 17828 9500 17834 9512
rect 17828 9472 19012 9500
rect 17828 9460 17834 9472
rect 9401 9435 9459 9441
rect 9401 9432 9413 9435
rect 8772 9404 9413 9432
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2130 9364 2136 9376
rect 2087 9336 2136 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9364 5503 9367
rect 5718 9364 5724 9376
rect 5491 9336 5724 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 7282 9324 7288 9376
rect 7340 9364 7346 9376
rect 7561 9367 7619 9373
rect 7561 9364 7573 9367
rect 7340 9336 7573 9364
rect 7340 9324 7346 9336
rect 7561 9333 7573 9336
rect 7607 9333 7619 9367
rect 7561 9327 7619 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 8772 9373 8800 9404
rect 9401 9401 9413 9404
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 13173 9435 13231 9441
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13532 9435 13590 9441
rect 13532 9432 13544 9435
rect 13219 9404 13544 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13532 9401 13544 9404
rect 13578 9432 13590 9435
rect 13722 9432 13728 9444
rect 13578 9404 13728 9432
rect 13578 9401 13590 9404
rect 13532 9395 13590 9401
rect 13722 9392 13728 9404
rect 13780 9392 13786 9444
rect 17497 9435 17555 9441
rect 17497 9401 17509 9435
rect 17543 9432 17555 9435
rect 17862 9432 17868 9444
rect 17543 9404 17868 9432
rect 17543 9401 17555 9404
rect 17497 9395 17555 9401
rect 17862 9392 17868 9404
rect 17920 9392 17926 9444
rect 18984 9376 19012 9472
rect 19260 9444 19288 9531
rect 19996 9500 20024 9596
rect 21910 9568 21916 9580
rect 21823 9540 21916 9568
rect 21910 9528 21916 9540
rect 21968 9568 21974 9580
rect 22646 9568 22652 9580
rect 21968 9540 22652 9568
rect 21968 9528 21974 9540
rect 22646 9528 22652 9540
rect 22704 9528 22710 9580
rect 23477 9571 23535 9577
rect 23477 9537 23489 9571
rect 23523 9568 23535 9571
rect 24578 9568 24584 9580
rect 23523 9540 24584 9568
rect 23523 9537 23535 9540
rect 23477 9531 23535 9537
rect 24578 9528 24584 9540
rect 24636 9528 24642 9580
rect 24688 9568 24716 9608
rect 26050 9596 26056 9608
rect 26108 9596 26114 9648
rect 27338 9636 27344 9648
rect 27299 9608 27344 9636
rect 27338 9596 27344 9608
rect 27396 9596 27402 9648
rect 24688 9540 24808 9568
rect 20349 9503 20407 9509
rect 20349 9500 20361 9503
rect 19996 9472 20361 9500
rect 20349 9469 20361 9472
rect 20395 9469 20407 9503
rect 20349 9463 20407 9469
rect 22094 9460 22100 9512
rect 22152 9500 22158 9512
rect 22465 9503 22523 9509
rect 22465 9500 22477 9503
rect 22152 9472 22477 9500
rect 22152 9460 22158 9472
rect 22465 9469 22477 9472
rect 22511 9500 22523 9503
rect 23382 9500 23388 9512
rect 22511 9472 23388 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 23382 9460 23388 9472
rect 23440 9460 23446 9512
rect 24670 9500 24676 9512
rect 24631 9472 24676 9500
rect 24670 9460 24676 9472
rect 24728 9460 24734 9512
rect 24780 9500 24808 9540
rect 27157 9503 27215 9509
rect 27157 9500 27169 9503
rect 24780 9472 27169 9500
rect 27157 9469 27169 9472
rect 27203 9500 27215 9503
rect 27709 9503 27767 9509
rect 27709 9500 27721 9503
rect 27203 9472 27721 9500
rect 27203 9469 27215 9472
rect 27157 9463 27215 9469
rect 27709 9469 27721 9472
rect 27755 9469 27767 9503
rect 27709 9463 27767 9469
rect 19242 9432 19248 9444
rect 19155 9404 19248 9432
rect 19242 9392 19248 9404
rect 19300 9432 19306 9444
rect 19705 9435 19763 9441
rect 19705 9432 19717 9435
rect 19300 9404 19717 9432
rect 19300 9392 19306 9404
rect 19705 9401 19717 9404
rect 19751 9432 19763 9435
rect 21545 9435 21603 9441
rect 19751 9404 20852 9432
rect 19751 9401 19763 9404
rect 19705 9395 19763 9401
rect 20824 9376 20852 9404
rect 21545 9401 21557 9435
rect 21591 9432 21603 9435
rect 22373 9435 22431 9441
rect 22373 9432 22385 9435
rect 21591 9404 22385 9432
rect 21591 9401 21603 9404
rect 21545 9395 21603 9401
rect 22373 9401 22385 9404
rect 22419 9432 22431 9435
rect 23474 9432 23480 9444
rect 22419 9404 23480 9432
rect 22419 9401 22431 9404
rect 22373 9395 22431 9401
rect 23474 9392 23480 9404
rect 23532 9392 23538 9444
rect 24578 9392 24584 9444
rect 24636 9432 24642 9444
rect 24918 9435 24976 9441
rect 24918 9432 24930 9435
rect 24636 9404 24930 9432
rect 24636 9392 24642 9404
rect 24918 9401 24930 9404
rect 24964 9401 24976 9435
rect 24918 9395 24976 9401
rect 8757 9367 8815 9373
rect 8757 9364 8769 9367
rect 8352 9336 8769 9364
rect 8352 9324 8358 9336
rect 8757 9333 8769 9336
rect 8803 9333 8815 9367
rect 8938 9364 8944 9376
rect 8899 9336 8944 9364
rect 8757 9327 8815 9333
rect 8938 9324 8944 9336
rect 8996 9324 9002 9376
rect 11517 9367 11575 9373
rect 11517 9333 11529 9367
rect 11563 9364 11575 9367
rect 11698 9364 11704 9376
rect 11563 9336 11704 9364
rect 11563 9333 11575 9336
rect 11517 9327 11575 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 18414 9364 18420 9376
rect 18375 9336 18420 9364
rect 18414 9324 18420 9336
rect 18472 9324 18478 9376
rect 18966 9364 18972 9376
rect 18927 9336 18972 9364
rect 18966 9324 18972 9336
rect 19024 9324 19030 9376
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 20806 9324 20812 9376
rect 20864 9364 20870 9376
rect 20901 9367 20959 9373
rect 20901 9364 20913 9367
rect 20864 9336 20913 9364
rect 20864 9324 20870 9336
rect 20901 9333 20913 9336
rect 20947 9333 20959 9367
rect 20901 9327 20959 9333
rect 22005 9367 22063 9373
rect 22005 9333 22017 9367
rect 22051 9364 22063 9367
rect 22186 9364 22192 9376
rect 22051 9336 22192 9364
rect 22051 9333 22063 9336
rect 22005 9327 22063 9333
rect 22186 9324 22192 9336
rect 22244 9324 22250 9376
rect 24210 9364 24216 9376
rect 24171 9336 24216 9364
rect 24210 9324 24216 9336
rect 24268 9324 24274 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 5074 9160 5080 9172
rect 4847 9132 5080 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 5074 9120 5080 9132
rect 5132 9120 5138 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7926 9160 7932 9172
rect 7699 9132 7932 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7926 9120 7932 9132
rect 7984 9120 7990 9172
rect 8113 9163 8171 9169
rect 8113 9129 8125 9163
rect 8159 9160 8171 9163
rect 8938 9160 8944 9172
rect 8159 9132 8944 9160
rect 8159 9129 8171 9132
rect 8113 9123 8171 9129
rect 8938 9120 8944 9132
rect 8996 9120 9002 9172
rect 9033 9163 9091 9169
rect 9033 9129 9045 9163
rect 9079 9160 9091 9163
rect 9306 9160 9312 9172
rect 9079 9132 9312 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9582 9120 9588 9172
rect 9640 9160 9646 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9640 9132 9689 9160
rect 9640 9120 9646 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 9677 9123 9735 9129
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 13262 9160 13268 9172
rect 11756 9132 13268 9160
rect 11756 9120 11762 9132
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 18601 9163 18659 9169
rect 18601 9129 18613 9163
rect 18647 9160 18659 9163
rect 18782 9160 18788 9172
rect 18647 9132 18788 9160
rect 18647 9129 18659 9132
rect 18601 9123 18659 9129
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 18969 9163 19027 9169
rect 18969 9129 18981 9163
rect 19015 9160 19027 9163
rect 19058 9160 19064 9172
rect 19015 9132 19064 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 19058 9120 19064 9132
rect 19116 9120 19122 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 26694 9160 26700 9172
rect 22152 9132 22197 9160
rect 26655 9132 26700 9160
rect 22152 9120 22158 9132
rect 26694 9120 26700 9132
rect 26752 9120 26758 9172
rect 15378 9052 15384 9104
rect 15436 9092 15442 9104
rect 15534 9095 15592 9101
rect 15534 9092 15546 9095
rect 15436 9064 15546 9092
rect 15436 9052 15442 9064
rect 15534 9061 15546 9064
rect 15580 9061 15592 9095
rect 15534 9055 15592 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2406 9024 2412 9036
rect 1443 8996 2412 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2406 8984 2412 8996
rect 2464 8984 2470 9036
rect 5718 9033 5724 9036
rect 5712 9024 5724 9033
rect 5679 8996 5724 9024
rect 5712 8987 5724 8996
rect 5718 8984 5724 8987
rect 5776 8984 5782 9036
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 7984 8996 9505 9024
rect 7984 8984 7990 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 10042 9024 10048 9036
rect 9493 8987 9551 8993
rect 9600 8996 10048 9024
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 5442 8956 5448 8968
rect 4120 8928 5448 8956
rect 4120 8916 4126 8928
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9600 8956 9628 8996
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 18414 9024 18420 9036
rect 10152 8996 18420 9024
rect 8996 8928 9628 8956
rect 8996 8916 9002 8928
rect 9674 8916 9680 8968
rect 9732 8956 9738 8968
rect 9950 8956 9956 8968
rect 9732 8928 9956 8956
rect 9732 8916 9738 8928
rect 9950 8916 9956 8928
rect 10008 8956 10014 8968
rect 10152 8965 10180 8996
rect 18414 8984 18420 8996
rect 18472 8984 18478 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 19061 9027 19119 9033
rect 19061 9024 19073 9027
rect 18748 8996 19073 9024
rect 18748 8984 18754 8996
rect 19061 8993 19073 8996
rect 19107 9024 19119 9027
rect 19334 9024 19340 9036
rect 19107 8996 19340 9024
rect 19107 8993 19119 8996
rect 19061 8987 19119 8993
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 23842 9024 23848 9036
rect 23803 8996 23848 9024
rect 23842 8984 23848 8996
rect 23900 8984 23906 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 10137 8959 10195 8965
rect 10137 8956 10149 8959
rect 10008 8928 10149 8956
rect 10008 8916 10014 8928
rect 10137 8925 10149 8928
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10244 8888 10272 8919
rect 14458 8916 14464 8968
rect 14516 8956 14522 8968
rect 15194 8956 15200 8968
rect 14516 8928 15200 8956
rect 14516 8916 14522 8928
rect 15194 8916 15200 8928
rect 15252 8956 15258 8968
rect 15289 8959 15347 8965
rect 15289 8956 15301 8959
rect 15252 8928 15301 8956
rect 15252 8916 15258 8928
rect 15289 8925 15301 8928
rect 15335 8925 15347 8959
rect 19242 8956 19248 8968
rect 19203 8928 19248 8956
rect 15289 8919 15347 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 23934 8956 23940 8968
rect 23895 8928 23940 8956
rect 23934 8916 23940 8928
rect 23992 8916 23998 8968
rect 24121 8959 24179 8965
rect 24121 8925 24133 8959
rect 24167 8956 24179 8959
rect 24167 8928 24624 8956
rect 24167 8925 24179 8928
rect 24121 8919 24179 8925
rect 10502 8888 10508 8900
rect 9916 8860 10508 8888
rect 9916 8848 9922 8860
rect 10502 8848 10508 8860
rect 10560 8848 10566 8900
rect 18322 8888 18328 8900
rect 18283 8860 18328 8888
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 24596 8832 24624 8928
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 6822 8820 6828 8832
rect 6783 8792 6828 8820
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 9180 8792 9321 8820
rect 9180 8780 9186 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9309 8783 9367 8789
rect 16298 8780 16304 8832
rect 16356 8820 16362 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 16356 8792 16681 8820
rect 16356 8780 16362 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 21177 8823 21235 8829
rect 21177 8789 21189 8823
rect 21223 8820 21235 8823
rect 21634 8820 21640 8832
rect 21223 8792 21640 8820
rect 21223 8789 21235 8792
rect 21177 8783 21235 8789
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 23474 8820 23480 8832
rect 23435 8792 23480 8820
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 24578 8780 24584 8832
rect 24636 8820 24642 8832
rect 24673 8823 24731 8829
rect 24673 8820 24685 8823
rect 24636 8792 24685 8820
rect 24636 8780 24642 8792
rect 24673 8789 24685 8792
rect 24719 8789 24731 8823
rect 24673 8783 24731 8789
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2406 8616 2412 8628
rect 2367 8588 2412 8616
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 4614 8616 4620 8628
rect 4575 8588 4620 8616
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8573 8619 8631 8625
rect 8573 8616 8585 8619
rect 7984 8588 8585 8616
rect 7984 8576 7990 8588
rect 8573 8585 8585 8588
rect 8619 8585 8631 8619
rect 10502 8616 10508 8628
rect 10463 8588 10508 8616
rect 8573 8579 8631 8585
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 14458 8616 14464 8628
rect 14419 8588 14464 8616
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8616 15255 8619
rect 15378 8616 15384 8628
rect 15243 8588 15384 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 18690 8616 18696 8628
rect 18651 8588 18696 8616
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19058 8616 19064 8628
rect 19019 8588 19064 8616
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19429 8619 19487 8625
rect 19429 8585 19441 8619
rect 19475 8616 19487 8619
rect 20806 8616 20812 8628
rect 19475 8588 20812 8616
rect 19475 8585 19487 8588
rect 19429 8579 19487 8585
rect 20806 8576 20812 8588
rect 20864 8576 20870 8628
rect 23842 8616 23848 8628
rect 23803 8588 23848 8616
rect 23842 8576 23848 8588
rect 23900 8576 23906 8628
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 1581 8551 1639 8557
rect 1581 8548 1593 8551
rect 1452 8520 1593 8548
rect 1452 8508 1458 8520
rect 1581 8517 1593 8520
rect 1627 8517 1639 8551
rect 1581 8511 1639 8517
rect 23290 8508 23296 8560
rect 23348 8548 23354 8560
rect 24029 8551 24087 8557
rect 24029 8548 24041 8551
rect 23348 8520 24041 8548
rect 23348 8508 23354 8520
rect 24029 8517 24041 8520
rect 24075 8517 24087 8551
rect 24029 8511 24087 8517
rect 2038 8480 2044 8492
rect 1412 8452 2044 8480
rect 1412 8421 1440 8452
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8480 4307 8483
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 4295 8452 5273 8480
rect 4295 8449 4307 8452
rect 4249 8443 4307 8449
rect 5261 8449 5273 8452
rect 5307 8480 5319 8483
rect 5718 8480 5724 8492
rect 5307 8452 5724 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 8938 8480 8944 8492
rect 7524 8452 8944 8480
rect 7524 8440 7530 8452
rect 8938 8440 8944 8452
rect 8996 8440 9002 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8480 14887 8483
rect 16206 8480 16212 8492
rect 14875 8452 16212 8480
rect 14875 8449 14887 8452
rect 14829 8443 14887 8449
rect 16206 8440 16212 8452
rect 16264 8440 16270 8492
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 24578 8480 24584 8492
rect 23523 8452 24584 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 24578 8440 24584 8452
rect 24636 8480 24642 8492
rect 26142 8480 26148 8492
rect 24636 8452 26148 8480
rect 24636 8440 24642 8452
rect 26142 8440 26148 8452
rect 26200 8440 26206 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 5169 8415 5227 8421
rect 5169 8412 5181 8415
rect 4672 8384 5181 8412
rect 4672 8372 4678 8384
rect 5169 8381 5181 8384
rect 5215 8381 5227 8415
rect 9122 8412 9128 8424
rect 5169 8375 5227 8381
rect 8404 8384 9128 8412
rect 5074 8344 5080 8356
rect 5035 8316 5080 8344
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 5500 8316 6193 8344
rect 5500 8304 5506 8316
rect 6181 8313 6193 8316
rect 6227 8344 6239 8347
rect 7282 8344 7288 8356
rect 6227 8316 7288 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4672 8248 4721 8276
rect 4672 8236 4678 8248
rect 4709 8245 4721 8248
rect 4755 8245 4767 8279
rect 4709 8239 4767 8245
rect 8294 8236 8300 8288
rect 8352 8276 8358 8288
rect 8404 8276 8432 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 16114 8412 16120 8424
rect 15611 8384 16120 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 20162 8412 20168 8424
rect 19392 8384 20168 8412
rect 19392 8372 19398 8384
rect 20162 8372 20168 8384
rect 20220 8412 20226 8424
rect 21085 8415 21143 8421
rect 21085 8412 21097 8415
rect 20220 8384 21097 8412
rect 20220 8372 20226 8384
rect 21085 8381 21097 8384
rect 21131 8412 21143 8415
rect 21361 8415 21419 8421
rect 21361 8412 21373 8415
rect 21131 8384 21373 8412
rect 21131 8381 21143 8384
rect 21085 8375 21143 8381
rect 21361 8381 21373 8384
rect 21407 8381 21419 8415
rect 21361 8375 21419 8381
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8412 24455 8415
rect 24670 8412 24676 8424
rect 24443 8384 24676 8412
rect 24443 8381 24455 8384
rect 24397 8375 24455 8381
rect 24670 8372 24676 8384
rect 24728 8412 24734 8424
rect 25409 8415 25467 8421
rect 25409 8412 25421 8415
rect 24728 8384 25421 8412
rect 24728 8372 24734 8384
rect 25409 8381 25421 8384
rect 25455 8381 25467 8415
rect 25409 8375 25467 8381
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 9370 8347 9428 8353
rect 9370 8344 9382 8347
rect 9272 8316 9382 8344
rect 9272 8304 9278 8316
rect 9370 8313 9382 8316
rect 9416 8313 9428 8347
rect 9370 8307 9428 8313
rect 23109 8347 23167 8353
rect 23109 8313 23121 8347
rect 23155 8344 23167 8347
rect 23934 8344 23940 8356
rect 23155 8316 23940 8344
rect 23155 8313 23167 8316
rect 23109 8307 23167 8313
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 24489 8347 24547 8353
rect 24489 8313 24501 8347
rect 24535 8344 24547 8347
rect 24854 8344 24860 8356
rect 24535 8316 24860 8344
rect 24535 8313 24547 8316
rect 24489 8307 24547 8313
rect 24854 8304 24860 8316
rect 24912 8344 24918 8356
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 24912 8316 25053 8344
rect 24912 8304 24918 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 26510 8304 26516 8356
rect 26568 8344 26574 8356
rect 26605 8347 26663 8353
rect 26605 8344 26617 8347
rect 26568 8316 26617 8344
rect 26568 8304 26574 8316
rect 26605 8313 26617 8316
rect 26651 8344 26663 8347
rect 26970 8344 26976 8356
rect 26651 8316 26976 8344
rect 26651 8313 26663 8316
rect 26605 8307 26663 8313
rect 26970 8304 26976 8316
rect 27028 8304 27034 8356
rect 15654 8276 15660 8288
rect 8352 8248 8445 8276
rect 15615 8248 15660 8276
rect 8352 8236 8358 8248
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 16022 8276 16028 8288
rect 15983 8248 16028 8276
rect 16022 8236 16028 8248
rect 16080 8236 16086 8288
rect 20901 8279 20959 8285
rect 20901 8245 20913 8279
rect 20947 8276 20959 8279
rect 21634 8276 21640 8288
rect 20947 8248 21640 8276
rect 20947 8245 20959 8248
rect 20901 8239 20959 8245
rect 21634 8236 21640 8248
rect 21692 8236 21698 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 1486 8032 1492 8084
rect 1544 8072 1550 8084
rect 1581 8075 1639 8081
rect 1581 8072 1593 8075
rect 1544 8044 1593 8072
rect 1544 8032 1550 8044
rect 1581 8041 1593 8044
rect 1627 8041 1639 8075
rect 1581 8035 1639 8041
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 4246 8072 4252 8084
rect 3660 8044 4252 8072
rect 3660 8032 3666 8044
rect 4246 8032 4252 8044
rect 4304 8072 4310 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4304 8044 4537 8072
rect 4304 8032 4310 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 9214 8072 9220 8084
rect 9175 8044 9220 8072
rect 4525 8035 4583 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 10321 8075 10379 8081
rect 10321 8041 10333 8075
rect 10367 8072 10379 8075
rect 10502 8072 10508 8084
rect 10367 8044 10508 8072
rect 10367 8041 10379 8044
rect 10321 8035 10379 8041
rect 10502 8032 10508 8044
rect 10560 8032 10566 8084
rect 23934 8032 23940 8084
rect 23992 8072 23998 8084
rect 24305 8075 24363 8081
rect 24305 8072 24317 8075
rect 23992 8044 24317 8072
rect 23992 8032 23998 8044
rect 24305 8041 24317 8044
rect 24351 8041 24363 8075
rect 24305 8035 24363 8041
rect 24394 8032 24400 8084
rect 24452 8072 24458 8084
rect 24673 8075 24731 8081
rect 24673 8072 24685 8075
rect 24452 8044 24685 8072
rect 24452 8032 24458 8044
rect 24673 8041 24685 8044
rect 24719 8041 24731 8075
rect 24673 8035 24731 8041
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25866 8072 25872 8084
rect 25004 8044 25872 8072
rect 25004 8032 25010 8044
rect 25866 8032 25872 8044
rect 25924 8072 25930 8084
rect 26145 8075 26203 8081
rect 26145 8072 26157 8075
rect 25924 8044 26157 8072
rect 25924 8032 25930 8044
rect 26145 8041 26157 8044
rect 26191 8041 26203 8075
rect 26694 8072 26700 8084
rect 26655 8044 26700 8072
rect 26145 8035 26203 8041
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 16206 7964 16212 8016
rect 16264 8013 16270 8016
rect 16264 8007 16328 8013
rect 16264 7973 16282 8007
rect 16316 7973 16328 8007
rect 16264 7967 16328 7973
rect 21260 8007 21318 8013
rect 21260 7973 21272 8007
rect 21306 8004 21318 8007
rect 21450 8004 21456 8016
rect 21306 7976 21456 8004
rect 21306 7973 21318 7976
rect 21260 7967 21318 7973
rect 16264 7964 16270 7967
rect 21450 7964 21456 7976
rect 21508 8004 21514 8016
rect 21910 8004 21916 8016
rect 21508 7976 21916 8004
rect 21508 7964 21514 7976
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 24121 8007 24179 8013
rect 24121 7973 24133 8007
rect 24167 8004 24179 8007
rect 24578 8004 24584 8016
rect 24167 7976 24584 8004
rect 24167 7973 24179 7976
rect 24121 7967 24179 7973
rect 24578 7964 24584 7976
rect 24636 7964 24642 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1946 7936 1952 7948
rect 1443 7908 1952 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1946 7896 1952 7908
rect 2004 7896 2010 7948
rect 11974 7945 11980 7948
rect 11968 7936 11980 7945
rect 11935 7908 11980 7936
rect 11968 7899 11980 7908
rect 11974 7896 11980 7899
rect 12032 7896 12038 7948
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15746 7936 15752 7948
rect 15252 7908 15752 7936
rect 15252 7896 15258 7908
rect 15746 7896 15752 7908
rect 15804 7936 15810 7948
rect 16025 7939 16083 7945
rect 16025 7936 16037 7939
rect 15804 7908 16037 7936
rect 15804 7896 15810 7908
rect 16025 7905 16037 7908
rect 16071 7905 16083 7939
rect 16025 7899 16083 7905
rect 18598 7896 18604 7948
rect 18656 7936 18662 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18656 7908 18705 7936
rect 18656 7896 18662 7908
rect 18693 7905 18705 7908
rect 18739 7936 18751 7939
rect 19242 7936 19248 7948
rect 18739 7908 19248 7936
rect 18739 7905 18751 7908
rect 18693 7899 18751 7905
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 20993 7939 21051 7945
rect 20993 7905 21005 7939
rect 21039 7936 21051 7939
rect 21634 7936 21640 7948
rect 21039 7908 21640 7936
rect 21039 7905 21051 7908
rect 20993 7899 21051 7905
rect 21634 7896 21640 7908
rect 21692 7896 21698 7948
rect 26510 7936 26516 7948
rect 26471 7908 26516 7936
rect 26510 7896 26516 7908
rect 26568 7896 26574 7948
rect 4338 7828 4344 7880
rect 4396 7868 4402 7880
rect 4614 7868 4620 7880
rect 4396 7840 4620 7868
rect 4396 7828 4402 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4798 7868 4804 7880
rect 4759 7840 4804 7868
rect 4798 7828 4804 7840
rect 4856 7828 4862 7880
rect 5261 7871 5319 7877
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5534 7868 5540 7880
rect 5307 7840 5540 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5534 7828 5540 7840
rect 5592 7868 5598 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5592 7840 5825 7868
rect 5592 7828 5598 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 11698 7868 11704 7880
rect 11659 7840 11704 7868
rect 5813 7831 5871 7837
rect 11698 7828 11704 7840
rect 11756 7828 11762 7880
rect 24118 7828 24124 7880
rect 24176 7868 24182 7880
rect 24765 7871 24823 7877
rect 24765 7868 24777 7871
rect 24176 7840 24777 7868
rect 24176 7828 24182 7840
rect 24765 7837 24777 7840
rect 24811 7837 24823 7871
rect 24765 7831 24823 7837
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 24995 7840 25452 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 15657 7803 15715 7809
rect 15657 7800 15669 7803
rect 12636 7772 15669 7800
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 1912 7704 2053 7732
rect 1912 7692 1918 7704
rect 2041 7701 2053 7704
rect 2087 7732 2099 7735
rect 3878 7732 3884 7744
rect 2087 7704 3884 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4154 7732 4160 7744
rect 4115 7704 4160 7732
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 9950 7732 9956 7744
rect 9911 7704 9956 7732
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 12434 7692 12440 7744
rect 12492 7732 12498 7744
rect 12636 7732 12664 7772
rect 15657 7769 15669 7772
rect 15703 7800 15715 7803
rect 16022 7800 16028 7812
rect 15703 7772 16028 7800
rect 15703 7769 15715 7772
rect 15657 7763 15715 7769
rect 16022 7760 16028 7772
rect 16080 7760 16086 7812
rect 18506 7800 18512 7812
rect 18467 7772 18512 7800
rect 18506 7760 18512 7772
rect 18564 7800 18570 7812
rect 19518 7800 19524 7812
rect 18564 7772 19524 7800
rect 18564 7760 18570 7772
rect 19518 7760 19524 7772
rect 19576 7760 19582 7812
rect 25424 7744 25452 7840
rect 13078 7732 13084 7744
rect 12492 7704 12664 7732
rect 13039 7704 13084 7732
rect 12492 7692 12498 7704
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 17402 7732 17408 7744
rect 17363 7704 17408 7732
rect 17402 7692 17408 7704
rect 17460 7692 17466 7744
rect 22370 7732 22376 7744
rect 22331 7704 22376 7732
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 25406 7732 25412 7744
rect 25367 7704 25412 7732
rect 25406 7692 25412 7704
rect 25464 7692 25470 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 4246 7528 4252 7540
rect 4207 7500 4252 7528
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9674 7528 9680 7540
rect 9272 7500 9680 7528
rect 9272 7488 9278 7500
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 15197 7531 15255 7537
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15654 7528 15660 7540
rect 15243 7500 15660 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15654 7488 15660 7500
rect 15712 7528 15718 7540
rect 15712 7500 16160 7528
rect 15712 7488 15718 7500
rect 3878 7392 3884 7404
rect 3791 7364 3884 7392
rect 3878 7352 3884 7364
rect 3936 7392 3942 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 3936 7364 4721 7392
rect 3936 7352 3942 7364
rect 4709 7361 4721 7364
rect 4755 7392 4767 7395
rect 4798 7392 4804 7404
rect 4755 7364 4804 7392
rect 4755 7361 4767 7364
rect 4709 7355 4767 7361
rect 4798 7352 4804 7364
rect 4856 7392 4862 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 4856 7364 5825 7392
rect 4856 7352 4862 7364
rect 5813 7361 5825 7364
rect 5859 7392 5871 7395
rect 6822 7392 6828 7404
rect 5859 7364 6828 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 11974 7392 11980 7404
rect 8352 7364 8397 7392
rect 11808 7364 11980 7392
rect 8352 7352 8358 7364
rect 1854 7333 1860 7336
rect 1581 7327 1639 7333
rect 1581 7293 1593 7327
rect 1627 7293 1639 7327
rect 1848 7324 1860 7333
rect 1815 7296 1860 7324
rect 1581 7287 1639 7293
rect 1848 7287 1860 7296
rect 1596 7256 1624 7287
rect 1854 7284 1860 7287
rect 1912 7284 1918 7336
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 2682 7256 2688 7268
rect 1596 7228 2688 7256
rect 1872 7200 1900 7228
rect 2682 7216 2688 7228
rect 2740 7216 2746 7268
rect 5074 7256 5080 7268
rect 4987 7228 5080 7256
rect 5074 7216 5080 7228
rect 5132 7256 5138 7268
rect 8205 7259 8263 7265
rect 5132 7228 5672 7256
rect 5132 7216 5138 7228
rect 5644 7200 5672 7228
rect 8205 7225 8217 7259
rect 8251 7256 8263 7259
rect 8542 7259 8600 7265
rect 8542 7256 8554 7259
rect 8251 7228 8554 7256
rect 8251 7225 8263 7228
rect 8205 7219 8263 7225
rect 8542 7225 8554 7228
rect 8588 7256 8600 7259
rect 9858 7256 9864 7268
rect 8588 7228 9864 7256
rect 8588 7225 8600 7228
rect 8542 7219 8600 7225
rect 9858 7216 9864 7228
rect 9916 7216 9922 7268
rect 1854 7148 1860 7200
rect 1912 7148 1918 7200
rect 2774 7148 2780 7200
rect 2832 7188 2838 7200
rect 2961 7191 3019 7197
rect 2961 7188 2973 7191
rect 2832 7160 2973 7188
rect 2832 7148 2838 7160
rect 2961 7157 2973 7160
rect 3007 7157 3019 7191
rect 5166 7188 5172 7200
rect 5127 7160 5172 7188
rect 2961 7151 3019 7157
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5626 7188 5632 7200
rect 5587 7160 5632 7188
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 11422 7188 11428 7200
rect 11383 7160 11428 7188
rect 11422 7148 11428 7160
rect 11480 7188 11486 7200
rect 11808 7197 11836 7364
rect 11974 7352 11980 7364
rect 12032 7392 12038 7404
rect 13262 7392 13268 7404
rect 12032 7364 13268 7392
rect 12032 7352 12038 7364
rect 13262 7352 13268 7364
rect 13320 7352 13326 7404
rect 16132 7401 16160 7500
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 16669 7531 16727 7537
rect 16669 7528 16681 7531
rect 16356 7500 16681 7528
rect 16356 7488 16362 7500
rect 16669 7497 16681 7500
rect 16715 7497 16727 7531
rect 18598 7528 18604 7540
rect 18559 7500 18604 7528
rect 16669 7491 16727 7497
rect 18598 7488 18604 7500
rect 18656 7488 18662 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 21450 7528 21456 7540
rect 21411 7500 21456 7528
rect 20901 7491 20959 7497
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 23477 7531 23535 7537
rect 23477 7497 23489 7531
rect 23523 7528 23535 7531
rect 23566 7528 23572 7540
rect 23523 7500 23572 7528
rect 23523 7497 23535 7500
rect 23477 7491 23535 7497
rect 23566 7488 23572 7500
rect 23624 7528 23630 7540
rect 24394 7528 24400 7540
rect 23624 7500 24400 7528
rect 23624 7488 23630 7500
rect 24394 7488 24400 7500
rect 24452 7488 24458 7540
rect 24581 7531 24639 7537
rect 24581 7497 24593 7531
rect 24627 7528 24639 7531
rect 24670 7528 24676 7540
rect 24627 7500 24676 7528
rect 24627 7497 24639 7500
rect 24581 7491 24639 7497
rect 24670 7488 24676 7500
rect 24728 7488 24734 7540
rect 26326 7488 26332 7540
rect 26384 7528 26390 7540
rect 27525 7531 27583 7537
rect 27525 7528 27537 7531
rect 26384 7500 27537 7528
rect 26384 7488 26390 7500
rect 27525 7497 27537 7500
rect 27571 7497 27583 7531
rect 27525 7491 27583 7497
rect 25774 7460 25780 7472
rect 24964 7432 25780 7460
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7392 16267 7395
rect 17402 7392 17408 7404
rect 16255 7364 17408 7392
rect 16255 7361 16267 7364
rect 16209 7355 16267 7361
rect 13081 7327 13139 7333
rect 13081 7293 13093 7327
rect 13127 7324 13139 7327
rect 13170 7324 13176 7336
rect 13127 7296 13176 7324
rect 13127 7293 13139 7296
rect 13081 7287 13139 7293
rect 13170 7284 13176 7296
rect 13228 7284 13234 7336
rect 15378 7284 15384 7336
rect 15436 7324 15442 7336
rect 16224 7324 16252 7355
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 22370 7392 22376 7404
rect 21836 7364 22376 7392
rect 19518 7324 19524 7336
rect 15436 7296 16252 7324
rect 19479 7296 19524 7324
rect 15436 7284 15442 7296
rect 19518 7284 19524 7296
rect 19576 7284 19582 7336
rect 12158 7256 12164 7268
rect 12119 7228 12164 7256
rect 12158 7216 12164 7228
rect 12216 7256 12222 7268
rect 12989 7259 13047 7265
rect 12989 7256 13001 7259
rect 12216 7228 13001 7256
rect 12216 7216 12222 7228
rect 12989 7225 13001 7228
rect 13035 7225 13047 7259
rect 15562 7256 15568 7268
rect 15475 7228 15568 7256
rect 12989 7219 13047 7225
rect 15562 7216 15568 7228
rect 15620 7256 15626 7268
rect 16025 7259 16083 7265
rect 16025 7256 16037 7259
rect 15620 7228 16037 7256
rect 15620 7216 15626 7228
rect 16025 7225 16037 7228
rect 16071 7256 16083 7259
rect 16390 7256 16396 7268
rect 16071 7228 16396 7256
rect 16071 7225 16083 7228
rect 16025 7219 16083 7225
rect 16390 7216 16396 7228
rect 16448 7216 16454 7268
rect 21836 7265 21864 7364
rect 22370 7352 22376 7364
rect 22428 7392 22434 7404
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 22428 7364 22569 7392
rect 22428 7352 22434 7364
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 24302 7352 24308 7404
rect 24360 7392 24366 7404
rect 24397 7395 24455 7401
rect 24397 7392 24409 7395
rect 24360 7364 24409 7392
rect 24360 7352 24366 7364
rect 24397 7361 24409 7364
rect 24443 7361 24455 7395
rect 24397 7355 24455 7361
rect 19429 7259 19487 7265
rect 19429 7225 19441 7259
rect 19475 7256 19487 7259
rect 19766 7259 19824 7265
rect 19766 7256 19778 7259
rect 19475 7228 19778 7256
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 19766 7225 19778 7228
rect 19812 7256 19824 7259
rect 21821 7259 21879 7265
rect 21821 7256 21833 7259
rect 19812 7228 21833 7256
rect 19812 7225 19824 7228
rect 19766 7219 19824 7225
rect 21821 7225 21833 7228
rect 21867 7225 21879 7259
rect 21821 7219 21879 7225
rect 22186 7216 22192 7268
rect 22244 7256 22250 7268
rect 22373 7259 22431 7265
rect 22373 7256 22385 7259
rect 22244 7228 22385 7256
rect 22244 7216 22250 7228
rect 22373 7225 22385 7228
rect 22419 7225 22431 7259
rect 24412 7256 24440 7355
rect 24964 7336 24992 7432
rect 25774 7420 25780 7432
rect 25832 7420 25838 7472
rect 25225 7395 25283 7401
rect 25225 7361 25237 7395
rect 25271 7392 25283 7395
rect 25406 7392 25412 7404
rect 25271 7364 25412 7392
rect 25271 7361 25283 7364
rect 25225 7355 25283 7361
rect 25406 7352 25412 7364
rect 25464 7392 25470 7404
rect 25464 7364 25728 7392
rect 25464 7352 25470 7364
rect 24946 7324 24952 7336
rect 24859 7296 24952 7324
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 25038 7256 25044 7268
rect 24412 7228 25044 7256
rect 22373 7219 22431 7225
rect 25038 7216 25044 7228
rect 25096 7216 25102 7268
rect 25700 7256 25728 7364
rect 25866 7352 25872 7404
rect 25924 7392 25930 7404
rect 26145 7395 26203 7401
rect 26145 7392 26157 7395
rect 25924 7364 26157 7392
rect 25924 7352 25930 7364
rect 26145 7361 26157 7364
rect 26191 7361 26203 7395
rect 26145 7355 26203 7361
rect 26390 7259 26448 7265
rect 26390 7256 26402 7259
rect 25700 7228 26402 7256
rect 25700 7200 25728 7228
rect 26390 7225 26402 7228
rect 26436 7225 26448 7259
rect 26390 7219 26448 7225
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 11480 7160 11805 7188
rect 11480 7148 11486 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 12618 7188 12624 7200
rect 12579 7160 12624 7188
rect 11793 7151 11851 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 14182 7188 14188 7200
rect 14143 7160 14188 7188
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 17586 7148 17592 7200
rect 17644 7188 17650 7200
rect 18049 7191 18107 7197
rect 18049 7188 18061 7191
rect 17644 7160 18061 7188
rect 17644 7148 17650 7160
rect 18049 7157 18061 7160
rect 18095 7157 18107 7191
rect 18049 7151 18107 7157
rect 20254 7148 20260 7200
rect 20312 7188 20318 7200
rect 22005 7191 22063 7197
rect 22005 7188 22017 7191
rect 20312 7160 22017 7188
rect 20312 7148 20318 7160
rect 22005 7157 22017 7160
rect 22051 7157 22063 7191
rect 22462 7188 22468 7200
rect 22423 7160 22468 7188
rect 22005 7151 22063 7157
rect 22462 7148 22468 7160
rect 22520 7148 22526 7200
rect 24118 7188 24124 7200
rect 24079 7160 24124 7188
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 25682 7188 25688 7200
rect 25643 7160 25688 7188
rect 25682 7148 25688 7160
rect 25740 7148 25746 7200
rect 25958 7188 25964 7200
rect 25919 7160 25964 7188
rect 25958 7148 25964 7160
rect 26016 7188 26022 7200
rect 26510 7188 26516 7200
rect 26016 7160 26516 7188
rect 26016 7148 26022 7160
rect 26510 7148 26516 7160
rect 26568 7148 26574 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 1946 6984 1952 6996
rect 1907 6956 1952 6984
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 2409 6987 2467 6993
rect 2409 6953 2421 6987
rect 2455 6984 2467 6987
rect 2682 6984 2688 6996
rect 2455 6956 2688 6984
rect 2455 6953 2467 6956
rect 2409 6947 2467 6953
rect 2682 6944 2688 6956
rect 2740 6944 2746 6996
rect 3418 6944 3424 6996
rect 3476 6984 3482 6996
rect 5718 6984 5724 6996
rect 3476 6956 5724 6984
rect 3476 6944 3482 6956
rect 5718 6944 5724 6956
rect 5776 6984 5782 6996
rect 6178 6984 6184 6996
rect 5776 6956 6184 6984
rect 5776 6944 5782 6956
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 11698 6984 11704 6996
rect 8352 6956 11704 6984
rect 8352 6944 8358 6956
rect 11698 6944 11704 6956
rect 11756 6944 11762 6996
rect 12989 6987 13047 6993
rect 12989 6953 13001 6987
rect 13035 6984 13047 6987
rect 13170 6984 13176 6996
rect 13035 6956 13176 6984
rect 13035 6953 13047 6956
rect 12989 6947 13047 6953
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 14182 6984 14188 6996
rect 13863 6956 14188 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 14182 6944 14188 6956
rect 14240 6944 14246 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15804 6956 16037 6984
rect 15804 6944 15810 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 19518 6984 19524 6996
rect 19479 6956 19524 6984
rect 16025 6947 16083 6953
rect 19518 6944 19524 6956
rect 19576 6944 19582 6996
rect 22097 6987 22155 6993
rect 22097 6953 22109 6987
rect 22143 6984 22155 6987
rect 22462 6984 22468 6996
rect 22143 6956 22468 6984
rect 22143 6953 22155 6956
rect 22097 6947 22155 6953
rect 22462 6944 22468 6956
rect 22520 6984 22526 6996
rect 22649 6987 22707 6993
rect 22649 6984 22661 6987
rect 22520 6956 22661 6984
rect 22520 6944 22526 6956
rect 22649 6953 22661 6956
rect 22695 6953 22707 6987
rect 22649 6947 22707 6953
rect 23017 6987 23075 6993
rect 23017 6953 23029 6987
rect 23063 6984 23075 6987
rect 23382 6984 23388 6996
rect 23063 6956 23388 6984
rect 23063 6953 23075 6956
rect 23017 6947 23075 6953
rect 23382 6944 23388 6956
rect 23440 6944 23446 6996
rect 25225 6987 25283 6993
rect 25225 6953 25237 6987
rect 25271 6984 25283 6987
rect 25498 6984 25504 6996
rect 25271 6956 25504 6984
rect 25271 6953 25283 6956
rect 25225 6947 25283 6953
rect 25498 6944 25504 6956
rect 25556 6944 25562 6996
rect 4338 6916 4344 6928
rect 4080 6888 4344 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 1762 6848 1768 6860
rect 1443 6820 1768 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 4080 6848 4108 6888
rect 4338 6876 4344 6888
rect 4396 6876 4402 6928
rect 4617 6919 4675 6925
rect 4617 6885 4629 6919
rect 4663 6916 4675 6919
rect 5074 6916 5080 6928
rect 4663 6888 5080 6916
rect 4663 6885 4675 6888
rect 4617 6879 4675 6885
rect 5074 6876 5080 6888
rect 5132 6876 5138 6928
rect 10045 6919 10103 6925
rect 10045 6916 10057 6919
rect 9600 6888 10057 6916
rect 6270 6848 6276 6860
rect 3927 6820 4108 6848
rect 6231 6820 6276 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 9490 6808 9496 6860
rect 9548 6848 9554 6860
rect 9600 6848 9628 6888
rect 10045 6885 10057 6888
rect 10091 6916 10103 6919
rect 13078 6916 13084 6928
rect 10091 6888 11100 6916
rect 10091 6885 10103 6888
rect 10045 6879 10103 6885
rect 9548 6820 9628 6848
rect 11072 6848 11100 6888
rect 12084 6888 13084 6916
rect 12084 6860 12112 6888
rect 11072 6820 11928 6848
rect 9548 6808 9554 6820
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4396 6752 4721 6780
rect 4396 6740 4402 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 6457 6783 6515 6789
rect 4856 6752 4901 6780
rect 4856 6740 4862 6752
rect 6457 6749 6469 6783
rect 6503 6780 6515 6783
rect 6822 6780 6828 6792
rect 6503 6752 6828 6780
rect 6503 6749 6515 6752
rect 6457 6743 6515 6749
rect 6822 6740 6828 6752
rect 6880 6740 6886 6792
rect 9674 6740 9680 6792
rect 9732 6740 9738 6792
rect 10134 6780 10140 6792
rect 10095 6752 10140 6780
rect 10134 6740 10140 6752
rect 10192 6740 10198 6792
rect 10229 6783 10287 6789
rect 10229 6749 10241 6783
rect 10275 6749 10287 6783
rect 10229 6743 10287 6749
rect 1578 6712 1584 6724
rect 1539 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 9692 6712 9720 6740
rect 10244 6712 10272 6743
rect 11900 6721 11928 6820
rect 12066 6808 12072 6860
rect 12124 6808 12130 6860
rect 12250 6848 12256 6860
rect 12211 6820 12256 6848
rect 12250 6808 12256 6820
rect 12308 6808 12314 6860
rect 12342 6780 12348 6792
rect 12303 6752 12348 6780
rect 12342 6740 12348 6752
rect 12400 6740 12406 6792
rect 12544 6789 12572 6888
rect 13078 6876 13084 6888
rect 13136 6876 13142 6928
rect 13262 6876 13268 6928
rect 13320 6916 13326 6928
rect 13320 6888 13860 6916
rect 13320 6876 13326 6888
rect 13832 6848 13860 6888
rect 21450 6876 21456 6928
rect 21508 6916 21514 6928
rect 21508 6888 22140 6916
rect 21508 6876 21514 6888
rect 22112 6860 22140 6888
rect 22186 6876 22192 6928
rect 22244 6916 22250 6928
rect 22373 6919 22431 6925
rect 22373 6916 22385 6919
rect 22244 6888 22385 6916
rect 22244 6876 22250 6888
rect 22373 6885 22385 6888
rect 22419 6885 22431 6919
rect 24946 6916 24952 6928
rect 22373 6879 22431 6885
rect 24872 6888 24952 6916
rect 13832 6820 14136 6848
rect 12529 6783 12587 6789
rect 12529 6749 12541 6783
rect 12575 6749 12587 6783
rect 13906 6780 13912 6792
rect 13867 6752 13912 6780
rect 12529 6743 12587 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14108 6789 14136 6820
rect 17586 6808 17592 6860
rect 17644 6848 17650 6860
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 17644 6820 17877 6848
rect 17644 6808 17650 6820
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 18506 6848 18512 6860
rect 18467 6820 18512 6848
rect 17865 6811 17923 6817
rect 18506 6808 18512 6820
rect 18564 6808 18570 6860
rect 22094 6808 22100 6860
rect 22152 6808 22158 6860
rect 23109 6851 23167 6857
rect 23109 6817 23121 6851
rect 23155 6848 23167 6851
rect 23290 6848 23296 6860
rect 23155 6820 23296 6848
rect 23155 6817 23167 6820
rect 23109 6811 23167 6817
rect 23290 6808 23296 6820
rect 23348 6808 23354 6860
rect 24670 6848 24676 6860
rect 24583 6820 24676 6848
rect 24670 6808 24676 6820
rect 24728 6848 24734 6860
rect 24872 6848 24900 6888
rect 24946 6876 24952 6888
rect 25004 6876 25010 6928
rect 24728 6820 24900 6848
rect 26513 6851 26571 6857
rect 24728 6808 24734 6820
rect 26513 6817 26525 6851
rect 26559 6848 26571 6851
rect 26602 6848 26608 6860
rect 26559 6820 26608 6848
rect 26559 6817 26571 6820
rect 26513 6811 26571 6817
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14458 6780 14464 6792
rect 14139 6752 14464 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 17678 6740 17684 6792
rect 17736 6780 17742 6792
rect 17957 6783 18015 6789
rect 17957 6780 17969 6783
rect 17736 6752 17969 6780
rect 17736 6740 17742 6752
rect 17957 6749 17969 6752
rect 18003 6749 18015 6783
rect 17957 6743 18015 6749
rect 18049 6783 18107 6789
rect 18049 6749 18061 6783
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 9692 6684 10272 6712
rect 11885 6715 11943 6721
rect 11885 6681 11897 6715
rect 11931 6681 11943 6715
rect 11885 6675 11943 6681
rect 17402 6672 17408 6724
rect 17460 6712 17466 6724
rect 18064 6712 18092 6743
rect 22646 6740 22652 6792
rect 22704 6780 22710 6792
rect 23201 6783 23259 6789
rect 23201 6780 23213 6783
rect 22704 6752 23213 6780
rect 22704 6740 22710 6752
rect 23201 6749 23213 6752
rect 23247 6749 23259 6783
rect 23201 6743 23259 6749
rect 24946 6740 24952 6792
rect 25004 6780 25010 6792
rect 25317 6783 25375 6789
rect 25317 6780 25329 6783
rect 25004 6752 25329 6780
rect 25004 6740 25010 6752
rect 25317 6749 25329 6752
rect 25363 6749 25375 6783
rect 25317 6743 25375 6749
rect 25501 6783 25559 6789
rect 25501 6749 25513 6783
rect 25547 6780 25559 6783
rect 25682 6780 25688 6792
rect 25547 6752 25688 6780
rect 25547 6749 25559 6752
rect 25501 6743 25559 6749
rect 25682 6740 25688 6752
rect 25740 6780 25746 6792
rect 25740 6752 26280 6780
rect 25740 6740 25746 6752
rect 18322 6712 18328 6724
rect 17460 6684 18328 6712
rect 17460 6672 17466 6684
rect 18322 6672 18328 6684
rect 18380 6672 18386 6724
rect 24854 6712 24860 6724
rect 24815 6684 24860 6712
rect 24854 6672 24860 6684
rect 24912 6672 24918 6724
rect 4249 6647 4307 6653
rect 4249 6613 4261 6647
rect 4295 6644 4307 6647
rect 4614 6644 4620 6656
rect 4295 6616 4620 6644
rect 4295 6613 4307 6616
rect 4249 6607 4307 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5810 6644 5816 6656
rect 5771 6616 5816 6644
rect 5810 6604 5816 6616
rect 5868 6604 5874 6656
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6644 7711 6647
rect 7926 6644 7932 6656
rect 7699 6616 7932 6644
rect 7699 6613 7711 6616
rect 7653 6607 7711 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 9766 6644 9772 6656
rect 9723 6616 9772 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 12250 6604 12256 6656
rect 12308 6644 12314 6656
rect 13449 6647 13507 6653
rect 13449 6644 13461 6647
rect 12308 6616 13461 6644
rect 12308 6604 12314 6616
rect 13449 6613 13461 6616
rect 13495 6613 13507 6647
rect 13449 6607 13507 6613
rect 15378 6604 15384 6656
rect 15436 6644 15442 6656
rect 15657 6647 15715 6653
rect 15657 6644 15669 6647
rect 15436 6616 15669 6644
rect 15436 6604 15442 6616
rect 15657 6613 15669 6616
rect 15703 6613 15715 6647
rect 15657 6607 15715 6613
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6644 16543 6647
rect 16850 6644 16856 6656
rect 16531 6616 16856 6644
rect 16531 6613 16543 6616
rect 16485 6607 16543 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17494 6644 17500 6656
rect 17455 6616 17500 6644
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6644 20131 6647
rect 20438 6644 20444 6656
rect 20119 6616 20444 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6644 21235 6647
rect 21634 6644 21640 6656
rect 21223 6616 21640 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21634 6604 21640 6616
rect 21692 6604 21698 6656
rect 26252 6653 26280 6752
rect 26694 6712 26700 6724
rect 26655 6684 26700 6712
rect 26694 6672 26700 6684
rect 26752 6672 26758 6724
rect 26237 6647 26295 6653
rect 26237 6613 26249 6647
rect 26283 6644 26295 6647
rect 26326 6644 26332 6656
rect 26283 6616 26332 6644
rect 26283 6613 26295 6616
rect 26237 6607 26295 6613
rect 26326 6604 26332 6616
rect 26384 6604 26390 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1673 6443 1731 6449
rect 1673 6409 1685 6443
rect 1719 6440 1731 6443
rect 1762 6440 1768 6452
rect 1719 6412 1768 6440
rect 1719 6409 1731 6412
rect 1673 6403 1731 6409
rect 1762 6400 1768 6412
rect 1820 6400 1826 6452
rect 3789 6443 3847 6449
rect 3789 6409 3801 6443
rect 3835 6440 3847 6443
rect 4798 6440 4804 6452
rect 3835 6412 4804 6440
rect 3835 6409 3847 6412
rect 3789 6403 3847 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5813 6443 5871 6449
rect 5813 6440 5825 6443
rect 5776 6412 5825 6440
rect 5776 6400 5782 6412
rect 5813 6409 5825 6412
rect 5859 6409 5871 6443
rect 6270 6440 6276 6452
rect 6231 6412 6276 6440
rect 5813 6403 5871 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 6641 6443 6699 6449
rect 6641 6409 6653 6443
rect 6687 6440 6699 6443
rect 6822 6440 6828 6452
rect 6687 6412 6828 6440
rect 6687 6409 6699 6412
rect 6641 6403 6699 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7374 6440 7380 6452
rect 7335 6412 7380 6440
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 9079 6412 10057 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 10045 6409 10057 6412
rect 10091 6440 10103 6443
rect 10134 6440 10140 6452
rect 10091 6412 10140 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6440 11667 6443
rect 12250 6440 12256 6452
rect 11655 6412 12256 6440
rect 11655 6409 11667 6412
rect 11609 6403 11667 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 12618 6440 12624 6452
rect 12400 6412 12624 6440
rect 12400 6400 12406 6412
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6440 13967 6443
rect 14182 6440 14188 6452
rect 13955 6412 14188 6440
rect 13955 6409 13967 6412
rect 13909 6403 13967 6409
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 17770 6440 17776 6452
rect 17731 6412 17776 6440
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 22094 6400 22100 6452
rect 22152 6440 22158 6452
rect 22646 6440 22652 6452
rect 22152 6412 22652 6440
rect 22152 6400 22158 6412
rect 22646 6400 22652 6412
rect 22704 6400 22710 6452
rect 23109 6443 23167 6449
rect 23109 6409 23121 6443
rect 23155 6440 23167 6443
rect 23290 6440 23296 6452
rect 23155 6412 23296 6440
rect 23155 6409 23167 6412
rect 23109 6403 23167 6409
rect 23290 6400 23296 6412
rect 23348 6400 23354 6452
rect 23474 6440 23480 6452
rect 23435 6412 23480 6440
rect 23474 6400 23480 6412
rect 23532 6400 23538 6452
rect 24854 6440 24860 6452
rect 24815 6412 24860 6440
rect 24854 6400 24860 6412
rect 24912 6400 24918 6452
rect 25317 6443 25375 6449
rect 25317 6409 25329 6443
rect 25363 6440 25375 6443
rect 25498 6440 25504 6452
rect 25363 6412 25504 6440
rect 25363 6409 25375 6412
rect 25317 6403 25375 6409
rect 25498 6400 25504 6412
rect 25556 6400 25562 6452
rect 25685 6443 25743 6449
rect 25685 6409 25697 6443
rect 25731 6440 25743 6443
rect 26326 6440 26332 6452
rect 25731 6412 26332 6440
rect 25731 6409 25743 6412
rect 25685 6403 25743 6409
rect 26326 6400 26332 6412
rect 26384 6400 26390 6452
rect 26602 6400 26608 6452
rect 26660 6440 26666 6452
rect 26973 6443 27031 6449
rect 26973 6440 26985 6443
rect 26660 6412 26985 6440
rect 26660 6400 26666 6412
rect 26973 6409 26985 6412
rect 27019 6409 27031 6443
rect 26973 6403 27031 6409
rect 3694 6332 3700 6384
rect 3752 6372 3758 6384
rect 4065 6375 4123 6381
rect 4065 6372 4077 6375
rect 3752 6344 4077 6372
rect 3752 6332 3758 6344
rect 4065 6341 4077 6344
rect 4111 6372 4123 6375
rect 5074 6372 5080 6384
rect 4111 6344 5080 6372
rect 4111 6341 4123 6344
rect 4065 6335 4123 6341
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 9674 6372 9680 6384
rect 9635 6344 9680 6372
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 17405 6375 17463 6381
rect 17405 6372 17417 6375
rect 13924 6344 17417 6372
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 4212 6276 4721 6304
rect 4212 6264 4218 6276
rect 4709 6273 4721 6276
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 4798 6264 4804 6316
rect 4856 6304 4862 6316
rect 5258 6304 5264 6316
rect 4856 6276 5264 6304
rect 4856 6264 4862 6276
rect 5258 6264 5264 6276
rect 5316 6264 5322 6316
rect 8110 6304 8116 6316
rect 8071 6276 8116 6304
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10597 6307 10655 6313
rect 10597 6304 10609 6307
rect 9916 6276 10609 6304
rect 9916 6264 9922 6276
rect 10597 6273 10609 6276
rect 10643 6304 10655 6307
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 10643 6276 11897 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 11885 6273 11897 6276
rect 11931 6304 11943 6307
rect 12066 6304 12072 6316
rect 11931 6276 12072 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 13924 6248 13952 6344
rect 17405 6341 17417 6344
rect 17451 6372 17463 6375
rect 17678 6372 17684 6384
rect 17451 6344 17684 6372
rect 17451 6341 17463 6344
rect 17405 6335 17463 6341
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 16942 6304 16948 6316
rect 16903 6276 16948 6304
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18380 6276 18613 6304
rect 18380 6264 18386 6276
rect 18601 6273 18613 6276
rect 18647 6304 18659 6307
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 18647 6276 19073 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 20438 6304 20444 6316
rect 20399 6276 20444 6304
rect 19061 6267 19119 6273
rect 20438 6264 20444 6276
rect 20496 6264 20502 6316
rect 20533 6307 20591 6313
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 1765 6239 1823 6245
rect 1765 6205 1777 6239
rect 1811 6236 1823 6239
rect 1854 6236 1860 6248
rect 1811 6208 1860 6236
rect 1811 6205 1823 6208
rect 1765 6199 1823 6205
rect 1854 6196 1860 6208
rect 1912 6196 1918 6248
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 8021 6239 8079 6245
rect 8021 6236 8033 6239
rect 7432 6208 8033 6236
rect 7432 6196 7438 6208
rect 8021 6205 8033 6208
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 13449 6239 13507 6245
rect 13449 6236 13461 6239
rect 12308 6208 13461 6236
rect 12308 6196 12314 6208
rect 13449 6205 13461 6208
rect 13495 6236 13507 6239
rect 13906 6236 13912 6248
rect 13495 6208 13912 6236
rect 13495 6205 13507 6208
rect 13449 6199 13507 6205
rect 13906 6196 13912 6208
rect 13964 6196 13970 6248
rect 15933 6239 15991 6245
rect 15933 6205 15945 6239
rect 15979 6236 15991 6239
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 15979 6208 16773 6236
rect 15979 6205 15991 6208
rect 15933 6199 15991 6205
rect 16761 6205 16773 6208
rect 16807 6236 16819 6239
rect 17494 6236 17500 6248
rect 16807 6208 17500 6236
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 17828 6208 18429 6236
rect 17828 6196 17834 6208
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 19889 6239 19947 6245
rect 18564 6208 18609 6236
rect 18564 6196 18570 6208
rect 19889 6205 19901 6239
rect 19935 6236 19947 6239
rect 19978 6236 19984 6248
rect 19935 6208 19984 6236
rect 19935 6205 19947 6208
rect 19889 6199 19947 6205
rect 19978 6196 19984 6208
rect 20036 6236 20042 6248
rect 20548 6236 20576 6267
rect 20036 6208 20576 6236
rect 26421 6239 26479 6245
rect 20036 6196 20042 6208
rect 26421 6205 26433 6239
rect 26467 6205 26479 6239
rect 26421 6199 26479 6205
rect 2038 6177 2044 6180
rect 2032 6168 2044 6177
rect 1951 6140 2044 6168
rect 2032 6131 2044 6140
rect 2096 6168 2102 6180
rect 2682 6168 2688 6180
rect 2096 6140 2688 6168
rect 2038 6128 2044 6131
rect 2096 6128 2102 6140
rect 2682 6128 2688 6140
rect 2740 6128 2746 6180
rect 10413 6171 10471 6177
rect 10413 6137 10425 6171
rect 10459 6168 10471 6171
rect 10778 6168 10784 6180
rect 10459 6140 10784 6168
rect 10459 6137 10471 6140
rect 10413 6131 10471 6137
rect 10778 6128 10784 6140
rect 10836 6168 10842 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10836 6140 11069 6168
rect 10836 6128 10842 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 16301 6171 16359 6177
rect 16301 6137 16313 6171
rect 16347 6168 16359 6171
rect 16482 6168 16488 6180
rect 16347 6140 16488 6168
rect 16347 6137 16359 6140
rect 16301 6131 16359 6137
rect 16482 6128 16488 6140
rect 16540 6168 16546 6180
rect 16942 6168 16948 6180
rect 16540 6140 16948 6168
rect 16540 6128 16546 6140
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 19521 6171 19579 6177
rect 19521 6137 19533 6171
rect 19567 6168 19579 6171
rect 20349 6171 20407 6177
rect 20349 6168 20361 6171
rect 19567 6140 20361 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 20349 6137 20361 6140
rect 20395 6168 20407 6171
rect 20530 6168 20536 6180
rect 20395 6140 20536 6168
rect 20395 6137 20407 6140
rect 20349 6131 20407 6137
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 26234 6168 26240 6180
rect 26195 6140 26240 6168
rect 26234 6128 26240 6140
rect 26292 6168 26298 6180
rect 26436 6168 26464 6199
rect 26292 6140 26464 6168
rect 26292 6128 26298 6140
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 3145 6103 3203 6109
rect 3145 6100 3157 6103
rect 3016 6072 3157 6100
rect 3016 6060 3022 6072
rect 3145 6069 3157 6072
rect 3191 6069 3203 6103
rect 4246 6100 4252 6112
rect 4207 6072 4252 6100
rect 3145 6063 3203 6069
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4614 6100 4620 6112
rect 4575 6072 4620 6100
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 7101 6103 7159 6109
rect 7101 6069 7113 6103
rect 7147 6100 7159 6103
rect 7190 6100 7196 6112
rect 7147 6072 7196 6100
rect 7147 6069 7159 6072
rect 7101 6063 7159 6069
rect 7190 6060 7196 6072
rect 7248 6060 7254 6112
rect 7561 6103 7619 6109
rect 7561 6069 7573 6103
rect 7607 6100 7619 6103
rect 7742 6100 7748 6112
rect 7607 6072 7748 6100
rect 7607 6069 7619 6072
rect 7561 6063 7619 6069
rect 7742 6060 7748 6072
rect 7800 6060 7806 6112
rect 7926 6100 7932 6112
rect 7887 6072 7932 6100
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 10502 6100 10508 6112
rect 9447 6072 10508 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 14277 6103 14335 6109
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14458 6100 14464 6112
rect 14323 6072 14464 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 16393 6103 16451 6109
rect 16393 6069 16405 6103
rect 16439 6100 16451 6103
rect 16574 6100 16580 6112
rect 16439 6072 16580 6100
rect 16439 6069 16451 6072
rect 16393 6063 16451 6069
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 16850 6100 16856 6112
rect 16811 6072 16856 6100
rect 16850 6060 16856 6072
rect 16908 6100 16914 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 16908 6072 18061 6100
rect 16908 6060 16914 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 19981 6103 20039 6109
rect 19981 6069 19993 6103
rect 20027 6100 20039 6103
rect 20714 6100 20720 6112
rect 20027 6072 20720 6100
rect 20027 6069 20039 6072
rect 19981 6063 20039 6069
rect 20714 6060 20720 6072
rect 20772 6060 20778 6112
rect 26602 6100 26608 6112
rect 26563 6072 26608 6100
rect 26602 6060 26608 6072
rect 26660 6060 26666 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2038 5896 2044 5908
rect 1999 5868 2044 5896
rect 2038 5856 2044 5868
rect 2096 5856 2102 5908
rect 2225 5899 2283 5905
rect 2225 5865 2237 5899
rect 2271 5896 2283 5899
rect 2774 5896 2780 5908
rect 2271 5868 2780 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3513 5899 3571 5905
rect 3513 5865 3525 5899
rect 3559 5896 3571 5899
rect 4614 5896 4620 5908
rect 3559 5868 4620 5896
rect 3559 5865 3571 5868
rect 3513 5859 3571 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5077 5899 5135 5905
rect 5077 5865 5089 5899
rect 5123 5896 5135 5899
rect 5442 5896 5448 5908
rect 5123 5868 5448 5896
rect 5123 5865 5135 5868
rect 5077 5859 5135 5865
rect 5442 5856 5448 5868
rect 5500 5896 5506 5908
rect 5810 5896 5816 5908
rect 5500 5868 5816 5896
rect 5500 5856 5506 5868
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 9490 5896 9496 5908
rect 9451 5868 9496 5896
rect 9490 5856 9496 5868
rect 9548 5856 9554 5908
rect 9858 5856 9864 5908
rect 9916 5896 9922 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 9916 5868 10057 5896
rect 9916 5856 9922 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 10045 5859 10103 5865
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 10735 5868 11253 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 11241 5865 11253 5868
rect 11287 5896 11299 5899
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 11287 5868 12357 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 12710 5896 12716 5908
rect 12492 5868 12716 5896
rect 12492 5856 12498 5868
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 17586 5896 17592 5908
rect 17547 5868 17592 5896
rect 17586 5856 17592 5868
rect 17644 5856 17650 5908
rect 18230 5896 18236 5908
rect 18191 5868 18236 5896
rect 18230 5856 18236 5868
rect 18288 5856 18294 5908
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 20901 5899 20959 5905
rect 20901 5896 20913 5899
rect 20496 5868 20913 5896
rect 20496 5856 20502 5868
rect 20901 5865 20913 5868
rect 20947 5865 20959 5899
rect 20901 5859 20959 5865
rect 21269 5899 21327 5905
rect 21269 5865 21281 5899
rect 21315 5896 21327 5899
rect 21726 5896 21732 5908
rect 21315 5868 21732 5896
rect 21315 5865 21327 5868
rect 21269 5859 21327 5865
rect 21726 5856 21732 5868
rect 21784 5896 21790 5908
rect 26970 5896 26976 5908
rect 21784 5868 26976 5896
rect 21784 5856 21790 5868
rect 26970 5856 26976 5868
rect 27028 5856 27034 5908
rect 3881 5831 3939 5837
rect 3881 5797 3893 5831
rect 3927 5828 3939 5831
rect 4154 5828 4160 5840
rect 3927 5800 4160 5828
rect 3927 5797 3939 5800
rect 3881 5791 3939 5797
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 4985 5831 5043 5837
rect 4985 5797 4997 5831
rect 5031 5828 5043 5831
rect 5166 5828 5172 5840
rect 5031 5800 5172 5828
rect 5031 5797 5043 5800
rect 4985 5791 5043 5797
rect 5166 5788 5172 5800
rect 5224 5788 5230 5840
rect 11146 5828 11152 5840
rect 11059 5800 11152 5828
rect 11146 5788 11152 5800
rect 11204 5828 11210 5840
rect 15010 5828 15016 5840
rect 11204 5800 15016 5828
rect 11204 5788 11210 5800
rect 15010 5788 15016 5800
rect 15068 5788 15074 5840
rect 15746 5828 15752 5840
rect 15304 5800 15752 5828
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 2406 5760 2412 5772
rect 1443 5732 2412 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 7926 5760 7932 5772
rect 7887 5732 7932 5760
rect 7926 5720 7932 5732
rect 7984 5720 7990 5772
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 13078 5760 13084 5772
rect 11756 5732 13084 5760
rect 11756 5720 11762 5732
rect 13078 5720 13084 5732
rect 13136 5760 13142 5772
rect 15304 5769 15332 5800
rect 15746 5788 15752 5800
rect 15804 5788 15810 5840
rect 17862 5788 17868 5840
rect 17920 5828 17926 5840
rect 17954 5828 17960 5840
rect 17920 5800 17960 5828
rect 17920 5788 17926 5800
rect 17954 5788 17960 5800
rect 18012 5828 18018 5840
rect 18141 5831 18199 5837
rect 18141 5828 18153 5831
rect 18012 5800 18153 5828
rect 18012 5788 18018 5800
rect 18141 5797 18153 5800
rect 18187 5828 18199 5831
rect 24118 5828 24124 5840
rect 18187 5800 24124 5828
rect 18187 5797 18199 5800
rect 18141 5791 18199 5797
rect 24118 5788 24124 5800
rect 24176 5828 24182 5840
rect 24176 5800 26556 5828
rect 24176 5788 24182 5800
rect 13725 5763 13783 5769
rect 13725 5760 13737 5763
rect 13136 5732 13737 5760
rect 13136 5720 13142 5732
rect 13725 5729 13737 5732
rect 13771 5729 13783 5763
rect 13725 5723 13783 5729
rect 15289 5763 15347 5769
rect 15289 5729 15301 5763
rect 15335 5729 15347 5763
rect 15289 5723 15347 5729
rect 15378 5720 15384 5772
rect 15436 5760 15442 5772
rect 15545 5763 15603 5769
rect 15545 5760 15557 5763
rect 15436 5732 15557 5760
rect 15436 5720 15442 5732
rect 15545 5729 15557 5732
rect 15591 5729 15603 5763
rect 22721 5763 22779 5769
rect 22721 5760 22733 5763
rect 15545 5723 15603 5729
rect 21468 5732 22733 5760
rect 1854 5652 1860 5704
rect 1912 5692 1918 5704
rect 2225 5695 2283 5701
rect 2225 5692 2237 5695
rect 1912 5664 2237 5692
rect 1912 5652 1918 5664
rect 2225 5661 2237 5664
rect 2271 5692 2283 5695
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2271 5664 2329 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 5258 5692 5264 5704
rect 5219 5664 5264 5692
rect 2317 5655 2375 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 8018 5692 8024 5704
rect 7979 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 11330 5692 11336 5704
rect 8168 5664 8213 5692
rect 11291 5664 11336 5692
rect 8168 5652 8174 5664
rect 11330 5652 11336 5664
rect 11388 5652 11394 5704
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 12805 5695 12863 5701
rect 12805 5692 12817 5695
rect 12768 5664 12817 5692
rect 12768 5652 12774 5664
rect 12805 5661 12817 5664
rect 12851 5661 12863 5695
rect 12805 5655 12863 5661
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5692 13047 5695
rect 13035 5664 13492 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 1578 5624 1584 5636
rect 1539 5596 1584 5624
rect 1578 5584 1584 5596
rect 1636 5584 1642 5636
rect 10778 5624 10784 5636
rect 10739 5596 10784 5624
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 4338 5556 4344 5568
rect 4299 5528 4344 5556
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4617 5559 4675 5565
rect 4617 5556 4629 5559
rect 4488 5528 4629 5556
rect 4488 5516 4494 5528
rect 4617 5525 4629 5528
rect 4663 5525 4675 5559
rect 7282 5556 7288 5568
rect 7243 5528 7288 5556
rect 4617 5519 4675 5525
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7558 5556 7564 5568
rect 7519 5528 7564 5556
rect 7558 5516 7564 5528
rect 7616 5516 7622 5568
rect 13464 5565 13492 5664
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 18785 5695 18843 5701
rect 18785 5692 18797 5695
rect 18380 5664 18797 5692
rect 18380 5652 18386 5664
rect 18785 5661 18797 5664
rect 18831 5661 18843 5695
rect 19794 5692 19800 5704
rect 19755 5664 19800 5692
rect 18785 5655 18843 5661
rect 19794 5652 19800 5664
rect 19852 5652 19858 5704
rect 20622 5652 20628 5704
rect 20680 5692 20686 5704
rect 21468 5701 21496 5732
rect 22721 5729 22733 5732
rect 22767 5729 22779 5763
rect 25314 5760 25320 5772
rect 25275 5732 25320 5760
rect 22721 5723 22779 5729
rect 25314 5720 25320 5732
rect 25372 5720 25378 5772
rect 26528 5769 26556 5800
rect 26513 5763 26571 5769
rect 26513 5729 26525 5763
rect 26559 5760 26571 5763
rect 27154 5760 27160 5772
rect 26559 5732 27160 5760
rect 26559 5729 26571 5732
rect 26513 5723 26571 5729
rect 27154 5720 27160 5732
rect 27212 5720 27218 5772
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 20680 5664 21373 5692
rect 20680 5652 20686 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 21361 5655 21419 5661
rect 21453 5695 21511 5701
rect 21453 5661 21465 5695
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 21468 5624 21496 5655
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 22094 5692 22100 5704
rect 21692 5664 22100 5692
rect 21692 5652 21698 5664
rect 22094 5652 22100 5664
rect 22152 5692 22158 5704
rect 22465 5695 22523 5701
rect 22465 5692 22477 5695
rect 22152 5664 22477 5692
rect 22152 5652 22158 5664
rect 22465 5661 22477 5664
rect 22511 5661 22523 5695
rect 22465 5655 22523 5661
rect 25498 5624 25504 5636
rect 20548 5596 21496 5624
rect 25459 5596 25504 5624
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13538 5556 13544 5568
rect 13495 5528 13544 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13538 5516 13544 5528
rect 13596 5516 13602 5568
rect 16482 5516 16488 5568
rect 16540 5556 16546 5568
rect 16669 5559 16727 5565
rect 16669 5556 16681 5559
rect 16540 5528 16681 5556
rect 16540 5516 16546 5528
rect 16669 5525 16681 5528
rect 16715 5525 16727 5559
rect 17770 5556 17776 5568
rect 17731 5528 17776 5556
rect 16669 5519 16727 5525
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 20438 5516 20444 5568
rect 20496 5556 20502 5568
rect 20548 5565 20576 5596
rect 25498 5584 25504 5596
rect 25556 5584 25562 5636
rect 20533 5559 20591 5565
rect 20533 5556 20545 5559
rect 20496 5528 20545 5556
rect 20496 5516 20502 5528
rect 20533 5525 20545 5528
rect 20579 5525 20591 5559
rect 20533 5519 20591 5525
rect 23566 5516 23572 5568
rect 23624 5556 23630 5568
rect 23845 5559 23903 5565
rect 23845 5556 23857 5559
rect 23624 5528 23857 5556
rect 23624 5516 23630 5528
rect 23845 5525 23857 5528
rect 23891 5525 23903 5559
rect 26694 5556 26700 5568
rect 26655 5528 26700 5556
rect 23845 5519 23903 5525
rect 26694 5516 26700 5528
rect 26752 5516 26758 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 2406 5352 2412 5364
rect 2367 5324 2412 5352
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 2958 5352 2964 5364
rect 2919 5324 2964 5352
rect 2958 5312 2964 5324
rect 3016 5312 3022 5364
rect 5077 5355 5135 5361
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5258 5352 5264 5364
rect 5123 5324 5264 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5258 5312 5264 5324
rect 5316 5312 5322 5364
rect 5442 5352 5448 5364
rect 5403 5324 5448 5352
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7926 5352 7932 5364
rect 7147 5324 7932 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 10502 5312 10508 5364
rect 10560 5352 10566 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10560 5324 10793 5352
rect 10560 5312 10566 5324
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 14458 5352 14464 5364
rect 14419 5324 14464 5352
rect 10781 5315 10839 5321
rect 14458 5312 14464 5324
rect 14516 5312 14522 5364
rect 15378 5352 15384 5364
rect 15339 5324 15384 5352
rect 15378 5312 15384 5324
rect 15436 5312 15442 5364
rect 17862 5352 17868 5364
rect 17823 5324 17868 5352
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18230 5352 18236 5364
rect 18012 5324 18236 5352
rect 18012 5312 18018 5324
rect 18230 5312 18236 5324
rect 18288 5312 18294 5364
rect 18322 5312 18328 5364
rect 18380 5352 18386 5364
rect 18601 5355 18659 5361
rect 18601 5352 18613 5355
rect 18380 5324 18613 5352
rect 18380 5312 18386 5324
rect 18601 5321 18613 5324
rect 18647 5321 18659 5355
rect 20346 5352 20352 5364
rect 20307 5324 20352 5352
rect 18601 5315 18659 5321
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 20530 5352 20536 5364
rect 20491 5324 20536 5352
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21726 5352 21732 5364
rect 21683 5324 21732 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 21726 5312 21732 5324
rect 21784 5312 21790 5364
rect 25133 5355 25191 5361
rect 25133 5321 25145 5355
rect 25179 5352 25191 5355
rect 25222 5352 25228 5364
rect 25179 5324 25228 5352
rect 25179 5321 25191 5324
rect 25133 5315 25191 5321
rect 25222 5312 25228 5324
rect 25280 5312 25286 5364
rect 26326 5312 26332 5364
rect 26384 5352 26390 5364
rect 26605 5355 26663 5361
rect 26605 5352 26617 5355
rect 26384 5324 26617 5352
rect 26384 5312 26390 5324
rect 26605 5321 26617 5324
rect 26651 5321 26663 5355
rect 27154 5352 27160 5364
rect 27115 5324 27160 5352
rect 26605 5315 26663 5321
rect 27154 5312 27160 5324
rect 27212 5312 27218 5364
rect 2038 5216 2044 5228
rect 1412 5188 2044 5216
rect 1412 5157 1440 5188
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2976 5216 3004 5312
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 11146 5284 11152 5296
rect 10735 5256 11152 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 11146 5244 11152 5256
rect 11204 5244 11210 5296
rect 16482 5244 16488 5296
rect 16540 5284 16546 5296
rect 16540 5256 16804 5284
rect 16540 5244 16546 5256
rect 9674 5216 9680 5228
rect 2976 5188 3188 5216
rect 9635 5188 9680 5216
rect 1397 5151 1455 5157
rect 1397 5117 1409 5151
rect 1443 5117 1455 5151
rect 1397 5111 1455 5117
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3053 5151 3111 5157
rect 3053 5148 3065 5151
rect 2832 5120 3065 5148
rect 2832 5108 2838 5120
rect 3053 5117 3065 5120
rect 3099 5117 3111 5151
rect 3160 5148 3188 5188
rect 9674 5176 9680 5188
rect 9732 5176 9738 5228
rect 10778 5176 10784 5228
rect 10836 5216 10842 5228
rect 11330 5216 11336 5228
rect 10836 5188 11336 5216
rect 10836 5176 10842 5188
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 13078 5216 13084 5228
rect 13039 5188 13084 5216
rect 13078 5176 13084 5188
rect 13136 5176 13142 5228
rect 15654 5176 15660 5228
rect 15712 5216 15718 5228
rect 16776 5225 16804 5256
rect 16669 5219 16727 5225
rect 16669 5216 16681 5219
rect 15712 5188 16681 5216
rect 15712 5176 15718 5188
rect 16669 5185 16681 5188
rect 16715 5185 16727 5219
rect 16669 5179 16727 5185
rect 16761 5219 16819 5225
rect 16761 5185 16773 5219
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20496 5188 21097 5216
rect 20496 5176 20502 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 3309 5151 3367 5157
rect 3309 5148 3321 5151
rect 3160 5120 3321 5148
rect 3053 5111 3111 5117
rect 3309 5117 3321 5120
rect 3355 5148 3367 5151
rect 3694 5148 3700 5160
rect 3355 5120 3700 5148
rect 3355 5117 3367 5120
rect 3309 5111 3367 5117
rect 3694 5108 3700 5120
rect 3752 5108 3758 5160
rect 7193 5151 7251 5157
rect 7193 5117 7205 5151
rect 7239 5148 7251 5151
rect 7282 5148 7288 5160
rect 7239 5120 7288 5148
rect 7239 5117 7251 5120
rect 7193 5111 7251 5117
rect 7282 5108 7288 5120
rect 7340 5108 7346 5160
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5148 15807 5151
rect 16577 5151 16635 5157
rect 16577 5148 16589 5151
rect 15795 5120 16589 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 16577 5117 16589 5120
rect 16623 5148 16635 5151
rect 17770 5148 17776 5160
rect 16623 5120 17776 5148
rect 16623 5117 16635 5120
rect 16577 5111 16635 5117
rect 17770 5108 17776 5120
rect 17828 5108 17834 5160
rect 20346 5108 20352 5160
rect 20404 5148 20410 5160
rect 20993 5151 21051 5157
rect 20993 5148 21005 5151
rect 20404 5120 21005 5148
rect 20404 5108 20410 5120
rect 20993 5117 21005 5120
rect 21039 5117 21051 5151
rect 20993 5111 21051 5117
rect 7438 5083 7496 5089
rect 7438 5080 7450 5083
rect 7208 5052 7450 5080
rect 7208 5024 7236 5052
rect 7438 5049 7450 5052
rect 7484 5080 7496 5083
rect 8110 5080 8116 5092
rect 7484 5052 8116 5080
rect 7484 5049 7496 5052
rect 7438 5043 7496 5049
rect 8110 5040 8116 5052
rect 8168 5080 8174 5092
rect 9125 5083 9183 5089
rect 9125 5080 9137 5083
rect 8168 5052 9137 5080
rect 8168 5040 8174 5052
rect 9125 5049 9137 5052
rect 9171 5049 9183 5083
rect 9125 5043 9183 5049
rect 11149 5083 11207 5089
rect 11149 5049 11161 5083
rect 11195 5080 11207 5083
rect 13348 5083 13406 5089
rect 11195 5052 11928 5080
rect 11195 5049 11207 5052
rect 11149 5043 11207 5049
rect 11900 5024 11928 5052
rect 13348 5049 13360 5083
rect 13394 5080 13406 5083
rect 13538 5080 13544 5092
rect 13394 5052 13544 5080
rect 13394 5049 13406 5052
rect 13348 5043 13406 5049
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 16117 5083 16175 5089
rect 16117 5049 16129 5083
rect 16163 5080 16175 5083
rect 16482 5080 16488 5092
rect 16163 5052 16488 5080
rect 16163 5049 16175 5052
rect 16117 5043 16175 5049
rect 16482 5040 16488 5052
rect 16540 5040 16546 5092
rect 20622 5080 20628 5092
rect 19996 5052 20628 5080
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 4433 5015 4491 5021
rect 4433 4981 4445 5015
rect 4479 5012 4491 5015
rect 4614 5012 4620 5024
rect 4479 4984 4620 5012
rect 4479 4981 4491 4984
rect 4433 4975 4491 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 7190 4972 7196 5024
rect 7248 4972 7254 5024
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 8573 5015 8631 5021
rect 8573 5012 8585 5015
rect 7708 4984 8585 5012
rect 7708 4972 7714 4984
rect 8573 4981 8585 4984
rect 8619 4981 8631 5015
rect 8573 4975 8631 4981
rect 10321 5015 10379 5021
rect 10321 4981 10333 5015
rect 10367 5012 10379 5015
rect 10778 5012 10784 5024
rect 10367 4984 10784 5012
rect 10367 4981 10379 4984
rect 10321 4975 10379 4981
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11241 5015 11299 5021
rect 11241 4981 11253 5015
rect 11287 5012 11299 5015
rect 11330 5012 11336 5024
rect 11287 4984 11336 5012
rect 11287 4981 11299 4984
rect 11241 4975 11299 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11882 5012 11888 5024
rect 11843 4984 11888 5012
rect 11882 4972 11888 4984
rect 11940 4972 11946 5024
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 12161 5015 12219 5021
rect 12161 5012 12173 5015
rect 12032 4984 12173 5012
rect 12032 4972 12038 4984
rect 12161 4981 12173 4984
rect 12207 5012 12219 5015
rect 12434 5012 12440 5024
rect 12207 4984 12440 5012
rect 12207 4981 12219 4984
rect 12161 4975 12219 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12710 5012 12716 5024
rect 12671 4984 12716 5012
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 16209 5015 16267 5021
rect 16209 4981 16221 5015
rect 16255 5012 16267 5015
rect 16298 5012 16304 5024
rect 16255 4984 16304 5012
rect 16255 4981 16267 4984
rect 16209 4975 16267 4981
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 19518 4972 19524 5024
rect 19576 5012 19582 5024
rect 19996 5021 20024 5052
rect 20622 5040 20628 5052
rect 20680 5040 20686 5092
rect 21100 5080 21128 5179
rect 25222 5148 25228 5160
rect 25183 5120 25228 5148
rect 25222 5108 25228 5120
rect 25280 5108 25286 5160
rect 21910 5080 21916 5092
rect 21100 5052 21916 5080
rect 21910 5040 21916 5052
rect 21968 5080 21974 5092
rect 22465 5083 22523 5089
rect 22465 5080 22477 5083
rect 21968 5052 22477 5080
rect 21968 5040 21974 5052
rect 22465 5049 22477 5052
rect 22511 5049 22523 5083
rect 25470 5083 25528 5089
rect 25470 5080 25482 5083
rect 22465 5043 22523 5049
rect 24872 5052 25482 5080
rect 24872 5024 24900 5052
rect 25470 5049 25482 5052
rect 25516 5049 25528 5083
rect 25470 5043 25528 5049
rect 19981 5015 20039 5021
rect 19981 5012 19993 5015
rect 19576 4984 19993 5012
rect 19576 4972 19582 4984
rect 19981 4981 19993 4984
rect 20027 4981 20039 5015
rect 19981 4975 20039 4981
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 20901 5015 20959 5021
rect 20901 5012 20913 5015
rect 20588 4984 20913 5012
rect 20588 4972 20594 4984
rect 20901 4981 20913 4984
rect 20947 4981 20959 5015
rect 22922 5012 22928 5024
rect 22883 4984 22928 5012
rect 20901 4975 20959 4981
rect 22922 4972 22928 4984
rect 22980 4972 22986 5024
rect 24765 5015 24823 5021
rect 24765 4981 24777 5015
rect 24811 5012 24823 5015
rect 24854 5012 24860 5024
rect 24811 4984 24860 5012
rect 24811 4981 24823 4984
rect 24765 4975 24823 4981
rect 24854 4972 24860 4984
rect 24912 4972 24918 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3053 4811 3111 4817
rect 3053 4808 3065 4811
rect 2832 4780 3065 4808
rect 2832 4768 2838 4780
rect 3053 4777 3065 4780
rect 3099 4808 3111 4811
rect 4154 4808 4160 4820
rect 3099 4780 4160 4808
rect 3099 4777 3111 4780
rect 3053 4771 3111 4777
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 4246 4768 4252 4820
rect 4304 4808 4310 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 4304 4780 4537 4808
rect 4304 4768 4310 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 5166 4808 5172 4820
rect 5127 4780 5172 4808
rect 4525 4771 4583 4777
rect 5166 4768 5172 4780
rect 5224 4768 5230 4820
rect 7558 4768 7564 4820
rect 7616 4808 7622 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7616 4780 7849 4808
rect 7616 4768 7622 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 10778 4808 10784 4820
rect 10739 4780 10784 4808
rect 7837 4771 7895 4777
rect 10778 4768 10784 4780
rect 10836 4768 10842 4820
rect 11241 4811 11299 4817
rect 11241 4777 11253 4811
rect 11287 4808 11299 4811
rect 11330 4808 11336 4820
rect 11287 4780 11336 4808
rect 11287 4777 11299 4780
rect 11241 4771 11299 4777
rect 11330 4768 11336 4780
rect 11388 4768 11394 4820
rect 11790 4808 11796 4820
rect 11751 4780 11796 4808
rect 11790 4768 11796 4780
rect 11848 4768 11854 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 11940 4780 12909 4808
rect 11940 4768 11946 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 12897 4771 12955 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 16209 4811 16267 4817
rect 16209 4808 16221 4811
rect 15712 4780 16221 4808
rect 15712 4768 15718 4780
rect 16209 4777 16221 4780
rect 16255 4777 16267 4811
rect 16574 4808 16580 4820
rect 16535 4780 16580 4808
rect 16209 4771 16267 4777
rect 16574 4768 16580 4780
rect 16632 4768 16638 4820
rect 19245 4811 19303 4817
rect 19245 4777 19257 4811
rect 19291 4808 19303 4811
rect 21361 4811 21419 4817
rect 21361 4808 21373 4811
rect 19291 4780 21373 4808
rect 19291 4777 19303 4780
rect 19245 4771 19303 4777
rect 21361 4777 21373 4780
rect 21407 4777 21419 4811
rect 21910 4808 21916 4820
rect 21871 4780 21916 4808
rect 21361 4771 21419 4777
rect 4430 4740 4436 4752
rect 4391 4712 4436 4740
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 7742 4740 7748 4752
rect 7703 4712 7748 4740
rect 7742 4700 7748 4712
rect 7800 4700 7806 4752
rect 11606 4700 11612 4752
rect 11664 4740 11670 4752
rect 11701 4743 11759 4749
rect 11701 4740 11713 4743
rect 11664 4712 11713 4740
rect 11664 4700 11670 4712
rect 11701 4709 11713 4712
rect 11747 4740 11759 4743
rect 12342 4740 12348 4752
rect 11747 4712 12348 4740
rect 11747 4709 11759 4712
rect 11701 4703 11759 4709
rect 12342 4700 12348 4712
rect 12400 4700 12406 4752
rect 15565 4743 15623 4749
rect 15565 4709 15577 4743
rect 15611 4740 15623 4743
rect 15746 4740 15752 4752
rect 15611 4712 15752 4740
rect 15611 4709 15623 4712
rect 15565 4703 15623 4709
rect 15746 4700 15752 4712
rect 15804 4700 15810 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 20530 4740 20536 4752
rect 19852 4712 20536 4740
rect 19852 4700 19858 4712
rect 20530 4700 20536 4712
rect 20588 4700 20594 4752
rect 20714 4700 20720 4752
rect 20772 4740 20778 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 20772 4712 21281 4740
rect 20772 4700 20778 4712
rect 21269 4709 21281 4712
rect 21315 4709 21327 4743
rect 21269 4703 21327 4709
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 2314 4632 2320 4684
rect 2372 4672 2378 4684
rect 2501 4675 2559 4681
rect 2501 4672 2513 4675
rect 2372 4644 2513 4672
rect 2372 4632 2378 4644
rect 2501 4641 2513 4644
rect 2547 4641 2559 4675
rect 13262 4672 13268 4684
rect 13223 4644 13268 4672
rect 2501 4635 2559 4641
rect 13262 4632 13268 4644
rect 13320 4632 13326 4684
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19886 4672 19892 4684
rect 19751 4644 19892 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 4617 4607 4675 4613
rect 4617 4604 4629 4607
rect 3752 4576 4629 4604
rect 3752 4564 3758 4576
rect 4617 4573 4629 4576
rect 4663 4573 4675 4607
rect 4617 4567 4675 4573
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7708 4576 7941 4604
rect 7708 4564 7714 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 8386 4604 8392 4616
rect 8347 4576 8392 4604
rect 7929 4567 7987 4573
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 11977 4607 12035 4613
rect 11977 4573 11989 4607
rect 12023 4604 12035 4607
rect 12158 4604 12164 4616
rect 12023 4576 12164 4604
rect 12023 4573 12035 4576
rect 11977 4567 12035 4573
rect 12158 4564 12164 4576
rect 12216 4604 12222 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 12216 4576 12449 4604
rect 12216 4564 12222 4576
rect 12437 4573 12449 4576
rect 12483 4604 12495 4607
rect 13538 4604 13544 4616
rect 12483 4576 13544 4604
rect 12483 4573 12495 4576
rect 12437 4567 12495 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 19426 4496 19432 4548
rect 19484 4536 19490 4548
rect 19628 4536 19656 4635
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 19978 4604 19984 4616
rect 19843 4576 19984 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 19978 4564 19984 4576
rect 20036 4564 20042 4616
rect 20622 4536 20628 4548
rect 19484 4508 20628 4536
rect 19484 4496 19490 4508
rect 20622 4496 20628 4508
rect 20680 4496 20686 4548
rect 21376 4536 21404 4771
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 25222 4768 25228 4820
rect 25280 4808 25286 4820
rect 25409 4811 25467 4817
rect 25409 4808 25421 4811
rect 25280 4780 25421 4808
rect 25280 4768 25286 4780
rect 25409 4777 25421 4780
rect 25455 4777 25467 4811
rect 25409 4771 25467 4777
rect 23566 4700 23572 4752
rect 23624 4740 23630 4752
rect 23722 4743 23780 4749
rect 23722 4740 23734 4743
rect 23624 4712 23734 4740
rect 23624 4700 23630 4712
rect 23722 4709 23734 4712
rect 23768 4709 23780 4743
rect 23722 4703 23780 4709
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 22094 4672 22100 4684
rect 21968 4644 22100 4672
rect 21968 4632 21974 4644
rect 22094 4632 22100 4644
rect 22152 4672 22158 4684
rect 22922 4672 22928 4684
rect 22152 4644 22928 4672
rect 22152 4632 22158 4644
rect 22922 4632 22928 4644
rect 22980 4672 22986 4684
rect 23477 4675 23535 4681
rect 23477 4672 23489 4675
rect 22980 4644 23489 4672
rect 22980 4632 22986 4644
rect 23477 4641 23489 4644
rect 23523 4672 23535 4675
rect 24302 4672 24308 4684
rect 23523 4644 24308 4672
rect 23523 4641 23535 4644
rect 23477 4635 23535 4641
rect 24302 4632 24308 4644
rect 24360 4632 24366 4684
rect 26510 4672 26516 4684
rect 26471 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4632 26574 4684
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4604 21603 4607
rect 21634 4604 21640 4616
rect 21591 4576 21640 4604
rect 21591 4573 21603 4576
rect 21545 4567 21603 4573
rect 21634 4564 21640 4576
rect 21692 4564 21698 4616
rect 22094 4536 22100 4548
rect 21376 4508 22100 4536
rect 22094 4496 22100 4508
rect 22152 4496 22158 4548
rect 24854 4536 24860 4548
rect 24815 4508 24860 4536
rect 24854 4496 24860 4508
rect 24912 4496 24918 4548
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 1670 4428 1676 4480
rect 1728 4468 1734 4480
rect 2685 4471 2743 4477
rect 2685 4468 2697 4471
rect 1728 4440 2697 4468
rect 1728 4428 1734 4440
rect 2685 4437 2697 4440
rect 2731 4437 2743 4471
rect 4062 4468 4068 4480
rect 4023 4440 4068 4468
rect 2685 4431 2743 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 6914 4468 6920 4480
rect 6875 4440 6920 4468
rect 6914 4428 6920 4440
rect 6972 4428 6978 4480
rect 7190 4468 7196 4480
rect 7151 4440 7196 4468
rect 7190 4428 7196 4440
rect 7248 4428 7254 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7377 4471 7435 4477
rect 7377 4468 7389 4471
rect 7340 4440 7389 4468
rect 7340 4428 7346 4440
rect 7377 4437 7389 4440
rect 7423 4437 7435 4471
rect 20898 4468 20904 4480
rect 20859 4440 20904 4468
rect 7377 4431 7435 4437
rect 20898 4428 20904 4440
rect 20956 4428 20962 4480
rect 26697 4471 26755 4477
rect 26697 4437 26709 4471
rect 26743 4468 26755 4471
rect 26786 4468 26792 4480
rect 26743 4440 26792 4468
rect 26743 4437 26755 4440
rect 26697 4431 26755 4437
rect 26786 4428 26792 4440
rect 26844 4428 26850 4480
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 4065 4267 4123 4273
rect 4065 4264 4077 4267
rect 3752 4236 4077 4264
rect 3752 4224 3758 4236
rect 4065 4233 4077 4236
rect 4111 4233 4123 4267
rect 4065 4227 4123 4233
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4433 4267 4491 4273
rect 4433 4264 4445 4267
rect 4304 4236 4445 4264
rect 4304 4224 4310 4236
rect 4433 4233 4445 4236
rect 4479 4233 4491 4267
rect 4433 4227 4491 4233
rect 7558 4224 7564 4276
rect 7616 4264 7622 4276
rect 7929 4267 7987 4273
rect 7929 4264 7941 4267
rect 7616 4236 7941 4264
rect 7616 4224 7622 4236
rect 7929 4233 7941 4236
rect 7975 4233 7987 4267
rect 7929 4227 7987 4233
rect 11425 4267 11483 4273
rect 11425 4233 11437 4267
rect 11471 4264 11483 4267
rect 11790 4264 11796 4276
rect 11471 4236 11796 4264
rect 11471 4233 11483 4236
rect 11425 4227 11483 4233
rect 11790 4224 11796 4236
rect 11848 4224 11854 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13633 4267 13691 4273
rect 13633 4264 13645 4267
rect 13596 4236 13645 4264
rect 13596 4224 13602 4236
rect 13633 4233 13645 4236
rect 13679 4233 13691 4267
rect 13633 4227 13691 4233
rect 15933 4267 15991 4273
rect 15933 4233 15945 4267
rect 15979 4264 15991 4267
rect 16298 4264 16304 4276
rect 15979 4236 16304 4264
rect 15979 4233 15991 4236
rect 15933 4227 15991 4233
rect 16298 4224 16304 4236
rect 16356 4224 16362 4276
rect 19061 4267 19119 4273
rect 19061 4233 19073 4267
rect 19107 4264 19119 4267
rect 19978 4264 19984 4276
rect 19107 4236 19984 4264
rect 19107 4233 19119 4236
rect 19061 4227 19119 4233
rect 19978 4224 19984 4236
rect 20036 4224 20042 4276
rect 23566 4224 23572 4276
rect 23624 4264 23630 4276
rect 23845 4267 23903 4273
rect 23845 4264 23857 4267
rect 23624 4236 23857 4264
rect 23624 4224 23630 4236
rect 23845 4233 23857 4236
rect 23891 4233 23903 4267
rect 24302 4264 24308 4276
rect 24215 4236 24308 4264
rect 23845 4227 23903 4233
rect 24302 4224 24308 4236
rect 24360 4264 24366 4276
rect 25222 4264 25228 4276
rect 24360 4236 25228 4264
rect 24360 4224 24366 4236
rect 25222 4224 25228 4236
rect 25280 4224 25286 4276
rect 26510 4224 26516 4276
rect 26568 4264 26574 4276
rect 26973 4267 27031 4273
rect 26973 4264 26985 4267
rect 26568 4236 26985 4264
rect 26568 4224 26574 4236
rect 26973 4233 26985 4236
rect 27019 4233 27031 4267
rect 26973 4227 27031 4233
rect 7742 4196 7748 4208
rect 6932 4168 7748 4196
rect 2314 4128 2320 4140
rect 2275 4100 2320 4128
rect 2314 4088 2320 4100
rect 2372 4128 2378 4140
rect 3786 4128 3792 4140
rect 2372 4100 3792 4128
rect 2372 4088 2378 4100
rect 3786 4088 3792 4100
rect 3844 4088 3850 4140
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4488 4100 4813 4128
rect 4488 4088 4494 4100
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 6932 4128 6960 4168
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 12989 4199 13047 4205
rect 12989 4165 13001 4199
rect 13035 4196 13047 4199
rect 13354 4196 13360 4208
rect 13035 4168 13360 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 13354 4156 13360 4168
rect 13412 4156 13418 4208
rect 6687 4100 6960 4128
rect 16316 4128 16344 4224
rect 19426 4196 19432 4208
rect 19352 4168 19432 4196
rect 16853 4131 16911 4137
rect 16853 4128 16865 4131
rect 16316 4100 16865 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 16853 4097 16865 4100
rect 16899 4097 16911 4131
rect 16853 4091 16911 4097
rect 16945 4131 17003 4137
rect 16945 4097 16957 4131
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 18693 4131 18751 4137
rect 18693 4097 18705 4131
rect 18739 4128 18751 4131
rect 19352 4128 19380 4168
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 19702 4128 19708 4140
rect 18739 4100 19380 4128
rect 19663 4100 19708 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4029 1455 4063
rect 1397 4023 1455 4029
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 3145 4063 3203 4069
rect 3145 4060 3157 4063
rect 2547 4032 3157 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 3145 4029 3157 4032
rect 3191 4060 3203 4063
rect 4890 4060 4896 4072
rect 3191 4032 4896 4060
rect 3191 4029 3203 4032
rect 3145 4023 3203 4029
rect 1412 3992 1440 4023
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6914 4020 6920 4032
rect 6972 4020 6978 4072
rect 7834 4020 7840 4072
rect 7892 4060 7898 4072
rect 8665 4063 8723 4069
rect 8665 4060 8677 4063
rect 7892 4032 8677 4060
rect 7892 4020 7898 4032
rect 8665 4029 8677 4032
rect 8711 4060 8723 4063
rect 9401 4063 9459 4069
rect 9401 4060 9413 4063
rect 8711 4032 9413 4060
rect 8711 4029 8723 4032
rect 8665 4023 8723 4029
rect 9401 4029 9413 4032
rect 9447 4029 9459 4063
rect 9401 4023 9459 4029
rect 16574 4020 16580 4072
rect 16632 4060 16638 4072
rect 16761 4063 16819 4069
rect 16761 4060 16773 4063
rect 16632 4032 16773 4060
rect 16632 4020 16638 4032
rect 16761 4029 16773 4032
rect 16807 4029 16819 4063
rect 16761 4023 16819 4029
rect 2038 3992 2044 4004
rect 1412 3964 2044 3992
rect 2038 3952 2044 3964
rect 2096 3952 2102 4004
rect 7101 3995 7159 4001
rect 7101 3961 7113 3995
rect 7147 3992 7159 3995
rect 7742 3992 7748 4004
rect 7147 3964 7748 3992
rect 7147 3961 7159 3964
rect 7101 3955 7159 3961
rect 7742 3952 7748 3964
rect 7800 3952 7806 4004
rect 8941 3995 8999 4001
rect 8941 3961 8953 3995
rect 8987 3992 8999 3995
rect 10594 3992 10600 4004
rect 8987 3964 10600 3992
rect 8987 3961 8999 3964
rect 8941 3955 8999 3961
rect 10594 3952 10600 3964
rect 10652 3952 10658 4004
rect 16301 3995 16359 4001
rect 16301 3961 16313 3995
rect 16347 3992 16359 3995
rect 16960 3992 16988 4091
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20438 4128 20444 4140
rect 20351 4100 20444 4128
rect 20438 4088 20444 4100
rect 20496 4088 20502 4140
rect 20993 4131 21051 4137
rect 20993 4097 21005 4131
rect 21039 4128 21051 4131
rect 21358 4128 21364 4140
rect 21039 4100 21364 4128
rect 21039 4097 21051 4100
rect 20993 4091 21051 4097
rect 21358 4088 21364 4100
rect 21416 4128 21422 4140
rect 21913 4131 21971 4137
rect 21913 4128 21925 4131
rect 21416 4100 21925 4128
rect 21416 4088 21422 4100
rect 21913 4097 21925 4100
rect 21959 4097 21971 4131
rect 21913 4091 21971 4097
rect 22002 4088 22008 4140
rect 22060 4128 22066 4140
rect 22060 4100 22105 4128
rect 22060 4088 22066 4100
rect 19429 4063 19487 4069
rect 19429 4029 19441 4063
rect 19475 4060 19487 4063
rect 20456 4060 20484 4088
rect 19475 4032 20484 4060
rect 19475 4029 19487 4032
rect 19429 4023 19487 4029
rect 20806 4020 20812 4072
rect 20864 4060 20870 4072
rect 21269 4063 21327 4069
rect 21269 4060 21281 4063
rect 20864 4032 21281 4060
rect 20864 4020 20870 4032
rect 21269 4029 21281 4032
rect 21315 4060 21327 4063
rect 21818 4060 21824 4072
rect 21315 4032 21824 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 22094 4020 22100 4072
rect 22152 4060 22158 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22152 4032 22477 4060
rect 22152 4020 22158 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 26421 4063 26479 4069
rect 26421 4060 26433 4063
rect 22465 4023 22523 4029
rect 26344 4032 26433 4060
rect 17678 3992 17684 4004
rect 16347 3964 17684 3992
rect 16347 3961 16359 3964
rect 16301 3955 16359 3961
rect 17678 3952 17684 3964
rect 17736 3952 17742 4004
rect 19702 3952 19708 4004
rect 19760 3992 19766 4004
rect 20257 3995 20315 4001
rect 20257 3992 20269 3995
rect 19760 3964 20269 3992
rect 19760 3952 19766 3964
rect 20257 3961 20269 3964
rect 20303 3992 20315 3995
rect 20438 3992 20444 4004
rect 20303 3964 20444 3992
rect 20303 3961 20315 3964
rect 20257 3955 20315 3961
rect 20438 3952 20444 3964
rect 20496 3952 20502 4004
rect 20622 3952 20628 4004
rect 20680 3992 20686 4004
rect 20680 3964 21496 3992
rect 20680 3952 20686 3964
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 2406 3884 2412 3936
rect 2464 3924 2470 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2464 3896 2697 3924
rect 2464 3884 2470 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 7558 3924 7564 3936
rect 7519 3896 7564 3924
rect 2685 3887 2743 3893
rect 7558 3884 7564 3896
rect 7616 3884 7622 3936
rect 10778 3884 10784 3936
rect 10836 3924 10842 3936
rect 11606 3924 11612 3936
rect 10836 3896 11612 3924
rect 10836 3884 10842 3896
rect 11606 3884 11612 3896
rect 11664 3924 11670 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11664 3896 11713 3924
rect 11664 3884 11670 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 12158 3924 12164 3936
rect 12119 3896 12164 3924
rect 11701 3887 11759 3893
rect 12158 3884 12164 3896
rect 12216 3884 12222 3936
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 13262 3924 13268 3936
rect 12308 3896 13268 3924
rect 12308 3884 12314 3896
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 16390 3924 16396 3936
rect 16351 3896 16396 3924
rect 16390 3884 16396 3896
rect 16448 3884 16454 3936
rect 19886 3924 19892 3936
rect 19847 3896 19892 3924
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 21468 3933 21496 3964
rect 26344 3936 26372 4032
rect 26421 4029 26433 4032
rect 26467 4029 26479 4063
rect 27522 4060 27528 4072
rect 27483 4032 27528 4060
rect 26421 4023 26479 4029
rect 27522 4020 27528 4032
rect 27580 4060 27586 4072
rect 28077 4063 28135 4069
rect 28077 4060 28089 4063
rect 27580 4032 28089 4060
rect 27580 4020 27586 4032
rect 28077 4029 28089 4032
rect 28123 4029 28135 4063
rect 28077 4023 28135 4029
rect 21453 3927 21511 3933
rect 20404 3896 20449 3924
rect 20404 3884 20410 3896
rect 21453 3893 21465 3927
rect 21499 3893 21511 3927
rect 26326 3924 26332 3936
rect 26287 3896 26332 3924
rect 21453 3887 21511 3893
rect 26326 3884 26332 3896
rect 26384 3884 26390 3936
rect 26602 3924 26608 3936
rect 26563 3896 26608 3924
rect 26602 3884 26608 3896
rect 26660 3884 26666 3936
rect 27706 3924 27712 3936
rect 27667 3896 27712 3924
rect 27706 3884 27712 3896
rect 27764 3884 27770 3936
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 2498 3680 2504 3732
rect 2556 3680 2562 3732
rect 3142 3720 3148 3732
rect 3103 3692 3148 3720
rect 3142 3680 3148 3692
rect 3200 3680 3206 3732
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4249 3723 4307 3729
rect 4249 3720 4261 3723
rect 4212 3692 4261 3720
rect 4212 3680 4218 3692
rect 4249 3689 4261 3692
rect 4295 3689 4307 3723
rect 4249 3683 4307 3689
rect 2516 3652 2544 3680
rect 1412 3624 2544 3652
rect 1412 3593 1440 3624
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 2501 3587 2559 3593
rect 2501 3553 2513 3587
rect 2547 3584 2559 3587
rect 2682 3584 2688 3596
rect 2547 3556 2688 3584
rect 2547 3553 2559 3556
rect 2501 3547 2559 3553
rect 2682 3544 2688 3556
rect 2740 3584 2746 3596
rect 2774 3584 2780 3596
rect 2740 3556 2780 3584
rect 2740 3544 2746 3556
rect 2774 3544 2780 3556
rect 2832 3544 2838 3596
rect 4264 3584 4292 3683
rect 7006 3680 7012 3732
rect 7064 3720 7070 3732
rect 7745 3723 7803 3729
rect 7745 3720 7757 3723
rect 7064 3692 7757 3720
rect 7064 3680 7070 3692
rect 7745 3689 7757 3692
rect 7791 3720 7803 3723
rect 8018 3720 8024 3732
rect 7791 3692 8024 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 12158 3680 12164 3732
rect 12216 3720 12222 3732
rect 12529 3723 12587 3729
rect 12529 3720 12541 3723
rect 12216 3692 12541 3720
rect 12216 3680 12222 3692
rect 12529 3689 12541 3692
rect 12575 3689 12587 3723
rect 17678 3720 17684 3732
rect 17639 3692 17684 3720
rect 12529 3683 12587 3689
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 19337 3723 19395 3729
rect 19337 3689 19349 3723
rect 19383 3720 19395 3723
rect 19886 3720 19892 3732
rect 19383 3692 19892 3720
rect 19383 3689 19395 3692
rect 19337 3683 19395 3689
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21634 3720 21640 3732
rect 21595 3692 21640 3720
rect 21634 3680 21640 3692
rect 21692 3680 21698 3732
rect 4614 3612 4620 3664
rect 4672 3661 4678 3664
rect 4672 3655 4736 3661
rect 4672 3621 4690 3655
rect 4724 3621 4736 3655
rect 11698 3652 11704 3664
rect 4672 3615 4736 3621
rect 11164 3624 11704 3652
rect 4672 3612 4678 3615
rect 4433 3587 4491 3593
rect 4433 3584 4445 3587
rect 4264 3556 4445 3584
rect 4433 3553 4445 3556
rect 4479 3553 4491 3587
rect 9858 3584 9864 3596
rect 9819 3556 9864 3584
rect 4433 3547 4491 3553
rect 9858 3544 9864 3556
rect 9916 3584 9922 3596
rect 11164 3593 11192 3624
rect 11698 3612 11704 3624
rect 11756 3612 11762 3664
rect 20254 3652 20260 3664
rect 19536 3624 20260 3652
rect 11422 3593 11428 3596
rect 10597 3587 10655 3593
rect 10597 3584 10609 3587
rect 9916 3556 10609 3584
rect 9916 3544 9922 3556
rect 10597 3553 10609 3556
rect 10643 3553 10655 3587
rect 10597 3547 10655 3553
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3553 11207 3587
rect 11416 3584 11428 3593
rect 11383 3556 11428 3584
rect 11149 3547 11207 3553
rect 11416 3547 11428 3556
rect 11422 3544 11428 3547
rect 11480 3544 11486 3596
rect 15746 3544 15752 3596
rect 15804 3584 15810 3596
rect 16298 3584 16304 3596
rect 15804 3556 16304 3584
rect 15804 3544 15810 3556
rect 16298 3544 16304 3556
rect 16356 3544 16362 3596
rect 16574 3593 16580 3596
rect 16568 3584 16580 3593
rect 16535 3556 16580 3584
rect 16568 3547 16580 3556
rect 16574 3544 16580 3547
rect 16632 3544 16638 3596
rect 19536 3593 19564 3624
rect 20254 3612 20260 3624
rect 20312 3612 20318 3664
rect 19521 3587 19579 3593
rect 19521 3553 19533 3587
rect 19567 3553 19579 3587
rect 19521 3547 19579 3553
rect 20070 3544 20076 3596
rect 20128 3584 20134 3596
rect 20806 3584 20812 3596
rect 20128 3556 20812 3584
rect 20128 3544 20134 3556
rect 20806 3544 20812 3556
rect 20864 3584 20870 3596
rect 20901 3587 20959 3593
rect 20901 3584 20913 3587
rect 20864 3556 20913 3584
rect 20864 3544 20870 3556
rect 20901 3553 20913 3556
rect 20947 3553 20959 3587
rect 23474 3584 23480 3596
rect 23435 3556 23480 3584
rect 20901 3547 20959 3553
rect 23474 3544 23480 3556
rect 23532 3544 23538 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7466 3516 7472 3528
rect 6604 3488 7472 3516
rect 6604 3476 6610 3488
rect 7466 3476 7472 3488
rect 7524 3516 7530 3528
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7524 3488 7849 3516
rect 7524 3476 7530 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 10134 3516 10140 3528
rect 10095 3488 10140 3516
rect 7929 3479 7987 3485
rect 7190 3448 7196 3460
rect 6288 3420 7196 3448
rect 6288 3392 6316 3420
rect 7190 3408 7196 3420
rect 7248 3448 7254 3460
rect 7944 3448 7972 3479
rect 10134 3476 10140 3488
rect 10192 3476 10198 3528
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3516 19855 3519
rect 20622 3516 20628 3528
rect 19843 3488 20628 3516
rect 19843 3485 19855 3488
rect 19797 3479 19855 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 21177 3519 21235 3525
rect 21177 3485 21189 3519
rect 21223 3516 21235 3519
rect 22002 3516 22008 3528
rect 21223 3488 22008 3516
rect 21223 3485 21235 3488
rect 21177 3479 21235 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 8386 3448 8392 3460
rect 7248 3420 8392 3448
rect 7248 3408 7254 3420
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 1578 3380 1584 3392
rect 1539 3352 1584 3380
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 2682 3380 2688 3392
rect 2643 3352 2688 3380
rect 2682 3340 2688 3352
rect 2740 3340 2746 3392
rect 5813 3383 5871 3389
rect 5813 3349 5825 3383
rect 5859 3380 5871 3383
rect 6270 3380 6276 3392
rect 5859 3352 6276 3380
rect 5859 3349 5871 3352
rect 5813 3343 5871 3349
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 7098 3380 7104 3392
rect 7059 3352 7104 3380
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7374 3380 7380 3392
rect 7335 3352 7380 3380
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 20254 3380 20260 3392
rect 20215 3352 20260 3380
rect 20254 3340 20260 3352
rect 20312 3340 20318 3392
rect 23658 3380 23664 3392
rect 23619 3352 23664 3380
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 26694 3380 26700 3392
rect 26655 3352 26700 3380
rect 26694 3340 26700 3352
rect 26752 3340 26758 3392
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2409 3179 2467 3185
rect 2409 3145 2421 3179
rect 2455 3176 2467 3179
rect 2498 3176 2504 3188
rect 2455 3148 2504 3176
rect 2455 3145 2467 3148
rect 2409 3139 2467 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 3786 3176 3792 3188
rect 2832 3148 2877 3176
rect 3747 3148 3792 3176
rect 2832 3136 2838 3148
rect 3786 3136 3792 3148
rect 3844 3136 3850 3188
rect 6914 3136 6920 3188
rect 6972 3176 6978 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 6972 3148 7021 3176
rect 6972 3136 6978 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 10781 3179 10839 3185
rect 10781 3176 10793 3179
rect 7009 3139 7067 3145
rect 7576 3148 10793 3176
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 5626 3108 5632 3120
rect 4387 3080 5632 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 5626 3068 5632 3080
rect 5684 3108 5690 3120
rect 5721 3111 5779 3117
rect 5721 3108 5733 3111
rect 5684 3080 5733 3108
rect 5684 3068 5690 3080
rect 5721 3077 5733 3080
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 2038 3040 2044 3052
rect 1412 3012 2044 3040
rect 1412 2981 1440 3012
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4672 3012 4905 3040
rect 4672 3000 4678 3012
rect 4893 3009 4905 3012
rect 4939 3040 4951 3043
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4939 3012 5365 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 6546 3040 6552 3052
rect 5592 3012 6552 3040
rect 5592 3000 5598 3012
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7576 3049 7604 3148
rect 10781 3145 10793 3148
rect 10827 3176 10839 3179
rect 11333 3179 11391 3185
rect 11333 3176 11345 3179
rect 10827 3148 11345 3176
rect 10827 3145 10839 3148
rect 10781 3139 10839 3145
rect 11333 3145 11345 3148
rect 11379 3176 11391 3179
rect 11422 3176 11428 3188
rect 11379 3148 11428 3176
rect 11379 3145 11391 3148
rect 11333 3139 11391 3145
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 11698 3176 11704 3188
rect 11659 3148 11704 3176
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 15344 3148 15485 3176
rect 15344 3136 15350 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 16574 3176 16580 3188
rect 16439 3148 16580 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 19058 3176 19064 3188
rect 19019 3148 19064 3176
rect 19058 3136 19064 3148
rect 19116 3136 19122 3188
rect 19334 3176 19340 3188
rect 19295 3148 19340 3176
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 19521 3179 19579 3185
rect 19521 3145 19533 3179
rect 19567 3176 19579 3179
rect 20254 3176 20260 3188
rect 19567 3148 20260 3176
rect 19567 3145 19579 3148
rect 19521 3139 19579 3145
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 22094 3136 22100 3188
rect 22152 3176 22158 3188
rect 22465 3179 22523 3185
rect 22465 3176 22477 3179
rect 22152 3148 22477 3176
rect 22152 3136 22158 3148
rect 22465 3145 22477 3148
rect 22511 3145 22523 3179
rect 24762 3176 24768 3188
rect 24723 3148 24768 3176
rect 22465 3139 22523 3145
rect 24762 3136 24768 3148
rect 24820 3136 24826 3188
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 27341 3179 27399 3185
rect 27341 3176 27353 3179
rect 26568 3148 27353 3176
rect 26568 3136 26574 3148
rect 27341 3145 27353 3148
rect 27387 3145 27399 3179
rect 27341 3139 27399 3145
rect 8018 3108 8024 3120
rect 7979 3080 8024 3108
rect 8018 3068 8024 3080
rect 8076 3068 8082 3120
rect 8386 3108 8392 3120
rect 8347 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3068 8450 3120
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16669 3111 16727 3117
rect 16669 3108 16681 3111
rect 16356 3080 16681 3108
rect 16356 3068 16362 3080
rect 16669 3077 16681 3080
rect 16715 3108 16727 3111
rect 17678 3108 17684 3120
rect 16715 3080 17684 3108
rect 16715 3077 16727 3080
rect 16669 3071 16727 3077
rect 17678 3068 17684 3080
rect 17736 3068 17742 3120
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7156 3012 7573 3040
rect 7156 3000 7162 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 20070 3040 20076 3052
rect 20031 3012 20076 3040
rect 7561 3003 7619 3009
rect 20070 3000 20076 3012
rect 20128 3040 20134 3052
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 20128 3012 20545 3040
rect 20128 3000 20134 3012
rect 20533 3009 20545 3012
rect 20579 3040 20591 3043
rect 20901 3043 20959 3049
rect 20901 3040 20913 3043
rect 20579 3012 20913 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 20901 3009 20913 3012
rect 20947 3040 20959 3043
rect 20947 3012 21220 3040
rect 20947 3009 20959 3012
rect 20901 3003 20959 3009
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 3053 2975 3111 2981
rect 3053 2941 3065 2975
rect 3099 2972 3111 2975
rect 3142 2972 3148 2984
rect 3099 2944 3148 2972
rect 3099 2941 3111 2944
rect 3053 2935 3111 2941
rect 3142 2932 3148 2944
rect 3200 2932 3206 2984
rect 3786 2932 3792 2984
rect 3844 2972 3850 2984
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 3844 2944 4721 2972
rect 3844 2932 3850 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 7282 2932 7288 2984
rect 7340 2972 7346 2984
rect 7377 2975 7435 2981
rect 7377 2972 7389 2975
rect 7340 2944 7389 2972
rect 7340 2932 7346 2944
rect 7377 2941 7389 2944
rect 7423 2972 7435 2975
rect 8757 2975 8815 2981
rect 8757 2972 8769 2975
rect 7423 2944 8769 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 8757 2941 8769 2944
rect 8803 2941 8815 2975
rect 8757 2935 8815 2941
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2972 9459 2975
rect 9490 2972 9496 2984
rect 9447 2944 9496 2972
rect 9447 2941 9459 2944
rect 9401 2935 9459 2941
rect 9490 2932 9496 2944
rect 9548 2972 9554 2984
rect 11698 2972 11704 2984
rect 9548 2944 11704 2972
rect 9548 2932 9554 2944
rect 11698 2932 11704 2944
rect 11756 2932 11762 2984
rect 14737 2975 14795 2981
rect 14737 2941 14749 2975
rect 14783 2972 14795 2975
rect 15286 2972 15292 2984
rect 14783 2944 15292 2972
rect 14783 2941 14795 2944
rect 14737 2935 14795 2941
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 17865 2975 17923 2981
rect 17865 2941 17877 2975
rect 17911 2972 17923 2975
rect 18230 2972 18236 2984
rect 17911 2944 18236 2972
rect 17911 2941 17923 2944
rect 17865 2935 17923 2941
rect 18230 2932 18236 2944
rect 18288 2932 18294 2984
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19889 2975 19947 2981
rect 19889 2972 19901 2975
rect 19116 2944 19901 2972
rect 19116 2932 19122 2944
rect 19889 2941 19901 2944
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 21085 2975 21143 2981
rect 21085 2941 21097 2975
rect 21131 2941 21143 2975
rect 21192 2972 21220 3012
rect 21341 2975 21399 2981
rect 21341 2972 21353 2975
rect 21192 2944 21353 2972
rect 21085 2935 21143 2941
rect 21341 2941 21353 2944
rect 21387 2941 21399 2975
rect 21341 2935 21399 2941
rect 24029 2975 24087 2981
rect 24029 2941 24041 2975
rect 24075 2972 24087 2975
rect 24762 2972 24768 2984
rect 24075 2944 24768 2972
rect 24075 2941 24087 2944
rect 24029 2935 24087 2941
rect 2038 2864 2044 2916
rect 2096 2904 2102 2916
rect 2590 2904 2596 2916
rect 2096 2876 2596 2904
rect 2096 2864 2102 2876
rect 2590 2864 2596 2876
rect 2648 2864 2654 2916
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2904 3387 2907
rect 4890 2904 4896 2916
rect 3375 2876 4896 2904
rect 3375 2873 3387 2876
rect 3329 2867 3387 2873
rect 4890 2864 4896 2876
rect 4948 2864 4954 2916
rect 6273 2907 6331 2913
rect 6273 2873 6285 2907
rect 6319 2904 6331 2907
rect 6914 2904 6920 2916
rect 6319 2876 6920 2904
rect 6319 2873 6331 2876
rect 6273 2867 6331 2873
rect 6914 2864 6920 2876
rect 6972 2904 6978 2916
rect 7469 2907 7527 2913
rect 7469 2904 7481 2907
rect 6972 2876 7481 2904
rect 6972 2864 6978 2876
rect 7469 2873 7481 2876
rect 7515 2873 7527 2907
rect 7469 2867 7527 2873
rect 7558 2864 7564 2916
rect 7616 2904 7622 2916
rect 9217 2907 9275 2913
rect 9217 2904 9229 2907
rect 7616 2876 9229 2904
rect 7616 2864 7622 2876
rect 9217 2873 9229 2876
rect 9263 2904 9275 2907
rect 9646 2907 9704 2913
rect 9646 2904 9658 2907
rect 9263 2876 9658 2904
rect 9263 2873 9275 2876
rect 9217 2867 9275 2873
rect 9646 2873 9658 2876
rect 9692 2873 9704 2907
rect 15010 2904 15016 2916
rect 14971 2876 15016 2904
rect 9646 2867 9704 2873
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 18509 2907 18567 2913
rect 18509 2873 18521 2907
rect 18555 2904 18567 2907
rect 19150 2904 19156 2916
rect 18555 2876 19156 2904
rect 18555 2873 18567 2876
rect 18509 2867 18567 2873
rect 19150 2864 19156 2876
rect 19208 2864 19214 2916
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19978 2904 19984 2916
rect 19392 2876 19984 2904
rect 19392 2864 19398 2876
rect 19978 2864 19984 2876
rect 20036 2864 20042 2916
rect 21100 2904 21128 2935
rect 24762 2932 24768 2944
rect 24820 2932 24826 2984
rect 26421 2975 26479 2981
rect 26421 2941 26433 2975
rect 26467 2972 26479 2975
rect 26878 2972 26884 2984
rect 26467 2944 26884 2972
rect 26467 2941 26479 2944
rect 26421 2935 26479 2941
rect 26878 2932 26884 2944
rect 26936 2972 26942 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26936 2944 26985 2972
rect 26936 2932 26942 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 27522 2972 27528 2984
rect 27483 2944 27528 2972
rect 26973 2935 27031 2941
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 28077 2975 28135 2981
rect 28077 2972 28089 2975
rect 27580 2944 28089 2972
rect 27580 2932 27586 2944
rect 28077 2941 28089 2944
rect 28123 2941 28135 2975
rect 28077 2935 28135 2941
rect 21450 2904 21456 2916
rect 21100 2876 21456 2904
rect 21450 2864 21456 2876
rect 21508 2904 21514 2916
rect 21910 2904 21916 2916
rect 21508 2876 21916 2904
rect 21508 2864 21514 2876
rect 21910 2864 21916 2876
rect 21968 2864 21974 2916
rect 24305 2907 24363 2913
rect 24305 2873 24317 2907
rect 24351 2904 24363 2907
rect 24854 2904 24860 2916
rect 24351 2876 24860 2904
rect 24351 2873 24363 2876
rect 24305 2867 24363 2873
rect 24854 2864 24860 2876
rect 24912 2864 24918 2916
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1452 2808 1593 2836
rect 1452 2796 1458 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 4249 2839 4307 2845
rect 4249 2805 4261 2839
rect 4295 2836 4307 2839
rect 4798 2836 4804 2848
rect 4295 2808 4804 2836
rect 4295 2805 4307 2808
rect 4249 2799 4307 2805
rect 4798 2796 4804 2808
rect 4856 2796 4862 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 23937 2839 23995 2845
rect 23937 2836 23949 2839
rect 23532 2808 23949 2836
rect 23532 2796 23538 2808
rect 23937 2805 23949 2808
rect 23983 2836 23995 2839
rect 25314 2836 25320 2848
rect 23983 2808 25320 2836
rect 23983 2805 23995 2808
rect 23937 2799 23995 2805
rect 25314 2796 25320 2808
rect 25372 2796 25378 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 27706 2836 27712 2848
rect 27667 2808 27712 2836
rect 27706 2796 27712 2808
rect 27764 2796 27770 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 3513 2635 3571 2641
rect 3513 2632 3525 2635
rect 2700 2604 3525 2632
rect 2700 2505 2728 2604
rect 3513 2601 3525 2604
rect 3559 2632 3571 2635
rect 4062 2632 4068 2644
rect 3559 2604 4068 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4614 2632 4620 2644
rect 4575 2604 4620 2632
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 5626 2632 5632 2644
rect 5587 2604 5632 2632
rect 5626 2592 5632 2604
rect 5684 2592 5690 2644
rect 6270 2632 6276 2644
rect 6231 2604 6276 2632
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 7009 2635 7067 2641
rect 7009 2632 7021 2635
rect 6972 2604 7021 2632
rect 6972 2592 6978 2604
rect 7009 2601 7021 2604
rect 7055 2601 7067 2635
rect 7374 2632 7380 2644
rect 7335 2604 7380 2632
rect 7009 2595 7067 2601
rect 7374 2592 7380 2604
rect 7432 2632 7438 2644
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 7432 2604 8401 2632
rect 7432 2592 7438 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 8389 2595 8447 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 17678 2632 17684 2644
rect 17639 2604 17684 2632
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 17770 2592 17776 2644
rect 17828 2632 17834 2644
rect 18049 2635 18107 2641
rect 18049 2632 18061 2635
rect 17828 2604 18061 2632
rect 17828 2592 17834 2604
rect 18049 2601 18061 2604
rect 18095 2601 18107 2635
rect 18049 2595 18107 2601
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 20070 2632 20076 2644
rect 19751 2604 20076 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 2958 2564 2964 2576
rect 2919 2536 2964 2564
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 7558 2564 7564 2576
rect 7392 2536 7564 2564
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 2685 2499 2743 2505
rect 2685 2465 2697 2499
rect 2731 2465 2743 2499
rect 2685 2459 2743 2465
rect 5077 2499 5135 2505
rect 5077 2465 5089 2499
rect 5123 2496 5135 2499
rect 5534 2496 5540 2508
rect 5123 2468 5540 2496
rect 5123 2465 5135 2468
rect 5077 2459 5135 2465
rect 1412 2428 1440 2459
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7392 2496 7420 2536
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 11514 2564 11520 2576
rect 11256 2536 11520 2564
rect 6779 2468 7420 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 2041 2431 2099 2437
rect 2041 2428 2053 2431
rect 1412 2400 2053 2428
rect 2041 2397 2053 2400
rect 2087 2428 2099 2431
rect 4338 2428 4344 2440
rect 2087 2400 4344 2428
rect 2087 2397 2099 2400
rect 2041 2391 2099 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6270 2428 6276 2440
rect 5859 2400 6276 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 6270 2388 6276 2400
rect 6328 2388 6334 2440
rect 7392 2428 7420 2468
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7515 2468 8033 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7392 2400 7573 2428
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 5169 2363 5227 2369
rect 5169 2329 5181 2363
rect 5215 2360 5227 2363
rect 7760 2360 7788 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 8021 2459 8079 2465
rect 9766 2456 9772 2468
rect 9824 2496 9830 2508
rect 11256 2505 11284 2536
rect 11514 2524 11520 2536
rect 11572 2564 11578 2576
rect 11977 2567 12035 2573
rect 11977 2564 11989 2567
rect 11572 2536 11989 2564
rect 11572 2524 11578 2536
rect 11977 2533 11989 2536
rect 12023 2533 12035 2567
rect 11977 2527 12035 2533
rect 10505 2499 10563 2505
rect 10505 2496 10517 2499
rect 9824 2468 10517 2496
rect 9824 2456 9830 2468
rect 10505 2465 10517 2468
rect 10551 2465 10563 2499
rect 10505 2459 10563 2465
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 13722 2456 13728 2508
rect 13780 2496 13786 2508
rect 13817 2499 13875 2505
rect 13817 2496 13829 2499
rect 13780 2468 13829 2496
rect 13780 2456 13786 2468
rect 13817 2465 13829 2468
rect 13863 2496 13875 2499
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 13863 2468 14565 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 16390 2496 16396 2508
rect 16303 2468 16396 2496
rect 14553 2459 14611 2465
rect 16390 2456 16396 2468
rect 16448 2496 16454 2508
rect 17129 2499 17187 2505
rect 17129 2496 17141 2499
rect 16448 2468 17141 2496
rect 16448 2456 16454 2468
rect 17129 2465 17141 2468
rect 17175 2465 17187 2499
rect 17696 2496 17724 2592
rect 18064 2564 18092 2595
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20162 2592 20168 2644
rect 20220 2632 20226 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 20220 2604 20269 2632
rect 20220 2592 20226 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 20806 2592 20812 2644
rect 20864 2632 20870 2644
rect 20901 2635 20959 2641
rect 20901 2632 20913 2635
rect 20864 2604 20913 2632
rect 20864 2592 20870 2604
rect 20901 2601 20913 2604
rect 20947 2601 20959 2635
rect 21450 2632 21456 2644
rect 21411 2604 21456 2632
rect 20901 2595 20959 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 24486 2592 24492 2644
rect 24544 2632 24550 2644
rect 24857 2635 24915 2641
rect 24857 2632 24869 2635
rect 24544 2604 24869 2632
rect 24544 2592 24550 2604
rect 24857 2601 24869 2604
rect 24903 2601 24915 2635
rect 25590 2632 25596 2644
rect 25551 2604 25596 2632
rect 24857 2595 24915 2601
rect 25590 2592 25596 2604
rect 25648 2592 25654 2644
rect 18570 2567 18628 2573
rect 18570 2564 18582 2567
rect 18064 2536 18582 2564
rect 18570 2533 18582 2536
rect 18616 2533 18628 2567
rect 18570 2527 18628 2533
rect 18325 2499 18383 2505
rect 18325 2496 18337 2499
rect 17696 2468 18337 2496
rect 17129 2459 17187 2465
rect 18325 2465 18337 2468
rect 18371 2465 18383 2499
rect 18325 2459 18383 2465
rect 21542 2456 21548 2508
rect 21600 2496 21606 2508
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21600 2468 21833 2496
rect 21600 2456 21606 2468
rect 21821 2465 21833 2468
rect 21867 2496 21879 2499
rect 22557 2499 22615 2505
rect 22557 2496 22569 2499
rect 21867 2468 22569 2496
rect 21867 2465 21879 2468
rect 21821 2459 21879 2465
rect 22557 2465 22569 2468
rect 22603 2465 22615 2499
rect 22557 2459 22615 2465
rect 24121 2499 24179 2505
rect 24121 2465 24133 2499
rect 24167 2496 24179 2499
rect 24504 2496 24532 2592
rect 24167 2468 24532 2496
rect 24167 2465 24179 2468
rect 24121 2459 24179 2465
rect 25314 2456 25320 2508
rect 25372 2496 25378 2508
rect 25409 2499 25467 2505
rect 25409 2496 25421 2499
rect 25372 2468 25421 2496
rect 25372 2456 25378 2468
rect 25409 2465 25421 2468
rect 25455 2496 25467 2499
rect 25961 2499 26019 2505
rect 25961 2496 25973 2499
rect 25455 2468 25973 2496
rect 25455 2465 25467 2468
rect 25409 2459 25467 2465
rect 25961 2465 25973 2468
rect 26007 2465 26019 2499
rect 26878 2496 26884 2508
rect 26839 2468 26884 2496
rect 25961 2459 26019 2465
rect 26878 2456 26884 2468
rect 26936 2496 26942 2508
rect 27433 2499 27491 2505
rect 27433 2496 27445 2499
rect 26936 2468 27445 2496
rect 26936 2456 26942 2468
rect 27433 2465 27445 2468
rect 27479 2465 27491 2499
rect 27433 2459 27491 2465
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9272 2400 9965 2428
rect 9272 2388 9278 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2428 11575 2431
rect 13446 2428 13452 2440
rect 11563 2400 13452 2428
rect 11563 2397 11575 2400
rect 11517 2391 11575 2397
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2428 14151 2431
rect 14918 2428 14924 2440
rect 14139 2400 14924 2428
rect 14139 2397 14151 2400
rect 14093 2391 14151 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 16669 2431 16727 2437
rect 16669 2397 16681 2431
rect 16715 2428 16727 2431
rect 17770 2428 17776 2440
rect 16715 2400 17776 2428
rect 16715 2397 16727 2400
rect 16669 2391 16727 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 22097 2431 22155 2437
rect 22097 2397 22109 2431
rect 22143 2428 22155 2431
rect 23474 2428 23480 2440
rect 22143 2400 23480 2428
rect 22143 2397 22155 2400
rect 22097 2391 22155 2397
rect 23474 2388 23480 2400
rect 23532 2388 23538 2440
rect 24397 2431 24455 2437
rect 24397 2397 24409 2431
rect 24443 2428 24455 2431
rect 26326 2428 26332 2440
rect 24443 2400 26332 2428
rect 24443 2397 24455 2400
rect 24397 2391 24455 2397
rect 26326 2388 26332 2400
rect 26384 2388 26390 2440
rect 5215 2332 7788 2360
rect 5215 2329 5227 2332
rect 5169 2323 5227 2329
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 3510 2252 3516 2304
rect 3568 2292 3574 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 3568 2264 4261 2292
rect 3568 2252 3574 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 27062 2292 27068 2304
rect 27023 2264 27068 2292
rect 4249 2255 4307 2261
rect 27062 2252 27068 2264
rect 27120 2252 27126 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3424 22244 3476 22296
rect 12164 22244 12216 22296
rect 2964 22108 3016 22160
rect 5816 22108 5868 22160
rect 20536 22108 20588 22160
rect 25412 22108 25464 22160
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 8300 21088 8352 21140
rect 21640 21088 21692 21140
rect 3700 20952 3752 21004
rect 10508 20952 10560 21004
rect 20812 20952 20864 21004
rect 4068 20748 4120 20800
rect 7656 20748 7708 20800
rect 23664 20791 23716 20800
rect 23664 20757 23673 20791
rect 23673 20757 23707 20791
rect 23707 20757 23716 20791
rect 23664 20748 23716 20757
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 1860 20587 1912 20596
rect 1860 20553 1869 20587
rect 1869 20553 1903 20587
rect 1903 20553 1912 20587
rect 1860 20544 1912 20553
rect 20812 20587 20864 20596
rect 20812 20553 20821 20587
rect 20821 20553 20855 20587
rect 20855 20553 20864 20587
rect 20812 20544 20864 20553
rect 28264 20544 28316 20596
rect 18328 20408 18380 20460
rect 23388 20408 23440 20460
rect 23664 20451 23716 20460
rect 23664 20417 23673 20451
rect 23673 20417 23707 20451
rect 23707 20417 23716 20451
rect 23664 20408 23716 20417
rect 2964 20383 3016 20392
rect 2964 20349 2973 20383
rect 2973 20349 3007 20383
rect 3007 20349 3016 20383
rect 2964 20340 3016 20349
rect 8484 20383 8536 20392
rect 8484 20349 8493 20383
rect 8493 20349 8527 20383
rect 8527 20349 8536 20383
rect 8484 20340 8536 20349
rect 13912 20383 13964 20392
rect 13912 20349 13921 20383
rect 13921 20349 13955 20383
rect 13955 20349 13964 20383
rect 13912 20340 13964 20349
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 19432 20383 19484 20392
rect 19432 20349 19441 20383
rect 19441 20349 19475 20383
rect 19475 20349 19484 20383
rect 19432 20340 19484 20349
rect 26424 20383 26476 20392
rect 26424 20349 26433 20383
rect 26433 20349 26467 20383
rect 26467 20349 26476 20383
rect 26424 20340 26476 20349
rect 4068 20272 4120 20324
rect 7104 20272 7156 20324
rect 14464 20272 14516 20324
rect 19708 20315 19760 20324
rect 19708 20281 19742 20315
rect 19742 20281 19760 20315
rect 19708 20272 19760 20281
rect 24676 20272 24728 20324
rect 2596 20204 2648 20256
rect 4344 20247 4396 20256
rect 4344 20213 4353 20247
rect 4353 20213 4387 20247
rect 4387 20213 4396 20247
rect 4344 20204 4396 20213
rect 6000 20204 6052 20256
rect 6828 20247 6880 20256
rect 6828 20213 6837 20247
rect 6837 20213 6871 20247
rect 6871 20213 6880 20247
rect 6828 20204 6880 20213
rect 6920 20204 6972 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 9864 20247 9916 20256
rect 9864 20213 9873 20247
rect 9873 20213 9907 20247
rect 9907 20213 9916 20247
rect 9864 20204 9916 20213
rect 15200 20204 15252 20256
rect 24860 20204 24912 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 1676 20000 1728 20052
rect 2412 20000 2464 20052
rect 6000 20043 6052 20052
rect 6000 20009 6009 20043
rect 6009 20009 6043 20043
rect 6043 20009 6052 20043
rect 6000 20000 6052 20009
rect 6920 20043 6972 20052
rect 6920 20009 6929 20043
rect 6929 20009 6963 20043
rect 6963 20009 6972 20043
rect 6920 20000 6972 20009
rect 7104 20043 7156 20052
rect 7104 20009 7113 20043
rect 7113 20009 7147 20043
rect 7147 20009 7156 20043
rect 7104 20000 7156 20009
rect 8484 20043 8536 20052
rect 8484 20009 8493 20043
rect 8493 20009 8527 20043
rect 8527 20009 8536 20043
rect 8484 20000 8536 20009
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 23204 20043 23256 20052
rect 23204 20009 23213 20043
rect 23213 20009 23247 20043
rect 23247 20009 23256 20043
rect 23204 20000 23256 20009
rect 26976 20043 27028 20052
rect 26976 20009 26985 20043
rect 26985 20009 27019 20043
rect 27019 20009 27028 20043
rect 26976 20000 27028 20009
rect 4896 19907 4948 19916
rect 4896 19873 4930 19907
rect 4930 19873 4948 19907
rect 4896 19864 4948 19873
rect 7472 19907 7524 19916
rect 7472 19873 7481 19907
rect 7481 19873 7515 19907
rect 7515 19873 7524 19907
rect 7472 19864 7524 19873
rect 10692 19932 10744 19984
rect 11612 19932 11664 19984
rect 10600 19907 10652 19916
rect 10600 19873 10609 19907
rect 10609 19873 10643 19907
rect 10643 19873 10652 19907
rect 10600 19864 10652 19873
rect 22100 19907 22152 19916
rect 22100 19873 22134 19907
rect 22134 19873 22152 19907
rect 26884 19907 26936 19916
rect 22100 19864 22152 19873
rect 26884 19873 26893 19907
rect 26893 19873 26927 19907
rect 26927 19873 26936 19907
rect 26884 19864 26936 19873
rect 7564 19839 7616 19848
rect 2964 19660 3016 19712
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 7748 19839 7800 19848
rect 7748 19805 7757 19839
rect 7757 19805 7791 19839
rect 7791 19805 7800 19839
rect 7748 19796 7800 19805
rect 16396 19796 16448 19848
rect 16488 19728 16540 19780
rect 17040 19796 17092 19848
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 25044 19839 25096 19848
rect 25044 19805 25053 19839
rect 25053 19805 25087 19839
rect 25087 19805 25096 19839
rect 25044 19796 25096 19805
rect 27068 19839 27120 19848
rect 24860 19728 24912 19780
rect 27068 19805 27077 19839
rect 27077 19805 27111 19839
rect 27111 19805 27120 19839
rect 27068 19796 27120 19805
rect 5356 19660 5408 19712
rect 11336 19660 11388 19712
rect 15660 19703 15712 19712
rect 15660 19669 15669 19703
rect 15669 19669 15703 19703
rect 15703 19669 15712 19703
rect 15660 19660 15712 19669
rect 15844 19660 15896 19712
rect 23848 19703 23900 19712
rect 23848 19669 23857 19703
rect 23857 19669 23891 19703
rect 23891 19669 23900 19703
rect 23848 19660 23900 19669
rect 24032 19660 24084 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 10692 19499 10744 19508
rect 10692 19465 10701 19499
rect 10701 19465 10735 19499
rect 10735 19465 10744 19499
rect 10692 19456 10744 19465
rect 14464 19499 14516 19508
rect 14464 19465 14473 19499
rect 14473 19465 14507 19499
rect 14507 19465 14516 19499
rect 14464 19456 14516 19465
rect 17040 19499 17092 19508
rect 17040 19465 17049 19499
rect 17049 19465 17083 19499
rect 17083 19465 17092 19499
rect 17040 19456 17092 19465
rect 23204 19456 23256 19508
rect 7472 19388 7524 19440
rect 7564 19252 7616 19304
rect 10600 19388 10652 19440
rect 24676 19456 24728 19508
rect 8484 19320 8536 19372
rect 15660 19320 15712 19372
rect 16028 19363 16080 19372
rect 16028 19329 16037 19363
rect 16037 19329 16071 19363
rect 16071 19329 16080 19363
rect 16028 19320 16080 19329
rect 21824 19320 21876 19372
rect 13084 19295 13136 19304
rect 13084 19261 13093 19295
rect 13093 19261 13127 19295
rect 13127 19261 13136 19295
rect 13084 19252 13136 19261
rect 13728 19252 13780 19304
rect 15844 19252 15896 19304
rect 4896 19184 4948 19236
rect 5724 19184 5776 19236
rect 13544 19184 13596 19236
rect 22008 19184 22060 19236
rect 23848 19320 23900 19372
rect 25044 19456 25096 19508
rect 26884 19499 26936 19508
rect 26884 19465 26893 19499
rect 26893 19465 26927 19499
rect 26927 19465 26936 19499
rect 26884 19456 26936 19465
rect 26976 19388 27028 19440
rect 27068 19320 27120 19372
rect 24032 19295 24084 19304
rect 24032 19261 24041 19295
rect 24041 19261 24075 19295
rect 24075 19261 24084 19295
rect 24032 19252 24084 19261
rect 23388 19184 23440 19236
rect 25596 19184 25648 19236
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 5448 19116 5500 19168
rect 7196 19159 7248 19168
rect 7196 19125 7205 19159
rect 7205 19125 7239 19159
rect 7239 19125 7248 19159
rect 7196 19116 7248 19125
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 16396 19116 16448 19168
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 20352 19159 20404 19168
rect 20352 19125 20361 19159
rect 20361 19125 20395 19159
rect 20395 19125 20404 19159
rect 20352 19116 20404 19125
rect 24492 19116 24544 19168
rect 25320 19159 25372 19168
rect 25320 19125 25329 19159
rect 25329 19125 25363 19159
rect 25363 19125 25372 19159
rect 25320 19116 25372 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 7564 18912 7616 18964
rect 7748 18912 7800 18964
rect 13084 18955 13136 18964
rect 13084 18921 13093 18955
rect 13093 18921 13127 18955
rect 13127 18921 13136 18955
rect 13084 18912 13136 18921
rect 14096 18912 14148 18964
rect 15568 18912 15620 18964
rect 16028 18955 16080 18964
rect 16028 18921 16037 18955
rect 16037 18921 16071 18955
rect 16071 18921 16080 18955
rect 16028 18912 16080 18921
rect 23848 18912 23900 18964
rect 25044 18955 25096 18964
rect 25044 18921 25053 18955
rect 25053 18921 25087 18955
rect 25087 18921 25096 18955
rect 25044 18912 25096 18921
rect 26884 18912 26936 18964
rect 10784 18844 10836 18896
rect 11336 18844 11388 18896
rect 2136 18776 2188 18828
rect 3792 18776 3844 18828
rect 4436 18776 4488 18828
rect 7656 18776 7708 18828
rect 10600 18776 10652 18828
rect 15844 18776 15896 18828
rect 18328 18776 18380 18828
rect 21272 18819 21324 18828
rect 21272 18785 21281 18819
rect 21281 18785 21315 18819
rect 21315 18785 21324 18819
rect 21272 18776 21324 18785
rect 21640 18776 21692 18828
rect 23756 18819 23808 18828
rect 23756 18785 23765 18819
rect 23765 18785 23799 18819
rect 23799 18785 23808 18819
rect 23756 18776 23808 18785
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 5264 18708 5316 18760
rect 7840 18751 7892 18760
rect 7840 18717 7849 18751
rect 7849 18717 7883 18751
rect 7883 18717 7892 18751
rect 7840 18708 7892 18717
rect 8484 18708 8536 18760
rect 13820 18708 13872 18760
rect 14372 18708 14424 18760
rect 15108 18708 15160 18760
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 16580 18751 16632 18760
rect 16580 18717 16589 18751
rect 16589 18717 16623 18751
rect 16623 18717 16632 18751
rect 18236 18751 18288 18760
rect 16580 18708 16632 18717
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 23848 18751 23900 18760
rect 23848 18717 23857 18751
rect 23857 18717 23891 18751
rect 23891 18717 23900 18751
rect 23848 18708 23900 18717
rect 23940 18751 23992 18760
rect 23940 18717 23949 18751
rect 23949 18717 23983 18751
rect 23983 18717 23992 18751
rect 23940 18708 23992 18717
rect 24768 18708 24820 18760
rect 1400 18572 1452 18624
rect 2044 18615 2096 18624
rect 2044 18581 2053 18615
rect 2053 18581 2087 18615
rect 2087 18581 2096 18615
rect 2044 18572 2096 18581
rect 2320 18615 2372 18624
rect 2320 18581 2329 18615
rect 2329 18581 2363 18615
rect 2363 18581 2372 18615
rect 2320 18572 2372 18581
rect 4620 18572 4672 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 9036 18615 9088 18624
rect 9036 18581 9045 18615
rect 9045 18581 9079 18615
rect 9079 18581 9088 18615
rect 9036 18572 9088 18581
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 13360 18572 13412 18624
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 19340 18572 19392 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 20812 18572 20864 18624
rect 25596 18615 25648 18624
rect 25596 18581 25605 18615
rect 25605 18581 25639 18615
rect 25639 18581 25648 18615
rect 25596 18572 25648 18581
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 3792 18411 3844 18420
rect 3792 18377 3801 18411
rect 3801 18377 3835 18411
rect 3835 18377 3844 18411
rect 3792 18368 3844 18377
rect 4804 18368 4856 18420
rect 6920 18368 6972 18420
rect 7656 18368 7708 18420
rect 10600 18368 10652 18420
rect 10784 18343 10836 18352
rect 2688 18232 2740 18284
rect 10784 18309 10793 18343
rect 10793 18309 10827 18343
rect 10827 18309 10836 18343
rect 10784 18300 10836 18309
rect 5080 18232 5132 18284
rect 5724 18232 5776 18284
rect 7748 18275 7800 18284
rect 7748 18241 7757 18275
rect 7757 18241 7791 18275
rect 7791 18241 7800 18275
rect 7748 18232 7800 18241
rect 8484 18232 8536 18284
rect 9312 18275 9364 18284
rect 9312 18241 9321 18275
rect 9321 18241 9355 18275
rect 9355 18241 9364 18275
rect 9312 18232 9364 18241
rect 1768 18164 1820 18216
rect 2320 18164 2372 18216
rect 4620 18207 4672 18216
rect 4620 18173 4629 18207
rect 4629 18173 4663 18207
rect 4663 18173 4672 18207
rect 4620 18164 4672 18173
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 9680 18164 9732 18216
rect 13084 18368 13136 18420
rect 13820 18368 13872 18420
rect 15844 18368 15896 18420
rect 16488 18411 16540 18420
rect 16488 18377 16497 18411
rect 16497 18377 16531 18411
rect 16531 18377 16540 18411
rect 16488 18368 16540 18377
rect 18236 18368 18288 18420
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 19248 18368 19300 18420
rect 21272 18411 21324 18420
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 23756 18411 23808 18420
rect 23756 18377 23765 18411
rect 23765 18377 23799 18411
rect 23799 18377 23808 18411
rect 23756 18368 23808 18377
rect 27068 18368 27120 18420
rect 14372 18343 14424 18352
rect 14372 18309 14381 18343
rect 14381 18309 14415 18343
rect 14415 18309 14424 18343
rect 14372 18300 14424 18309
rect 14464 18300 14516 18352
rect 15016 18232 15068 18284
rect 15568 18300 15620 18352
rect 21640 18343 21692 18352
rect 21640 18309 21649 18343
rect 21649 18309 21683 18343
rect 21683 18309 21692 18343
rect 21640 18300 21692 18309
rect 22008 18300 22060 18352
rect 23940 18300 23992 18352
rect 15844 18232 15896 18284
rect 16580 18232 16632 18284
rect 18328 18232 18380 18284
rect 20260 18232 20312 18284
rect 12440 18207 12492 18216
rect 12440 18173 12449 18207
rect 12449 18173 12483 18207
rect 12483 18173 12492 18207
rect 20076 18207 20128 18216
rect 12440 18164 12492 18173
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20352 18164 20404 18216
rect 24676 18232 24728 18284
rect 25780 18164 25832 18216
rect 26148 18207 26200 18216
rect 26148 18173 26157 18207
rect 26157 18173 26191 18207
rect 26191 18173 26200 18207
rect 26148 18164 26200 18173
rect 2044 18096 2096 18148
rect 2504 18096 2556 18148
rect 7840 18096 7892 18148
rect 4252 18071 4304 18080
rect 4252 18037 4261 18071
rect 4261 18037 4295 18071
rect 4295 18037 4304 18071
rect 4252 18028 4304 18037
rect 4344 18028 4396 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 13452 18096 13504 18148
rect 20536 18096 20588 18148
rect 8760 18028 8812 18080
rect 9588 18028 9640 18080
rect 13544 18028 13596 18080
rect 14556 18028 14608 18080
rect 15292 18071 15344 18080
rect 15292 18037 15301 18071
rect 15301 18037 15335 18071
rect 15335 18037 15344 18071
rect 15292 18028 15344 18037
rect 18328 18071 18380 18080
rect 18328 18037 18337 18071
rect 18337 18037 18371 18071
rect 18371 18037 18380 18071
rect 18328 18028 18380 18037
rect 20628 18028 20680 18080
rect 24124 18071 24176 18080
rect 24124 18037 24133 18071
rect 24133 18037 24167 18071
rect 24167 18037 24176 18071
rect 24124 18028 24176 18037
rect 24216 18071 24268 18080
rect 24216 18037 24225 18071
rect 24225 18037 24259 18071
rect 24259 18037 24268 18071
rect 24216 18028 24268 18037
rect 25044 18028 25096 18080
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 2136 17824 2188 17876
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 4712 17867 4764 17876
rect 4712 17833 4721 17867
rect 4721 17833 4755 17867
rect 4755 17833 4764 17867
rect 4712 17824 4764 17833
rect 7472 17824 7524 17876
rect 9680 17867 9732 17876
rect 9680 17833 9689 17867
rect 9689 17833 9723 17867
rect 9723 17833 9732 17867
rect 9680 17824 9732 17833
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 13728 17867 13780 17876
rect 12440 17824 12492 17833
rect 13728 17833 13737 17867
rect 13737 17833 13771 17867
rect 13771 17833 13780 17867
rect 13728 17824 13780 17833
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 20720 17824 20772 17876
rect 22560 17824 22612 17876
rect 23848 17824 23900 17876
rect 26240 17867 26292 17876
rect 26240 17833 26249 17867
rect 26249 17833 26283 17867
rect 26283 17833 26292 17867
rect 26240 17824 26292 17833
rect 7840 17799 7892 17808
rect 7840 17765 7849 17799
rect 7849 17765 7883 17799
rect 7883 17765 7892 17799
rect 7840 17756 7892 17765
rect 17316 17756 17368 17808
rect 24032 17756 24084 17808
rect 1676 17688 1728 17740
rect 4068 17688 4120 17740
rect 7932 17688 7984 17740
rect 8024 17688 8076 17740
rect 10416 17688 10468 17740
rect 15660 17731 15712 17740
rect 15660 17697 15669 17731
rect 15669 17697 15703 17731
rect 15703 17697 15712 17731
rect 15660 17688 15712 17697
rect 20628 17688 20680 17740
rect 21824 17688 21876 17740
rect 24308 17731 24360 17740
rect 24308 17697 24317 17731
rect 24317 17697 24351 17731
rect 24351 17697 24360 17731
rect 24308 17688 24360 17697
rect 2320 17620 2372 17672
rect 2688 17620 2740 17672
rect 4160 17552 4212 17604
rect 5264 17620 5316 17672
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8576 17663 8628 17672
rect 8576 17629 8585 17663
rect 8585 17629 8619 17663
rect 8619 17629 8628 17663
rect 10140 17663 10192 17672
rect 8576 17620 8628 17629
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 10784 17620 10836 17672
rect 15568 17620 15620 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 17224 17620 17276 17672
rect 16580 17552 16632 17604
rect 20168 17620 20220 17672
rect 20812 17620 20864 17672
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 24400 17663 24452 17672
rect 21456 17620 21508 17629
rect 24400 17629 24409 17663
rect 24409 17629 24443 17663
rect 24443 17629 24452 17663
rect 24400 17620 24452 17629
rect 24676 17756 24728 17808
rect 26516 17731 26568 17740
rect 26516 17697 26525 17731
rect 26525 17697 26559 17731
rect 26559 17697 26568 17731
rect 26516 17688 26568 17697
rect 1492 17484 1544 17536
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 16856 17527 16908 17536
rect 16856 17493 16865 17527
rect 16865 17493 16899 17527
rect 16899 17493 16908 17527
rect 16856 17484 16908 17493
rect 18880 17484 18932 17536
rect 21272 17484 21324 17536
rect 25044 17527 25096 17536
rect 25044 17493 25053 17527
rect 25053 17493 25087 17527
rect 25087 17493 25096 17527
rect 25044 17484 25096 17493
rect 26884 17484 26936 17536
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 4068 17323 4120 17332
rect 1676 17280 1728 17289
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 8484 17280 8536 17332
rect 10784 17323 10836 17332
rect 10784 17289 10793 17323
rect 10793 17289 10827 17323
rect 10827 17289 10836 17323
rect 10784 17280 10836 17289
rect 14556 17323 14608 17332
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 2320 17144 2372 17196
rect 4712 17144 4764 17196
rect 5356 17212 5408 17264
rect 6184 17144 6236 17196
rect 8576 17144 8628 17196
rect 9404 17144 9456 17196
rect 10784 17144 10836 17196
rect 15016 17280 15068 17332
rect 15660 17280 15712 17332
rect 18236 17323 18288 17332
rect 18236 17289 18245 17323
rect 18245 17289 18279 17323
rect 18279 17289 18288 17323
rect 18236 17280 18288 17289
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 22560 17323 22612 17332
rect 22560 17289 22569 17323
rect 22569 17289 22603 17323
rect 22603 17289 22612 17323
rect 22560 17280 22612 17289
rect 26516 17323 26568 17332
rect 26516 17289 26525 17323
rect 26525 17289 26559 17323
rect 26559 17289 26568 17323
rect 26516 17280 26568 17289
rect 24308 17212 24360 17264
rect 24952 17212 25004 17264
rect 25320 17212 25372 17264
rect 15844 17144 15896 17196
rect 18328 17144 18380 17196
rect 19064 17187 19116 17196
rect 19064 17153 19073 17187
rect 19073 17153 19107 17187
rect 19107 17153 19116 17187
rect 19064 17144 19116 17153
rect 20628 17187 20680 17196
rect 20628 17153 20637 17187
rect 20637 17153 20671 17187
rect 20671 17153 20680 17187
rect 20628 17144 20680 17153
rect 25044 17187 25096 17196
rect 25044 17153 25053 17187
rect 25053 17153 25087 17187
rect 25087 17153 25096 17187
rect 25044 17144 25096 17153
rect 1860 17076 1912 17128
rect 2688 17076 2740 17128
rect 4252 17076 4304 17128
rect 16856 17076 16908 17128
rect 18236 17076 18288 17128
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 23940 17076 23992 17128
rect 24860 17076 24912 17128
rect 9864 17008 9916 17060
rect 17224 17008 17276 17060
rect 17868 17008 17920 17060
rect 21456 17008 21508 17060
rect 24400 17008 24452 17060
rect 2228 16940 2280 16992
rect 4712 16940 4764 16992
rect 8024 16983 8076 16992
rect 8024 16949 8033 16983
rect 8033 16949 8067 16983
rect 8067 16949 8076 16983
rect 8024 16940 8076 16949
rect 8852 16983 8904 16992
rect 8852 16949 8861 16983
rect 8861 16949 8895 16983
rect 8895 16949 8904 16983
rect 8852 16940 8904 16949
rect 9128 16940 9180 16992
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 15476 16983 15528 16992
rect 15476 16949 15485 16983
rect 15485 16949 15519 16983
rect 15519 16949 15528 16983
rect 15476 16940 15528 16949
rect 16580 16983 16632 16992
rect 16580 16949 16589 16983
rect 16589 16949 16623 16983
rect 16623 16949 16632 16983
rect 16580 16940 16632 16949
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 18420 16983 18472 16992
rect 18420 16949 18429 16983
rect 18429 16949 18463 16983
rect 18463 16949 18472 16983
rect 18420 16940 18472 16949
rect 20444 16983 20496 16992
rect 20444 16949 20453 16983
rect 20453 16949 20487 16983
rect 20487 16949 20496 16983
rect 20444 16940 20496 16949
rect 21640 16940 21692 16992
rect 24308 16983 24360 16992
rect 24308 16949 24317 16983
rect 24317 16949 24351 16983
rect 24351 16949 24360 16983
rect 24860 16983 24912 16992
rect 24308 16940 24360 16949
rect 24860 16949 24869 16983
rect 24869 16949 24903 16983
rect 24903 16949 24912 16983
rect 24860 16940 24912 16949
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2320 16779 2372 16788
rect 2320 16745 2329 16779
rect 2329 16745 2363 16779
rect 2363 16745 2372 16779
rect 2320 16736 2372 16745
rect 6184 16779 6236 16788
rect 6184 16745 6193 16779
rect 6193 16745 6227 16779
rect 6227 16745 6236 16779
rect 6184 16736 6236 16745
rect 9680 16779 9732 16788
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 13452 16736 13504 16788
rect 15476 16736 15528 16788
rect 5080 16711 5132 16720
rect 5080 16677 5114 16711
rect 5114 16677 5132 16711
rect 5080 16668 5132 16677
rect 10324 16668 10376 16720
rect 15292 16668 15344 16720
rect 19340 16668 19392 16720
rect 20444 16668 20496 16720
rect 1584 16600 1636 16652
rect 2688 16600 2740 16652
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 4160 16600 4212 16652
rect 9128 16643 9180 16652
rect 9128 16609 9137 16643
rect 9137 16609 9171 16643
rect 9171 16609 9180 16643
rect 9128 16600 9180 16609
rect 12348 16643 12400 16652
rect 12348 16609 12357 16643
rect 12357 16609 12391 16643
rect 12391 16609 12400 16643
rect 12348 16600 12400 16609
rect 12440 16600 12492 16652
rect 13728 16600 13780 16652
rect 4804 16575 4856 16584
rect 1768 16464 1820 16516
rect 2136 16464 2188 16516
rect 4804 16541 4813 16575
rect 4813 16541 4847 16575
rect 4847 16541 4856 16575
rect 4804 16532 4856 16541
rect 9864 16532 9916 16584
rect 10784 16532 10836 16584
rect 15568 16600 15620 16652
rect 18420 16600 18472 16652
rect 21272 16779 21324 16788
rect 21272 16745 21281 16779
rect 21281 16745 21315 16779
rect 21315 16745 21324 16779
rect 21272 16736 21324 16745
rect 24032 16779 24084 16788
rect 24032 16745 24041 16779
rect 24041 16745 24075 16779
rect 24075 16745 24084 16779
rect 24032 16736 24084 16745
rect 24400 16736 24452 16788
rect 21548 16668 21600 16720
rect 25412 16668 25464 16720
rect 21364 16643 21416 16652
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 16580 16532 16632 16584
rect 16672 16532 16724 16584
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 24768 16600 24820 16652
rect 17868 16464 17920 16516
rect 20168 16532 20220 16584
rect 21640 16532 21692 16584
rect 25044 16575 25096 16584
rect 25044 16541 25053 16575
rect 25053 16541 25087 16575
rect 25087 16541 25096 16575
rect 25044 16532 25096 16541
rect 19340 16464 19392 16516
rect 24676 16396 24728 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 1584 16192 1636 16244
rect 2504 16192 2556 16244
rect 4160 16192 4212 16244
rect 5080 16192 5132 16244
rect 6276 16192 6328 16244
rect 9404 16235 9456 16244
rect 2136 16056 2188 16108
rect 9404 16201 9413 16235
rect 9413 16201 9447 16235
rect 9447 16201 9456 16235
rect 9404 16192 9456 16201
rect 12348 16192 12400 16244
rect 13728 16192 13780 16244
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 16672 16192 16724 16244
rect 17868 16235 17920 16244
rect 17868 16201 17877 16235
rect 17877 16201 17911 16235
rect 17911 16201 17920 16235
rect 17868 16192 17920 16201
rect 18880 16192 18932 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 21272 16192 21324 16244
rect 24216 16192 24268 16244
rect 24768 16192 24820 16244
rect 21364 16167 21416 16176
rect 4804 15988 4856 16040
rect 5448 15988 5500 16040
rect 6828 16031 6880 16040
rect 6828 15997 6837 16031
rect 6837 15997 6871 16031
rect 6871 15997 6880 16031
rect 6828 15988 6880 15997
rect 9680 16056 9732 16108
rect 21364 16133 21373 16167
rect 21373 16133 21407 16167
rect 21407 16133 21416 16167
rect 21364 16124 21416 16133
rect 12256 16056 12308 16108
rect 16580 16056 16632 16108
rect 19064 16099 19116 16108
rect 19064 16065 19073 16099
rect 19073 16065 19107 16099
rect 19107 16065 19116 16099
rect 19064 16056 19116 16065
rect 21640 16056 21692 16108
rect 24952 16099 25004 16108
rect 24952 16065 24961 16099
rect 24961 16065 24995 16099
rect 24995 16065 25004 16099
rect 24952 16056 25004 16065
rect 25044 16056 25096 16108
rect 25688 16056 25740 16108
rect 9588 15988 9640 16040
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 16396 15988 16448 16040
rect 24400 15988 24452 16040
rect 25504 15988 25556 16040
rect 25964 15988 26016 16040
rect 2688 15920 2740 15972
rect 10232 15920 10284 15972
rect 11888 15963 11940 15972
rect 8208 15895 8260 15904
rect 8208 15861 8217 15895
rect 8217 15861 8251 15895
rect 8251 15861 8260 15895
rect 8208 15852 8260 15861
rect 9864 15852 9916 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 11888 15929 11897 15963
rect 11897 15929 11931 15963
rect 11931 15929 11940 15963
rect 11888 15920 11940 15929
rect 15384 15963 15436 15972
rect 15384 15929 15393 15963
rect 15393 15929 15427 15963
rect 15427 15929 15436 15963
rect 15384 15920 15436 15929
rect 15292 15852 15344 15904
rect 24860 15920 24912 15972
rect 25044 15920 25096 15972
rect 18788 15895 18840 15904
rect 18788 15861 18797 15895
rect 18797 15861 18831 15895
rect 18831 15861 18840 15895
rect 18788 15852 18840 15861
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 24124 15895 24176 15904
rect 24124 15861 24133 15895
rect 24133 15861 24167 15895
rect 24167 15861 24176 15895
rect 24124 15852 24176 15861
rect 24676 15895 24728 15904
rect 24676 15861 24685 15895
rect 24685 15861 24719 15895
rect 24719 15861 24728 15895
rect 24676 15852 24728 15861
rect 25688 15895 25740 15904
rect 25688 15861 25697 15895
rect 25697 15861 25731 15895
rect 25731 15861 25740 15895
rect 25688 15852 25740 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 2228 15648 2280 15700
rect 11888 15648 11940 15700
rect 12256 15648 12308 15700
rect 18880 15691 18932 15700
rect 18880 15657 18889 15691
rect 18889 15657 18923 15691
rect 18923 15657 18932 15691
rect 18880 15648 18932 15657
rect 24952 15691 25004 15700
rect 24952 15657 24961 15691
rect 24961 15657 24995 15691
rect 24995 15657 25004 15691
rect 24952 15648 25004 15657
rect 25504 15648 25556 15700
rect 25964 15691 26016 15700
rect 25964 15657 25973 15691
rect 25973 15657 26007 15691
rect 26007 15657 26016 15691
rect 25964 15648 26016 15657
rect 2136 15623 2188 15632
rect 2136 15589 2145 15623
rect 2145 15589 2179 15623
rect 2179 15589 2188 15623
rect 2136 15580 2188 15589
rect 15200 15580 15252 15632
rect 17960 15580 18012 15632
rect 19340 15623 19392 15632
rect 19340 15589 19349 15623
rect 19349 15589 19383 15623
rect 19383 15589 19392 15623
rect 19340 15580 19392 15589
rect 21640 15580 21692 15632
rect 7288 15555 7340 15564
rect 2228 15487 2280 15496
rect 2228 15453 2237 15487
rect 2237 15453 2271 15487
rect 2271 15453 2280 15487
rect 2228 15444 2280 15453
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 9680 15555 9732 15564
rect 9680 15521 9689 15555
rect 9689 15521 9723 15555
rect 9723 15521 9732 15555
rect 9680 15512 9732 15521
rect 9956 15555 10008 15564
rect 9956 15521 9990 15555
rect 9990 15521 10008 15555
rect 9956 15512 10008 15521
rect 18604 15512 18656 15564
rect 19248 15555 19300 15564
rect 19248 15521 19257 15555
rect 19257 15521 19291 15555
rect 19291 15521 19300 15555
rect 19248 15512 19300 15521
rect 21824 15512 21876 15564
rect 24952 15512 25004 15564
rect 25228 15512 25280 15564
rect 26516 15555 26568 15564
rect 26516 15521 26525 15555
rect 26525 15521 26559 15555
rect 26559 15521 26568 15555
rect 26516 15512 26568 15521
rect 2504 15444 2556 15496
rect 3056 15444 3108 15496
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 19616 15444 19668 15496
rect 2688 15308 2740 15360
rect 6828 15308 6880 15360
rect 7656 15308 7708 15360
rect 12808 15308 12860 15360
rect 16672 15351 16724 15360
rect 16672 15317 16681 15351
rect 16681 15317 16715 15351
rect 16715 15317 16724 15351
rect 16672 15308 16724 15317
rect 19064 15308 19116 15360
rect 20720 15308 20772 15360
rect 23388 15351 23440 15360
rect 23388 15317 23397 15351
rect 23397 15317 23431 15351
rect 23431 15317 23440 15351
rect 23388 15308 23440 15317
rect 24584 15351 24636 15360
rect 24584 15317 24593 15351
rect 24593 15317 24627 15351
rect 24627 15317 24636 15351
rect 24584 15308 24636 15317
rect 25412 15308 25464 15360
rect 26792 15308 26844 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 7288 15104 7340 15156
rect 9588 15104 9640 15156
rect 9680 15104 9732 15156
rect 12164 15147 12216 15156
rect 12164 15113 12173 15147
rect 12173 15113 12207 15147
rect 12207 15113 12216 15147
rect 12164 15104 12216 15113
rect 15200 15147 15252 15156
rect 15200 15113 15209 15147
rect 15209 15113 15243 15147
rect 15243 15113 15252 15147
rect 15200 15104 15252 15113
rect 18604 15147 18656 15156
rect 18604 15113 18613 15147
rect 18613 15113 18647 15147
rect 18647 15113 18656 15147
rect 18604 15104 18656 15113
rect 18696 15104 18748 15156
rect 19340 15147 19392 15156
rect 19340 15113 19349 15147
rect 19349 15113 19383 15147
rect 19383 15113 19392 15147
rect 19340 15104 19392 15113
rect 19708 15104 19760 15156
rect 20720 15104 20772 15156
rect 21640 15104 21692 15156
rect 26516 15147 26568 15156
rect 26516 15113 26525 15147
rect 26525 15113 26559 15147
rect 26559 15113 26568 15147
rect 26516 15104 26568 15113
rect 2228 15036 2280 15088
rect 15292 15036 15344 15088
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 16396 14968 16448 15020
rect 16672 14968 16724 15020
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 2228 14832 2280 14884
rect 2872 14832 2924 14884
rect 8208 14900 8260 14952
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 8300 14764 8352 14816
rect 9956 14900 10008 14952
rect 12624 14900 12676 14952
rect 12164 14832 12216 14884
rect 12900 14900 12952 14952
rect 15660 14900 15712 14952
rect 19340 14900 19392 14952
rect 19524 14943 19576 14952
rect 19524 14909 19533 14943
rect 19533 14909 19567 14943
rect 19567 14909 19576 14943
rect 19524 14900 19576 14909
rect 11888 14764 11940 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 12808 14764 12860 14816
rect 15752 14764 15804 14816
rect 19616 14832 19668 14884
rect 16488 14764 16540 14816
rect 21824 14764 21876 14816
rect 23940 14764 23992 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 2228 14603 2280 14612
rect 2228 14569 2237 14603
rect 2237 14569 2271 14603
rect 2271 14569 2280 14603
rect 2228 14560 2280 14569
rect 2688 14560 2740 14612
rect 8300 14603 8352 14612
rect 8300 14569 8309 14603
rect 8309 14569 8343 14603
rect 8343 14569 8352 14603
rect 8300 14560 8352 14569
rect 9588 14560 9640 14612
rect 11888 14603 11940 14612
rect 11888 14569 11897 14603
rect 11897 14569 11931 14603
rect 11931 14569 11940 14603
rect 11888 14560 11940 14569
rect 16580 14560 16632 14612
rect 19524 14560 19576 14612
rect 2136 14492 2188 14544
rect 5448 14492 5500 14544
rect 15292 14492 15344 14544
rect 2780 14424 2832 14476
rect 5080 14424 5132 14476
rect 9036 14467 9088 14476
rect 9036 14433 9045 14467
rect 9045 14433 9079 14467
rect 9079 14433 9088 14467
rect 9036 14424 9088 14433
rect 13728 14424 13780 14476
rect 16672 14492 16724 14544
rect 18788 14492 18840 14544
rect 16396 14467 16448 14476
rect 16396 14433 16430 14467
rect 16430 14433 16448 14467
rect 16396 14424 16448 14433
rect 19340 14424 19392 14476
rect 21824 14560 21876 14612
rect 23388 14492 23440 14544
rect 21732 14467 21784 14476
rect 21732 14433 21766 14467
rect 21766 14433 21784 14467
rect 21732 14424 21784 14433
rect 23296 14424 23348 14476
rect 10784 14356 10836 14408
rect 12348 14356 12400 14408
rect 13544 14399 13596 14408
rect 13544 14365 13553 14399
rect 13553 14365 13587 14399
rect 13587 14365 13596 14399
rect 13544 14356 13596 14365
rect 23940 14399 23992 14408
rect 23940 14365 23949 14399
rect 23949 14365 23983 14399
rect 23983 14365 23992 14399
rect 23940 14356 23992 14365
rect 25044 14356 25096 14408
rect 25780 14356 25832 14408
rect 4988 14220 5040 14272
rect 7656 14220 7708 14272
rect 8576 14220 8628 14272
rect 11060 14220 11112 14272
rect 11520 14263 11572 14272
rect 11520 14229 11529 14263
rect 11529 14229 11563 14263
rect 11563 14229 11572 14263
rect 11520 14220 11572 14229
rect 12624 14263 12676 14272
rect 12624 14229 12633 14263
rect 12633 14229 12667 14263
rect 12667 14229 12676 14263
rect 12624 14220 12676 14229
rect 12808 14220 12860 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 19616 14263 19668 14272
rect 19616 14229 19625 14263
rect 19625 14229 19659 14263
rect 19659 14229 19668 14263
rect 19616 14220 19668 14229
rect 23296 14220 23348 14272
rect 25872 14220 25924 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 5080 14016 5132 14068
rect 7656 14016 7708 14068
rect 10784 14059 10836 14068
rect 10784 14025 10793 14059
rect 10793 14025 10827 14059
rect 10827 14025 10836 14059
rect 10784 14016 10836 14025
rect 11888 14016 11940 14068
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 19616 14016 19668 14068
rect 21824 14059 21876 14068
rect 21824 14025 21833 14059
rect 21833 14025 21867 14059
rect 21867 14025 21876 14059
rect 21824 14016 21876 14025
rect 4068 13948 4120 14000
rect 8208 13991 8260 14000
rect 8208 13957 8217 13991
rect 8217 13957 8251 13991
rect 8251 13957 8260 13991
rect 8208 13948 8260 13957
rect 2872 13812 2924 13864
rect 4436 13812 4488 13864
rect 8300 13880 8352 13932
rect 11980 13948 12032 14000
rect 12348 13880 12400 13932
rect 12440 13880 12492 13932
rect 21732 13948 21784 14000
rect 23940 13948 23992 14000
rect 27436 13991 27488 14000
rect 16396 13923 16448 13932
rect 16396 13889 16405 13923
rect 16405 13889 16439 13923
rect 16439 13889 16448 13923
rect 27436 13957 27445 13991
rect 27445 13957 27479 13991
rect 27479 13957 27488 13991
rect 27436 13948 27488 13957
rect 16396 13880 16448 13889
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 7472 13812 7524 13864
rect 2780 13744 2832 13796
rect 4252 13787 4304 13796
rect 4252 13753 4261 13787
rect 4261 13753 4295 13787
rect 4295 13753 4304 13787
rect 4252 13744 4304 13753
rect 1768 13719 1820 13728
rect 1768 13685 1777 13719
rect 1777 13685 1811 13719
rect 1811 13685 1820 13719
rect 1768 13676 1820 13685
rect 4344 13719 4396 13728
rect 4344 13685 4353 13719
rect 4353 13685 4387 13719
rect 4387 13685 4396 13719
rect 4344 13676 4396 13685
rect 4988 13744 5040 13796
rect 8392 13744 8444 13796
rect 9036 13744 9088 13796
rect 10784 13744 10836 13796
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 13728 13812 13780 13864
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 11060 13744 11112 13796
rect 11336 13744 11388 13796
rect 15292 13787 15344 13796
rect 15292 13753 15301 13787
rect 15301 13753 15335 13787
rect 15335 13753 15344 13787
rect 15292 13744 15344 13753
rect 16304 13744 16356 13796
rect 5632 13676 5684 13728
rect 8208 13676 8260 13728
rect 9588 13676 9640 13728
rect 12256 13676 12308 13728
rect 13544 13676 13596 13728
rect 15660 13676 15712 13728
rect 18788 13812 18840 13864
rect 25504 13880 25556 13932
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 26056 13880 26108 13889
rect 19524 13855 19576 13864
rect 19524 13821 19558 13855
rect 19558 13821 19576 13855
rect 19524 13812 19576 13821
rect 23296 13812 23348 13864
rect 19432 13744 19484 13796
rect 17592 13676 17644 13728
rect 25872 13719 25924 13728
rect 25872 13685 25881 13719
rect 25881 13685 25915 13719
rect 25915 13685 25924 13719
rect 25872 13676 25924 13685
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 1768 13515 1820 13524
rect 1768 13481 1777 13515
rect 1777 13481 1811 13515
rect 1811 13481 1820 13515
rect 1768 13472 1820 13481
rect 2872 13515 2924 13524
rect 2872 13481 2881 13515
rect 2881 13481 2915 13515
rect 2915 13481 2924 13515
rect 2872 13472 2924 13481
rect 4528 13472 4580 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 10784 13515 10836 13524
rect 10784 13481 10793 13515
rect 10793 13481 10827 13515
rect 10827 13481 10836 13515
rect 10784 13472 10836 13481
rect 11336 13472 11388 13524
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 13728 13472 13780 13524
rect 19340 13472 19392 13524
rect 26056 13515 26108 13524
rect 26056 13481 26065 13515
rect 26065 13481 26099 13515
rect 26099 13481 26108 13515
rect 26056 13472 26108 13481
rect 2964 13404 3016 13456
rect 15200 13404 15252 13456
rect 15752 13447 15804 13456
rect 15752 13413 15761 13447
rect 15761 13413 15795 13447
rect 15795 13413 15804 13447
rect 15752 13404 15804 13413
rect 16672 13404 16724 13456
rect 19432 13404 19484 13456
rect 3332 13336 3384 13388
rect 4160 13336 4212 13388
rect 7840 13379 7892 13388
rect 2504 13311 2556 13320
rect 2504 13277 2513 13311
rect 2513 13277 2547 13311
rect 2547 13277 2556 13311
rect 2504 13268 2556 13277
rect 4344 13268 4396 13320
rect 7840 13345 7849 13379
rect 7849 13345 7883 13379
rect 7883 13345 7892 13379
rect 7840 13336 7892 13345
rect 7932 13379 7984 13388
rect 7932 13345 7941 13379
rect 7941 13345 7975 13379
rect 7975 13345 7984 13379
rect 7932 13336 7984 13345
rect 11244 13336 11296 13388
rect 17224 13379 17276 13388
rect 17224 13345 17233 13379
rect 17233 13345 17267 13379
rect 17267 13345 17276 13379
rect 17224 13336 17276 13345
rect 19984 13336 20036 13388
rect 22928 13336 22980 13388
rect 5080 13268 5132 13320
rect 7564 13268 7616 13320
rect 7748 13268 7800 13320
rect 8116 13311 8168 13320
rect 8116 13277 8125 13311
rect 8125 13277 8159 13311
rect 8159 13277 8168 13311
rect 8116 13268 8168 13277
rect 11704 13311 11756 13320
rect 11704 13277 11713 13311
rect 11713 13277 11747 13311
rect 11747 13277 11756 13311
rect 11704 13268 11756 13277
rect 12072 13268 12124 13320
rect 12624 13268 12676 13320
rect 16488 13268 16540 13320
rect 17408 13268 17460 13320
rect 17592 13268 17644 13320
rect 22284 13268 22336 13320
rect 23388 13268 23440 13320
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4160 13132 4212 13184
rect 15752 13132 15804 13184
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 24216 13175 24268 13184
rect 24216 13141 24225 13175
rect 24225 13141 24259 13175
rect 24259 13141 24268 13175
rect 24216 13132 24268 13141
rect 25780 13175 25832 13184
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 2964 12971 3016 12980
rect 2964 12937 2973 12971
rect 2973 12937 3007 12971
rect 3007 12937 3016 12971
rect 2964 12928 3016 12937
rect 4528 12928 4580 12980
rect 5080 12971 5132 12980
rect 5080 12937 5089 12971
rect 5089 12937 5123 12971
rect 5123 12937 5132 12971
rect 5080 12928 5132 12937
rect 7564 12971 7616 12980
rect 7564 12937 7573 12971
rect 7573 12937 7607 12971
rect 7607 12937 7616 12971
rect 7564 12928 7616 12937
rect 7840 12971 7892 12980
rect 7840 12937 7849 12971
rect 7849 12937 7883 12971
rect 7883 12937 7892 12971
rect 7840 12928 7892 12937
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 572 12860 624 12912
rect 7012 12860 7064 12912
rect 8116 12860 8168 12912
rect 2320 12835 2372 12844
rect 2320 12801 2329 12835
rect 2329 12801 2363 12835
rect 2363 12801 2372 12835
rect 2320 12792 2372 12801
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3884 12792 3936 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 16488 12928 16540 12980
rect 17592 12971 17644 12980
rect 17592 12937 17601 12971
rect 17601 12937 17635 12971
rect 17635 12937 17644 12971
rect 17592 12928 17644 12937
rect 22284 12928 22336 12980
rect 23388 12928 23440 12980
rect 22008 12860 22060 12912
rect 22928 12860 22980 12912
rect 24952 12860 25004 12912
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 19064 12792 19116 12844
rect 19432 12792 19484 12844
rect 25872 12792 25924 12844
rect 4160 12724 4212 12776
rect 8576 12767 8628 12776
rect 8576 12733 8585 12767
rect 8585 12733 8619 12767
rect 8619 12733 8628 12767
rect 8576 12724 8628 12733
rect 11244 12767 11296 12776
rect 11244 12733 11253 12767
rect 11253 12733 11287 12767
rect 11287 12733 11296 12767
rect 11244 12724 11296 12733
rect 11704 12767 11756 12776
rect 11704 12733 11713 12767
rect 11713 12733 11747 12767
rect 11747 12733 11756 12767
rect 11704 12724 11756 12733
rect 17224 12724 17276 12776
rect 2320 12656 2372 12708
rect 2780 12656 2832 12708
rect 3792 12656 3844 12708
rect 2044 12588 2096 12640
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 3976 12588 4028 12640
rect 8944 12656 8996 12708
rect 15016 12699 15068 12708
rect 15016 12665 15025 12699
rect 15025 12665 15059 12699
rect 15059 12665 15068 12699
rect 15016 12656 15068 12665
rect 16580 12656 16632 12708
rect 17408 12656 17460 12708
rect 18880 12656 18932 12708
rect 24216 12724 24268 12776
rect 25780 12724 25832 12776
rect 24400 12656 24452 12708
rect 9956 12631 10008 12640
rect 9956 12597 9965 12631
rect 9965 12597 9999 12631
rect 9999 12597 10008 12631
rect 9956 12588 10008 12597
rect 14740 12631 14792 12640
rect 14740 12597 14749 12631
rect 14749 12597 14783 12631
rect 14783 12597 14792 12631
rect 14740 12588 14792 12597
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 17224 12588 17276 12640
rect 17684 12588 17736 12640
rect 19616 12588 19668 12640
rect 20444 12588 20496 12640
rect 24584 12631 24636 12640
rect 24584 12597 24593 12631
rect 24593 12597 24627 12631
rect 24627 12597 24636 12631
rect 24584 12588 24636 12597
rect 25412 12588 25464 12640
rect 25688 12631 25740 12640
rect 25688 12597 25697 12631
rect 25697 12597 25731 12631
rect 25731 12597 25740 12631
rect 25688 12588 25740 12597
rect 26148 12631 26200 12640
rect 26148 12597 26157 12631
rect 26157 12597 26191 12631
rect 26191 12597 26200 12631
rect 26148 12588 26200 12597
rect 26332 12588 26384 12640
rect 26516 12588 26568 12640
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 1860 12384 1912 12436
rect 4344 12427 4396 12436
rect 4344 12393 4353 12427
rect 4353 12393 4387 12427
rect 4387 12393 4396 12427
rect 4344 12384 4396 12393
rect 7656 12427 7708 12436
rect 7656 12393 7665 12427
rect 7665 12393 7699 12427
rect 7699 12393 7708 12427
rect 7656 12384 7708 12393
rect 8576 12427 8628 12436
rect 8576 12393 8585 12427
rect 8585 12393 8619 12427
rect 8619 12393 8628 12427
rect 8576 12384 8628 12393
rect 15108 12427 15160 12436
rect 15108 12393 15117 12427
rect 15117 12393 15151 12427
rect 15151 12393 15160 12427
rect 15108 12384 15160 12393
rect 19524 12384 19576 12436
rect 20444 12384 20496 12436
rect 22376 12384 22428 12436
rect 23204 12427 23256 12436
rect 23204 12393 23213 12427
rect 23213 12393 23247 12427
rect 23247 12393 23256 12427
rect 23204 12384 23256 12393
rect 24216 12384 24268 12436
rect 24768 12427 24820 12436
rect 24768 12393 24777 12427
rect 24777 12393 24811 12427
rect 24811 12393 24820 12427
rect 24768 12384 24820 12393
rect 25504 12384 25556 12436
rect 25872 12384 25924 12436
rect 26332 12384 26384 12436
rect 15752 12359 15804 12368
rect 15752 12325 15761 12359
rect 15761 12325 15795 12359
rect 15795 12325 15804 12359
rect 15752 12316 15804 12325
rect 15844 12316 15896 12368
rect 16488 12316 16540 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 6552 12291 6604 12300
rect 2780 12248 2832 12257
rect 6552 12257 6586 12291
rect 6586 12257 6604 12291
rect 6552 12248 6604 12257
rect 11244 12291 11296 12300
rect 11244 12257 11253 12291
rect 11253 12257 11287 12291
rect 11287 12257 11296 12291
rect 11244 12248 11296 12257
rect 15200 12248 15252 12300
rect 18052 12248 18104 12300
rect 19064 12316 19116 12368
rect 18972 12248 19024 12300
rect 21272 12291 21324 12300
rect 21272 12257 21281 12291
rect 21281 12257 21315 12291
rect 21315 12257 21324 12291
rect 21272 12248 21324 12257
rect 22836 12248 22888 12300
rect 23112 12291 23164 12300
rect 23112 12257 23121 12291
rect 23121 12257 23155 12291
rect 23155 12257 23164 12291
rect 23112 12248 23164 12257
rect 24308 12248 24360 12300
rect 26608 12316 26660 12368
rect 25412 12248 25464 12300
rect 2136 12223 2188 12232
rect 2136 12189 2145 12223
rect 2145 12189 2179 12223
rect 2179 12189 2188 12223
rect 2136 12180 2188 12189
rect 2412 12180 2464 12232
rect 5172 12180 5224 12232
rect 5540 12180 5592 12232
rect 10784 12180 10836 12232
rect 12348 12180 12400 12232
rect 15016 12180 15068 12232
rect 15384 12180 15436 12232
rect 15476 12180 15528 12232
rect 21364 12223 21416 12232
rect 21364 12189 21373 12223
rect 21373 12189 21407 12223
rect 21407 12189 21416 12223
rect 21364 12180 21416 12189
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 23388 12223 23440 12232
rect 21456 12180 21508 12189
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 24860 12223 24912 12232
rect 24860 12189 24869 12223
rect 24869 12189 24903 12223
rect 24903 12189 24912 12223
rect 27160 12223 27212 12232
rect 24860 12180 24912 12189
rect 27160 12189 27169 12223
rect 27169 12189 27203 12223
rect 27203 12189 27212 12223
rect 27160 12180 27212 12189
rect 2688 12112 2740 12164
rect 19708 12155 19760 12164
rect 19708 12121 19717 12155
rect 19717 12121 19751 12155
rect 19751 12121 19760 12155
rect 19708 12112 19760 12121
rect 24584 12112 24636 12164
rect 26148 12112 26200 12164
rect 3056 12044 3108 12096
rect 3884 12044 3936 12096
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 10048 12044 10100 12096
rect 15292 12087 15344 12096
rect 15292 12053 15301 12087
rect 15301 12053 15335 12087
rect 15335 12053 15344 12087
rect 15292 12044 15344 12053
rect 16304 12087 16356 12096
rect 16304 12053 16313 12087
rect 16313 12053 16347 12087
rect 16347 12053 16356 12087
rect 16304 12044 16356 12053
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 20904 12087 20956 12096
rect 20904 12053 20913 12087
rect 20913 12053 20947 12087
rect 20947 12053 20956 12087
rect 20904 12044 20956 12053
rect 22008 12087 22060 12096
rect 22008 12053 22017 12087
rect 22017 12053 22051 12087
rect 22051 12053 22060 12087
rect 22008 12044 22060 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 7656 11883 7708 11892
rect 7656 11849 7665 11883
rect 7665 11849 7699 11883
rect 7699 11849 7708 11883
rect 7656 11840 7708 11849
rect 8484 11840 8536 11892
rect 9956 11840 10008 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14832 11840 14884 11892
rect 19524 11840 19576 11892
rect 21272 11840 21324 11892
rect 23112 11840 23164 11892
rect 4252 11704 4304 11756
rect 5080 11704 5132 11756
rect 6460 11704 6512 11756
rect 8208 11772 8260 11824
rect 21916 11772 21968 11824
rect 24676 11840 24728 11892
rect 24860 11840 24912 11892
rect 11244 11747 11296 11756
rect 11244 11713 11253 11747
rect 11253 11713 11287 11747
rect 11287 11713 11296 11747
rect 11244 11704 11296 11713
rect 16396 11747 16448 11756
rect 16396 11713 16405 11747
rect 16405 11713 16439 11747
rect 16439 11713 16448 11747
rect 16396 11704 16448 11713
rect 19708 11704 19760 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 20720 11704 20772 11756
rect 22008 11747 22060 11756
rect 5172 11679 5224 11688
rect 2044 11568 2096 11620
rect 5172 11645 5181 11679
rect 5181 11645 5215 11679
rect 5215 11645 5224 11679
rect 5172 11636 5224 11645
rect 6552 11636 6604 11688
rect 7748 11636 7800 11688
rect 8208 11679 8260 11688
rect 8208 11645 8217 11679
rect 8217 11645 8251 11679
rect 8251 11645 8260 11679
rect 8208 11636 8260 11645
rect 10048 11679 10100 11688
rect 10048 11645 10057 11679
rect 10057 11645 10091 11679
rect 10091 11645 10100 11679
rect 10048 11636 10100 11645
rect 13820 11636 13872 11688
rect 15660 11636 15712 11688
rect 16304 11636 16356 11688
rect 18972 11636 19024 11688
rect 20352 11636 20404 11688
rect 20904 11636 20956 11688
rect 22008 11713 22017 11747
rect 22017 11713 22051 11747
rect 22051 11713 22060 11747
rect 22008 11704 22060 11713
rect 24308 11747 24360 11756
rect 24308 11713 24317 11747
rect 24317 11713 24351 11747
rect 24351 11713 24360 11747
rect 24308 11704 24360 11713
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 25780 11840 25832 11892
rect 25412 11772 25464 11824
rect 27160 11772 27212 11824
rect 25688 11636 25740 11688
rect 26516 11679 26568 11688
rect 26516 11645 26525 11679
rect 26525 11645 26559 11679
rect 26559 11645 26568 11679
rect 26516 11636 26568 11645
rect 2780 11568 2832 11620
rect 5264 11611 5316 11620
rect 5264 11577 5273 11611
rect 5273 11577 5307 11611
rect 5307 11577 5316 11611
rect 5264 11568 5316 11577
rect 10600 11568 10652 11620
rect 15200 11568 15252 11620
rect 18144 11568 18196 11620
rect 21732 11568 21784 11620
rect 24952 11611 25004 11620
rect 24952 11577 24961 11611
rect 24961 11577 24995 11611
rect 24995 11577 25004 11611
rect 24952 11568 25004 11577
rect 26148 11568 26200 11620
rect 3056 11543 3108 11552
rect 3056 11509 3065 11543
rect 3065 11509 3099 11543
rect 3099 11509 3108 11543
rect 3056 11500 3108 11509
rect 4252 11543 4304 11552
rect 4252 11509 4261 11543
rect 4261 11509 4295 11543
rect 4295 11509 4304 11543
rect 4252 11500 4304 11509
rect 4804 11543 4856 11552
rect 4804 11509 4813 11543
rect 4813 11509 4847 11543
rect 4847 11509 4856 11543
rect 4804 11500 4856 11509
rect 5540 11500 5592 11552
rect 7380 11543 7432 11552
rect 7380 11509 7389 11543
rect 7389 11509 7423 11543
rect 7423 11509 7432 11543
rect 7380 11500 7432 11509
rect 7840 11543 7892 11552
rect 7840 11509 7849 11543
rect 7849 11509 7883 11543
rect 7883 11509 7892 11543
rect 7840 11500 7892 11509
rect 10784 11500 10836 11552
rect 12348 11500 12400 11552
rect 15384 11500 15436 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 18328 11543 18380 11552
rect 18328 11509 18337 11543
rect 18337 11509 18371 11543
rect 18371 11509 18380 11543
rect 18328 11500 18380 11509
rect 18788 11543 18840 11552
rect 18788 11509 18797 11543
rect 18797 11509 18831 11543
rect 18831 11509 18840 11543
rect 18788 11500 18840 11509
rect 20076 11500 20128 11552
rect 20168 11500 20220 11552
rect 22836 11500 22888 11552
rect 23388 11543 23440 11552
rect 23388 11509 23397 11543
rect 23397 11509 23431 11543
rect 23431 11509 23440 11543
rect 23388 11500 23440 11509
rect 24768 11500 24820 11552
rect 26516 11500 26568 11552
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2412 11339 2464 11348
rect 2044 11296 2096 11305
rect 2412 11305 2421 11339
rect 2421 11305 2455 11339
rect 2455 11305 2464 11339
rect 2412 11296 2464 11305
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 4804 11296 4856 11348
rect 7380 11296 7432 11348
rect 10048 11296 10100 11348
rect 10600 11339 10652 11348
rect 10600 11305 10609 11339
rect 10609 11305 10643 11339
rect 10643 11305 10652 11339
rect 10600 11296 10652 11305
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18328 11296 18380 11348
rect 20168 11296 20220 11348
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 21364 11339 21416 11348
rect 21364 11305 21373 11339
rect 21373 11305 21407 11339
rect 21407 11305 21416 11339
rect 21364 11296 21416 11305
rect 22836 11339 22888 11348
rect 22836 11305 22845 11339
rect 22845 11305 22879 11339
rect 22879 11305 22888 11339
rect 22836 11296 22888 11305
rect 23204 11339 23256 11348
rect 23204 11305 23213 11339
rect 23213 11305 23247 11339
rect 23247 11305 23256 11339
rect 23204 11296 23256 11305
rect 24952 11339 25004 11348
rect 24952 11305 24961 11339
rect 24961 11305 24995 11339
rect 24995 11305 25004 11339
rect 24952 11296 25004 11305
rect 25688 11296 25740 11348
rect 26700 11339 26752 11348
rect 26700 11305 26709 11339
rect 26709 11305 26743 11339
rect 26743 11305 26752 11339
rect 26700 11296 26752 11305
rect 2136 11228 2188 11280
rect 1492 11160 1544 11212
rect 2504 11203 2556 11212
rect 2504 11169 2513 11203
rect 2513 11169 2547 11203
rect 2547 11169 2556 11203
rect 9588 11228 9640 11280
rect 12256 11228 12308 11280
rect 16028 11271 16080 11280
rect 16028 11237 16037 11271
rect 16037 11237 16071 11271
rect 16071 11237 16080 11271
rect 16028 11228 16080 11237
rect 18052 11271 18104 11280
rect 18052 11237 18061 11271
rect 18061 11237 18095 11271
rect 18095 11237 18104 11271
rect 18052 11228 18104 11237
rect 21456 11228 21508 11280
rect 25044 11228 25096 11280
rect 2504 11160 2556 11169
rect 3884 11160 3936 11212
rect 5816 11160 5868 11212
rect 8208 11203 8260 11212
rect 8208 11169 8217 11203
rect 8217 11169 8251 11203
rect 8251 11169 8260 11203
rect 8208 11160 8260 11169
rect 10508 11160 10560 11212
rect 10876 11160 10928 11212
rect 12992 11160 13044 11212
rect 15844 11160 15896 11212
rect 16304 11160 16356 11212
rect 17960 11160 18012 11212
rect 21364 11160 21416 11212
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 6276 11135 6328 11144
rect 1584 11067 1636 11076
rect 1584 11033 1593 11067
rect 1593 11033 1627 11067
rect 1627 11033 1636 11067
rect 1584 11024 1636 11033
rect 4344 11024 4396 11076
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 8024 11092 8076 11144
rect 8484 11135 8536 11144
rect 8484 11101 8493 11135
rect 8493 11101 8527 11135
rect 8527 11101 8536 11135
rect 8484 11092 8536 11101
rect 11060 11135 11112 11144
rect 11060 11101 11069 11135
rect 11069 11101 11103 11135
rect 11103 11101 11112 11135
rect 11060 11092 11112 11101
rect 12900 11135 12952 11144
rect 7748 11024 7800 11076
rect 10600 11024 10652 11076
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 12348 11024 12400 11076
rect 16396 11092 16448 11144
rect 18604 11135 18656 11144
rect 18604 11101 18613 11135
rect 18613 11101 18647 11135
rect 18647 11101 18656 11135
rect 18604 11092 18656 11101
rect 18972 11092 19024 11144
rect 20812 11092 20864 11144
rect 21824 11135 21876 11144
rect 21824 11101 21833 11135
rect 21833 11101 21867 11135
rect 21867 11101 21876 11135
rect 21824 11092 21876 11101
rect 22008 11135 22060 11144
rect 22008 11101 22017 11135
rect 22017 11101 22051 11135
rect 22051 11101 22060 11135
rect 22008 11092 22060 11101
rect 4896 10956 4948 11008
rect 8668 10956 8720 11008
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14280 10956 14332 10965
rect 14740 10956 14792 11008
rect 20720 11024 20772 11076
rect 25136 11024 25188 11076
rect 26148 11067 26200 11076
rect 26148 11033 26157 11067
rect 26157 11033 26191 11067
rect 26191 11033 26200 11067
rect 26148 11024 26200 11033
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 16580 10956 16632 11008
rect 17868 10956 17920 11008
rect 19156 10999 19208 11008
rect 19156 10965 19165 10999
rect 19165 10965 19199 10999
rect 19199 10965 19208 10999
rect 19156 10956 19208 10965
rect 24216 10956 24268 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 1492 10752 1544 10804
rect 5080 10752 5132 10804
rect 5724 10752 5776 10804
rect 6460 10752 6512 10804
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 12900 10752 12952 10804
rect 13268 10795 13320 10804
rect 13268 10761 13277 10795
rect 13277 10761 13311 10795
rect 13311 10761 13320 10795
rect 13268 10752 13320 10761
rect 15844 10752 15896 10804
rect 16304 10795 16356 10804
rect 16304 10761 16313 10795
rect 16313 10761 16347 10795
rect 16347 10761 16356 10795
rect 16304 10752 16356 10761
rect 5908 10727 5960 10736
rect 5908 10693 5917 10727
rect 5917 10693 5951 10727
rect 5951 10693 5960 10727
rect 5908 10684 5960 10693
rect 7932 10684 7984 10736
rect 8300 10684 8352 10736
rect 12992 10727 13044 10736
rect 12992 10693 13001 10727
rect 13001 10693 13035 10727
rect 13035 10693 13044 10727
rect 14740 10727 14792 10736
rect 12992 10684 13044 10693
rect 14740 10693 14749 10727
rect 14749 10693 14783 10727
rect 14783 10693 14792 10727
rect 14740 10684 14792 10693
rect 3976 10616 4028 10668
rect 7564 10616 7616 10668
rect 2688 10548 2740 10600
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 7656 10548 7708 10600
rect 8392 10616 8444 10668
rect 8668 10659 8720 10668
rect 8668 10625 8677 10659
rect 8677 10625 8711 10659
rect 8711 10625 8720 10659
rect 8668 10616 8720 10625
rect 8944 10616 8996 10668
rect 9864 10616 9916 10668
rect 14280 10616 14332 10668
rect 15476 10659 15528 10668
rect 15476 10625 15485 10659
rect 15485 10625 15519 10659
rect 15519 10625 15528 10659
rect 15476 10616 15528 10625
rect 18788 10752 18840 10804
rect 18604 10684 18656 10736
rect 18972 10659 19024 10668
rect 18972 10625 18981 10659
rect 18981 10625 19015 10659
rect 19015 10625 19024 10659
rect 22008 10752 22060 10804
rect 22284 10795 22336 10804
rect 22284 10761 22293 10795
rect 22293 10761 22327 10795
rect 22327 10761 22336 10795
rect 22284 10752 22336 10761
rect 26516 10752 26568 10804
rect 21364 10727 21416 10736
rect 21364 10693 21373 10727
rect 21373 10693 21407 10727
rect 21407 10693 21416 10727
rect 21364 10684 21416 10693
rect 21732 10659 21784 10668
rect 18972 10616 19024 10625
rect 21732 10625 21741 10659
rect 21741 10625 21775 10659
rect 21775 10625 21784 10659
rect 21732 10616 21784 10625
rect 24584 10616 24636 10668
rect 15568 10548 15620 10600
rect 18604 10548 18656 10600
rect 19156 10548 19208 10600
rect 26424 10591 26476 10600
rect 2136 10480 2188 10532
rect 3056 10480 3108 10532
rect 4160 10480 4212 10532
rect 4988 10523 5040 10532
rect 4988 10489 4997 10523
rect 4997 10489 5031 10523
rect 5031 10489 5040 10523
rect 4988 10480 5040 10489
rect 8024 10480 8076 10532
rect 8576 10523 8628 10532
rect 8576 10489 8585 10523
rect 8585 10489 8619 10523
rect 8619 10489 8628 10523
rect 8576 10480 8628 10489
rect 11060 10480 11112 10532
rect 15384 10523 15436 10532
rect 15384 10489 15393 10523
rect 15393 10489 15427 10523
rect 15427 10489 15436 10523
rect 15384 10480 15436 10489
rect 26424 10557 26433 10591
rect 26433 10557 26467 10591
rect 26467 10557 26476 10591
rect 26424 10548 26476 10557
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 24308 10523 24360 10532
rect 24308 10489 24317 10523
rect 24317 10489 24351 10523
rect 24351 10489 24360 10523
rect 24308 10480 24360 10489
rect 4528 10455 4580 10464
rect 4528 10421 4537 10455
rect 4537 10421 4571 10455
rect 4571 10421 4580 10455
rect 4528 10412 4580 10421
rect 6184 10455 6236 10464
rect 6184 10421 6193 10455
rect 6193 10421 6227 10455
rect 6227 10421 6236 10455
rect 6184 10412 6236 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 9220 10455 9272 10464
rect 9220 10421 9229 10455
rect 9229 10421 9263 10455
rect 9263 10421 9272 10455
rect 10140 10455 10192 10464
rect 9220 10412 9272 10421
rect 10140 10421 10149 10455
rect 10149 10421 10183 10455
rect 10183 10421 10192 10455
rect 10140 10412 10192 10421
rect 10232 10455 10284 10464
rect 10232 10421 10241 10455
rect 10241 10421 10275 10455
rect 10275 10421 10284 10455
rect 10876 10455 10928 10464
rect 10232 10412 10284 10421
rect 10876 10421 10885 10455
rect 10885 10421 10919 10455
rect 10919 10421 10928 10455
rect 10876 10412 10928 10421
rect 11612 10412 11664 10464
rect 14924 10455 14976 10464
rect 14924 10421 14933 10455
rect 14933 10421 14967 10455
rect 14967 10421 14976 10455
rect 14924 10412 14976 10421
rect 17868 10455 17920 10464
rect 17868 10421 17877 10455
rect 17877 10421 17911 10455
rect 17911 10421 17920 10455
rect 17868 10412 17920 10421
rect 18788 10455 18840 10464
rect 18788 10421 18797 10455
rect 18797 10421 18831 10455
rect 18831 10421 18840 10455
rect 18788 10412 18840 10421
rect 23480 10412 23532 10464
rect 24216 10455 24268 10464
rect 24216 10421 24225 10455
rect 24225 10421 24259 10455
rect 24259 10421 24268 10455
rect 24216 10412 24268 10421
rect 26608 10455 26660 10464
rect 26608 10421 26617 10455
rect 26617 10421 26651 10455
rect 26651 10421 26660 10455
rect 26608 10412 26660 10421
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 2136 10251 2188 10260
rect 2136 10217 2145 10251
rect 2145 10217 2179 10251
rect 2179 10217 2188 10251
rect 2136 10208 2188 10217
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 4344 10251 4396 10260
rect 4344 10217 4353 10251
rect 4353 10217 4387 10251
rect 4387 10217 4396 10251
rect 4344 10208 4396 10217
rect 4804 10208 4856 10260
rect 4988 10251 5040 10260
rect 4988 10217 4997 10251
rect 4997 10217 5031 10251
rect 5031 10217 5040 10251
rect 4988 10208 5040 10217
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 7748 10208 7800 10260
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 12348 10208 12400 10260
rect 15292 10208 15344 10260
rect 15660 10208 15712 10260
rect 18512 10208 18564 10260
rect 22008 10208 22060 10260
rect 24216 10208 24268 10260
rect 8300 10140 8352 10192
rect 9588 10140 9640 10192
rect 18972 10140 19024 10192
rect 23664 10140 23716 10192
rect 8944 10072 8996 10124
rect 11152 10072 11204 10124
rect 14924 10072 14976 10124
rect 15752 10072 15804 10124
rect 18052 10072 18104 10124
rect 18696 10115 18748 10124
rect 18696 10081 18705 10115
rect 18705 10081 18739 10115
rect 18739 10081 18748 10115
rect 18696 10072 18748 10081
rect 20812 10072 20864 10124
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 7472 10004 7524 10056
rect 8116 10004 8168 10056
rect 8852 10004 8904 10056
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 2412 9936 2464 9988
rect 7288 9936 7340 9988
rect 1584 9911 1636 9920
rect 1584 9877 1593 9911
rect 1593 9877 1627 9911
rect 1627 9877 1636 9911
rect 1584 9868 1636 9877
rect 2688 9868 2740 9920
rect 9864 9911 9916 9920
rect 9864 9877 9873 9911
rect 9873 9877 9907 9911
rect 9907 9877 9916 9911
rect 9864 9868 9916 9877
rect 15384 10004 15436 10056
rect 18328 10004 18380 10056
rect 11704 9868 11756 9920
rect 13728 9868 13780 9920
rect 14280 9868 14332 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 19248 9868 19300 9920
rect 23572 10004 23624 10056
rect 24216 10047 24268 10056
rect 24216 10013 24225 10047
rect 24225 10013 24259 10047
rect 24259 10013 24268 10047
rect 24216 10004 24268 10013
rect 24584 10004 24636 10056
rect 21640 9868 21692 9920
rect 23388 9868 23440 9920
rect 24860 9911 24912 9920
rect 24860 9877 24869 9911
rect 24869 9877 24903 9911
rect 24903 9877 24912 9911
rect 24860 9868 24912 9877
rect 26792 9868 26844 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 2688 9664 2740 9716
rect 3976 9707 4028 9716
rect 3976 9673 3985 9707
rect 3985 9673 4019 9707
rect 4019 9673 4028 9707
rect 3976 9664 4028 9673
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 8300 9664 8352 9716
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 15660 9707 15712 9716
rect 15660 9673 15669 9707
rect 15669 9673 15703 9707
rect 15703 9673 15712 9707
rect 15660 9664 15712 9673
rect 15752 9664 15804 9716
rect 18604 9707 18656 9716
rect 18604 9673 18613 9707
rect 18613 9673 18647 9707
rect 18647 9673 18656 9707
rect 18604 9664 18656 9673
rect 23664 9664 23716 9716
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 4068 9503 4120 9512
rect 4068 9469 4077 9503
rect 4077 9469 4111 9503
rect 4111 9469 4120 9503
rect 4068 9460 4120 9469
rect 9864 9528 9916 9580
rect 11152 9528 11204 9580
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 18420 9528 18472 9580
rect 18880 9528 18932 9580
rect 19708 9596 19760 9648
rect 19984 9639 20036 9648
rect 19984 9605 19993 9639
rect 19993 9605 20027 9639
rect 20027 9605 20036 9639
rect 19984 9596 20036 9605
rect 26516 9664 26568 9716
rect 26056 9639 26108 9648
rect 7932 9460 7984 9512
rect 9312 9503 9364 9512
rect 9312 9469 9321 9503
rect 9321 9469 9355 9503
rect 9355 9469 9364 9503
rect 9312 9460 9364 9469
rect 10048 9460 10100 9512
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 2136 9324 2188 9376
rect 5724 9324 5776 9376
rect 7288 9324 7340 9376
rect 8300 9324 8352 9376
rect 13728 9392 13780 9444
rect 17868 9392 17920 9444
rect 21916 9571 21968 9580
rect 21916 9537 21925 9571
rect 21925 9537 21959 9571
rect 21959 9537 21968 9571
rect 22652 9571 22704 9580
rect 21916 9528 21968 9537
rect 22652 9537 22661 9571
rect 22661 9537 22695 9571
rect 22695 9537 22704 9571
rect 22652 9528 22704 9537
rect 24584 9528 24636 9580
rect 26056 9605 26065 9639
rect 26065 9605 26099 9639
rect 26099 9605 26108 9639
rect 26056 9596 26108 9605
rect 27344 9639 27396 9648
rect 27344 9605 27353 9639
rect 27353 9605 27387 9639
rect 27387 9605 27396 9639
rect 27344 9596 27396 9605
rect 22100 9460 22152 9512
rect 23388 9460 23440 9512
rect 24676 9503 24728 9512
rect 24676 9469 24685 9503
rect 24685 9469 24719 9503
rect 24719 9469 24728 9503
rect 24676 9460 24728 9469
rect 19248 9392 19300 9444
rect 23480 9392 23532 9444
rect 24584 9392 24636 9444
rect 8944 9367 8996 9376
rect 8944 9333 8953 9367
rect 8953 9333 8987 9367
rect 8987 9333 8996 9367
rect 8944 9324 8996 9333
rect 11704 9324 11756 9376
rect 18420 9367 18472 9376
rect 18420 9333 18429 9367
rect 18429 9333 18463 9367
rect 18463 9333 18472 9367
rect 18420 9324 18472 9333
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 20812 9324 20864 9376
rect 22192 9324 22244 9376
rect 24216 9367 24268 9376
rect 24216 9333 24225 9367
rect 24225 9333 24259 9367
rect 24259 9333 24268 9367
rect 24216 9324 24268 9333
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 5080 9120 5132 9172
rect 7932 9120 7984 9172
rect 8944 9120 8996 9172
rect 9312 9120 9364 9172
rect 9588 9120 9640 9172
rect 11704 9120 11756 9172
rect 13268 9163 13320 9172
rect 13268 9129 13277 9163
rect 13277 9129 13311 9163
rect 13311 9129 13320 9163
rect 13268 9120 13320 9129
rect 18788 9120 18840 9172
rect 19064 9120 19116 9172
rect 22100 9163 22152 9172
rect 22100 9129 22109 9163
rect 22109 9129 22143 9163
rect 22143 9129 22152 9163
rect 26700 9163 26752 9172
rect 22100 9120 22152 9129
rect 26700 9129 26709 9163
rect 26709 9129 26743 9163
rect 26743 9129 26752 9163
rect 26700 9120 26752 9129
rect 15384 9052 15436 9104
rect 2412 8984 2464 9036
rect 5724 9027 5776 9036
rect 5724 8993 5758 9027
rect 5758 8993 5776 9027
rect 5724 8984 5776 8993
rect 7932 8984 7984 9036
rect 10048 9027 10100 9036
rect 4068 8916 4120 8968
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 8944 8916 8996 8968
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 9680 8916 9732 8968
rect 9956 8916 10008 8968
rect 18420 8984 18472 9036
rect 18696 8984 18748 9036
rect 19340 8984 19392 9036
rect 23848 9027 23900 9036
rect 23848 8993 23857 9027
rect 23857 8993 23891 9027
rect 23891 8993 23900 9027
rect 23848 8984 23900 8993
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 9864 8848 9916 8900
rect 14464 8916 14516 8968
rect 15200 8916 15252 8968
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 23940 8959 23992 8968
rect 23940 8925 23949 8959
rect 23949 8925 23983 8959
rect 23983 8925 23992 8959
rect 23940 8916 23992 8925
rect 10508 8848 10560 8900
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 6828 8823 6880 8832
rect 6828 8789 6837 8823
rect 6837 8789 6871 8823
rect 6871 8789 6880 8823
rect 6828 8780 6880 8789
rect 9128 8780 9180 8832
rect 16304 8780 16356 8832
rect 21640 8780 21692 8832
rect 23480 8823 23532 8832
rect 23480 8789 23489 8823
rect 23489 8789 23523 8823
rect 23523 8789 23532 8823
rect 23480 8780 23532 8789
rect 24584 8780 24636 8832
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 4620 8619 4672 8628
rect 4620 8585 4629 8619
rect 4629 8585 4663 8619
rect 4663 8585 4672 8619
rect 4620 8576 4672 8585
rect 7932 8576 7984 8628
rect 10508 8619 10560 8628
rect 10508 8585 10517 8619
rect 10517 8585 10551 8619
rect 10551 8585 10560 8619
rect 10508 8576 10560 8585
rect 14464 8619 14516 8628
rect 14464 8585 14473 8619
rect 14473 8585 14507 8619
rect 14507 8585 14516 8619
rect 14464 8576 14516 8585
rect 15384 8576 15436 8628
rect 18696 8619 18748 8628
rect 18696 8585 18705 8619
rect 18705 8585 18739 8619
rect 18739 8585 18748 8619
rect 18696 8576 18748 8585
rect 19064 8619 19116 8628
rect 19064 8585 19073 8619
rect 19073 8585 19107 8619
rect 19107 8585 19116 8619
rect 19064 8576 19116 8585
rect 20812 8576 20864 8628
rect 23848 8619 23900 8628
rect 23848 8585 23857 8619
rect 23857 8585 23891 8619
rect 23891 8585 23900 8619
rect 23848 8576 23900 8585
rect 1400 8508 1452 8560
rect 23296 8508 23348 8560
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 7472 8440 7524 8492
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 24584 8483 24636 8492
rect 24584 8449 24593 8483
rect 24593 8449 24627 8483
rect 24627 8449 24636 8483
rect 24584 8440 24636 8449
rect 26148 8440 26200 8492
rect 4620 8372 4672 8424
rect 9128 8415 9180 8424
rect 5080 8347 5132 8356
rect 5080 8313 5089 8347
rect 5089 8313 5123 8347
rect 5123 8313 5132 8347
rect 5080 8304 5132 8313
rect 5448 8304 5500 8356
rect 7288 8304 7340 8356
rect 4620 8236 4672 8288
rect 8300 8279 8352 8288
rect 8300 8245 8309 8279
rect 8309 8245 8343 8279
rect 8343 8245 8352 8279
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 19340 8372 19392 8424
rect 20168 8372 20220 8424
rect 24676 8372 24728 8424
rect 9220 8304 9272 8356
rect 23940 8304 23992 8356
rect 24860 8304 24912 8356
rect 26516 8304 26568 8356
rect 26976 8304 27028 8356
rect 15660 8279 15712 8288
rect 8300 8236 8352 8245
rect 15660 8245 15669 8279
rect 15669 8245 15703 8279
rect 15703 8245 15712 8279
rect 15660 8236 15712 8245
rect 16028 8279 16080 8288
rect 16028 8245 16037 8279
rect 16037 8245 16071 8279
rect 16071 8245 16080 8279
rect 16028 8236 16080 8245
rect 21640 8236 21692 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 1492 8032 1544 8084
rect 3608 8032 3660 8084
rect 4252 8032 4304 8084
rect 9220 8075 9272 8084
rect 9220 8041 9229 8075
rect 9229 8041 9263 8075
rect 9263 8041 9272 8075
rect 9220 8032 9272 8041
rect 10508 8032 10560 8084
rect 23940 8032 23992 8084
rect 24400 8032 24452 8084
rect 24952 8032 25004 8084
rect 25872 8032 25924 8084
rect 26700 8075 26752 8084
rect 26700 8041 26709 8075
rect 26709 8041 26743 8075
rect 26743 8041 26752 8075
rect 26700 8032 26752 8041
rect 16212 7964 16264 8016
rect 21456 7964 21508 8016
rect 21916 7964 21968 8016
rect 24584 7964 24636 8016
rect 1952 7896 2004 7948
rect 11980 7939 12032 7948
rect 11980 7905 12014 7939
rect 12014 7905 12032 7939
rect 11980 7896 12032 7905
rect 15200 7896 15252 7948
rect 15752 7896 15804 7948
rect 18604 7896 18656 7948
rect 19248 7896 19300 7948
rect 21640 7896 21692 7948
rect 26516 7939 26568 7948
rect 26516 7905 26525 7939
rect 26525 7905 26559 7939
rect 26559 7905 26568 7939
rect 26516 7896 26568 7905
rect 4344 7828 4396 7880
rect 4620 7871 4672 7880
rect 4620 7837 4629 7871
rect 4629 7837 4663 7871
rect 4663 7837 4672 7871
rect 4620 7828 4672 7837
rect 4804 7871 4856 7880
rect 4804 7837 4813 7871
rect 4813 7837 4847 7871
rect 4847 7837 4856 7871
rect 4804 7828 4856 7837
rect 5540 7828 5592 7880
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 24124 7828 24176 7880
rect 1860 7692 1912 7744
rect 3884 7692 3936 7744
rect 4160 7735 4212 7744
rect 4160 7701 4169 7735
rect 4169 7701 4203 7735
rect 4203 7701 4212 7735
rect 4160 7692 4212 7701
rect 9956 7735 10008 7744
rect 9956 7701 9965 7735
rect 9965 7701 9999 7735
rect 9999 7701 10008 7735
rect 9956 7692 10008 7701
rect 12440 7692 12492 7744
rect 16028 7760 16080 7812
rect 18512 7803 18564 7812
rect 18512 7769 18521 7803
rect 18521 7769 18555 7803
rect 18555 7769 18564 7803
rect 18512 7760 18564 7769
rect 19524 7760 19576 7812
rect 13084 7735 13136 7744
rect 13084 7701 13093 7735
rect 13093 7701 13127 7735
rect 13127 7701 13136 7735
rect 13084 7692 13136 7701
rect 17408 7735 17460 7744
rect 17408 7701 17417 7735
rect 17417 7701 17451 7735
rect 17451 7701 17460 7735
rect 17408 7692 17460 7701
rect 22376 7735 22428 7744
rect 22376 7701 22385 7735
rect 22385 7701 22419 7735
rect 22419 7701 22428 7735
rect 22376 7692 22428 7701
rect 25412 7735 25464 7744
rect 25412 7701 25421 7735
rect 25421 7701 25455 7735
rect 25455 7701 25464 7735
rect 25412 7692 25464 7701
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 9220 7488 9272 7540
rect 9680 7531 9732 7540
rect 9680 7497 9689 7531
rect 9689 7497 9723 7531
rect 9723 7497 9732 7531
rect 9680 7488 9732 7497
rect 15660 7488 15712 7540
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4804 7352 4856 7404
rect 6828 7352 6880 7404
rect 8300 7395 8352 7404
rect 8300 7361 8309 7395
rect 8309 7361 8343 7395
rect 8343 7361 8352 7395
rect 8300 7352 8352 7361
rect 1860 7327 1912 7336
rect 1860 7293 1894 7327
rect 1894 7293 1912 7327
rect 1860 7284 1912 7293
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 2688 7216 2740 7268
rect 5080 7259 5132 7268
rect 5080 7225 5089 7259
rect 5089 7225 5123 7259
rect 5123 7225 5132 7259
rect 5080 7216 5132 7225
rect 9864 7216 9916 7268
rect 1860 7148 1912 7200
rect 2780 7148 2832 7200
rect 5172 7191 5224 7200
rect 5172 7157 5181 7191
rect 5181 7157 5215 7191
rect 5215 7157 5224 7191
rect 5172 7148 5224 7157
rect 5632 7191 5684 7200
rect 5632 7157 5641 7191
rect 5641 7157 5675 7191
rect 5675 7157 5684 7191
rect 5632 7148 5684 7157
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11980 7352 12032 7404
rect 13268 7395 13320 7404
rect 13268 7361 13277 7395
rect 13277 7361 13311 7395
rect 13311 7361 13320 7395
rect 13268 7352 13320 7361
rect 16304 7488 16356 7540
rect 18604 7531 18656 7540
rect 18604 7497 18613 7531
rect 18613 7497 18647 7531
rect 18647 7497 18656 7531
rect 18604 7488 18656 7497
rect 20812 7488 20864 7540
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 23572 7488 23624 7540
rect 24400 7488 24452 7540
rect 24676 7488 24728 7540
rect 26332 7488 26384 7540
rect 13176 7284 13228 7336
rect 15384 7284 15436 7336
rect 17408 7352 17460 7404
rect 19524 7327 19576 7336
rect 19524 7293 19533 7327
rect 19533 7293 19567 7327
rect 19567 7293 19576 7327
rect 19524 7284 19576 7293
rect 12164 7259 12216 7268
rect 12164 7225 12173 7259
rect 12173 7225 12207 7259
rect 12207 7225 12216 7259
rect 12164 7216 12216 7225
rect 15568 7259 15620 7268
rect 15568 7225 15577 7259
rect 15577 7225 15611 7259
rect 15611 7225 15620 7259
rect 15568 7216 15620 7225
rect 16396 7216 16448 7268
rect 22376 7352 22428 7404
rect 24308 7352 24360 7404
rect 22192 7216 22244 7268
rect 25780 7420 25832 7472
rect 25412 7352 25464 7404
rect 24952 7327 25004 7336
rect 24952 7293 24961 7327
rect 24961 7293 24995 7327
rect 24995 7293 25004 7327
rect 24952 7284 25004 7293
rect 25044 7259 25096 7268
rect 25044 7225 25053 7259
rect 25053 7225 25087 7259
rect 25087 7225 25096 7259
rect 25044 7216 25096 7225
rect 25872 7352 25924 7404
rect 11428 7148 11480 7157
rect 12624 7191 12676 7200
rect 12624 7157 12633 7191
rect 12633 7157 12667 7191
rect 12667 7157 12676 7191
rect 12624 7148 12676 7157
rect 14188 7191 14240 7200
rect 14188 7157 14197 7191
rect 14197 7157 14231 7191
rect 14231 7157 14240 7191
rect 14188 7148 14240 7157
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 17592 7148 17644 7200
rect 20260 7148 20312 7200
rect 22468 7191 22520 7200
rect 22468 7157 22477 7191
rect 22477 7157 22511 7191
rect 22511 7157 22520 7191
rect 22468 7148 22520 7157
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 25688 7191 25740 7200
rect 25688 7157 25697 7191
rect 25697 7157 25731 7191
rect 25731 7157 25740 7191
rect 25688 7148 25740 7157
rect 25964 7191 26016 7200
rect 25964 7157 25973 7191
rect 25973 7157 26007 7191
rect 26007 7157 26016 7191
rect 25964 7148 26016 7157
rect 26516 7148 26568 7200
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 1952 6987 2004 6996
rect 1952 6953 1961 6987
rect 1961 6953 1995 6987
rect 1995 6953 2004 6987
rect 1952 6944 2004 6953
rect 2688 6944 2740 6996
rect 3424 6944 3476 6996
rect 5724 6944 5776 6996
rect 6184 6987 6236 6996
rect 6184 6953 6193 6987
rect 6193 6953 6227 6987
rect 6227 6953 6236 6987
rect 6184 6944 6236 6953
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 11704 6987 11756 6996
rect 8300 6944 8352 6953
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 13176 6944 13228 6996
rect 14188 6944 14240 6996
rect 15752 6944 15804 6996
rect 19524 6987 19576 6996
rect 19524 6953 19533 6987
rect 19533 6953 19567 6987
rect 19567 6953 19576 6987
rect 19524 6944 19576 6953
rect 22468 6944 22520 6996
rect 23388 6944 23440 6996
rect 25504 6944 25556 6996
rect 1768 6808 1820 6860
rect 4344 6876 4396 6928
rect 5080 6876 5132 6928
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 9496 6808 9548 6860
rect 4344 6740 4396 6792
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 6828 6740 6880 6792
rect 9680 6740 9732 6792
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 1584 6715 1636 6724
rect 1584 6681 1593 6715
rect 1593 6681 1627 6715
rect 1627 6681 1636 6715
rect 1584 6672 1636 6681
rect 12072 6808 12124 6860
rect 12256 6851 12308 6860
rect 12256 6817 12265 6851
rect 12265 6817 12299 6851
rect 12299 6817 12308 6851
rect 12256 6808 12308 6817
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 13084 6876 13136 6928
rect 13268 6876 13320 6928
rect 21456 6876 21508 6928
rect 22192 6876 22244 6928
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 17592 6808 17644 6860
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 22100 6808 22152 6860
rect 23296 6808 23348 6860
rect 24676 6851 24728 6860
rect 24676 6817 24685 6851
rect 24685 6817 24719 6851
rect 24719 6817 24728 6851
rect 24952 6876 25004 6928
rect 24676 6808 24728 6817
rect 26608 6808 26660 6860
rect 14464 6740 14516 6792
rect 17684 6740 17736 6792
rect 17408 6672 17460 6724
rect 22652 6740 22704 6792
rect 24952 6740 25004 6792
rect 25688 6740 25740 6792
rect 18328 6672 18380 6724
rect 24860 6715 24912 6724
rect 24860 6681 24869 6715
rect 24869 6681 24903 6715
rect 24903 6681 24912 6715
rect 24860 6672 24912 6681
rect 4620 6604 4672 6656
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 7932 6604 7984 6656
rect 9772 6604 9824 6656
rect 12256 6604 12308 6656
rect 15384 6604 15436 6656
rect 16856 6604 16908 6656
rect 17500 6647 17552 6656
rect 17500 6613 17509 6647
rect 17509 6613 17543 6647
rect 17543 6613 17552 6647
rect 17500 6604 17552 6613
rect 20444 6604 20496 6656
rect 21640 6604 21692 6656
rect 26700 6715 26752 6724
rect 26700 6681 26709 6715
rect 26709 6681 26743 6715
rect 26743 6681 26752 6715
rect 26700 6672 26752 6681
rect 26332 6604 26384 6656
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1768 6400 1820 6452
rect 4804 6400 4856 6452
rect 5724 6400 5776 6452
rect 6276 6443 6328 6452
rect 6276 6409 6285 6443
rect 6285 6409 6319 6443
rect 6319 6409 6328 6443
rect 6276 6400 6328 6409
rect 6828 6400 6880 6452
rect 7380 6443 7432 6452
rect 7380 6409 7389 6443
rect 7389 6409 7423 6443
rect 7423 6409 7432 6443
rect 7380 6400 7432 6409
rect 10140 6400 10192 6452
rect 12256 6400 12308 6452
rect 12348 6400 12400 6452
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 14188 6400 14240 6452
rect 17776 6443 17828 6452
rect 17776 6409 17785 6443
rect 17785 6409 17819 6443
rect 17819 6409 17828 6443
rect 17776 6400 17828 6409
rect 22100 6400 22152 6452
rect 22652 6443 22704 6452
rect 22652 6409 22661 6443
rect 22661 6409 22695 6443
rect 22695 6409 22704 6443
rect 22652 6400 22704 6409
rect 23296 6400 23348 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 24860 6443 24912 6452
rect 24860 6409 24869 6443
rect 24869 6409 24903 6443
rect 24903 6409 24912 6443
rect 24860 6400 24912 6409
rect 25504 6400 25556 6452
rect 26332 6400 26384 6452
rect 26608 6400 26660 6452
rect 3700 6332 3752 6384
rect 5080 6332 5132 6384
rect 9680 6375 9732 6384
rect 9680 6341 9689 6375
rect 9689 6341 9723 6375
rect 9723 6341 9732 6375
rect 9680 6332 9732 6341
rect 4160 6264 4212 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 5264 6307 5316 6316
rect 4804 6264 4856 6273
rect 5264 6273 5273 6307
rect 5273 6273 5307 6307
rect 5307 6273 5316 6307
rect 5264 6264 5316 6273
rect 8116 6307 8168 6316
rect 8116 6273 8125 6307
rect 8125 6273 8159 6307
rect 8159 6273 8168 6307
rect 8116 6264 8168 6273
rect 9864 6264 9916 6316
rect 12072 6264 12124 6316
rect 17684 6332 17736 6384
rect 16948 6307 17000 6316
rect 16948 6273 16957 6307
rect 16957 6273 16991 6307
rect 16991 6273 17000 6307
rect 16948 6264 17000 6273
rect 18328 6264 18380 6316
rect 20444 6307 20496 6316
rect 20444 6273 20453 6307
rect 20453 6273 20487 6307
rect 20487 6273 20496 6307
rect 20444 6264 20496 6273
rect 1860 6196 1912 6248
rect 7380 6196 7432 6248
rect 12256 6196 12308 6248
rect 13912 6196 13964 6248
rect 17500 6196 17552 6248
rect 17776 6196 17828 6248
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 19984 6196 20036 6248
rect 2044 6171 2096 6180
rect 2044 6137 2078 6171
rect 2078 6137 2096 6171
rect 2044 6128 2096 6137
rect 2688 6128 2740 6180
rect 10784 6128 10836 6180
rect 16488 6128 16540 6180
rect 16948 6128 17000 6180
rect 20536 6128 20588 6180
rect 26240 6171 26292 6180
rect 26240 6137 26249 6171
rect 26249 6137 26283 6171
rect 26283 6137 26292 6171
rect 26240 6128 26292 6137
rect 2964 6060 3016 6112
rect 4252 6103 4304 6112
rect 4252 6069 4261 6103
rect 4261 6069 4295 6103
rect 4295 6069 4304 6103
rect 4252 6060 4304 6069
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 7196 6060 7248 6112
rect 7748 6060 7800 6112
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 14464 6060 14516 6112
rect 16580 6060 16632 6112
rect 16856 6103 16908 6112
rect 16856 6069 16865 6103
rect 16865 6069 16899 6103
rect 16899 6069 16908 6103
rect 16856 6060 16908 6069
rect 20720 6060 20772 6112
rect 26608 6103 26660 6112
rect 26608 6069 26617 6103
rect 26617 6069 26651 6103
rect 26651 6069 26660 6103
rect 26608 6060 26660 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2044 5899 2096 5908
rect 2044 5865 2053 5899
rect 2053 5865 2087 5899
rect 2087 5865 2096 5899
rect 2044 5856 2096 5865
rect 2780 5856 2832 5908
rect 4620 5856 4672 5908
rect 5448 5856 5500 5908
rect 5816 5856 5868 5908
rect 9496 5899 9548 5908
rect 9496 5865 9505 5899
rect 9505 5865 9539 5899
rect 9539 5865 9548 5899
rect 9496 5856 9548 5865
rect 9864 5856 9916 5908
rect 12440 5856 12492 5908
rect 12716 5899 12768 5908
rect 12716 5865 12725 5899
rect 12725 5865 12759 5899
rect 12759 5865 12768 5899
rect 12716 5856 12768 5865
rect 17592 5899 17644 5908
rect 17592 5865 17601 5899
rect 17601 5865 17635 5899
rect 17635 5865 17644 5899
rect 17592 5856 17644 5865
rect 18236 5899 18288 5908
rect 18236 5865 18245 5899
rect 18245 5865 18279 5899
rect 18279 5865 18288 5899
rect 18236 5856 18288 5865
rect 20444 5856 20496 5908
rect 21732 5856 21784 5908
rect 26976 5856 27028 5908
rect 4160 5788 4212 5840
rect 5172 5788 5224 5840
rect 11152 5831 11204 5840
rect 11152 5797 11161 5831
rect 11161 5797 11195 5831
rect 11195 5797 11204 5831
rect 11152 5788 11204 5797
rect 15016 5788 15068 5840
rect 2412 5720 2464 5772
rect 7932 5763 7984 5772
rect 7932 5729 7941 5763
rect 7941 5729 7975 5763
rect 7975 5729 7984 5763
rect 7932 5720 7984 5729
rect 11704 5720 11756 5772
rect 13084 5720 13136 5772
rect 15752 5788 15804 5840
rect 17868 5788 17920 5840
rect 17960 5788 18012 5840
rect 24124 5788 24176 5840
rect 15384 5720 15436 5772
rect 1860 5652 1912 5704
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 8024 5695 8076 5704
rect 8024 5661 8033 5695
rect 8033 5661 8067 5695
rect 8067 5661 8076 5695
rect 8024 5652 8076 5661
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 11336 5695 11388 5704
rect 8116 5652 8168 5661
rect 11336 5661 11345 5695
rect 11345 5661 11379 5695
rect 11379 5661 11388 5695
rect 11336 5652 11388 5661
rect 12716 5652 12768 5704
rect 1584 5627 1636 5636
rect 1584 5593 1593 5627
rect 1593 5593 1627 5627
rect 1627 5593 1636 5627
rect 1584 5584 1636 5593
rect 10784 5627 10836 5636
rect 10784 5593 10793 5627
rect 10793 5593 10827 5627
rect 10827 5593 10836 5627
rect 10784 5584 10836 5593
rect 4344 5559 4396 5568
rect 4344 5525 4353 5559
rect 4353 5525 4387 5559
rect 4387 5525 4396 5559
rect 4344 5516 4396 5525
rect 4436 5516 4488 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 7564 5559 7616 5568
rect 7564 5525 7573 5559
rect 7573 5525 7607 5559
rect 7607 5525 7616 5559
rect 7564 5516 7616 5525
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 19800 5695 19852 5704
rect 19800 5661 19809 5695
rect 19809 5661 19843 5695
rect 19843 5661 19852 5695
rect 19800 5652 19852 5661
rect 20628 5652 20680 5704
rect 25320 5763 25372 5772
rect 25320 5729 25329 5763
rect 25329 5729 25363 5763
rect 25363 5729 25372 5763
rect 25320 5720 25372 5729
rect 27160 5720 27212 5772
rect 21640 5652 21692 5704
rect 22100 5652 22152 5704
rect 25504 5627 25556 5636
rect 13544 5516 13596 5568
rect 16488 5516 16540 5568
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 20444 5516 20496 5568
rect 25504 5593 25513 5627
rect 25513 5593 25547 5627
rect 25547 5593 25556 5627
rect 25504 5584 25556 5593
rect 23572 5516 23624 5568
rect 26700 5559 26752 5568
rect 26700 5525 26709 5559
rect 26709 5525 26743 5559
rect 26743 5525 26752 5559
rect 26700 5516 26752 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 2412 5355 2464 5364
rect 2412 5321 2421 5355
rect 2421 5321 2455 5355
rect 2455 5321 2464 5355
rect 2412 5312 2464 5321
rect 2964 5355 3016 5364
rect 2964 5321 2973 5355
rect 2973 5321 3007 5355
rect 3007 5321 3016 5355
rect 2964 5312 3016 5321
rect 5264 5312 5316 5364
rect 5448 5355 5500 5364
rect 5448 5321 5457 5355
rect 5457 5321 5491 5355
rect 5491 5321 5500 5355
rect 5448 5312 5500 5321
rect 7932 5312 7984 5364
rect 10508 5312 10560 5364
rect 14464 5355 14516 5364
rect 14464 5321 14473 5355
rect 14473 5321 14507 5355
rect 14507 5321 14516 5355
rect 14464 5312 14516 5321
rect 15384 5355 15436 5364
rect 15384 5321 15393 5355
rect 15393 5321 15427 5355
rect 15427 5321 15436 5355
rect 15384 5312 15436 5321
rect 17868 5355 17920 5364
rect 17868 5321 17877 5355
rect 17877 5321 17911 5355
rect 17911 5321 17920 5355
rect 17868 5312 17920 5321
rect 17960 5312 18012 5364
rect 18236 5355 18288 5364
rect 18236 5321 18245 5355
rect 18245 5321 18279 5355
rect 18279 5321 18288 5355
rect 18236 5312 18288 5321
rect 18328 5312 18380 5364
rect 20352 5355 20404 5364
rect 20352 5321 20361 5355
rect 20361 5321 20395 5355
rect 20395 5321 20404 5355
rect 20352 5312 20404 5321
rect 20536 5355 20588 5364
rect 20536 5321 20545 5355
rect 20545 5321 20579 5355
rect 20579 5321 20588 5355
rect 20536 5312 20588 5321
rect 21732 5312 21784 5364
rect 25228 5312 25280 5364
rect 26332 5312 26384 5364
rect 27160 5355 27212 5364
rect 27160 5321 27169 5355
rect 27169 5321 27203 5355
rect 27203 5321 27212 5355
rect 27160 5312 27212 5321
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 11152 5244 11204 5296
rect 16488 5244 16540 5296
rect 9680 5219 9732 5228
rect 2780 5108 2832 5160
rect 9680 5185 9689 5219
rect 9689 5185 9723 5219
rect 9723 5185 9732 5219
rect 9680 5176 9732 5185
rect 10784 5176 10836 5228
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 15660 5176 15712 5228
rect 20444 5176 20496 5228
rect 3700 5108 3752 5160
rect 7288 5108 7340 5160
rect 17776 5108 17828 5160
rect 20352 5108 20404 5160
rect 8116 5040 8168 5092
rect 13544 5040 13596 5092
rect 16488 5040 16540 5092
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 4620 4972 4672 5024
rect 7196 4972 7248 5024
rect 7656 4972 7708 5024
rect 10784 4972 10836 5024
rect 11336 4972 11388 5024
rect 11888 5015 11940 5024
rect 11888 4981 11897 5015
rect 11897 4981 11931 5015
rect 11931 4981 11940 5015
rect 11888 4972 11940 4981
rect 11980 4972 12032 5024
rect 12440 4972 12492 5024
rect 12716 5015 12768 5024
rect 12716 4981 12725 5015
rect 12725 4981 12759 5015
rect 12759 4981 12768 5015
rect 12716 4972 12768 4981
rect 16304 4972 16356 5024
rect 19524 4972 19576 5024
rect 20628 5040 20680 5092
rect 25228 5151 25280 5160
rect 25228 5117 25237 5151
rect 25237 5117 25271 5151
rect 25271 5117 25280 5151
rect 25228 5108 25280 5117
rect 21916 5083 21968 5092
rect 21916 5049 21925 5083
rect 21925 5049 21959 5083
rect 21959 5049 21968 5083
rect 21916 5040 21968 5049
rect 20536 4972 20588 5024
rect 22928 5015 22980 5024
rect 22928 4981 22937 5015
rect 22937 4981 22971 5015
rect 22971 4981 22980 5015
rect 22928 4972 22980 4981
rect 24860 4972 24912 5024
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 2780 4768 2832 4820
rect 4160 4768 4212 4820
rect 4252 4768 4304 4820
rect 5172 4811 5224 4820
rect 5172 4777 5181 4811
rect 5181 4777 5215 4811
rect 5215 4777 5224 4811
rect 5172 4768 5224 4777
rect 7564 4768 7616 4820
rect 10784 4811 10836 4820
rect 10784 4777 10793 4811
rect 10793 4777 10827 4811
rect 10827 4777 10836 4811
rect 10784 4768 10836 4777
rect 11336 4811 11388 4820
rect 11336 4777 11345 4811
rect 11345 4777 11379 4811
rect 11379 4777 11388 4811
rect 11336 4768 11388 4777
rect 11796 4811 11848 4820
rect 11796 4777 11805 4811
rect 11805 4777 11839 4811
rect 11839 4777 11848 4811
rect 11796 4768 11848 4777
rect 11888 4768 11940 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 15660 4768 15712 4820
rect 16580 4811 16632 4820
rect 16580 4777 16589 4811
rect 16589 4777 16623 4811
rect 16623 4777 16632 4811
rect 16580 4768 16632 4777
rect 21916 4811 21968 4820
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 7748 4743 7800 4752
rect 7748 4709 7757 4743
rect 7757 4709 7791 4743
rect 7791 4709 7800 4743
rect 7748 4700 7800 4709
rect 11612 4700 11664 4752
rect 12348 4700 12400 4752
rect 15752 4700 15804 4752
rect 19800 4700 19852 4752
rect 20536 4743 20588 4752
rect 20536 4709 20545 4743
rect 20545 4709 20579 4743
rect 20579 4709 20588 4743
rect 20536 4700 20588 4709
rect 20720 4700 20772 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 2320 4632 2372 4684
rect 13268 4675 13320 4684
rect 13268 4641 13277 4675
rect 13277 4641 13311 4675
rect 13311 4641 13320 4675
rect 13268 4632 13320 4641
rect 3700 4564 3752 4616
rect 7656 4564 7708 4616
rect 8392 4607 8444 4616
rect 8392 4573 8401 4607
rect 8401 4573 8435 4607
rect 8435 4573 8444 4607
rect 8392 4564 8444 4573
rect 12164 4564 12216 4616
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 19432 4496 19484 4548
rect 19892 4632 19944 4684
rect 19984 4564 20036 4616
rect 20628 4496 20680 4548
rect 21916 4777 21925 4811
rect 21925 4777 21959 4811
rect 21959 4777 21968 4811
rect 21916 4768 21968 4777
rect 25228 4768 25280 4820
rect 23572 4700 23624 4752
rect 21916 4632 21968 4684
rect 22100 4632 22152 4684
rect 22928 4632 22980 4684
rect 24308 4632 24360 4684
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 21640 4564 21692 4616
rect 22100 4496 22152 4548
rect 24860 4539 24912 4548
rect 24860 4505 24869 4539
rect 24869 4505 24903 4539
rect 24903 4505 24912 4539
rect 24860 4496 24912 4505
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 1676 4428 1728 4480
rect 4068 4471 4120 4480
rect 4068 4437 4077 4471
rect 4077 4437 4111 4471
rect 4111 4437 4120 4471
rect 4068 4428 4120 4437
rect 6920 4471 6972 4480
rect 6920 4437 6929 4471
rect 6929 4437 6963 4471
rect 6963 4437 6972 4471
rect 6920 4428 6972 4437
rect 7196 4471 7248 4480
rect 7196 4437 7205 4471
rect 7205 4437 7239 4471
rect 7239 4437 7248 4471
rect 7196 4428 7248 4437
rect 7288 4428 7340 4480
rect 20904 4471 20956 4480
rect 20904 4437 20913 4471
rect 20913 4437 20947 4471
rect 20947 4437 20956 4471
rect 20904 4428 20956 4437
rect 26792 4428 26844 4480
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 3700 4224 3752 4276
rect 4252 4224 4304 4276
rect 7564 4224 7616 4276
rect 11796 4224 11848 4276
rect 13544 4224 13596 4276
rect 16304 4224 16356 4276
rect 19984 4224 20036 4276
rect 23572 4224 23624 4276
rect 24308 4267 24360 4276
rect 24308 4233 24317 4267
rect 24317 4233 24351 4267
rect 24351 4233 24360 4267
rect 24308 4224 24360 4233
rect 25228 4224 25280 4276
rect 26516 4224 26568 4276
rect 2320 4131 2372 4140
rect 2320 4097 2329 4131
rect 2329 4097 2363 4131
rect 2363 4097 2372 4131
rect 2320 4088 2372 4097
rect 3792 4088 3844 4140
rect 4436 4088 4488 4140
rect 7748 4156 7800 4208
rect 13360 4156 13412 4208
rect 19432 4156 19484 4208
rect 19708 4131 19760 4140
rect 4896 4020 4948 4072
rect 6920 4020 6972 4072
rect 7840 4020 7892 4072
rect 16580 4020 16632 4072
rect 2044 3995 2096 4004
rect 2044 3961 2053 3995
rect 2053 3961 2087 3995
rect 2087 3961 2096 3995
rect 2044 3952 2096 3961
rect 7748 3952 7800 4004
rect 10600 3952 10652 4004
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 20444 4131 20496 4140
rect 20444 4097 20453 4131
rect 20453 4097 20487 4131
rect 20487 4097 20496 4131
rect 20444 4088 20496 4097
rect 21364 4088 21416 4140
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 20812 4020 20864 4072
rect 21824 4063 21876 4072
rect 21824 4029 21833 4063
rect 21833 4029 21867 4063
rect 21867 4029 21876 4063
rect 21824 4020 21876 4029
rect 22100 4020 22152 4072
rect 17684 3952 17736 4004
rect 19708 3952 19760 4004
rect 20444 3952 20496 4004
rect 20628 3952 20680 4004
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 2412 3884 2464 3936
rect 7564 3927 7616 3936
rect 7564 3893 7573 3927
rect 7573 3893 7607 3927
rect 7607 3893 7616 3927
rect 7564 3884 7616 3893
rect 10784 3884 10836 3936
rect 11612 3884 11664 3936
rect 12164 3927 12216 3936
rect 12164 3893 12173 3927
rect 12173 3893 12207 3927
rect 12207 3893 12216 3927
rect 12164 3884 12216 3893
rect 12256 3884 12308 3936
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 16396 3927 16448 3936
rect 16396 3893 16405 3927
rect 16405 3893 16439 3927
rect 16439 3893 16448 3927
rect 16396 3884 16448 3893
rect 19892 3927 19944 3936
rect 19892 3893 19901 3927
rect 19901 3893 19935 3927
rect 19935 3893 19944 3927
rect 19892 3884 19944 3893
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 27528 4063 27580 4072
rect 27528 4029 27537 4063
rect 27537 4029 27571 4063
rect 27571 4029 27580 4063
rect 27528 4020 27580 4029
rect 20352 3884 20404 3893
rect 26332 3927 26384 3936
rect 26332 3893 26341 3927
rect 26341 3893 26375 3927
rect 26375 3893 26384 3927
rect 26332 3884 26384 3893
rect 26608 3927 26660 3936
rect 26608 3893 26617 3927
rect 26617 3893 26651 3927
rect 26651 3893 26660 3927
rect 26608 3884 26660 3893
rect 27712 3927 27764 3936
rect 27712 3893 27721 3927
rect 27721 3893 27755 3927
rect 27755 3893 27764 3927
rect 27712 3884 27764 3893
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 2504 3680 2556 3732
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 4160 3680 4212 3732
rect 2688 3544 2740 3596
rect 2780 3544 2832 3596
rect 7012 3680 7064 3732
rect 8024 3680 8076 3732
rect 12164 3680 12216 3732
rect 17684 3723 17736 3732
rect 17684 3689 17693 3723
rect 17693 3689 17727 3723
rect 17727 3689 17736 3723
rect 17684 3680 17736 3689
rect 19892 3680 19944 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 21640 3723 21692 3732
rect 21640 3689 21649 3723
rect 21649 3689 21683 3723
rect 21683 3689 21692 3723
rect 21640 3680 21692 3689
rect 4620 3612 4672 3664
rect 9864 3587 9916 3596
rect 9864 3553 9873 3587
rect 9873 3553 9907 3587
rect 9907 3553 9916 3587
rect 11704 3612 11756 3664
rect 9864 3544 9916 3553
rect 11428 3587 11480 3596
rect 11428 3553 11462 3587
rect 11462 3553 11480 3587
rect 11428 3544 11480 3553
rect 15752 3544 15804 3596
rect 16304 3587 16356 3596
rect 16304 3553 16313 3587
rect 16313 3553 16347 3587
rect 16347 3553 16356 3587
rect 16304 3544 16356 3553
rect 16580 3587 16632 3596
rect 16580 3553 16614 3587
rect 16614 3553 16632 3587
rect 16580 3544 16632 3553
rect 20260 3612 20312 3664
rect 20076 3544 20128 3596
rect 20812 3544 20864 3596
rect 23480 3587 23532 3596
rect 23480 3553 23489 3587
rect 23489 3553 23523 3587
rect 23523 3553 23532 3587
rect 23480 3544 23532 3553
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 6552 3476 6604 3528
rect 7472 3476 7524 3528
rect 10140 3519 10192 3528
rect 7196 3408 7248 3460
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 20628 3476 20680 3528
rect 22008 3476 22060 3528
rect 8392 3408 8444 3460
rect 1584 3383 1636 3392
rect 1584 3349 1593 3383
rect 1593 3349 1627 3383
rect 1627 3349 1636 3383
rect 1584 3340 1636 3349
rect 2688 3383 2740 3392
rect 2688 3349 2697 3383
rect 2697 3349 2731 3383
rect 2731 3349 2740 3383
rect 2688 3340 2740 3349
rect 6276 3340 6328 3392
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 20260 3383 20312 3392
rect 20260 3349 20269 3383
rect 20269 3349 20303 3383
rect 20303 3349 20312 3383
rect 20260 3340 20312 3349
rect 23664 3383 23716 3392
rect 23664 3349 23673 3383
rect 23673 3349 23707 3383
rect 23707 3349 23716 3383
rect 23664 3340 23716 3349
rect 26700 3383 26752 3392
rect 26700 3349 26709 3383
rect 26709 3349 26743 3383
rect 26743 3349 26752 3383
rect 26700 3340 26752 3349
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2504 3136 2556 3188
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 3792 3179 3844 3188
rect 2780 3136 2832 3145
rect 3792 3145 3801 3179
rect 3801 3145 3835 3179
rect 3835 3145 3844 3179
rect 3792 3136 3844 3145
rect 6920 3136 6972 3188
rect 5632 3068 5684 3120
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 4620 3000 4672 3052
rect 5540 3000 5592 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 7104 3000 7156 3052
rect 11428 3136 11480 3188
rect 11704 3179 11756 3188
rect 11704 3145 11713 3179
rect 11713 3145 11747 3179
rect 11747 3145 11756 3179
rect 11704 3136 11756 3145
rect 15292 3136 15344 3188
rect 16580 3136 16632 3188
rect 19064 3179 19116 3188
rect 19064 3145 19073 3179
rect 19073 3145 19107 3179
rect 19107 3145 19116 3179
rect 19064 3136 19116 3145
rect 19340 3179 19392 3188
rect 19340 3145 19349 3179
rect 19349 3145 19383 3179
rect 19383 3145 19392 3179
rect 19340 3136 19392 3145
rect 20260 3136 20312 3188
rect 22100 3136 22152 3188
rect 24768 3179 24820 3188
rect 24768 3145 24777 3179
rect 24777 3145 24811 3179
rect 24811 3145 24820 3179
rect 24768 3136 24820 3145
rect 26516 3136 26568 3188
rect 8024 3111 8076 3120
rect 8024 3077 8033 3111
rect 8033 3077 8067 3111
rect 8067 3077 8076 3111
rect 8024 3068 8076 3077
rect 8392 3111 8444 3120
rect 8392 3077 8401 3111
rect 8401 3077 8435 3111
rect 8435 3077 8444 3111
rect 8392 3068 8444 3077
rect 16304 3068 16356 3120
rect 17684 3068 17736 3120
rect 20076 3043 20128 3052
rect 20076 3009 20085 3043
rect 20085 3009 20119 3043
rect 20119 3009 20128 3043
rect 20076 3000 20128 3009
rect 3148 2932 3200 2984
rect 3792 2932 3844 2984
rect 7288 2932 7340 2984
rect 9496 2932 9548 2984
rect 11704 2932 11756 2984
rect 15292 2932 15344 2984
rect 18236 2975 18288 2984
rect 18236 2941 18245 2975
rect 18245 2941 18279 2975
rect 18279 2941 18288 2975
rect 18236 2932 18288 2941
rect 19064 2932 19116 2984
rect 2044 2864 2096 2916
rect 2596 2864 2648 2916
rect 4896 2864 4948 2916
rect 6920 2864 6972 2916
rect 7564 2864 7616 2916
rect 15016 2907 15068 2916
rect 15016 2873 15025 2907
rect 15025 2873 15059 2907
rect 15059 2873 15068 2907
rect 15016 2864 15068 2873
rect 19156 2864 19208 2916
rect 19340 2864 19392 2916
rect 19984 2907 20036 2916
rect 19984 2873 19993 2907
rect 19993 2873 20027 2907
rect 20027 2873 20036 2907
rect 19984 2864 20036 2873
rect 24768 2932 24820 2984
rect 26884 2932 26936 2984
rect 27528 2975 27580 2984
rect 27528 2941 27537 2975
rect 27537 2941 27571 2975
rect 27571 2941 27580 2975
rect 27528 2932 27580 2941
rect 21456 2864 21508 2916
rect 21916 2864 21968 2916
rect 24860 2864 24912 2916
rect 1400 2796 1452 2848
rect 4804 2839 4856 2848
rect 4804 2805 4813 2839
rect 4813 2805 4847 2839
rect 4847 2805 4856 2839
rect 4804 2796 4856 2805
rect 23480 2796 23532 2848
rect 25320 2796 25372 2848
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 27712 2839 27764 2848
rect 27712 2805 27721 2839
rect 27721 2805 27755 2839
rect 27755 2805 27764 2839
rect 27712 2796 27764 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 4068 2592 4120 2644
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 5632 2635 5684 2644
rect 5632 2601 5641 2635
rect 5641 2601 5675 2635
rect 5675 2601 5684 2635
rect 5632 2592 5684 2601
rect 6276 2635 6328 2644
rect 6276 2601 6285 2635
rect 6285 2601 6319 2635
rect 6319 2601 6328 2635
rect 6276 2592 6328 2601
rect 6920 2592 6972 2644
rect 7380 2635 7432 2644
rect 7380 2601 7389 2635
rect 7389 2601 7423 2635
rect 7423 2601 7432 2635
rect 7380 2592 7432 2601
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 17684 2635 17736 2644
rect 17684 2601 17693 2635
rect 17693 2601 17727 2635
rect 17727 2601 17736 2635
rect 17684 2592 17736 2601
rect 17776 2592 17828 2644
rect 2964 2567 3016 2576
rect 2964 2533 2973 2567
rect 2973 2533 3007 2567
rect 3007 2533 3016 2567
rect 2964 2524 3016 2533
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 7564 2524 7616 2576
rect 4344 2388 4396 2440
rect 6276 2388 6328 2440
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 11520 2524 11572 2576
rect 9772 2456 9824 2465
rect 13728 2456 13780 2508
rect 16396 2499 16448 2508
rect 16396 2465 16405 2499
rect 16405 2465 16439 2499
rect 16439 2465 16448 2499
rect 16396 2456 16448 2465
rect 20076 2592 20128 2644
rect 20168 2592 20220 2644
rect 20812 2592 20864 2644
rect 21456 2635 21508 2644
rect 21456 2601 21465 2635
rect 21465 2601 21499 2635
rect 21499 2601 21508 2635
rect 21456 2592 21508 2601
rect 24492 2592 24544 2644
rect 25596 2635 25648 2644
rect 25596 2601 25605 2635
rect 25605 2601 25639 2635
rect 25639 2601 25648 2635
rect 25596 2592 25648 2601
rect 21548 2456 21600 2508
rect 25320 2456 25372 2508
rect 26884 2499 26936 2508
rect 26884 2465 26893 2499
rect 26893 2465 26927 2499
rect 26927 2465 26936 2499
rect 26884 2456 26936 2465
rect 9220 2388 9272 2440
rect 13452 2388 13504 2440
rect 14924 2388 14976 2440
rect 17776 2388 17828 2440
rect 23480 2388 23532 2440
rect 26332 2388 26384 2440
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 3516 2252 3568 2304
rect 27068 2295 27120 2304
rect 27068 2261 27077 2295
rect 27077 2261 27111 2295
rect 27111 2261 27120 2295
rect 27068 2252 27120 2261
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 1674 23520 1730 24000
rect 3422 23624 3478 23633
rect 3422 23559 3478 23568
rect 1688 20058 1716 23520
rect 2962 22400 3018 22409
rect 2962 22335 3018 22344
rect 2976 22166 3004 22335
rect 3436 22302 3464 23559
rect 4986 23520 5042 24000
rect 8298 23520 8354 24000
rect 11610 23520 11666 24000
rect 14922 23520 14978 24000
rect 18326 23520 18382 24000
rect 21638 23520 21694 24000
rect 24950 23520 25006 24000
rect 25134 23624 25190 23633
rect 25134 23559 25190 23568
rect 4158 23080 4214 23089
rect 4158 23015 4214 23024
rect 3424 22296 3476 22302
rect 3424 22238 3476 22244
rect 2964 22160 3016 22166
rect 2964 22102 3016 22108
rect 4066 21856 4122 21865
rect 4066 21791 4122 21800
rect 3698 21312 3754 21321
rect 3698 21247 3754 21256
rect 3712 21010 3740 21247
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 4080 20806 4108 21791
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 1858 20632 1914 20641
rect 1858 20567 1860 20576
rect 1912 20567 1914 20576
rect 1860 20538 1912 20544
rect 3422 20496 3478 20505
rect 3422 20431 3478 20440
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 2596 20256 2648 20262
rect 2596 20198 2648 20204
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2136 18828 2188 18834
rect 2136 18770 2188 18776
rect 1400 18624 1452 18630
rect 1400 18566 1452 18572
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 570 16416 626 16425
rect 570 16351 626 16360
rect 584 12918 612 16351
rect 572 12912 624 12918
rect 572 12854 624 12860
rect 1412 11121 1440 18566
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 13274 1532 17478
rect 1596 16658 1624 18255
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1688 17338 1716 17682
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1596 16250 1624 16594
rect 1780 16522 1808 18158
rect 2056 18154 2084 18566
rect 2148 18193 2176 18770
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2332 18222 2360 18566
rect 2320 18216 2372 18222
rect 2134 18184 2190 18193
rect 2044 18148 2096 18154
rect 2320 18158 2372 18164
rect 2134 18119 2190 18128
rect 2044 18090 2096 18096
rect 2148 17882 2176 18119
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2332 17202 2360 17614
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 1872 16794 1900 17070
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 2136 16516 2188 16522
rect 2136 16458 2188 16464
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2148 16114 2176 16458
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 2134 16008 2190 16017
rect 2134 15943 2190 15952
rect 2148 15638 2176 15943
rect 2240 15706 2268 16934
rect 2318 16824 2374 16833
rect 2318 16759 2320 16768
rect 2372 16759 2374 16768
rect 2320 16730 2372 16736
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2136 15632 2188 15638
rect 2136 15574 2188 15580
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1768 13728 1820 13734
rect 1768 13670 1820 13676
rect 1780 13530 1808 13670
rect 1768 13524 1820 13530
rect 1768 13466 1820 13472
rect 1504 13246 1716 13274
rect 1490 11520 1546 11529
rect 1490 11455 1546 11464
rect 1504 11218 1532 11455
rect 1492 11212 1544 11218
rect 1492 11154 1544 11160
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1504 10810 1532 11154
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1596 10441 1624 11018
rect 1582 10432 1638 10441
rect 1582 10367 1638 10376
rect 1584 9920 1636 9926
rect 1582 9888 1584 9897
rect 1636 9888 1638 9897
rect 1582 9823 1638 9832
rect 1584 9376 1636 9382
rect 1582 9344 1584 9353
rect 1636 9344 1638 9353
rect 1582 9279 1638 9288
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1412 7449 1440 8502
rect 1504 8090 1532 8599
rect 1596 8129 1624 8774
rect 1582 8120 1638 8129
rect 1492 8084 1544 8090
rect 1582 8055 1638 8064
rect 1492 8026 1544 8032
rect 1398 7440 1454 7449
rect 1398 7375 1454 7384
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6730 1624 6831
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1688 6361 1716 13246
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12442 1900 13126
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 1964 12345 1992 14758
rect 2148 14550 2176 15574
rect 2228 15496 2280 15502
rect 2228 15438 2280 15444
rect 2240 15094 2268 15438
rect 2228 15088 2280 15094
rect 2228 15030 2280 15036
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 14618 2268 14826
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 2148 13433 2176 14486
rect 2134 13424 2190 13433
rect 2134 13359 2190 13368
rect 2318 12880 2374 12889
rect 2318 12815 2320 12824
rect 2372 12815 2374 12824
rect 2320 12786 2372 12792
rect 2424 12730 2452 19994
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2516 16590 2544 18090
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2516 16250 2544 16526
rect 2504 16244 2556 16250
rect 2504 16186 2556 16192
rect 2516 15502 2544 16186
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2516 12850 2544 13262
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2320 12708 2372 12714
rect 2424 12702 2544 12730
rect 2320 12650 2372 12656
rect 2044 12640 2096 12646
rect 2096 12588 2176 12594
rect 2044 12582 2176 12588
rect 2056 12566 2176 12582
rect 1950 12336 2006 12345
rect 1950 12271 2006 12280
rect 1964 11121 1992 12271
rect 2148 12238 2176 12566
rect 2332 12345 2360 12650
rect 2318 12336 2374 12345
rect 2318 12271 2374 12280
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2056 11354 2084 11562
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2148 11286 2176 12174
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 1950 11112 2006 11121
rect 1950 11047 2006 11056
rect 2136 10532 2188 10538
rect 2136 10474 2188 10480
rect 2148 10266 2176 10474
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1766 10024 1822 10033
rect 1766 9959 1822 9968
rect 1780 6866 1808 9959
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2042 8528 2098 8537
rect 2042 8463 2044 8472
rect 2096 8463 2098 8472
rect 2044 8434 2096 8440
rect 2148 8401 2176 9318
rect 2134 8392 2190 8401
rect 2134 8327 2190 8336
rect 1952 7948 2004 7954
rect 1952 7890 2004 7896
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7342 1900 7686
rect 1860 7336 1912 7342
rect 1964 7313 1992 7890
rect 1860 7278 1912 7284
rect 1950 7304 2006 7313
rect 1950 7239 2006 7248
rect 1860 7200 1912 7206
rect 1860 7142 1912 7148
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1780 6458 1808 6802
rect 1768 6452 1820 6458
rect 1768 6394 1820 6400
rect 1674 6352 1730 6361
rect 1674 6287 1730 6296
rect 1872 6254 1900 7142
rect 1964 7002 1992 7239
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1860 6248 1912 6254
rect 1860 6190 1912 6196
rect 1872 5710 1900 6190
rect 2044 6180 2096 6186
rect 2044 6122 2096 6128
rect 2056 5914 2084 6122
rect 2044 5908 2096 5914
rect 2044 5850 2096 5856
rect 1860 5704 1912 5710
rect 1582 5672 1638 5681
rect 1860 5646 1912 5652
rect 1582 5607 1584 5616
rect 1636 5607 1638 5616
rect 1584 5578 1636 5584
rect 2042 5264 2098 5273
rect 2042 5199 2044 5208
rect 2096 5199 2098 5208
rect 2044 5170 2096 5176
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 5030 1624 5063
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 2332 4690 2360 12271
rect 2412 12232 2464 12238
rect 2516 12209 2544 12702
rect 2412 12174 2464 12180
rect 2502 12200 2558 12209
rect 2424 11393 2452 12174
rect 2502 12135 2558 12144
rect 2410 11384 2466 11393
rect 2410 11319 2412 11328
rect 2464 11319 2466 11328
rect 2412 11290 2464 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2516 10266 2544 11154
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2424 9722 2452 9930
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2410 9072 2466 9081
rect 2410 9007 2412 9016
rect 2464 9007 2466 9016
rect 2412 8978 2464 8984
rect 2424 8634 2452 8978
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2410 5808 2466 5817
rect 2410 5743 2412 5752
rect 2464 5743 2466 5752
rect 2412 5714 2464 5720
rect 2424 5370 2452 5714
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 2320 4684 2372 4690
rect 2320 4626 2372 4632
rect 1412 4593 1440 4626
rect 1398 4584 1454 4593
rect 1398 4519 1454 4528
rect 1950 4584 2006 4593
rect 1950 4519 2006 4528
rect 1584 4480 1636 4486
rect 1582 4448 1584 4457
rect 1676 4480 1728 4486
rect 1636 4448 1638 4457
rect 1676 4422 1728 4428
rect 1582 4383 1638 4392
rect 1584 3936 1636 3942
rect 1582 3904 1584 3913
rect 1636 3904 1638 3913
rect 1582 3839 1638 3848
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 662 3224 718 3233
rect 662 3159 718 3168
rect 676 480 704 3159
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 2145 1440 2790
rect 1596 2689 1624 3334
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1398 2136 1454 2145
rect 1398 2071 1454 2080
rect 1596 1465 1624 2246
rect 1582 1456 1638 1465
rect 1582 1391 1638 1400
rect 1688 921 1716 4422
rect 1964 3738 1992 4519
rect 2332 4146 2360 4626
rect 2502 4176 2558 4185
rect 2320 4140 2372 4146
rect 2502 4111 2558 4120
rect 2320 4082 2372 4088
rect 2042 4040 2098 4049
rect 2042 3975 2044 3984
rect 2096 3975 2098 3984
rect 2044 3946 2096 3952
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 2042 3088 2098 3097
rect 2042 3023 2044 3032
rect 2096 3023 2098 3032
rect 2044 2994 2096 3000
rect 2044 2916 2096 2922
rect 2044 2858 2096 2864
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 2056 480 2084 2858
rect 662 0 718 480
rect 2042 0 2098 480
rect 2424 377 2452 3878
rect 2516 3738 2544 4111
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2516 3194 2544 3674
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2608 2922 2636 20198
rect 2976 19718 3004 20334
rect 2964 19712 3016 19718
rect 2964 19654 3016 19660
rect 3146 19408 3202 19417
rect 3146 19343 3202 19352
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2700 17678 2728 18226
rect 3160 17785 3188 19343
rect 3146 17776 3202 17785
rect 3146 17711 3202 17720
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2700 17134 2728 17478
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2686 16960 2742 16969
rect 2686 16895 2742 16904
rect 2700 16658 2728 16895
rect 2688 16652 2740 16658
rect 2688 16594 2740 16600
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15366 2728 15914
rect 3056 15496 3108 15502
rect 3056 15438 3108 15444
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 15026 2728 15302
rect 3068 15162 3096 15438
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2700 14618 2728 14962
rect 2872 14884 2924 14890
rect 2872 14826 2924 14832
rect 2884 14793 2912 14826
rect 2870 14784 2926 14793
rect 2870 14719 2926 14728
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2780 14476 2832 14482
rect 2780 14418 2832 14424
rect 2792 13802 2820 14418
rect 2962 14104 3018 14113
rect 2962 14039 3018 14048
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13796 2832 13802
rect 2780 13738 2832 13744
rect 2884 13530 2912 13806
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 13462 3004 14039
rect 2964 13456 3016 13462
rect 2964 13398 3016 13404
rect 2976 13297 3004 13398
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 2962 13288 3018 13297
rect 2962 13223 3018 13232
rect 2976 12986 3004 13223
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12594 2820 12650
rect 3344 12646 3372 13330
rect 2700 12566 2820 12594
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 2700 12170 2728 12566
rect 3344 12481 3372 12582
rect 3330 12472 3386 12481
rect 3330 12407 3386 12416
rect 2778 12336 2834 12345
rect 2778 12271 2780 12280
rect 2832 12271 2834 12280
rect 2780 12242 2832 12248
rect 2688 12164 2740 12170
rect 2688 12106 2740 12112
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 2780 11620 2832 11626
rect 2700 11354 2728 11591
rect 2780 11562 2832 11568
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2792 11234 2820 11562
rect 3068 11558 3096 12038
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2700 11206 2820 11234
rect 2700 10606 2728 11206
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 9926 2728 10542
rect 3068 10538 3096 11494
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2700 9722 2728 9862
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2700 7274 2728 9658
rect 2688 7268 2740 7274
rect 2688 7210 2740 7216
rect 2700 7002 2728 7210
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2792 6361 2820 7142
rect 3436 7002 3464 20431
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 4080 20097 4108 20266
rect 3882 20088 3938 20097
rect 3882 20023 3938 20032
rect 4066 20088 4122 20097
rect 4066 20023 4122 20032
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3804 18426 3832 18770
rect 3792 18420 3844 18426
rect 3792 18362 3844 18368
rect 3514 17640 3570 17649
rect 3514 17575 3570 17584
rect 3528 10577 3556 17575
rect 3698 15872 3754 15881
rect 3698 15807 3754 15816
rect 3606 13424 3662 13433
rect 3606 13359 3662 13368
rect 3514 10568 3570 10577
rect 3514 10503 3570 10512
rect 3620 8090 3648 13359
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3424 6996 3476 7002
rect 3424 6938 3476 6944
rect 3712 6390 3740 15807
rect 3896 13433 3924 20023
rect 4172 18737 4200 23015
rect 5000 20641 5028 23520
rect 5816 22160 5868 22166
rect 5816 22102 5868 22108
rect 4986 20632 5042 20641
rect 4986 20567 5042 20576
rect 4344 20256 4396 20262
rect 4344 20198 4396 20204
rect 4158 18728 4214 18737
rect 4158 18663 4214 18672
rect 4356 18170 4384 20198
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4908 19242 4936 19858
rect 5356 19712 5408 19718
rect 5408 19660 5488 19666
rect 5356 19654 5488 19660
rect 5368 19638 5488 19654
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 5460 19174 5488 19638
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 4448 18834 4476 19110
rect 4526 18864 4582 18873
rect 4436 18828 4488 18834
rect 4526 18799 4582 18808
rect 4436 18770 4488 18776
rect 4356 18142 4476 18170
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4080 17338 4108 17682
rect 4160 17604 4212 17610
rect 4160 17546 4212 17552
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4172 16658 4200 17546
rect 4264 17134 4292 18022
rect 4356 17882 4384 18022
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4252 17128 4304 17134
rect 4252 17070 4304 17076
rect 4160 16652 4212 16658
rect 4160 16594 4212 16600
rect 4172 16250 4200 16594
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4250 15328 4306 15337
rect 4250 15263 4306 15272
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3882 13424 3938 13433
rect 4080 13410 4108 13942
rect 4264 13802 4292 15263
rect 4448 13870 4476 18142
rect 4436 13864 4488 13870
rect 4436 13806 4488 13812
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4080 13394 4200 13410
rect 4080 13388 4212 13394
rect 4080 13382 4160 13388
rect 3882 13359 3938 13368
rect 4160 13330 4212 13336
rect 4356 13326 4384 13670
rect 4540 13530 4568 18799
rect 4804 18760 4856 18766
rect 4710 18728 4766 18737
rect 4804 18702 4856 18708
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4710 18663 4766 18672
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4632 18222 4660 18566
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4724 17882 4752 18663
rect 4816 18426 4844 18702
rect 4804 18420 4856 18426
rect 4804 18362 4856 18368
rect 4816 18193 4844 18362
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 4802 18184 4858 18193
rect 4802 18119 4858 18128
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4724 17202 4752 17818
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 3804 12714 3832 13126
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3896 12102 3924 12786
rect 4172 12782 4200 13126
rect 4160 12776 4212 12782
rect 4160 12718 4212 12724
rect 3976 12640 4028 12646
rect 4028 12588 4108 12594
rect 3976 12582 4108 12588
rect 3988 12566 4108 12582
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11218 3924 12038
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3976 10668 4028 10674
rect 3976 10610 4028 10616
rect 3988 9722 4016 10610
rect 4080 10554 4108 12566
rect 4356 12442 4384 13262
rect 4540 12986 4568 13466
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 4540 12753 4568 12922
rect 4526 12744 4582 12753
rect 4526 12679 4582 12688
rect 4344 12436 4396 12442
rect 4344 12378 4396 12384
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4264 11558 4292 11698
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11393 4292 11494
rect 4250 11384 4306 11393
rect 4250 11319 4306 11328
rect 4618 11112 4674 11121
rect 4344 11076 4396 11082
rect 4618 11047 4674 11056
rect 4344 11018 4396 11024
rect 4080 10538 4200 10554
rect 4080 10532 4212 10538
rect 4080 10526 4160 10532
rect 4160 10474 4212 10480
rect 4356 10266 4384 11018
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4344 10260 4396 10266
rect 4344 10202 4396 10208
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 8974 4108 9454
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3896 7410 3924 7686
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3700 6384 3752 6390
rect 2778 6352 2834 6361
rect 3700 6326 3752 6332
rect 4172 6322 4200 7686
rect 4264 7546 4292 8026
rect 4344 7880 4396 7886
rect 4344 7822 4396 7828
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4356 6934 4384 7822
rect 4344 6928 4396 6934
rect 4344 6870 4396 6876
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 2778 6287 2834 6296
rect 4160 6316 4212 6322
rect 2792 6202 2820 6287
rect 4160 6258 4212 6264
rect 2700 6186 2820 6202
rect 2688 6180 2820 6186
rect 2740 6174 2820 6180
rect 2688 6122 2740 6128
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2780 5908 2832 5914
rect 2780 5850 2832 5856
rect 2792 5166 2820 5850
rect 2976 5370 3004 6054
rect 4172 5846 4200 6258
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3146 5672 3202 5681
rect 3146 5607 3202 5616
rect 2964 5364 3016 5370
rect 2964 5306 3016 5312
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 2792 4826 2820 5102
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3160 3738 3188 5607
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 3712 4622 3740 5102
rect 4264 4826 4292 6054
rect 4356 5574 4384 6734
rect 4540 5681 4568 10406
rect 4632 8634 4660 11047
rect 4724 9897 4752 16934
rect 5092 16726 5120 18226
rect 5276 18086 5304 18702
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5276 17678 5304 18022
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17270 5396 17478
rect 5356 17264 5408 17270
rect 5356 17206 5408 17212
rect 5080 16720 5132 16726
rect 5080 16662 5132 16668
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4816 16046 4844 16526
rect 5092 16250 5120 16662
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 5460 16046 5488 19110
rect 5736 18290 5764 19178
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 4804 16040 4856 16046
rect 4804 15982 4856 15988
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5722 14784 5778 14793
rect 5722 14719 5778 14728
rect 5448 14544 5500 14550
rect 5448 14486 5500 14492
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 4988 14272 5040 14278
rect 4988 14214 5040 14220
rect 5000 13802 5028 14214
rect 5092 14074 5120 14418
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5460 13870 5488 14486
rect 5448 13864 5500 13870
rect 5446 13832 5448 13841
rect 5500 13832 5502 13841
rect 4988 13796 5040 13802
rect 5446 13767 5502 13776
rect 4988 13738 5040 13744
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11354 4844 11494
rect 4804 11348 4856 11354
rect 4804 11290 4856 11296
rect 4816 10266 4844 11290
rect 5000 11200 5028 13738
rect 5632 13728 5684 13734
rect 5632 13670 5684 13676
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5092 12986 5120 13262
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5092 11762 5120 12922
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5184 11694 5212 12174
rect 5172 11688 5224 11694
rect 5172 11630 5224 11636
rect 5262 11656 5318 11665
rect 5262 11591 5264 11600
rect 5316 11591 5318 11600
rect 5264 11562 5316 11568
rect 5552 11558 5580 12174
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5000 11172 5212 11200
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10606 4936 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 10266 5028 10474
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4710 9888 4766 9897
rect 4710 9823 4766 9832
rect 4710 9752 4766 9761
rect 4710 9687 4766 9696
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4632 8430 4660 8570
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7886 4660 8230
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4632 6118 4660 6598
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4632 5914 4660 6054
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4526 5672 4582 5681
rect 4526 5607 4582 5616
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4252 4820 4304 4826
rect 4252 4762 4304 4768
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 3712 4282 3740 4558
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 2686 3632 2742 3641
rect 2686 3567 2688 3576
rect 2740 3567 2742 3576
rect 2780 3596 2832 3602
rect 2688 3538 2740 3544
rect 2780 3538 2832 3544
rect 2688 3392 2740 3398
rect 2686 3360 2688 3369
rect 2740 3360 2742 3369
rect 2686 3295 2742 3304
rect 2792 3194 2820 3538
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 3160 2990 3188 3674
rect 3804 3194 3832 4082
rect 3792 3188 3844 3194
rect 3792 3130 3844 3136
rect 3804 2990 3832 3130
rect 3148 2984 3200 2990
rect 3148 2926 3200 2932
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2962 2816 3018 2825
rect 2962 2751 3018 2760
rect 2976 2582 3004 2751
rect 4080 2650 4108 4422
rect 4172 3738 4200 4762
rect 4264 4282 4292 4762
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4356 3505 4384 5510
rect 4448 4758 4476 5510
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4448 4146 4476 4694
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4632 3670 4660 4966
rect 4620 3664 4672 3670
rect 4724 3641 4752 9687
rect 5092 9178 5120 10746
rect 5184 10305 5212 11172
rect 5170 10296 5226 10305
rect 5170 10231 5226 10240
rect 5184 9761 5212 10231
rect 5170 9752 5226 9761
rect 5170 9687 5226 9696
rect 5552 9602 5580 11494
rect 5644 10441 5672 13670
rect 5736 10810 5764 14719
rect 5828 11218 5856 22102
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 8312 21146 8340 23520
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 8300 21140 8352 21146
rect 8300 21082 8352 21088
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 7656 20800 7708 20806
rect 7656 20742 7708 20748
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6826 20360 6882 20369
rect 6826 20295 6882 20304
rect 7104 20324 7156 20330
rect 6840 20262 6868 20295
rect 7104 20266 7156 20272
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6920 20256 6972 20262
rect 6920 20198 6972 20204
rect 6012 20097 6040 20198
rect 5998 20088 6054 20097
rect 6932 20058 6960 20198
rect 7116 20058 7144 20266
rect 5998 20023 6000 20032
rect 6052 20023 6054 20032
rect 6920 20052 6972 20058
rect 6000 19994 6052 20000
rect 6920 19994 6972 20000
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 6932 18426 6960 19994
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7484 19446 7512 19858
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7576 19310 7604 19790
rect 7564 19304 7616 19310
rect 7564 19246 7616 19252
rect 7196 19168 7248 19174
rect 7196 19110 7248 19116
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6196 16794 6224 17138
rect 6184 16788 6236 16794
rect 6236 16748 6316 16776
rect 6184 16730 6236 16736
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6288 16250 6316 16748
rect 6276 16244 6328 16250
rect 6276 16186 6328 16192
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6840 15366 6868 15982
rect 6828 15360 6880 15366
rect 6828 15302 6880 15308
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 7208 14940 7236 19110
rect 7576 18970 7604 19246
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7668 18873 7696 20742
rect 8484 20392 8536 20398
rect 8484 20334 8536 20340
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7746 19952 7802 19961
rect 7746 19887 7802 19896
rect 7760 19854 7788 19887
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7760 18970 7788 19790
rect 8404 19394 8432 20198
rect 8496 20058 8524 20334
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 8484 20052 8536 20058
rect 8484 19994 8536 20000
rect 9876 19961 9904 20198
rect 9862 19952 9918 19961
rect 9862 19887 9918 19896
rect 8404 19378 8524 19394
rect 8404 19372 8536 19378
rect 8404 19366 8484 19372
rect 8484 19314 8536 19320
rect 8496 19174 8524 19314
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7654 18864 7710 18873
rect 7654 18799 7656 18808
rect 7708 18799 7710 18808
rect 7656 18770 7708 18776
rect 7668 18426 7696 18770
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18290 7788 18906
rect 8496 18766 8524 19110
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 7852 18465 7880 18702
rect 7838 18456 7894 18465
rect 7894 18414 7972 18442
rect 7838 18391 7894 18400
rect 7748 18284 7800 18290
rect 7748 18226 7800 18232
rect 7840 18148 7892 18154
rect 7840 18090 7892 18096
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7484 17882 7512 18022
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7852 17814 7880 18090
rect 7840 17808 7892 17814
rect 7840 17750 7892 17756
rect 7944 17746 7972 18414
rect 8496 18290 8524 18702
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 9036 18624 9088 18630
rect 9036 18566 9088 18572
rect 8484 18284 8536 18290
rect 8536 18244 8616 18272
rect 8484 18226 8536 18232
rect 7932 17740 7984 17746
rect 7932 17682 7984 17688
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8036 17649 8064 17682
rect 8588 17678 8616 18244
rect 8772 18086 8800 18566
rect 9048 18222 9076 18566
rect 9310 18320 9366 18329
rect 9310 18255 9312 18264
rect 9364 18255 9366 18264
rect 9312 18226 9364 18232
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9600 17762 9628 18022
rect 9692 17882 9720 18158
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9600 17734 9720 17762
rect 8484 17672 8536 17678
rect 8022 17640 8078 17649
rect 8484 17614 8536 17620
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8022 17575 8078 17584
rect 8036 16998 8064 17575
rect 8496 17338 8524 17614
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8588 17202 8616 17614
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 8024 16992 8076 16998
rect 8022 16960 8024 16969
rect 8852 16992 8904 16998
rect 8076 16960 8078 16969
rect 8852 16934 8904 16940
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8022 16895 8078 16904
rect 8208 15904 8260 15910
rect 8208 15846 8260 15852
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 15162 7328 15506
rect 7656 15360 7708 15366
rect 7656 15302 7708 15308
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7668 14958 7696 15302
rect 8220 14958 8248 15846
rect 8864 15473 8892 16934
rect 9140 16697 9168 16934
rect 9126 16688 9182 16697
rect 9126 16623 9128 16632
rect 9180 16623 9182 16632
rect 9128 16594 9180 16600
rect 9416 16250 9444 17138
rect 9692 16794 9720 17734
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10140 17672 10192 17678
rect 10060 17632 10140 17660
rect 9864 17060 9916 17066
rect 9864 17002 9916 17008
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9876 16590 9904 17002
rect 10060 16998 10088 17632
rect 10140 17614 10192 17620
rect 10428 17105 10456 17682
rect 10230 17096 10286 17105
rect 10230 17031 10286 17040
rect 10414 17096 10470 17105
rect 10414 17031 10470 17040
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 8850 15464 8906 15473
rect 8850 15399 8906 15408
rect 7656 14952 7708 14958
rect 6274 14920 6330 14929
rect 7208 14912 7328 14940
rect 6274 14855 6330 14864
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 5816 11212 5868 11218
rect 5816 11154 5868 11160
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5828 10690 5856 11154
rect 6288 11150 6316 14855
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11150 6500 11698
rect 6564 11694 6592 12242
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5908 10736 5960 10742
rect 5906 10704 5908 10713
rect 5960 10704 5962 10713
rect 5828 10662 5906 10690
rect 6288 10690 6316 11086
rect 6472 10810 6500 11086
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 5906 10639 5962 10648
rect 6196 10662 6316 10690
rect 6196 10470 6224 10662
rect 6184 10464 6236 10470
rect 5630 10432 5686 10441
rect 6184 10406 6236 10412
rect 5630 10367 5686 10376
rect 6196 10033 6224 10406
rect 6182 10024 6238 10033
rect 6182 9959 6238 9968
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5460 9574 5580 9602
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5092 8362 5120 9114
rect 5460 8974 5488 9574
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 9042 5764 9318
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8362 5488 8910
rect 5736 8498 5764 8978
rect 7024 8945 7052 12854
rect 7194 12472 7250 12481
rect 7194 12407 7250 12416
rect 7102 9616 7158 9625
rect 7102 9551 7158 9560
rect 7010 8936 7066 8945
rect 7010 8871 7066 8880
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4816 7410 4844 7822
rect 5092 7426 5120 8298
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4908 7398 5120 7426
rect 4816 6798 4844 7346
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 6458 4844 6734
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4802 6352 4858 6361
rect 4802 6287 4804 6296
rect 4856 6287 4858 6296
rect 4804 6258 4856 6264
rect 4908 4078 4936 7398
rect 5552 7342 5580 7822
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 6840 7410 6868 8774
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 5540 7336 5592 7342
rect 5078 7304 5134 7313
rect 5540 7278 5592 7284
rect 6182 7304 6238 7313
rect 5078 7239 5080 7248
rect 5132 7239 5134 7248
rect 6182 7239 6238 7248
rect 5080 7210 5132 7216
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5080 6928 5132 6934
rect 5080 6870 5132 6876
rect 5092 6390 5120 6870
rect 5080 6384 5132 6390
rect 5078 6352 5080 6361
rect 5132 6352 5134 6361
rect 5078 6287 5134 6296
rect 5184 5846 5212 7142
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5184 4826 5212 5782
rect 5276 5710 5304 6258
rect 5644 6225 5672 7142
rect 6196 7002 6224 7239
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 5736 6458 5764 6938
rect 6274 6896 6330 6905
rect 6274 6831 6276 6840
rect 6328 6831 6330 6840
rect 6276 6802 6328 6808
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5630 6216 5686 6225
rect 5630 6151 5686 6160
rect 5828 5914 5856 6598
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 6288 6458 6316 6802
rect 6840 6798 6868 7346
rect 6828 6792 6880 6798
rect 6828 6734 6880 6740
rect 6840 6458 6868 6734
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5276 5370 5304 5646
rect 5460 5370 5488 5850
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 4896 4072 4948 4078
rect 6288 4049 6316 6394
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6932 4078 6960 4422
rect 6920 4072 6972 4078
rect 4896 4014 4948 4020
rect 6274 4040 6330 4049
rect 4802 3904 4858 3913
rect 4802 3839 4858 3848
rect 4620 3606 4672 3612
rect 4710 3632 4766 3641
rect 4342 3496 4398 3505
rect 4342 3431 4398 3440
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 4356 2446 4384 3431
rect 4632 3058 4660 3606
rect 4710 3567 4766 3576
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4632 2650 4660 2994
rect 4816 2854 4844 3839
rect 4908 3777 4936 4014
rect 6920 4014 6972 4020
rect 6274 3975 6330 3984
rect 4894 3768 4950 3777
rect 4894 3703 4950 3712
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5632 3120 5684 3126
rect 5538 3088 5594 3097
rect 5632 3062 5684 3068
rect 5538 3023 5540 3032
rect 5592 3023 5594 3032
rect 5540 2994 5592 3000
rect 4896 2916 4948 2922
rect 4896 2858 4948 2864
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 480 3556 2246
rect 4908 480 4936 2858
rect 5644 2650 5672 3062
rect 6288 2650 6316 3334
rect 6564 3058 6592 3470
rect 6932 3194 6960 4014
rect 7024 3738 7052 8871
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3641 7144 9551
rect 7208 9466 7236 12407
rect 7300 10169 7328 14912
rect 8208 14952 8260 14958
rect 7656 14894 7708 14900
rect 8128 14912 8208 14940
rect 7668 14278 7696 14894
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 14074 7696 14214
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7654 13832 7710 13841
rect 7484 13530 7512 13806
rect 7654 13767 7710 13776
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7470 13424 7526 13433
rect 7470 13359 7526 13368
rect 7484 13025 7512 13359
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7470 13016 7526 13025
rect 7576 12986 7604 13262
rect 7470 12951 7526 12960
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7576 12889 7604 12922
rect 7562 12880 7618 12889
rect 7562 12815 7618 12824
rect 7668 12442 7696 13767
rect 7930 13424 7986 13433
rect 7840 13388 7892 13394
rect 7930 13359 7932 13368
rect 7840 13330 7892 13336
rect 7984 13359 7986 13368
rect 7932 13330 7984 13336
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7760 12730 7788 13262
rect 7852 12986 7880 13330
rect 8128 13326 8156 14912
rect 8208 14894 8260 14900
rect 8300 14816 8352 14822
rect 8300 14758 8352 14764
rect 8312 14618 8340 14758
rect 8864 14657 8892 15399
rect 9600 15162 9628 15982
rect 9692 15570 9720 16050
rect 9876 15910 9904 16526
rect 10060 16017 10088 16934
rect 10046 16008 10102 16017
rect 10244 15978 10272 17031
rect 10428 16998 10456 17031
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 16833 10456 16934
rect 10414 16824 10470 16833
rect 10414 16759 10470 16768
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10046 15943 10102 15952
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10336 15910 10364 16662
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9692 15162 9720 15506
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 8850 14648 8906 14657
rect 8300 14612 8352 14618
rect 9600 14618 9628 15098
rect 8850 14583 8906 14592
rect 9588 14612 9640 14618
rect 8300 14554 8352 14560
rect 9588 14554 9640 14560
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 13841 8248 13942
rect 8312 13938 8340 14554
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8206 13832 8262 13841
rect 8206 13767 8262 13776
rect 8392 13796 8444 13802
rect 8392 13738 8444 13744
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13320 8168 13326
rect 8220 13297 8248 13670
rect 8116 13262 8168 13268
rect 8206 13288 8262 13297
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7852 12832 7880 12922
rect 8128 12918 8156 13262
rect 8206 13223 8262 13232
rect 8116 12912 8168 12918
rect 8404 12889 8432 13738
rect 8116 12854 8168 12860
rect 8390 12880 8446 12889
rect 7852 12804 7972 12832
rect 8390 12815 8446 12824
rect 7760 12702 7880 12730
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11898 7696 12378
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7852 11642 7880 12702
rect 7944 12345 7972 12804
rect 7930 12336 7986 12345
rect 7930 12271 7986 12280
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8220 11830 8248 12038
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8220 11694 8248 11766
rect 8208 11688 8260 11694
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 11354 7420 11494
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7760 11082 7788 11630
rect 7852 11614 7972 11642
rect 8208 11630 8260 11636
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 11076 7800 11082
rect 7748 11018 7800 11024
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7286 10160 7342 10169
rect 7286 10095 7342 10104
rect 7300 9994 7328 10095
rect 7484 10062 7512 10406
rect 7576 10266 7604 10610
rect 7656 10600 7708 10606
rect 7654 10568 7656 10577
rect 7708 10568 7710 10577
rect 7654 10503 7710 10512
rect 7760 10266 7788 11018
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7288 9988 7340 9994
rect 7288 9930 7340 9936
rect 7208 9438 7512 9466
rect 7288 9376 7340 9382
rect 7288 9318 7340 9324
rect 7300 8362 7328 9318
rect 7484 8498 7512 9438
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7378 8392 7434 8401
rect 7288 8356 7340 8362
rect 7378 8327 7434 8336
rect 7288 8298 7340 8304
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7208 5030 7236 6054
rect 7300 5574 7328 8298
rect 7392 6458 7420 8327
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7392 6254 7420 6394
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5166 7328 5510
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7196 5024 7248 5030
rect 7196 4966 7248 4972
rect 7208 4486 7236 4966
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7102 3632 7158 3641
rect 7102 3567 7158 3576
rect 7208 3466 7236 4422
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 7116 3058 7144 3334
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7300 2990 7328 4422
rect 7484 3534 7512 8434
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7564 5568 7616 5574
rect 7564 5510 7616 5516
rect 7576 4826 7604 5510
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7576 4282 7604 4762
rect 7668 4622 7696 4966
rect 7760 4758 7788 6054
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7564 3936 7616 3942
rect 7668 3924 7696 4558
rect 7760 4214 7788 4694
rect 7748 4208 7800 4214
rect 7748 4150 7800 4156
rect 7852 4078 7880 11494
rect 7944 10742 7972 11614
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 8036 10538 8064 11086
rect 8220 10810 8248 11154
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8300 10736 8352 10742
rect 8220 10684 8300 10690
rect 8220 10678 8352 10684
rect 8220 10662 8340 10678
rect 8404 10674 8432 12815
rect 8588 12782 8616 14214
rect 9048 13802 9076 14418
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 9588 13728 9640 13734
rect 9640 13676 9720 13682
rect 9588 13670 9720 13676
rect 9600 13654 9720 13670
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8588 12442 8616 12718
rect 8944 12708 8996 12714
rect 8944 12650 8996 12656
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8496 11150 8524 11834
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8668 11008 8720 11014
rect 8574 10976 8630 10985
rect 8668 10950 8720 10956
rect 8574 10911 8630 10920
rect 8392 10668 8444 10674
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 9518 7972 10406
rect 8036 10266 8064 10474
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9722 8156 9998
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 9178 7972 9454
rect 8220 9330 8248 10662
rect 8392 10610 8444 10616
rect 8588 10577 8616 10911
rect 8680 10674 8708 10950
rect 8956 10674 8984 12650
rect 9310 12336 9366 12345
rect 9310 12271 9366 12280
rect 8668 10668 8720 10674
rect 8944 10668 8996 10674
rect 8668 10610 8720 10616
rect 8864 10628 8944 10656
rect 8574 10568 8630 10577
rect 8574 10503 8576 10512
rect 8628 10503 8630 10512
rect 8576 10474 8628 10480
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8312 9722 8340 10134
rect 8864 10062 8892 10628
rect 8944 10610 8996 10616
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10305 9260 10406
rect 9218 10296 9274 10305
rect 9218 10231 9274 10240
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8956 9382 8984 10066
rect 9324 9518 9352 12271
rect 9588 11280 9640 11286
rect 9586 11248 9588 11257
rect 9640 11248 9642 11257
rect 9586 11183 9642 11192
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9312 9512 9364 9518
rect 9312 9454 9364 9460
rect 8300 9376 8352 9382
rect 8220 9324 8300 9330
rect 8220 9318 8352 9324
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8220 9302 8340 9318
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7944 9042 7972 9114
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7944 8634 7972 8978
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6118 7972 6598
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 7932 6112 7984 6118
rect 7930 6080 7932 6089
rect 7984 6080 7986 6089
rect 7930 6015 7986 6024
rect 7932 5772 7984 5778
rect 7932 5714 7984 5720
rect 7944 5681 7972 5714
rect 8128 5710 8156 6258
rect 8024 5704 8076 5710
rect 7930 5672 7986 5681
rect 8024 5646 8076 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7930 5607 7986 5616
rect 7944 5370 7972 5607
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 8036 4593 8064 5646
rect 8128 5098 8156 5646
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8022 4584 8078 4593
rect 8022 4519 8078 4528
rect 7840 4072 7892 4078
rect 7840 4014 7892 4020
rect 7748 4004 7800 4010
rect 7748 3946 7800 3952
rect 7616 3896 7696 3924
rect 7564 3878 7616 3884
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6366 2816 6422 2825
rect 6366 2751 6422 2760
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 5538 2544 5594 2553
rect 5538 2479 5540 2488
rect 5592 2479 5594 2488
rect 5540 2450 5592 2456
rect 6288 2446 6316 2586
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6380 480 6408 2751
rect 6932 2650 6960 2858
rect 7392 2650 7420 3334
rect 7576 2922 7604 3878
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 7576 2582 7604 2858
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7760 480 7788 3946
rect 8220 3913 8248 9302
rect 8956 9178 8984 9318
rect 9324 9178 9352 9454
rect 9600 9178 9628 10134
rect 8944 9172 8996 9178
rect 8944 9114 8996 9120
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9588 9172 9640 9178
rect 9588 9114 9640 9120
rect 9692 8974 9720 13654
rect 9876 11121 9904 15846
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 9968 14958 9996 15506
rect 10336 15065 10364 15846
rect 10322 15056 10378 15065
rect 10322 14991 10378 15000
rect 9956 14952 10008 14958
rect 9956 14894 10008 14900
rect 10336 14793 10364 14991
rect 10322 14784 10378 14793
rect 10322 14719 10378 14728
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9968 11898 9996 12582
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10060 11694 10088 12038
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10060 11354 10088 11630
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10520 11218 10548 20946
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 11624 19990 11652 23520
rect 12164 22296 12216 22302
rect 12164 22238 12216 22244
rect 10692 19984 10744 19990
rect 10692 19926 10744 19932
rect 11612 19984 11664 19990
rect 11612 19926 11664 19932
rect 10600 19916 10652 19922
rect 10600 19858 10652 19864
rect 10612 19446 10640 19858
rect 10704 19514 10732 19926
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10600 19440 10652 19446
rect 10600 19382 10652 19388
rect 10612 18834 10640 19382
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 11348 18902 11376 19654
rect 10784 18896 10836 18902
rect 10784 18838 10836 18844
rect 11336 18896 11388 18902
rect 11336 18838 11388 18844
rect 10600 18828 10652 18834
rect 10600 18770 10652 18776
rect 10612 18426 10640 18770
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10796 18358 10824 18838
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 10784 18352 10836 18358
rect 12084 18329 12112 18566
rect 10784 18294 10836 18300
rect 12070 18320 12126 18329
rect 10796 17678 10824 18294
rect 12070 18255 12126 18264
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10784 17672 10836 17678
rect 10784 17614 10836 17620
rect 10796 17338 10824 17614
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10796 17202 10824 17274
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 10796 16590 10824 17138
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10784 16584 10836 16590
rect 10784 16526 10836 16532
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 11900 15706 11928 15914
rect 11888 15700 11940 15706
rect 11888 15642 11940 15648
rect 11900 14906 11928 15642
rect 12176 15162 12204 22238
rect 14936 20505 14964 23520
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 14922 20496 14978 20505
rect 18340 20466 18368 23520
rect 20536 22160 20588 22166
rect 20536 22102 20588 22108
rect 14922 20431 14978 20440
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 13912 20392 13964 20398
rect 16672 20392 16724 20398
rect 13912 20334 13964 20340
rect 16670 20360 16672 20369
rect 19432 20392 19484 20398
rect 16724 20360 16726 20369
rect 13924 20058 13952 20334
rect 14464 20324 14516 20330
rect 19432 20334 19484 20340
rect 19706 20360 19762 20369
rect 16670 20295 16726 20304
rect 14464 20266 14516 20272
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 13728 19304 13780 19310
rect 13924 19258 13952 19994
rect 14476 19514 14504 20266
rect 15200 20256 15252 20262
rect 15200 20198 15252 20204
rect 14464 19508 14516 19514
rect 14464 19450 14516 19456
rect 13780 19252 13952 19258
rect 13728 19246 13952 19252
rect 13096 18970 13124 19246
rect 13544 19236 13596 19242
rect 13740 19230 13952 19246
rect 13544 19178 13596 19184
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 13096 18426 13124 18906
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12452 17882 12480 18158
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12452 17762 12480 17818
rect 12360 17734 12480 17762
rect 12360 16658 12388 17734
rect 12348 16652 12400 16658
rect 12268 16612 12348 16640
rect 12268 16114 12296 16612
rect 12348 16594 12400 16600
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12348 16244 12400 16250
rect 12452 16232 12480 16594
rect 12714 16552 12770 16561
rect 12714 16487 12770 16496
rect 12400 16204 12480 16232
rect 12348 16186 12400 16192
rect 12256 16108 12308 16114
rect 12256 16050 12308 16056
rect 12268 15706 12296 16050
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12164 15156 12216 15162
rect 12164 15098 12216 15104
rect 11900 14878 12020 14906
rect 12176 14890 12204 15098
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11900 14618 11928 14758
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 14074 10824 14350
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10782 13832 10838 13841
rect 11072 13802 11100 14214
rect 10782 13767 10784 13776
rect 10836 13767 10838 13776
rect 11060 13796 11112 13802
rect 10784 13738 10836 13744
rect 11060 13738 11112 13744
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 10796 13530 10824 13738
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 11348 13530 11376 13738
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11256 12782 11284 13330
rect 11426 13016 11482 13025
rect 11426 12951 11482 12960
rect 11244 12776 11296 12782
rect 11242 12744 11244 12753
rect 11440 12753 11468 12951
rect 11296 12744 11298 12753
rect 11426 12744 11482 12753
rect 11298 12702 11376 12730
rect 11242 12679 11298 12688
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10796 11937 10824 12174
rect 10782 11928 10838 11937
rect 10782 11863 10838 11872
rect 10600 11620 10652 11626
rect 10600 11562 10652 11568
rect 10612 11354 10640 11562
rect 10796 11558 10824 11863
rect 11256 11762 11284 12242
rect 11348 11801 11376 12702
rect 11426 12679 11482 12688
rect 11334 11792 11390 11801
rect 11244 11756 11296 11762
rect 11334 11727 11390 11736
rect 11244 11698 11296 11704
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 9862 11112 9918 11121
rect 9862 11047 9918 11056
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9876 9926 9904 10610
rect 10138 10568 10194 10577
rect 10138 10503 10194 10512
rect 10152 10470 10180 10503
rect 10140 10464 10192 10470
rect 10232 10464 10284 10470
rect 10140 10406 10192 10412
rect 10230 10432 10232 10441
rect 10284 10432 10286 10441
rect 10230 10367 10286 10376
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9876 9586 9904 9862
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 8956 8498 8984 8910
rect 9876 8906 9904 9522
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9042 10088 9454
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9140 8430 9168 8774
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 8300 8288 8352 8294
rect 8300 8230 8352 8236
rect 8312 7410 8340 8230
rect 9232 8090 9260 8298
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9232 7546 9260 8026
rect 9968 7750 9996 8910
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8312 7002 8340 7346
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9508 5914 9536 6802
rect 9692 6798 9720 7482
rect 9864 7268 9916 7274
rect 9864 7210 9916 7216
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6390 9720 6734
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9678 6080 9734 6089
rect 9678 6015 9734 6024
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9692 5234 9720 6015
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 8392 4616 8444 4622
rect 8390 4584 8392 4593
rect 8444 4584 8446 4593
rect 8390 4519 8446 4528
rect 8206 3904 8262 3913
rect 8206 3839 8262 3848
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8036 3126 8064 3674
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8404 3126 8432 3402
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 9496 2984 9548 2990
rect 9496 2926 9548 2932
rect 9508 2650 9536 2926
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9784 2514 9812 6598
rect 9876 6322 9904 7210
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9876 5914 9904 6258
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9862 3632 9918 3641
rect 9862 3567 9864 3576
rect 9916 3567 9918 3576
rect 9864 3538 9916 3544
rect 9968 2553 9996 7686
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6458 10180 6734
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10152 3233 10180 3470
rect 10138 3224 10194 3233
rect 10138 3159 10194 3168
rect 10244 2961 10272 10367
rect 10612 10062 10640 11018
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10520 8634 10548 8842
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10520 8090 10548 8570
rect 10796 8401 10824 11494
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10888 10470 10916 11154
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10538 11100 11086
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 10782 8392 10838 8401
rect 10782 8327 10838 8336
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5370 10548 6054
rect 10796 5642 10824 6122
rect 10888 5658 10916 10406
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11152 10124 11204 10130
rect 11152 10066 11204 10072
rect 11164 9586 11192 10066
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 11152 5840 11204 5846
rect 11152 5782 11204 5788
rect 10966 5672 11022 5681
rect 10784 5636 10836 5642
rect 10888 5630 10966 5658
rect 10966 5607 11022 5616
rect 10784 5578 10836 5584
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 11164 5302 11192 5782
rect 11336 5704 11388 5710
rect 11440 5692 11468 7142
rect 11388 5664 11468 5692
rect 11336 5646 11388 5652
rect 11152 5296 11204 5302
rect 11152 5238 11204 5244
rect 11348 5234 11376 5646
rect 10784 5228 10836 5234
rect 10784 5170 10836 5176
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 10796 5030 10824 5170
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 10796 4826 10824 4966
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 11348 4826 11376 4966
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 11336 4820 11388 4826
rect 11336 4762 11388 4768
rect 10600 4004 10652 4010
rect 10600 3946 10652 3952
rect 10230 2952 10286 2961
rect 10230 2887 10286 2896
rect 9954 2544 10010 2553
rect 9772 2508 9824 2514
rect 9954 2479 10010 2488
rect 9772 2450 9824 2456
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9232 480 9260 2382
rect 10612 480 10640 3946
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10796 3777 10824 3878
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10782 3768 10838 3777
rect 10956 3760 11252 3780
rect 10782 3703 10838 3712
rect 11428 3596 11480 3602
rect 11428 3538 11480 3544
rect 11440 3194 11468 3538
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 11532 2582 11560 14214
rect 11900 14074 11928 14554
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11992 14006 12020 14878
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12360 14414 12388 16186
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 12360 13938 12388 14350
rect 12452 13938 12480 14758
rect 12636 14278 12664 14894
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12256 13728 12308 13734
rect 12256 13670 12308 13676
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11716 12782 11744 13262
rect 12084 12986 12112 13262
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11610 12064 11666 12073
rect 11610 11999 11666 12008
rect 11624 10470 11652 11999
rect 12268 11286 12296 13670
rect 12452 13530 12480 13874
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12636 13326 12664 14214
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12622 12336 12678 12345
rect 12622 12271 12678 12280
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12360 11558 12388 12174
rect 12636 11937 12664 12271
rect 12622 11928 12678 11937
rect 12622 11863 12678 11872
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12256 11280 12308 11286
rect 12254 11248 12256 11257
rect 12308 11248 12310 11257
rect 12254 11183 12310 11192
rect 12268 11157 12296 11183
rect 12360 11082 12388 11494
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11624 5817 11652 10406
rect 12360 10266 12388 11018
rect 12348 10260 12400 10266
rect 12348 10202 12400 10208
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11716 9382 11744 9862
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11716 9178 11744 9318
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 7886 11744 9114
rect 11794 8392 11850 8401
rect 11794 8327 11850 8336
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11716 7002 11744 7822
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 11610 5808 11666 5817
rect 11716 5778 11744 6938
rect 11610 5743 11666 5752
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11612 4752 11664 4758
rect 11612 4694 11664 4700
rect 11624 3942 11652 4694
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11716 3670 11744 5714
rect 11808 4826 11836 8327
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 11992 7410 12020 7890
rect 12440 7744 12492 7750
rect 12440 7686 12492 7692
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 12162 7304 12218 7313
rect 12162 7239 12164 7248
rect 12216 7239 12218 7248
rect 12164 7210 12216 7216
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12084 6322 12112 6802
rect 12268 6662 12296 6802
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6458 12296 6598
rect 12360 6458 12388 6734
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12162 6352 12218 6361
rect 12072 6316 12124 6322
rect 12452 6338 12480 7686
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 6458 12664 7142
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12162 6287 12218 6296
rect 12360 6310 12480 6338
rect 12072 6258 12124 6264
rect 12176 6089 12204 6287
rect 12256 6248 12308 6254
rect 12254 6216 12256 6225
rect 12308 6216 12310 6225
rect 12254 6151 12310 6160
rect 12162 6080 12218 6089
rect 12162 6015 12218 6024
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11900 4826 11928 4966
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11808 4282 11836 4762
rect 11796 4276 11848 4282
rect 11796 4218 11848 4224
rect 11992 4185 12020 4966
rect 12360 4758 12388 6310
rect 12728 5914 12756 16487
rect 12990 15464 13046 15473
rect 12990 15399 13046 15408
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 12820 14929 12848 15302
rect 12900 14952 12952 14958
rect 12806 14920 12862 14929
rect 12900 14894 12952 14900
rect 12806 14855 12862 14864
rect 12820 14822 12848 14855
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13870 12848 14214
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12912 11937 12940 14894
rect 12898 11928 12954 11937
rect 12898 11863 12954 11872
rect 13004 11370 13032 15399
rect 12820 11342 13032 11370
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12452 5030 12480 5850
rect 12820 5794 12848 11342
rect 12992 11212 13044 11218
rect 12992 11154 13044 11160
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12912 10810 12940 11086
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 13004 10742 13032 11154
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 12992 10736 13044 10742
rect 12992 10678 13044 10684
rect 13280 9586 13308 10746
rect 13372 9761 13400 18566
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13464 16794 13492 18090
rect 13556 18086 13584 19178
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 13820 18760 13872 18766
rect 13740 18708 13820 18714
rect 13740 18702 13872 18708
rect 13740 18686 13860 18702
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13740 17882 13768 18686
rect 13832 18426 13860 18686
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 14108 17882 14136 18906
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14384 18358 14412 18702
rect 14476 18358 14504 19450
rect 15212 18850 15240 20198
rect 19444 20058 19472 20334
rect 19706 20295 19708 20304
rect 19760 20295 19762 20304
rect 19708 20266 19760 20272
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15672 19378 15700 19654
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15856 19310 15884 19654
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15844 19304 15896 19310
rect 15844 19246 15896 19252
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18970 15608 19110
rect 16040 18970 16068 19314
rect 16408 19174 16436 19790
rect 16488 19780 16540 19786
rect 16488 19722 16540 19728
rect 16500 19258 16528 19722
rect 17052 19514 17080 19790
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 16500 19230 16620 19258
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 16028 18964 16080 18970
rect 16028 18906 16080 18912
rect 15120 18822 15240 18850
rect 15120 18766 15148 18822
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 15028 18290 15056 18566
rect 15016 18284 15068 18290
rect 15016 18226 15068 18232
rect 14556 18080 14608 18086
rect 14556 18022 14608 18028
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14568 17338 14596 18022
rect 15028 17338 15056 18226
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 14646 17096 14702 17105
rect 14646 17031 14702 17040
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13464 16697 13492 16730
rect 13450 16688 13506 16697
rect 13450 16623 13506 16632
rect 13728 16652 13780 16658
rect 13728 16594 13780 16600
rect 13740 16250 13768 16594
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 14660 16046 14688 17031
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 15212 15638 15240 18822
rect 15844 18828 15896 18834
rect 15844 18770 15896 18776
rect 15856 18737 15884 18770
rect 16592 18766 16620 19230
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16488 18760 16540 18766
rect 15842 18728 15898 18737
rect 16488 18702 16540 18708
rect 16580 18760 16632 18766
rect 16580 18702 16632 18708
rect 15842 18663 15898 18672
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15580 18358 15608 18566
rect 15856 18426 15884 18663
rect 16500 18601 16528 18702
rect 16486 18592 16542 18601
rect 15956 18524 16252 18544
rect 16486 18527 16542 18536
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16500 18426 16528 18527
rect 15844 18420 15896 18426
rect 15844 18362 15896 18368
rect 16488 18420 16540 18426
rect 16488 18362 16540 18368
rect 15568 18352 15620 18358
rect 15568 18294 15620 18300
rect 16592 18290 16620 18702
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17882 15332 18022
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15658 17776 15714 17785
rect 15658 17711 15660 17720
rect 15712 17711 15714 17720
rect 15660 17682 15712 17688
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15488 16794 15516 16934
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15304 15910 15332 16662
rect 15488 16250 15516 16730
rect 15580 16658 15608 17614
rect 15672 17338 15700 17682
rect 15856 17678 15884 18226
rect 16684 18193 16712 19110
rect 18328 18828 18380 18834
rect 18328 18770 18380 18776
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 18248 18426 18276 18702
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18340 18290 18368 18770
rect 19444 18714 19472 19994
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 19260 18686 19472 18714
rect 19260 18426 19288 18686
rect 19340 18624 19392 18630
rect 19340 18566 19392 18572
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 16670 18184 16726 18193
rect 16670 18119 16726 18128
rect 18340 18086 18368 18226
rect 18328 18080 18380 18086
rect 18328 18022 18380 18028
rect 17316 17808 17368 17814
rect 17316 17750 17368 17756
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15476 16244 15528 16250
rect 15672 16232 15700 17274
rect 15856 17202 15884 17614
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16394 17504 16450 17513
rect 15956 17436 16252 17456
rect 16394 17439 16450 17448
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15844 17196 15896 17202
rect 15844 17138 15896 17144
rect 16026 16688 16082 16697
rect 16026 16623 16082 16632
rect 16040 16590 16068 16623
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15672 16204 15884 16232
rect 15476 16186 15528 16192
rect 15382 16008 15438 16017
rect 15382 15943 15384 15952
rect 15436 15943 15438 15952
rect 15384 15914 15436 15920
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15200 15632 15252 15638
rect 15200 15574 15252 15580
rect 15304 15586 15332 15846
rect 15212 15162 15240 15574
rect 15304 15558 15424 15586
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 15094 15332 15438
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15304 14550 15332 15030
rect 15292 14544 15344 14550
rect 15292 14486 15344 14492
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 13544 14408 13596 14414
rect 13544 14350 13596 14356
rect 13556 13734 13584 14350
rect 13740 13870 13768 14418
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13740 13530 13768 13806
rect 15292 13796 15344 13802
rect 15292 13738 15344 13744
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 14830 12880 14886 12889
rect 14830 12815 14886 12824
rect 14740 12640 14792 12646
rect 14740 12582 14792 12588
rect 13818 12200 13874 12209
rect 13818 12135 13874 12144
rect 13832 11898 13860 12135
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13832 11694 13860 11834
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 14752 11014 14780 12582
rect 14844 11898 14872 12815
rect 15014 12744 15070 12753
rect 15212 12730 15240 13398
rect 15014 12679 15016 12688
rect 15068 12679 15070 12688
rect 15120 12702 15240 12730
rect 15016 12650 15068 12656
rect 15120 12442 15148 12702
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15212 12306 15240 12582
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15016 12232 15068 12238
rect 15304 12186 15332 13738
rect 15396 12238 15424 15558
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15672 14278 15700 14894
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15568 13864 15620 13870
rect 15672 13841 15700 14214
rect 15568 13806 15620 13812
rect 15658 13832 15714 13841
rect 15474 13696 15530 13705
rect 15474 13631 15530 13640
rect 15488 12617 15516 13631
rect 15474 12608 15530 12617
rect 15474 12543 15530 12552
rect 15016 12174 15068 12180
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14292 10674 14320 10950
rect 14752 10742 14780 10950
rect 14740 10736 14792 10742
rect 14740 10678 14792 10684
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14292 9926 14320 10610
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14936 10130 14964 10406
rect 14924 10124 14976 10130
rect 14924 10066 14976 10072
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 13358 9752 13414 9761
rect 13358 9687 13414 9696
rect 13634 9752 13690 9761
rect 13634 9687 13690 9696
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 9178 13308 9522
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 6934 13124 7686
rect 13174 7440 13230 7449
rect 13174 7375 13230 7384
rect 13268 7404 13320 7410
rect 13188 7342 13216 7375
rect 13268 7346 13320 7352
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 13188 7002 13216 7278
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 12728 5766 12848 5794
rect 13084 5772 13136 5778
rect 12728 5710 12756 5766
rect 13084 5714 13136 5720
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 12728 5030 12756 5646
rect 13096 5234 13124 5714
rect 13188 5273 13216 6938
rect 13280 6934 13308 7346
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13174 5264 13230 5273
rect 13084 5228 13136 5234
rect 13174 5199 13230 5208
rect 13084 5170 13136 5176
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12348 4752 12400 4758
rect 12348 4694 12400 4700
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11978 4176 12034 4185
rect 11978 4111 12034 4120
rect 12176 3942 12204 4558
rect 12164 3936 12216 3942
rect 12164 3878 12216 3884
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12176 3738 12204 3878
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 11704 3664 11756 3670
rect 11704 3606 11756 3612
rect 11716 3194 11744 3606
rect 12268 3505 12296 3878
rect 12728 3505 12756 4966
rect 13372 4826 13400 6967
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13556 5098 13584 5510
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13280 4049 13308 4626
rect 13372 4214 13400 4762
rect 13556 4622 13584 5034
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13556 4282 13584 4558
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13266 4040 13322 4049
rect 13266 3975 13322 3984
rect 13280 3942 13308 3975
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13648 3890 13676 9687
rect 13740 9450 13768 9862
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14476 8634 14504 8910
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 7002 14228 7142
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13924 6254 13952 6734
rect 14200 6458 14228 6938
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14476 6118 14504 6734
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5370 14504 6054
rect 15028 5953 15056 12174
rect 15212 12158 15332 12186
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 15212 12073 15240 12158
rect 15292 12096 15344 12102
rect 15198 12064 15254 12073
rect 15292 12038 15344 12044
rect 15198 11999 15254 12008
rect 15198 11928 15254 11937
rect 15198 11863 15254 11872
rect 15212 11626 15240 11863
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15304 10266 15332 12038
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 10538 15424 11494
rect 15488 10674 15516 12174
rect 15580 11778 15608 13806
rect 15658 13767 15714 13776
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15672 12850 15700 13670
rect 15764 13462 15792 14758
rect 15752 13456 15804 13462
rect 15752 13398 15804 13404
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15764 12374 15792 13126
rect 15856 12374 15884 16204
rect 16408 16046 16436 17439
rect 16592 16998 16620 17546
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 17134 16896 17478
rect 16856 17128 16908 17134
rect 16670 17096 16726 17105
rect 16856 17070 16908 17076
rect 17236 17066 17264 17614
rect 16670 17031 16726 17040
rect 17224 17060 17276 17066
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16592 16590 16620 16934
rect 16684 16590 16712 17031
rect 17224 17002 17276 17008
rect 17328 16998 17356 17750
rect 18234 17640 18290 17649
rect 18234 17575 18290 17584
rect 18248 17338 18276 17575
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18248 17134 18276 17274
rect 18340 17202 18368 18022
rect 18328 17196 18380 17202
rect 18328 17138 18380 17144
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 17868 17060 17920 17066
rect 17868 17002 17920 17008
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16592 16114 16620 16526
rect 16684 16250 16712 16526
rect 16672 16244 16724 16250
rect 16724 16204 16804 16232
rect 16672 16186 16724 16192
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16684 15026 16712 15302
rect 16396 15020 16448 15026
rect 16396 14962 16448 14968
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 16408 14482 16436 14962
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16302 14376 16358 14385
rect 16302 14311 16358 14320
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16316 13802 16344 14311
rect 16408 13938 16436 14418
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16500 13433 16528 14758
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16488 13320 16540 13326
rect 16592 13308 16620 14554
rect 16672 14544 16724 14550
rect 16672 14486 16724 14492
rect 16684 13462 16712 14486
rect 16672 13456 16724 13462
rect 16672 13398 16724 13404
rect 16540 13280 16620 13308
rect 16488 13262 16540 13268
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 16488 12980 16540 12986
rect 16408 12940 16488 12968
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15580 11750 15792 11778
rect 15660 11688 15712 11694
rect 15660 11630 15712 11636
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15476 10668 15528 10674
rect 15476 10610 15528 10616
rect 15580 10606 15608 10950
rect 15568 10600 15620 10606
rect 15568 10542 15620 10548
rect 15384 10532 15436 10538
rect 15384 10474 15436 10480
rect 15672 10418 15700 11630
rect 15764 10985 15792 11750
rect 16316 11694 16344 12038
rect 16408 11762 16436 12940
rect 16592 12968 16620 13280
rect 16540 12940 16620 12968
rect 16488 12922 16540 12928
rect 16580 12708 16632 12714
rect 16580 12650 16632 12656
rect 16488 12368 16540 12374
rect 16488 12310 16540 12316
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16304 11688 16356 11694
rect 16304 11630 16356 11636
rect 16026 11520 16082 11529
rect 16026 11455 16082 11464
rect 16040 11286 16068 11455
rect 16316 11393 16344 11630
rect 16302 11384 16358 11393
rect 16302 11319 16358 11328
rect 16028 11280 16080 11286
rect 16028 11222 16080 11228
rect 15844 11212 15896 11218
rect 15844 11154 15896 11160
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 15750 10976 15806 10985
rect 15750 10911 15806 10920
rect 15580 10390 15700 10418
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15212 7954 15240 8910
rect 15200 7948 15252 7954
rect 15200 7890 15252 7896
rect 15014 5944 15070 5953
rect 15014 5879 15070 5888
rect 15028 5846 15056 5879
rect 15016 5840 15068 5846
rect 15016 5782 15068 5788
rect 14464 5364 14516 5370
rect 14464 5306 14516 5312
rect 13648 3862 13768 3890
rect 12254 3496 12310 3505
rect 12254 3431 12310 3440
rect 12714 3496 12770 3505
rect 12714 3431 12770 3440
rect 12070 3224 12126 3233
rect 11704 3188 11756 3194
rect 12070 3159 12126 3168
rect 11704 3130 11756 3136
rect 11716 2990 11744 3130
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 12084 480 12112 3159
rect 13740 2514 13768 3862
rect 15304 3194 15332 9862
rect 15396 9722 15424 9998
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15396 9110 15424 9658
rect 15384 9104 15436 9110
rect 15580 9081 15608 10390
rect 15764 10305 15792 10911
rect 15856 10810 15884 11154
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16316 10810 16344 11154
rect 16408 11150 16436 11698
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 15750 10296 15806 10305
rect 15660 10260 15712 10266
rect 15750 10231 15806 10240
rect 16394 10296 16450 10305
rect 16394 10231 16450 10240
rect 15660 10202 15712 10208
rect 15672 9722 15700 10202
rect 15752 10124 15804 10130
rect 15752 10066 15804 10072
rect 15764 9722 15792 10066
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15384 9046 15436 9052
rect 15566 9072 15622 9081
rect 15396 8634 15424 9046
rect 15566 9007 15622 9016
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 16316 8514 16344 8774
rect 16224 8498 16344 8514
rect 16212 8492 16344 8498
rect 16264 8486 16344 8492
rect 16408 8514 16436 10231
rect 16500 8673 16528 12310
rect 16592 11014 16620 12650
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16486 8664 16542 8673
rect 16486 8599 16542 8608
rect 16408 8486 16528 8514
rect 16212 8434 16264 8440
rect 16120 8424 16172 8430
rect 16118 8392 16120 8401
rect 16172 8392 16174 8401
rect 16118 8327 16174 8336
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 16028 8288 16080 8294
rect 16028 8230 16080 8236
rect 15672 7546 15700 8230
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7857 15792 7890
rect 15750 7848 15806 7857
rect 16040 7818 16068 8230
rect 16224 8022 16252 8434
rect 16212 8016 16264 8022
rect 16212 7958 16264 7964
rect 16224 7834 16252 7958
rect 15750 7783 15806 7792
rect 16028 7812 16080 7818
rect 15660 7540 15712 7546
rect 15660 7482 15712 7488
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15396 6662 15424 7278
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15580 7041 15608 7210
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15566 7032 15622 7041
rect 15566 6967 15622 6976
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15396 5778 15424 6598
rect 15384 5772 15436 5778
rect 15384 5714 15436 5720
rect 15396 5370 15424 5714
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15672 5234 15700 7142
rect 15764 7002 15792 7783
rect 16224 7806 16344 7834
rect 16028 7754 16080 7760
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16316 7546 16344 7806
rect 16394 7576 16450 7585
rect 16304 7540 16356 7546
rect 16394 7511 16450 7520
rect 16304 7482 16356 7488
rect 16408 7274 16436 7511
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 15752 6996 15804 7002
rect 15752 6938 15804 6944
rect 15764 5846 15792 6938
rect 16500 6633 16528 8486
rect 16776 7449 16804 16204
rect 17328 15337 17356 16934
rect 17880 16640 17908 17002
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18432 16658 18460 16934
rect 18420 16652 18472 16658
rect 17880 16612 18000 16640
rect 17868 16516 17920 16522
rect 17868 16458 17920 16464
rect 17880 16250 17908 16458
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17972 15638 18000 16612
rect 18420 16594 18472 16600
rect 17960 15632 18012 15638
rect 17960 15574 18012 15580
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18616 15337 18644 15506
rect 17314 15328 17370 15337
rect 17314 15263 17370 15272
rect 18602 15328 18658 15337
rect 18602 15263 18658 15272
rect 18616 15162 18644 15263
rect 18708 15162 18736 18362
rect 18892 17542 18920 17573
rect 18880 17536 18932 17542
rect 18878 17504 18880 17513
rect 18932 17504 18934 17513
rect 18878 17439 18934 17448
rect 18786 17232 18842 17241
rect 18786 17167 18842 17176
rect 18800 17134 18828 17167
rect 18892 17134 18920 17439
rect 19064 17196 19116 17202
rect 19064 17138 19116 17144
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18892 16250 18920 16526
rect 18880 16244 18932 16250
rect 18880 16186 18932 16192
rect 19076 16114 19104 17138
rect 19352 16726 19380 18566
rect 20272 18290 20300 18566
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20364 18222 20392 19110
rect 20076 18216 20128 18222
rect 20074 18184 20076 18193
rect 20352 18216 20404 18222
rect 20128 18184 20130 18193
rect 20352 18158 20404 18164
rect 20074 18119 20130 18128
rect 20364 17882 20392 18158
rect 20548 18154 20576 22102
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 21652 21146 21680 23520
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20824 20602 20852 20946
rect 23664 20800 23716 20806
rect 23664 20742 23716 20748
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20824 20505 20852 20538
rect 20810 20496 20866 20505
rect 23676 20466 23704 20742
rect 20810 20431 20866 20440
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23202 20360 23258 20369
rect 23202 20295 23258 20304
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 23216 20058 23244 20295
rect 23204 20052 23256 20058
rect 23204 19994 23256 20000
rect 22100 19916 22152 19922
rect 22100 19858 22152 19864
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21836 19378 21864 19790
rect 21824 19372 21876 19378
rect 21824 19314 21876 19320
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21640 18828 21692 18834
rect 21640 18770 21692 18776
rect 21284 18737 21312 18770
rect 21270 18728 21326 18737
rect 21270 18663 21326 18672
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20536 18148 20588 18154
rect 20536 18090 20588 18096
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20640 17898 20668 18022
rect 20640 17882 20760 17898
rect 20352 17876 20404 17882
rect 20640 17876 20772 17882
rect 20640 17870 20720 17876
rect 20352 17818 20404 17824
rect 20720 17818 20772 17824
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20180 17338 20208 17614
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 20640 17202 20668 17682
rect 20824 17678 20852 18566
rect 21284 18426 21312 18663
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21652 18358 21680 18770
rect 21640 18352 21692 18358
rect 21638 18320 21640 18329
rect 21692 18320 21694 18329
rect 21638 18255 21694 18264
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21836 17746 21864 19314
rect 22112 19258 22140 19858
rect 23216 19514 23244 19994
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 22020 19242 22140 19258
rect 23400 19242 23428 20402
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 24032 19712 24084 19718
rect 24032 19654 24084 19660
rect 23860 19378 23888 19654
rect 23848 19372 23900 19378
rect 23848 19314 23900 19320
rect 22008 19236 22140 19242
rect 22060 19230 22140 19236
rect 23388 19236 23440 19242
rect 22008 19178 22060 19184
rect 23388 19178 23440 19184
rect 22020 18358 22048 19178
rect 23860 18970 23888 19314
rect 24044 19310 24072 19654
rect 24688 19514 24716 20266
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24872 19786 24900 20198
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24872 19666 24900 19722
rect 24780 19638 24900 19666
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23662 18864 23718 18873
rect 23662 18799 23718 18808
rect 23756 18828 23808 18834
rect 23570 18592 23626 18601
rect 23570 18527 23626 18536
rect 22008 18352 22060 18358
rect 22008 18294 22060 18300
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 21824 17740 21876 17746
rect 21824 17682 21876 17688
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20456 16726 20484 16934
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21284 16794 21312 17478
rect 21468 17066 21496 17614
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21640 16992 21692 16998
rect 21640 16934 21692 16940
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 19340 16720 19392 16726
rect 19340 16662 19392 16668
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 19352 16522 19380 16662
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 19338 16280 19394 16289
rect 20180 16250 20208 16526
rect 21284 16250 21312 16730
rect 21548 16720 21600 16726
rect 21548 16662 21600 16668
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 19338 16215 19394 16224
rect 20168 16244 20220 16250
rect 19064 16108 19116 16114
rect 19064 16050 19116 16056
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18800 15609 18828 15846
rect 18892 15706 18920 15846
rect 18880 15700 18932 15706
rect 18880 15642 18932 15648
rect 18786 15600 18842 15609
rect 18786 15535 18842 15544
rect 19076 15366 19104 16050
rect 19352 15638 19380 16215
rect 20168 16186 20220 16192
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21376 16182 21404 16594
rect 21364 16176 21416 16182
rect 21364 16118 21416 16124
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 19340 15632 19392 15638
rect 19340 15574 19392 15580
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19260 15473 19288 15506
rect 19246 15464 19302 15473
rect 19246 15399 19302 15408
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 19352 15162 19380 15574
rect 19616 15496 19668 15502
rect 19616 15438 19668 15444
rect 18604 15156 18656 15162
rect 18604 15098 18656 15104
rect 18696 15156 18748 15162
rect 19340 15156 19392 15162
rect 18748 15116 18828 15144
rect 18696 15098 18748 15104
rect 18800 14550 18828 15116
rect 19340 15098 19392 15104
rect 19340 14952 19392 14958
rect 19340 14894 19392 14900
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 18788 14544 18840 14550
rect 18694 14512 18750 14521
rect 18788 14486 18840 14492
rect 18694 14447 18750 14456
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17236 12782 17264 13330
rect 17604 13326 17632 13670
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17236 12646 17264 12718
rect 17420 12714 17448 13262
rect 17604 12986 17632 13262
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17408 12708 17460 12714
rect 17408 12650 17460 12656
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17696 12424 17724 12582
rect 17696 12396 17816 12424
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11257 16896 11494
rect 16854 11248 16910 11257
rect 16854 11183 16910 11192
rect 17222 10840 17278 10849
rect 17222 10775 17278 10784
rect 17236 10577 17264 10775
rect 17222 10568 17278 10577
rect 17222 10503 17278 10512
rect 17788 9518 17816 12396
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18064 11286 18092 12242
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11626 18184 12038
rect 18144 11620 18196 11626
rect 18144 11562 18196 11568
rect 18156 11354 18184 11562
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18340 11354 18368 11494
rect 18144 11348 18196 11354
rect 18144 11290 18196 11296
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 11098 18000 11154
rect 17880 11070 18000 11098
rect 18604 11144 18656 11150
rect 18604 11086 18656 11092
rect 17880 11014 17908 11070
rect 17868 11008 17920 11014
rect 17868 10950 17920 10956
rect 17880 10470 17908 10950
rect 18616 10742 18644 11086
rect 18604 10736 18656 10742
rect 18524 10684 18604 10690
rect 18524 10678 18656 10684
rect 18524 10662 18644 10678
rect 17868 10464 17920 10470
rect 17868 10406 17920 10412
rect 17880 10169 17908 10406
rect 18524 10266 18552 10662
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 17866 10160 17922 10169
rect 17866 10095 17922 10104
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 9330 17908 9386
rect 18064 9330 18092 10066
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 17880 9302 18092 9330
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 16762 7440 16818 7449
rect 17420 7410 17448 7686
rect 16762 7375 16818 7384
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17420 6730 17448 7346
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17774 7168 17830 7177
rect 17604 6866 17632 7142
rect 17774 7103 17830 7112
rect 17592 6860 17644 6866
rect 17592 6802 17644 6808
rect 17408 6724 17460 6730
rect 17408 6666 17460 6672
rect 16856 6656 16908 6662
rect 16486 6624 16542 6633
rect 15956 6556 16252 6576
rect 16856 6598 16908 6604
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 16486 6559 16542 6568
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16488 6180 16540 6186
rect 16488 6122 16540 6128
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15672 4826 15700 5170
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15764 4758 15792 5782
rect 16500 5574 16528 6122
rect 16868 6118 16896 6598
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 16960 6186 16988 6258
rect 17512 6254 17540 6598
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16856 6112 16908 6118
rect 16856 6054 16908 6060
rect 16488 5568 16540 5574
rect 16488 5510 16540 5516
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 16500 5302 16528 5510
rect 16488 5296 16540 5302
rect 16488 5238 16540 5244
rect 16500 5098 16528 5238
rect 16488 5092 16540 5098
rect 16488 5034 16540 5040
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 15752 4752 15804 4758
rect 15752 4694 15804 4700
rect 15764 3602 15792 4694
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 16316 4282 16344 4966
rect 16304 4276 16356 4282
rect 16304 4218 16356 4224
rect 16396 3936 16448 3942
rect 16396 3878 16448 3884
rect 16500 3890 16528 5034
rect 16592 4826 16620 6054
rect 17604 5914 17632 6802
rect 17696 6798 17724 6829
rect 17684 6792 17736 6798
rect 17682 6760 17684 6769
rect 17736 6760 17738 6769
rect 17682 6695 17738 6704
rect 17696 6390 17724 6695
rect 17788 6458 17816 7103
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17788 6254 17816 6394
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17958 6080 18014 6089
rect 17958 6015 18014 6024
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17972 5846 18000 6015
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17788 5166 17816 5510
rect 17880 5370 17908 5782
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 16592 4078 16620 4762
rect 16580 4072 16632 4078
rect 17972 4049 18000 5306
rect 18064 4593 18092 9302
rect 18340 8945 18368 9998
rect 18616 9722 18644 10542
rect 18708 10130 18736 14447
rect 18800 14074 18828 14486
rect 19352 14482 19380 14894
rect 19536 14618 19564 14894
rect 19628 14890 19656 15438
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20732 15162 20760 15302
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 19616 14884 19668 14890
rect 19616 14826 19668 14832
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18800 13870 18828 14010
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 19154 13696 19210 13705
rect 19154 13631 19210 13640
rect 19168 13025 19196 13631
rect 19352 13530 19380 14418
rect 19628 14278 19656 14826
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19628 14074 19656 14214
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19432 13796 19484 13802
rect 19432 13738 19484 13744
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19444 13462 19472 13738
rect 19432 13456 19484 13462
rect 19338 13424 19394 13433
rect 19432 13398 19484 13404
rect 19338 13359 19394 13368
rect 19154 13016 19210 13025
rect 19154 12951 19210 12960
rect 18970 12880 19026 12889
rect 18970 12815 18972 12824
rect 19024 12815 19026 12824
rect 19064 12844 19116 12850
rect 18972 12786 19024 12792
rect 19064 12786 19116 12792
rect 18878 12744 18934 12753
rect 18878 12679 18880 12688
rect 18932 12679 18934 12688
rect 18880 12650 18932 12656
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 10810 18828 11494
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18788 10464 18840 10470
rect 18788 10406 18840 10412
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 9382 18460 9522
rect 18420 9376 18472 9382
rect 18420 9318 18472 9324
rect 18432 9042 18460 9318
rect 18800 9178 18828 10406
rect 18892 9586 18920 12650
rect 19076 12374 19104 12786
rect 19064 12368 19116 12374
rect 19064 12310 19116 12316
rect 18972 12300 19024 12306
rect 18972 12242 19024 12248
rect 18984 11694 19012 12242
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18984 11150 19012 11630
rect 18972 11144 19024 11150
rect 19168 11098 19196 12951
rect 18972 11086 19024 11092
rect 18984 10674 19012 11086
rect 19076 11070 19196 11098
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18984 10198 19012 10610
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18984 9081 19012 9318
rect 19076 9178 19104 11070
rect 19156 11008 19208 11014
rect 19156 10950 19208 10956
rect 19168 10606 19196 10950
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 19260 9450 19288 9862
rect 19248 9444 19300 9450
rect 19248 9386 19300 9392
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18970 9072 19026 9081
rect 18420 9036 18472 9042
rect 18420 8978 18472 8984
rect 18696 9036 18748 9042
rect 18970 9007 19026 9016
rect 18696 8978 18748 8984
rect 18326 8936 18382 8945
rect 18326 8871 18328 8880
rect 18380 8871 18382 8880
rect 18328 8842 18380 8848
rect 18340 6848 18368 8842
rect 18708 8634 18736 8978
rect 19076 8634 19104 9114
rect 19260 8974 19288 9386
rect 19352 9042 19380 13359
rect 19444 12850 19472 13398
rect 19432 12844 19484 12850
rect 19432 12786 19484 12792
rect 19430 12608 19486 12617
rect 19430 12543 19486 12552
rect 19444 11778 19472 12543
rect 19536 12442 19564 13806
rect 19616 12640 19668 12646
rect 19720 12617 19748 15098
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19996 12889 20024 13330
rect 19982 12880 20038 12889
rect 19982 12815 20038 12824
rect 19616 12582 19668 12588
rect 19706 12608 19762 12617
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19536 11898 19564 12378
rect 19628 12152 19656 12582
rect 19706 12543 19762 12552
rect 19708 12164 19760 12170
rect 19628 12124 19708 12152
rect 19708 12106 19760 12112
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19444 11750 19656 11778
rect 19720 11762 19748 12106
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18510 7848 18566 7857
rect 18510 7783 18512 7792
rect 18564 7783 18566 7792
rect 18512 7754 18564 7760
rect 18616 7546 18644 7890
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18510 7440 18566 7449
rect 18510 7375 18566 7384
rect 18524 6905 18552 7375
rect 18510 6896 18566 6905
rect 18340 6820 18460 6848
rect 18510 6831 18512 6840
rect 18328 6724 18380 6730
rect 18328 6666 18380 6672
rect 18234 6352 18290 6361
rect 18340 6322 18368 6666
rect 18234 6287 18290 6296
rect 18328 6316 18380 6322
rect 18248 5914 18276 6287
rect 18328 6258 18380 6264
rect 18236 5908 18288 5914
rect 18236 5850 18288 5856
rect 18248 5370 18276 5850
rect 18340 5710 18368 6258
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 5370 18368 5646
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18050 4584 18106 4593
rect 18050 4519 18106 4528
rect 16580 4014 16632 4020
rect 17958 4040 18014 4049
rect 17684 4004 17736 4010
rect 17958 3975 18014 3984
rect 18234 4040 18290 4049
rect 18234 3975 18290 3984
rect 17684 3946 17736 3952
rect 15752 3596 15804 3602
rect 15752 3538 15804 3544
rect 16304 3596 16356 3602
rect 16304 3538 16356 3544
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15304 2990 15332 3130
rect 16316 3126 16344 3538
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15028 2825 15056 2858
rect 15014 2816 15070 2825
rect 15014 2751 15070 2760
rect 16302 2816 16358 2825
rect 16302 2751 16358 2760
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 13464 480 13492 2382
rect 14936 480 14964 2382
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 480 16344 2751
rect 16408 2514 16436 3878
rect 16500 3862 16620 3890
rect 16592 3602 16620 3862
rect 17696 3738 17724 3946
rect 17684 3732 17736 3738
rect 17736 3692 17816 3720
rect 17684 3674 17736 3680
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16592 3194 16620 3538
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17696 2650 17724 3062
rect 17788 2650 17816 3692
rect 18248 2990 18276 3975
rect 18432 3913 18460 6820
rect 18564 6831 18566 6840
rect 18512 6802 18564 6808
rect 18524 6254 18552 6802
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18418 3904 18474 3913
rect 18418 3839 18474 3848
rect 19076 3194 19104 8570
rect 19352 8514 19380 8978
rect 19352 8486 19472 8514
rect 19340 8424 19392 8430
rect 19260 8372 19340 8378
rect 19260 8366 19392 8372
rect 19260 8350 19380 8366
rect 19260 7954 19288 8350
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19444 6338 19472 8486
rect 19628 8401 19656 11750
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19996 9654 20024 12815
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20456 12442 20484 12582
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20258 12336 20314 12345
rect 20258 12271 20314 12280
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 19524 7812 19576 7818
rect 19524 7754 19576 7760
rect 19536 7342 19564 7754
rect 19524 7336 19576 7342
rect 19524 7278 19576 7284
rect 19536 7002 19564 7278
rect 19524 6996 19576 7002
rect 19524 6938 19576 6944
rect 19628 6497 19656 8327
rect 19614 6488 19670 6497
rect 19614 6423 19670 6432
rect 19352 6310 19472 6338
rect 19352 3194 19380 6310
rect 19524 5024 19576 5030
rect 19524 4966 19576 4972
rect 19536 4593 19564 4966
rect 19522 4584 19578 4593
rect 19432 4548 19484 4554
rect 19522 4519 19578 4528
rect 19432 4490 19484 4496
rect 19444 4214 19472 4490
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19720 4146 19748 9590
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19812 4758 19840 5646
rect 19800 4752 19852 4758
rect 19996 4729 20024 6190
rect 19800 4694 19852 4700
rect 19982 4720 20038 4729
rect 19892 4684 19944 4690
rect 19982 4655 20038 4664
rect 19892 4626 19944 4632
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19720 4010 19748 4082
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19904 3942 19932 4626
rect 19996 4622 20024 4655
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 4282 20024 4558
rect 19984 4276 20036 4282
rect 19984 4218 20036 4224
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19904 3738 19932 3878
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 20088 3602 20116 11494
rect 20180 11354 20208 11494
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 20180 8430 20208 9318
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20272 7936 20300 12271
rect 20456 11762 20484 12378
rect 21272 12300 21324 12306
rect 21272 12242 21324 12248
rect 20904 12096 20956 12102
rect 20904 12038 20956 12044
rect 20718 11928 20774 11937
rect 20718 11863 20774 11872
rect 20732 11762 20760 11863
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20352 11688 20404 11694
rect 20732 11665 20760 11698
rect 20916 11694 20944 12038
rect 21284 11898 21312 12242
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 20904 11688 20956 11694
rect 20352 11630 20404 11636
rect 20718 11656 20774 11665
rect 20364 11354 20392 11630
rect 20904 11630 20956 11636
rect 20718 11591 20774 11600
rect 20718 11520 20774 11529
rect 20718 11455 20774 11464
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20732 11082 20760 11455
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20810 11384 20866 11393
rect 20956 11376 21252 11396
rect 21376 11354 21404 12174
rect 20810 11319 20866 11328
rect 21364 11348 21416 11354
rect 20824 11150 20852 11319
rect 21364 11290 21416 11296
rect 21468 11286 21496 12174
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 21364 11212 21416 11218
rect 21364 11154 21416 11160
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 21376 10742 21404 11154
rect 21364 10736 21416 10742
rect 21362 10704 21364 10713
rect 21416 10704 21418 10713
rect 21362 10639 21418 10648
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20824 9382 20852 10066
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20824 8634 20852 9318
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 21362 9072 21418 9081
rect 21362 9007 21418 9016
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20272 7908 20392 7936
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20272 3670 20300 7142
rect 20364 5370 20392 7908
rect 20824 7546 20852 8570
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20456 6322 20484 6598
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 5914 20484 6258
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20444 5568 20496 5574
rect 20444 5510 20496 5516
rect 20352 5364 20404 5370
rect 20352 5306 20404 5312
rect 20364 5166 20392 5306
rect 20456 5234 20484 5510
rect 20548 5370 20576 6122
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20456 4146 20484 5170
rect 20640 5098 20668 5646
rect 20628 5092 20680 5098
rect 20628 5034 20680 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 20548 4758 20576 4966
rect 20732 4758 20760 6054
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 20536 4752 20588 4758
rect 20536 4694 20588 4700
rect 20720 4752 20772 4758
rect 20720 4694 20772 4700
rect 20628 4548 20680 4554
rect 20628 4490 20680 4496
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 20640 4010 20668 4490
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20628 4004 20680 4010
rect 20628 3946 20680 3952
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20260 3664 20312 3670
rect 20180 3612 20260 3618
rect 20180 3606 20312 3612
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 20180 3590 20300 3606
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19076 2990 19104 3130
rect 18236 2984 18288 2990
rect 18236 2926 18288 2932
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19352 2922 19380 3130
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 19156 2916 19208 2922
rect 19156 2858 19208 2864
rect 19340 2916 19392 2922
rect 19340 2858 19392 2864
rect 19984 2916 20036 2922
rect 19984 2858 20036 2864
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17788 480 17816 2382
rect 19168 480 19196 2858
rect 19996 2553 20024 2858
rect 20088 2650 20116 2994
rect 20180 2650 20208 3590
rect 20364 3482 20392 3878
rect 20456 3641 20484 3946
rect 20732 3738 20760 4694
rect 20904 4480 20956 4486
rect 20904 4422 20956 4428
rect 20812 4072 20864 4078
rect 20916 4049 20944 4422
rect 21376 4146 21404 9007
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21468 7546 21496 7958
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21468 6934 21496 7482
rect 21456 6928 21508 6934
rect 21456 6870 21508 6876
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 20812 4014 20864 4020
rect 20902 4040 20958 4049
rect 20824 3913 20852 4014
rect 20902 3975 20958 3984
rect 20810 3904 20866 3913
rect 20810 3839 20866 3848
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20442 3632 20498 3641
rect 20442 3567 20498 3576
rect 20812 3596 20864 3602
rect 20812 3538 20864 3544
rect 20272 3454 20392 3482
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20272 3398 20300 3454
rect 20260 3392 20312 3398
rect 20260 3334 20312 3340
rect 20272 3194 20300 3334
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20168 2644 20220 2650
rect 20168 2586 20220 2592
rect 19982 2544 20038 2553
rect 19982 2479 20038 2488
rect 20640 480 20668 3470
rect 20824 2650 20852 3538
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 21468 2650 21496 2858
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21560 2514 21588 16662
rect 21652 16590 21680 16934
rect 21640 16584 21692 16590
rect 21640 16526 21692 16532
rect 21652 16114 21680 16526
rect 21640 16108 21692 16114
rect 21640 16050 21692 16056
rect 21652 15638 21680 16050
rect 21640 15632 21692 15638
rect 21640 15574 21692 15580
rect 21652 15162 21680 15574
rect 21836 15570 21864 17682
rect 22572 17338 22600 17818
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 21824 15564 21876 15570
rect 21824 15506 21876 15512
rect 21640 15156 21692 15162
rect 21640 15098 21692 15104
rect 21836 14822 21864 15506
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 21824 14816 21876 14822
rect 21824 14758 21876 14764
rect 21836 14618 21864 14758
rect 21824 14612 21876 14618
rect 21824 14554 21876 14560
rect 21732 14476 21784 14482
rect 21732 14418 21784 14424
rect 21744 14006 21772 14418
rect 21836 14074 21864 14554
rect 23400 14550 23428 15302
rect 23388 14544 23440 14550
rect 23388 14486 23440 14492
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23308 14278 23336 14418
rect 23296 14272 23348 14278
rect 23296 14214 23348 14220
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 21732 14000 21784 14006
rect 21732 13942 21784 13948
rect 23308 13870 23336 14214
rect 23296 13864 23348 13870
rect 23296 13806 23348 13812
rect 22282 13424 22338 13433
rect 22282 13359 22338 13368
rect 22928 13388 22980 13394
rect 22296 13326 22324 13359
rect 22928 13330 22980 13336
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22006 13016 22062 13025
rect 22296 12986 22324 13262
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22006 12951 22062 12960
rect 22284 12980 22336 12986
rect 22020 12918 22048 12951
rect 22284 12922 22336 12928
rect 22008 12912 22060 12918
rect 22008 12854 22060 12860
rect 22388 12442 22416 13126
rect 22940 12918 22968 13330
rect 22928 12912 22980 12918
rect 22926 12880 22928 12889
rect 22980 12880 22982 12889
rect 22926 12815 22982 12824
rect 22834 12744 22890 12753
rect 22834 12679 22890 12688
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22848 12306 22876 12679
rect 23204 12436 23256 12442
rect 23204 12378 23256 12384
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 23112 12300 23164 12306
rect 23112 12242 23164 12248
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21916 11824 21968 11830
rect 21916 11766 21968 11772
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21744 10674 21772 11562
rect 21822 11384 21878 11393
rect 21822 11319 21878 11328
rect 21836 11150 21864 11319
rect 21824 11144 21876 11150
rect 21824 11086 21876 11092
rect 21928 10996 21956 11766
rect 22020 11762 22048 12038
rect 23124 11898 23152 12242
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 22008 11756 22060 11762
rect 22008 11698 22060 11704
rect 22020 11150 22048 11698
rect 22836 11552 22888 11558
rect 22836 11494 22888 11500
rect 22282 11384 22338 11393
rect 22848 11354 22876 11494
rect 23216 11354 23244 12378
rect 23308 12322 23336 13806
rect 23400 13326 23428 14486
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23400 12986 23428 13262
rect 23388 12980 23440 12986
rect 23388 12922 23440 12928
rect 23308 12294 23428 12322
rect 23400 12238 23428 12294
rect 23388 12232 23440 12238
rect 23388 12174 23440 12180
rect 23400 11558 23428 12174
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 22282 11319 22338 11328
rect 22836 11348 22888 11354
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21836 10968 21956 10996
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 21652 9489 21680 9862
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 21652 8838 21680 9415
rect 21836 9081 21864 10968
rect 22020 10810 22048 11086
rect 22296 10810 22324 11319
rect 22836 11290 22888 11296
rect 23204 11348 23256 11354
rect 23204 11290 23256 11296
rect 22008 10804 22060 10810
rect 22008 10746 22060 10752
rect 22284 10804 22336 10810
rect 22284 10746 22336 10752
rect 22020 10266 22048 10746
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 23388 9920 23440 9926
rect 23388 9862 23440 9868
rect 22650 9616 22706 9625
rect 21916 9580 21968 9586
rect 22650 9551 22652 9560
rect 21916 9522 21968 9528
rect 22704 9551 22706 9560
rect 22652 9522 22704 9528
rect 21822 9072 21878 9081
rect 21822 9007 21878 9016
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21652 8294 21680 8774
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21652 7954 21680 8230
rect 21928 8022 21956 9522
rect 23400 9518 23428 9862
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 22112 9178 22140 9454
rect 23492 9450 23520 10406
rect 23584 10062 23612 18527
rect 23676 10198 23704 18799
rect 23756 18770 23808 18776
rect 23768 18426 23796 18770
rect 23848 18760 23900 18766
rect 23848 18702 23900 18708
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23756 18420 23808 18426
rect 23756 18362 23808 18368
rect 23860 17882 23888 18702
rect 23952 18358 23980 18702
rect 23940 18352 23992 18358
rect 23940 18294 23992 18300
rect 24124 18080 24176 18086
rect 24124 18022 24176 18028
rect 24216 18080 24268 18086
rect 24216 18022 24268 18028
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 24032 17808 24084 17814
rect 24032 17750 24084 17756
rect 23938 17504 23994 17513
rect 23938 17439 23994 17448
rect 23952 17134 23980 17439
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 24044 16794 24072 17750
rect 24136 17241 24164 18022
rect 24122 17232 24178 17241
rect 24122 17167 24178 17176
rect 24032 16788 24084 16794
rect 24032 16730 24084 16736
rect 24228 16250 24256 18022
rect 24308 17740 24360 17746
rect 24308 17682 24360 17688
rect 24320 17270 24348 17682
rect 24400 17672 24452 17678
rect 24400 17614 24452 17620
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24412 17066 24440 17614
rect 24400 17060 24452 17066
rect 24400 17002 24452 17008
rect 24308 16992 24360 16998
rect 24308 16934 24360 16940
rect 24216 16244 24268 16250
rect 24216 16186 24268 16192
rect 24124 15904 24176 15910
rect 24124 15846 24176 15852
rect 24136 15337 24164 15846
rect 24320 15609 24348 16934
rect 24412 16794 24440 17002
rect 24400 16788 24452 16794
rect 24400 16730 24452 16736
rect 24400 16040 24452 16046
rect 24400 15982 24452 15988
rect 24306 15600 24362 15609
rect 24306 15535 24362 15544
rect 24122 15328 24178 15337
rect 24122 15263 24178 15272
rect 23940 14816 23992 14822
rect 23940 14758 23992 14764
rect 23952 14414 23980 14758
rect 23940 14408 23992 14414
rect 23940 14350 23992 14356
rect 23952 14006 23980 14350
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 24216 13184 24268 13190
rect 24216 13126 24268 13132
rect 24228 12782 24256 13126
rect 24216 12776 24268 12782
rect 24216 12718 24268 12724
rect 24228 12442 24256 12718
rect 24320 12594 24348 15535
rect 24412 14929 24440 15982
rect 24398 14920 24454 14929
rect 24398 14855 24454 14864
rect 24412 12714 24440 14855
rect 24400 12708 24452 12714
rect 24400 12650 24452 12656
rect 24320 12566 24440 12594
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24320 11801 24348 12242
rect 24306 11792 24362 11801
rect 24306 11727 24308 11736
rect 24360 11727 24362 11736
rect 24308 11698 24360 11704
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24228 10470 24256 10950
rect 24306 10568 24362 10577
rect 24306 10503 24308 10512
rect 24360 10503 24362 10512
rect 24308 10474 24360 10480
rect 24216 10464 24268 10470
rect 24216 10406 24268 10412
rect 24228 10266 24256 10406
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 23664 10192 23716 10198
rect 23664 10134 23716 10140
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23676 9722 23704 10134
rect 24216 10056 24268 10062
rect 24216 9998 24268 10004
rect 23664 9716 23716 9722
rect 23664 9658 23716 9664
rect 23480 9444 23532 9450
rect 23480 9386 23532 9392
rect 24228 9382 24256 9998
rect 22192 9376 22244 9382
rect 22192 9318 22244 9324
rect 24216 9376 24268 9382
rect 24216 9318 24268 9324
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 21640 7948 21692 7954
rect 21640 7890 21692 7896
rect 21652 6662 21680 7890
rect 22204 7274 22232 9318
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23296 8560 23348 8566
rect 23296 8502 23348 8508
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22388 7410 22416 7686
rect 22376 7404 22428 7410
rect 22376 7346 22428 7352
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22204 6934 22232 7210
rect 22468 7200 22520 7206
rect 22468 7142 22520 7148
rect 22480 7002 22508 7142
rect 22468 6996 22520 7002
rect 22468 6938 22520 6944
rect 22192 6928 22244 6934
rect 22192 6870 22244 6876
rect 23308 6866 23336 8502
rect 23492 7018 23520 8774
rect 23860 8673 23888 8978
rect 23940 8968 23992 8974
rect 23940 8910 23992 8916
rect 23846 8664 23902 8673
rect 23846 8599 23848 8608
rect 23900 8599 23902 8608
rect 23848 8570 23900 8576
rect 23952 8362 23980 8910
rect 24228 8537 24256 9318
rect 24214 8528 24270 8537
rect 24214 8463 24270 8472
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23952 8090 23980 8298
rect 24412 8242 24440 12566
rect 24320 8214 24440 8242
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 23572 7540 23624 7546
rect 23572 7482 23624 7488
rect 23584 7449 23612 7482
rect 23570 7440 23626 7449
rect 23570 7375 23626 7384
rect 24136 7206 24164 7822
rect 24320 7585 24348 8214
rect 24398 8120 24454 8129
rect 24398 8055 24400 8064
rect 24452 8055 24454 8064
rect 24400 8026 24452 8032
rect 24306 7576 24362 7585
rect 24412 7546 24440 8026
rect 24306 7511 24362 7520
rect 24400 7540 24452 7546
rect 24320 7410 24348 7511
rect 24400 7482 24452 7488
rect 24308 7404 24360 7410
rect 24308 7346 24360 7352
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23400 7002 23520 7018
rect 23388 6996 23520 7002
rect 23440 6990 23520 6996
rect 23388 6938 23440 6944
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 23296 6860 23348 6866
rect 23296 6802 23348 6808
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 21652 5710 21680 6598
rect 22112 6458 22140 6802
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 6458 22692 6734
rect 23308 6458 23336 6802
rect 23492 6458 23520 6990
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21744 5409 21772 5850
rect 24136 5846 24164 7142
rect 24124 5840 24176 5846
rect 24124 5782 24176 5788
rect 22100 5704 22152 5710
rect 22100 5646 22152 5652
rect 21730 5400 21786 5409
rect 21730 5335 21732 5344
rect 21784 5335 21786 5344
rect 21732 5306 21784 5312
rect 21744 5275 21772 5306
rect 21916 5092 21968 5098
rect 21916 5034 21968 5040
rect 21928 4826 21956 5034
rect 21916 4820 21968 4826
rect 21968 4780 22048 4808
rect 21916 4762 21968 4768
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 21640 4616 21692 4622
rect 21638 4584 21640 4593
rect 21692 4584 21694 4593
rect 21638 4519 21694 4528
rect 21652 3738 21680 4519
rect 21824 4072 21876 4078
rect 21822 4040 21824 4049
rect 21876 4040 21878 4049
rect 21822 3975 21878 3984
rect 21640 3732 21692 3738
rect 21640 3674 21692 3680
rect 21928 2922 21956 4626
rect 22020 4146 22048 4780
rect 22112 4690 22140 5646
rect 23572 5568 23624 5574
rect 23572 5510 23624 5516
rect 22928 5024 22980 5030
rect 22928 4966 22980 4972
rect 22940 4690 22968 4966
rect 23584 4758 23612 5510
rect 23572 4752 23624 4758
rect 23570 4720 23572 4729
rect 23624 4720 23626 4729
rect 22100 4684 22152 4690
rect 22100 4626 22152 4632
rect 22928 4684 22980 4690
rect 23570 4655 23626 4664
rect 24308 4684 24360 4690
rect 22928 4626 22980 4632
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 22020 3618 22048 4082
rect 22112 4078 22140 4490
rect 23584 4282 23612 4655
rect 24308 4626 24360 4632
rect 24320 4282 24348 4626
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 24308 4276 24360 4282
rect 24308 4218 24360 4224
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22020 3590 22140 3618
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 21916 2916 21968 2922
rect 21916 2858 21968 2864
rect 21548 2508 21600 2514
rect 21548 2450 21600 2456
rect 22020 480 22048 3470
rect 22112 3194 22140 3590
rect 23480 3596 23532 3602
rect 23480 3538 23532 3544
rect 22100 3188 22152 3194
rect 22100 3130 22152 3136
rect 23492 2854 23520 3538
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23676 3097 23704 3334
rect 23662 3088 23718 3097
rect 23662 3023 23718 3032
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 24504 2650 24532 19110
rect 24688 18290 24716 19450
rect 24780 18766 24808 19638
rect 24768 18760 24820 18766
rect 24768 18702 24820 18708
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24688 17814 24716 18226
rect 24676 17808 24728 17814
rect 24676 17750 24728 17756
rect 24964 17270 24992 23520
rect 25044 19848 25096 19854
rect 25044 19790 25096 19796
rect 25056 19514 25084 19790
rect 25044 19508 25096 19514
rect 25044 19450 25096 19456
rect 25056 18970 25084 19450
rect 25044 18964 25096 18970
rect 25044 18906 25096 18912
rect 25044 18080 25096 18086
rect 25044 18022 25096 18028
rect 25056 17542 25084 18022
rect 25044 17536 25096 17542
rect 25044 17478 25096 17484
rect 24952 17264 25004 17270
rect 24952 17206 25004 17212
rect 25056 17202 25084 17478
rect 25044 17196 25096 17202
rect 25044 17138 25096 17144
rect 24860 17128 24912 17134
rect 24860 17070 24912 17076
rect 24872 16998 24900 17070
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24768 16652 24820 16658
rect 24768 16594 24820 16600
rect 24674 16552 24730 16561
rect 24674 16487 24730 16496
rect 24688 16454 24716 16487
rect 24676 16448 24728 16454
rect 24676 16390 24728 16396
rect 24688 15910 24716 16390
rect 24780 16289 24808 16594
rect 24766 16280 24822 16289
rect 24766 16215 24768 16224
rect 24820 16215 24822 16224
rect 24768 16186 24820 16192
rect 24780 16155 24808 16186
rect 24872 15978 24900 16934
rect 25056 16590 25084 17138
rect 25044 16584 25096 16590
rect 25044 16526 25096 16532
rect 25056 16114 25084 16526
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24860 15972 24912 15978
rect 24860 15914 24912 15920
rect 24676 15904 24728 15910
rect 24676 15846 24728 15852
rect 24582 15464 24638 15473
rect 24582 15399 24638 15408
rect 24596 15366 24624 15399
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24688 14657 24716 15846
rect 24964 15706 24992 16050
rect 25044 15972 25096 15978
rect 25044 15914 25096 15920
rect 24952 15700 25004 15706
rect 24952 15642 25004 15648
rect 24952 15564 25004 15570
rect 24952 15506 25004 15512
rect 24674 14648 24730 14657
rect 24674 14583 24730 14592
rect 24766 13968 24822 13977
rect 24766 13903 24822 13912
rect 24584 12640 24636 12646
rect 24584 12582 24636 12588
rect 24596 12170 24624 12582
rect 24780 12442 24808 13903
rect 24964 13002 24992 15506
rect 25056 14414 25084 15914
rect 25044 14408 25096 14414
rect 25044 14350 25096 14356
rect 25042 13832 25098 13841
rect 25042 13767 25098 13776
rect 24872 12974 24992 13002
rect 24768 12436 24820 12442
rect 24688 12396 24768 12424
rect 24584 12164 24636 12170
rect 24584 12106 24636 12112
rect 24688 11898 24716 12396
rect 24768 12378 24820 12384
rect 24766 12336 24822 12345
rect 24872 12322 24900 12974
rect 24952 12912 25004 12918
rect 24952 12854 25004 12860
rect 24822 12294 24900 12322
rect 24766 12271 24822 12280
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24872 11898 24900 12174
rect 24676 11892 24728 11898
rect 24676 11834 24728 11840
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24964 11626 24992 12854
rect 25056 11762 25084 13767
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24768 11552 24820 11558
rect 24768 11494 24820 11500
rect 24584 10668 24636 10674
rect 24584 10610 24636 10616
rect 24596 10062 24624 10610
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24596 9586 24624 9998
rect 24584 9580 24636 9586
rect 24584 9522 24636 9528
rect 24596 9450 24624 9522
rect 24676 9512 24728 9518
rect 24674 9480 24676 9489
rect 24728 9480 24730 9489
rect 24584 9444 24636 9450
rect 24674 9415 24730 9424
rect 24584 9386 24636 9392
rect 24596 8838 24624 9386
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24596 8498 24624 8774
rect 24584 8492 24636 8498
rect 24584 8434 24636 8440
rect 24596 8022 24624 8434
rect 24676 8424 24728 8430
rect 24676 8366 24728 8372
rect 24584 8016 24636 8022
rect 24584 7958 24636 7964
rect 24688 7546 24716 8366
rect 24676 7540 24728 7546
rect 24676 7482 24728 7488
rect 24676 6860 24728 6866
rect 24676 6802 24728 6808
rect 24688 6361 24716 6802
rect 24674 6352 24730 6361
rect 24674 6287 24730 6296
rect 24780 3194 24808 11494
rect 24964 11354 24992 11562
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 25056 11286 25084 11698
rect 25044 11280 25096 11286
rect 25044 11222 25096 11228
rect 25148 11082 25176 23559
rect 28262 23520 28318 24000
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25424 22166 25452 23015
rect 25412 22160 25464 22166
rect 25412 22102 25464 22108
rect 26974 21856 27030 21865
rect 25956 21788 26252 21808
rect 26974 21791 27030 21800
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25226 21312 25282 21321
rect 25226 21247 25282 21256
rect 25240 15570 25268 21247
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25686 20496 25742 20505
rect 25686 20431 25742 20440
rect 25410 19408 25466 19417
rect 25410 19343 25466 19352
rect 25320 19168 25372 19174
rect 25320 19110 25372 19116
rect 25332 18873 25360 19110
rect 25318 18864 25374 18873
rect 25318 18799 25374 18808
rect 25424 18601 25452 19343
rect 25596 19236 25648 19242
rect 25596 19178 25648 19184
rect 25502 18864 25558 18873
rect 25502 18799 25558 18808
rect 25410 18592 25466 18601
rect 25410 18527 25466 18536
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25228 15564 25280 15570
rect 25228 15506 25280 15512
rect 25226 15464 25282 15473
rect 25226 15399 25282 15408
rect 25136 11076 25188 11082
rect 25136 11018 25188 11024
rect 25240 10849 25268 15399
rect 25226 10840 25282 10849
rect 25226 10775 25282 10784
rect 24860 9920 24912 9926
rect 24860 9862 24912 9868
rect 24872 9489 24900 9862
rect 24858 9480 24914 9489
rect 24914 9438 24992 9466
rect 24858 9415 24914 9424
rect 24860 8356 24912 8362
rect 24860 8298 24912 8304
rect 24872 6730 24900 8298
rect 24964 8090 24992 9438
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 24964 6934 24992 7278
rect 25044 7268 25096 7274
rect 25044 7210 25096 7216
rect 25056 7041 25084 7210
rect 25042 7032 25098 7041
rect 25042 6967 25098 6976
rect 24952 6928 25004 6934
rect 24952 6870 25004 6876
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 25332 6746 25360 17206
rect 25412 16720 25464 16726
rect 25412 16662 25464 16668
rect 25424 15366 25452 16662
rect 25516 16046 25544 18799
rect 25608 18630 25636 19178
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25608 18329 25636 18566
rect 25594 18320 25650 18329
rect 25594 18255 25650 18264
rect 25700 16538 25728 20431
rect 26424 20392 26476 20398
rect 26424 20334 26476 20340
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 25608 16510 25728 16538
rect 25504 16040 25556 16046
rect 25504 15982 25556 15988
rect 25504 15700 25556 15706
rect 25504 15642 25556 15648
rect 25412 15360 25464 15366
rect 25412 15302 25464 15308
rect 25424 12753 25452 15302
rect 25516 13938 25544 15642
rect 25504 13932 25556 13938
rect 25504 13874 25556 13880
rect 25502 13424 25558 13433
rect 25502 13359 25558 13368
rect 25410 12744 25466 12753
rect 25410 12679 25466 12688
rect 25412 12640 25464 12646
rect 25412 12582 25464 12588
rect 25424 12306 25452 12582
rect 25516 12442 25544 13359
rect 25504 12436 25556 12442
rect 25504 12378 25556 12384
rect 25502 12336 25558 12345
rect 25412 12300 25464 12306
rect 25502 12271 25558 12280
rect 25412 12242 25464 12248
rect 25424 11830 25452 12242
rect 25412 11824 25464 11830
rect 25412 11766 25464 11772
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25424 7410 25452 7686
rect 25412 7404 25464 7410
rect 25412 7346 25464 7352
rect 25516 7002 25544 12271
rect 25504 6996 25556 7002
rect 25504 6938 25556 6944
rect 24860 6724 24912 6730
rect 24860 6666 24912 6672
rect 24858 6488 24914 6497
rect 24964 6474 24992 6734
rect 25332 6718 25452 6746
rect 25318 6624 25374 6633
rect 25318 6559 25374 6568
rect 24914 6446 24992 6474
rect 24858 6423 24860 6432
rect 24912 6423 24914 6432
rect 24860 6394 24912 6400
rect 25332 5778 25360 6559
rect 25320 5772 25372 5778
rect 25320 5714 25372 5720
rect 25332 5386 25360 5714
rect 25240 5370 25360 5386
rect 25228 5364 25360 5370
rect 25280 5358 25360 5364
rect 25228 5306 25280 5312
rect 25228 5160 25280 5166
rect 25228 5102 25280 5108
rect 24860 5024 24912 5030
rect 24860 4966 24912 4972
rect 24872 4593 24900 4966
rect 25240 4826 25268 5102
rect 25228 4820 25280 4826
rect 25228 4762 25280 4768
rect 24858 4584 24914 4593
rect 24858 4519 24860 4528
rect 24912 4519 24914 4528
rect 24860 4490 24912 4496
rect 25240 4282 25268 4762
rect 25228 4276 25280 4282
rect 25228 4218 25280 4224
rect 24768 3188 24820 3194
rect 24768 3130 24820 3136
rect 24780 2990 24808 3130
rect 24768 2984 24820 2990
rect 24768 2926 24820 2932
rect 24860 2916 24912 2922
rect 24860 2858 24912 2864
rect 24492 2644 24544 2650
rect 24492 2586 24544 2592
rect 23480 2440 23532 2446
rect 23480 2382 23532 2388
rect 23492 480 23520 2382
rect 24872 480 24900 2858
rect 25332 2854 25360 2885
rect 25320 2848 25372 2854
rect 25424 2802 25452 6718
rect 25516 6458 25544 6938
rect 25608 6769 25636 16510
rect 25792 16266 25820 18158
rect 26160 17898 26188 18158
rect 26160 17882 26280 17898
rect 26160 17876 26292 17882
rect 26160 17870 26240 17876
rect 26240 17818 26292 17824
rect 25870 17640 25926 17649
rect 25870 17575 25926 17584
rect 25700 16238 25820 16266
rect 25700 16114 25728 16238
rect 25778 16144 25834 16153
rect 25688 16108 25740 16114
rect 25778 16079 25834 16088
rect 25688 16050 25740 16056
rect 25688 15904 25740 15910
rect 25688 15846 25740 15852
rect 25700 13841 25728 15846
rect 25792 14521 25820 16079
rect 25778 14512 25834 14521
rect 25778 14447 25834 14456
rect 25780 14408 25832 14414
rect 25884 14385 25912 17575
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25964 16040 26016 16046
rect 25964 15982 26016 15988
rect 25976 15706 26004 15982
rect 25964 15700 26016 15706
rect 25964 15642 26016 15648
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25780 14350 25832 14356
rect 25870 14376 25926 14385
rect 25686 13832 25742 13841
rect 25686 13767 25742 13776
rect 25792 13433 25820 14350
rect 25870 14311 25926 14320
rect 25872 14272 25924 14278
rect 25872 14214 25924 14220
rect 25884 13734 25912 14214
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26056 13932 26108 13938
rect 26056 13874 26108 13880
rect 25872 13728 25924 13734
rect 25872 13670 25924 13676
rect 25778 13424 25834 13433
rect 25778 13359 25834 13368
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 12782 25820 13126
rect 25884 12850 25912 13670
rect 26068 13530 26096 13874
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25872 12844 25924 12850
rect 25872 12786 25924 12792
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 25688 12640 25740 12646
rect 25688 12582 25740 12588
rect 25700 11694 25728 12582
rect 25792 11898 25820 12718
rect 26148 12640 26200 12646
rect 26148 12582 26200 12588
rect 26332 12640 26384 12646
rect 26332 12582 26384 12588
rect 25872 12436 25924 12442
rect 25872 12378 25924 12384
rect 25780 11892 25832 11898
rect 25780 11834 25832 11840
rect 25688 11688 25740 11694
rect 25688 11630 25740 11636
rect 25700 11354 25728 11630
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25884 8242 25912 12378
rect 26160 12170 26188 12582
rect 26344 12442 26372 12582
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 26148 12164 26200 12170
rect 26148 12106 26200 12112
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 26160 11082 26188 11562
rect 26148 11076 26200 11082
rect 26148 11018 26200 11024
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 26436 10826 26464 20334
rect 26988 20058 27016 21791
rect 28276 20602 28304 23520
rect 28264 20596 28316 20602
rect 28264 20538 28316 20544
rect 26976 20052 27028 20058
rect 26976 19994 27028 20000
rect 26884 19916 26936 19922
rect 26884 19858 26936 19864
rect 26896 19514 26924 19858
rect 26884 19508 26936 19514
rect 26884 19450 26936 19456
rect 26896 18970 26924 19450
rect 26988 19446 27016 19994
rect 27068 19848 27120 19854
rect 27068 19790 27120 19796
rect 26976 19440 27028 19446
rect 26976 19382 27028 19388
rect 26884 18964 26936 18970
rect 26884 18906 26936 18912
rect 26514 18728 26570 18737
rect 26514 18663 26570 18672
rect 26528 17746 26556 18663
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26528 17338 26556 17682
rect 26884 17536 26936 17542
rect 26884 17478 26936 17484
rect 26516 17332 26568 17338
rect 26516 17274 26568 17280
rect 26514 17232 26570 17241
rect 26514 17167 26570 17176
rect 26528 15570 26556 17167
rect 26516 15564 26568 15570
rect 26516 15506 26568 15512
rect 26528 15162 26556 15506
rect 26792 15360 26844 15366
rect 26792 15302 26844 15308
rect 26516 15156 26568 15162
rect 26516 15098 26568 15104
rect 26516 12640 26568 12646
rect 26516 12582 26568 12588
rect 26528 11694 26556 12582
rect 26608 12368 26660 12374
rect 26608 12310 26660 12316
rect 26516 11688 26568 11694
rect 26516 11630 26568 11636
rect 26516 11552 26568 11558
rect 26620 11506 26648 12310
rect 26698 11656 26754 11665
rect 26698 11591 26754 11600
rect 26568 11500 26648 11506
rect 26516 11494 26648 11500
rect 26528 11478 26648 11494
rect 26528 11257 26556 11478
rect 26712 11354 26740 11591
rect 26700 11348 26752 11354
rect 26700 11290 26752 11296
rect 26514 11248 26570 11257
rect 26514 11183 26516 11192
rect 26568 11183 26570 11192
rect 26516 11154 26568 11160
rect 26344 10798 26464 10826
rect 26528 10810 26556 11154
rect 26516 10804 26568 10810
rect 26344 10418 26372 10798
rect 26516 10746 26568 10752
rect 26422 10704 26478 10713
rect 26422 10639 26478 10648
rect 26436 10606 26464 10639
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26608 10464 26660 10470
rect 26606 10432 26608 10441
rect 26660 10432 26662 10441
rect 26344 10390 26464 10418
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26056 9648 26108 9654
rect 26054 9616 26056 9625
rect 26108 9616 26110 9625
rect 26054 9551 26110 9560
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 26160 8378 26188 8434
rect 26160 8350 26280 8378
rect 26252 8276 26280 8350
rect 26252 8248 26372 8276
rect 25792 8214 25912 8242
rect 25792 7478 25820 8214
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25780 7472 25832 7478
rect 25780 7414 25832 7420
rect 25884 7410 25912 8026
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26344 7546 26372 8248
rect 26332 7540 26384 7546
rect 26332 7482 26384 7488
rect 25872 7404 25924 7410
rect 25872 7346 25924 7352
rect 25688 7200 25740 7206
rect 25964 7200 26016 7206
rect 25688 7142 25740 7148
rect 25962 7168 25964 7177
rect 26016 7168 26018 7177
rect 25700 6798 25728 7142
rect 25962 7103 26018 7112
rect 25688 6792 25740 6798
rect 25594 6760 25650 6769
rect 25688 6734 25740 6740
rect 25594 6695 25650 6704
rect 26332 6656 26384 6662
rect 26332 6598 26384 6604
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26344 6458 26372 6598
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 26332 6452 26384 6458
rect 26332 6394 26384 6400
rect 26238 6216 26294 6225
rect 26238 6151 26240 6160
rect 26292 6151 26294 6160
rect 26240 6122 26292 6128
rect 25502 5672 25558 5681
rect 25502 5607 25504 5616
rect 25556 5607 25558 5616
rect 25504 5578 25556 5584
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26344 5370 26372 6394
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26332 3936 26384 3942
rect 26332 3878 26384 3884
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26344 2961 26372 3878
rect 26436 3777 26464 10390
rect 26606 10367 26662 10376
rect 26514 10160 26570 10169
rect 26514 10095 26516 10104
rect 26568 10095 26570 10104
rect 26516 10066 26568 10072
rect 26528 9722 26556 10066
rect 26804 10010 26832 15302
rect 26896 11121 26924 17478
rect 26882 11112 26938 11121
rect 26882 11047 26938 11056
rect 26988 10577 27016 19382
rect 27080 19378 27108 19790
rect 27068 19372 27120 19378
rect 27068 19314 27120 19320
rect 27080 18426 27108 19314
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 27436 14000 27488 14006
rect 27436 13942 27488 13948
rect 27448 13841 27476 13942
rect 27434 13832 27490 13841
rect 27434 13767 27490 13776
rect 27160 12232 27212 12238
rect 27160 12174 27212 12180
rect 27172 11830 27200 12174
rect 27160 11824 27212 11830
rect 27160 11766 27212 11772
rect 27526 11792 27582 11801
rect 27526 11727 27582 11736
rect 27540 10606 27568 11727
rect 27528 10600 27580 10606
rect 26974 10568 27030 10577
rect 27528 10542 27580 10548
rect 26974 10503 27030 10512
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 26804 9982 26924 10010
rect 26792 9920 26844 9926
rect 26792 9862 26844 9868
rect 26516 9716 26568 9722
rect 26516 9658 26568 9664
rect 26698 9344 26754 9353
rect 26698 9279 26754 9288
rect 26712 9178 26740 9279
rect 26700 9172 26752 9178
rect 26700 9114 26752 9120
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8362 26556 8978
rect 26698 8664 26754 8673
rect 26698 8599 26754 8608
rect 26606 8528 26662 8537
rect 26606 8463 26662 8472
rect 26516 8356 26568 8362
rect 26516 8298 26568 8304
rect 26516 7948 26568 7954
rect 26516 7890 26568 7896
rect 26528 7206 26556 7890
rect 26516 7200 26568 7206
rect 26516 7142 26568 7148
rect 26620 6866 26648 8463
rect 26712 8090 26740 8599
rect 26804 8129 26832 9862
rect 26790 8120 26846 8129
rect 26700 8084 26752 8090
rect 26790 8055 26846 8064
rect 26700 8026 26752 8032
rect 26698 7440 26754 7449
rect 26698 7375 26754 7384
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26620 6458 26648 6802
rect 26712 6730 26740 7375
rect 26790 7032 26846 7041
rect 26790 6967 26846 6976
rect 26700 6724 26752 6730
rect 26700 6666 26752 6672
rect 26608 6452 26660 6458
rect 26608 6394 26660 6400
rect 26514 6352 26570 6361
rect 26514 6287 26570 6296
rect 26528 4690 26556 6287
rect 26608 6112 26660 6118
rect 26608 6054 26660 6060
rect 26620 5137 26648 6054
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 26528 4282 26556 4626
rect 26516 4276 26568 4282
rect 26516 4218 26568 4224
rect 26608 3936 26660 3942
rect 26712 3913 26740 5510
rect 26804 4570 26832 6967
rect 26896 6361 26924 9982
rect 27344 9648 27396 9654
rect 27342 9616 27344 9625
rect 27396 9616 27398 9625
rect 27342 9551 27398 9560
rect 26976 8356 27028 8362
rect 26976 8298 27028 8304
rect 26882 6352 26938 6361
rect 26882 6287 26938 6296
rect 26988 5914 27016 8298
rect 27724 6905 27752 10406
rect 27710 6896 27766 6905
rect 27710 6831 27766 6840
rect 26976 5908 27028 5914
rect 26976 5850 27028 5856
rect 27160 5772 27212 5778
rect 27160 5714 27212 5720
rect 27172 5370 27200 5714
rect 27160 5364 27212 5370
rect 27160 5306 27212 5312
rect 26804 4542 26924 4570
rect 26792 4480 26844 4486
rect 26792 4422 26844 4428
rect 26608 3878 26660 3884
rect 26698 3904 26754 3913
rect 26422 3768 26478 3777
rect 26422 3703 26478 3712
rect 26514 3632 26570 3641
rect 26514 3567 26516 3576
rect 26568 3567 26570 3576
rect 26516 3538 26568 3544
rect 26528 3194 26556 3538
rect 26620 3369 26648 3878
rect 26698 3839 26754 3848
rect 26700 3392 26752 3398
rect 26606 3360 26662 3369
rect 26700 3334 26752 3340
rect 26606 3295 26662 3304
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26330 2952 26386 2961
rect 26330 2887 26386 2896
rect 26608 2848 26660 2854
rect 25372 2796 25452 2802
rect 25320 2790 25452 2796
rect 25332 2774 25452 2790
rect 25594 2816 25650 2825
rect 25332 2514 25360 2774
rect 26608 2790 26660 2796
rect 25594 2751 25650 2760
rect 25608 2650 25636 2751
rect 25596 2644 25648 2650
rect 25596 2586 25648 2592
rect 25320 2508 25372 2514
rect 25320 2450 25372 2456
rect 26332 2440 26384 2446
rect 26332 2382 26384 2388
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 26344 480 26372 2382
rect 26620 1465 26648 2790
rect 26712 2145 26740 3334
rect 26698 2136 26754 2145
rect 26698 2071 26754 2080
rect 26606 1456 26662 1465
rect 26606 1391 26662 1400
rect 2410 368 2466 377
rect 2410 303 2466 312
rect 3514 0 3570 480
rect 4894 0 4950 480
rect 6366 0 6422 480
rect 7746 0 7802 480
rect 9218 0 9274 480
rect 10598 0 10654 480
rect 12070 0 12126 480
rect 13450 0 13506 480
rect 14922 0 14978 480
rect 16302 0 16358 480
rect 17774 0 17830 480
rect 19154 0 19210 480
rect 20626 0 20682 480
rect 22006 0 22062 480
rect 23478 0 23534 480
rect 24858 0 24914 480
rect 26330 0 26386 480
rect 26804 377 26832 4422
rect 26896 2990 26924 4542
rect 27710 4448 27766 4457
rect 27710 4383 27766 4392
rect 27528 4072 27580 4078
rect 27526 4040 27528 4049
rect 27580 4040 27582 4049
rect 27526 3975 27582 3984
rect 27724 3942 27752 4383
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 27618 3768 27674 3777
rect 27618 3703 27674 3712
rect 27526 3496 27582 3505
rect 27526 3431 27582 3440
rect 27540 2990 27568 3431
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 26882 2544 26938 2553
rect 27632 2530 27660 3703
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 29182 2816 29238 2825
rect 27724 2689 27752 2790
rect 29182 2751 29238 2760
rect 27710 2680 27766 2689
rect 27710 2615 27766 2624
rect 27632 2502 27752 2530
rect 26882 2479 26884 2488
rect 26936 2479 26938 2488
rect 26884 2450 26936 2456
rect 27068 2304 27120 2310
rect 27068 2246 27120 2252
rect 27080 921 27108 2246
rect 27066 912 27122 921
rect 27066 847 27122 856
rect 27724 480 27752 2502
rect 29196 480 29224 2751
rect 26790 368 26846 377
rect 26790 303 26846 312
rect 27710 0 27766 480
rect 29182 0 29238 480
<< via2 >>
rect 3422 23568 3478 23624
rect 2962 22344 3018 22400
rect 25134 23568 25190 23624
rect 4158 23024 4214 23080
rect 4066 21800 4122 21856
rect 3698 21256 3754 21312
rect 1858 20596 1914 20632
rect 1858 20576 1860 20596
rect 1860 20576 1912 20596
rect 1912 20576 1914 20596
rect 3422 20440 3478 20496
rect 570 16360 626 16416
rect 1582 18264 1638 18320
rect 2134 18128 2190 18184
rect 2134 15952 2190 16008
rect 2318 16788 2374 16824
rect 2318 16768 2320 16788
rect 2320 16768 2372 16788
rect 2372 16768 2374 16788
rect 1490 11464 1546 11520
rect 1398 11056 1454 11112
rect 1582 10376 1638 10432
rect 1582 9868 1584 9888
rect 1584 9868 1636 9888
rect 1636 9868 1638 9888
rect 1582 9832 1638 9868
rect 1582 9324 1584 9344
rect 1584 9324 1636 9344
rect 1636 9324 1638 9344
rect 1582 9288 1638 9324
rect 1490 8608 1546 8664
rect 1582 8064 1638 8120
rect 1398 7384 1454 7440
rect 1582 6840 1638 6896
rect 2134 13368 2190 13424
rect 2318 12844 2374 12880
rect 2318 12824 2320 12844
rect 2320 12824 2372 12844
rect 2372 12824 2374 12844
rect 1950 12280 2006 12336
rect 2318 12280 2374 12336
rect 1950 11056 2006 11112
rect 1766 9968 1822 10024
rect 2042 8492 2098 8528
rect 2042 8472 2044 8492
rect 2044 8472 2096 8492
rect 2096 8472 2098 8492
rect 2134 8336 2190 8392
rect 1950 7248 2006 7304
rect 1674 6296 1730 6352
rect 1582 5636 1638 5672
rect 1582 5616 1584 5636
rect 1584 5616 1636 5636
rect 1636 5616 1638 5636
rect 2042 5228 2098 5264
rect 2042 5208 2044 5228
rect 2044 5208 2096 5228
rect 2096 5208 2098 5228
rect 1582 5072 1638 5128
rect 2502 12144 2558 12200
rect 2410 11348 2466 11384
rect 2410 11328 2412 11348
rect 2412 11328 2464 11348
rect 2464 11328 2466 11348
rect 2410 9036 2466 9072
rect 2410 9016 2412 9036
rect 2412 9016 2464 9036
rect 2464 9016 2466 9036
rect 2410 5772 2466 5808
rect 2410 5752 2412 5772
rect 2412 5752 2464 5772
rect 2464 5752 2466 5772
rect 1398 4528 1454 4584
rect 1950 4528 2006 4584
rect 1582 4428 1584 4448
rect 1584 4428 1636 4448
rect 1636 4428 1638 4448
rect 1582 4392 1638 4428
rect 1582 3884 1584 3904
rect 1584 3884 1636 3904
rect 1636 3884 1638 3904
rect 1582 3848 1638 3884
rect 662 3168 718 3224
rect 1582 2624 1638 2680
rect 1398 2080 1454 2136
rect 1582 1400 1638 1456
rect 2502 4120 2558 4176
rect 2042 4004 2098 4040
rect 2042 3984 2044 4004
rect 2044 3984 2096 4004
rect 2096 3984 2098 4004
rect 2042 3052 2098 3088
rect 2042 3032 2044 3052
rect 2044 3032 2096 3052
rect 2096 3032 2098 3052
rect 1674 856 1730 912
rect 3146 19352 3202 19408
rect 3146 17720 3202 17776
rect 2686 16904 2742 16960
rect 2870 14728 2926 14784
rect 2962 14048 3018 14104
rect 2962 13232 3018 13288
rect 3330 12416 3386 12472
rect 2778 12300 2834 12336
rect 2778 12280 2780 12300
rect 2780 12280 2832 12300
rect 2832 12280 2834 12300
rect 2686 11600 2742 11656
rect 3882 20032 3938 20088
rect 4066 20032 4122 20088
rect 3514 17584 3570 17640
rect 3698 15816 3754 15872
rect 3606 13368 3662 13424
rect 3514 10512 3570 10568
rect 4986 20576 5042 20632
rect 4158 18672 4214 18728
rect 4526 18808 4582 18864
rect 4250 15272 4306 15328
rect 3882 13368 3938 13424
rect 4710 18672 4766 18728
rect 4802 18128 4858 18184
rect 4526 12688 4582 12744
rect 4250 11328 4306 11384
rect 4618 11056 4674 11112
rect 2778 6296 2834 6352
rect 3146 5616 3202 5672
rect 5722 14728 5778 14784
rect 5446 13812 5448 13832
rect 5448 13812 5500 13832
rect 5500 13812 5502 13832
rect 5446 13776 5502 13812
rect 5262 11620 5318 11656
rect 5262 11600 5264 11620
rect 5264 11600 5316 11620
rect 5316 11600 5318 11620
rect 4710 9832 4766 9888
rect 4710 9696 4766 9752
rect 4526 5616 4582 5672
rect 2686 3596 2742 3632
rect 2686 3576 2688 3596
rect 2688 3576 2740 3596
rect 2740 3576 2742 3596
rect 2686 3340 2688 3360
rect 2688 3340 2740 3360
rect 2740 3340 2742 3360
rect 2686 3304 2742 3340
rect 2962 2760 3018 2816
rect 5170 10240 5226 10296
rect 5170 9696 5226 9752
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 6826 20304 6882 20360
rect 5998 20052 6054 20088
rect 5998 20032 6000 20052
rect 6000 20032 6052 20052
rect 6052 20032 6054 20052
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 7746 19896 7802 19952
rect 9862 19896 9918 19952
rect 7654 18828 7710 18864
rect 7654 18808 7656 18828
rect 7656 18808 7708 18828
rect 7708 18808 7710 18828
rect 7838 18400 7894 18456
rect 9310 18284 9366 18320
rect 9310 18264 9312 18284
rect 9312 18264 9364 18284
rect 9364 18264 9366 18284
rect 8022 17584 8078 17640
rect 8022 16940 8024 16960
rect 8024 16940 8076 16960
rect 8076 16940 8078 16960
rect 8022 16904 8078 16940
rect 9126 16652 9182 16688
rect 9126 16632 9128 16652
rect 9128 16632 9180 16652
rect 9180 16632 9182 16652
rect 10230 17040 10286 17096
rect 10414 17040 10470 17096
rect 8850 15408 8906 15464
rect 6274 14864 6330 14920
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5906 10684 5908 10704
rect 5908 10684 5960 10704
rect 5960 10684 5962 10704
rect 5906 10648 5962 10684
rect 5630 10376 5686 10432
rect 6182 9968 6238 10024
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 7194 12416 7250 12472
rect 7102 9560 7158 9616
rect 7010 8880 7066 8936
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 4802 6316 4858 6352
rect 4802 6296 4804 6316
rect 4804 6296 4856 6316
rect 4856 6296 4858 6316
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 5078 7268 5134 7304
rect 5078 7248 5080 7268
rect 5080 7248 5132 7268
rect 5132 7248 5134 7268
rect 6182 7248 6238 7304
rect 5078 6332 5080 6352
rect 5080 6332 5132 6352
rect 5132 6332 5134 6352
rect 5078 6296 5134 6332
rect 6274 6860 6330 6896
rect 6274 6840 6276 6860
rect 6276 6840 6328 6860
rect 6328 6840 6330 6860
rect 5630 6160 5686 6216
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 4802 3848 4858 3904
rect 4342 3440 4398 3496
rect 4710 3576 4766 3632
rect 6274 3984 6330 4040
rect 4894 3712 4950 3768
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 5538 3052 5594 3088
rect 5538 3032 5540 3052
rect 5540 3032 5592 3052
rect 5592 3032 5594 3052
rect 7654 13776 7710 13832
rect 7470 13368 7526 13424
rect 7470 12960 7526 13016
rect 7562 12824 7618 12880
rect 7930 13388 7986 13424
rect 7930 13368 7932 13388
rect 7932 13368 7984 13388
rect 7984 13368 7986 13388
rect 10046 15952 10102 16008
rect 10414 16768 10470 16824
rect 8850 14592 8906 14648
rect 8206 13776 8262 13832
rect 8206 13232 8262 13288
rect 8390 12824 8446 12880
rect 7930 12280 7986 12336
rect 7286 10104 7342 10160
rect 7654 10548 7656 10568
rect 7656 10548 7708 10568
rect 7708 10548 7710 10568
rect 7654 10512 7710 10548
rect 7378 8336 7434 8392
rect 7102 3576 7158 3632
rect 8574 10920 8630 10976
rect 9310 12280 9366 12336
rect 8574 10532 8630 10568
rect 8574 10512 8576 10532
rect 8576 10512 8628 10532
rect 8628 10512 8630 10532
rect 9218 10240 9274 10296
rect 9586 11228 9588 11248
rect 9588 11228 9640 11248
rect 9640 11228 9642 11248
rect 9586 11192 9642 11228
rect 7930 6060 7932 6080
rect 7932 6060 7984 6080
rect 7984 6060 7986 6080
rect 7930 6024 7986 6060
rect 7930 5616 7986 5672
rect 8022 4528 8078 4584
rect 6366 2760 6422 2816
rect 5538 2508 5594 2544
rect 5538 2488 5540 2508
rect 5540 2488 5592 2508
rect 5592 2488 5594 2508
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 10322 15000 10378 15056
rect 10322 14728 10378 14784
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 12070 18264 12126 18320
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 14922 20440 14978 20496
rect 16670 20340 16672 20360
rect 16672 20340 16724 20360
rect 16724 20340 16726 20360
rect 16670 20304 16726 20340
rect 12714 16496 12770 16552
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10782 13796 10838 13832
rect 10782 13776 10784 13796
rect 10784 13776 10836 13796
rect 10836 13776 10838 13796
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 11426 12960 11482 13016
rect 11242 12724 11244 12744
rect 11244 12724 11296 12744
rect 11296 12724 11298 12744
rect 11242 12688 11298 12724
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10782 11872 10838 11928
rect 11426 12688 11482 12744
rect 11334 11736 11390 11792
rect 9862 11056 9918 11112
rect 10138 10512 10194 10568
rect 10230 10412 10232 10432
rect 10232 10412 10284 10432
rect 10284 10412 10286 10432
rect 10230 10376 10286 10412
rect 9678 6024 9734 6080
rect 8390 4564 8392 4584
rect 8392 4564 8444 4584
rect 8444 4564 8446 4584
rect 8390 4528 8446 4564
rect 8206 3848 8262 3904
rect 9862 3596 9918 3632
rect 9862 3576 9864 3596
rect 9864 3576 9916 3596
rect 9916 3576 9918 3596
rect 10138 3168 10194 3224
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10782 8336 10838 8392
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10966 5616 11022 5672
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10230 2896 10286 2952
rect 9954 2488 10010 2544
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 10782 3712 10838 3768
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 11610 12008 11666 12064
rect 12622 12280 12678 12336
rect 12622 11872 12678 11928
rect 12254 11228 12256 11248
rect 12256 11228 12308 11248
rect 12308 11228 12310 11248
rect 12254 11192 12310 11228
rect 11794 8336 11850 8392
rect 11610 5752 11666 5808
rect 12162 7268 12218 7304
rect 12162 7248 12164 7268
rect 12164 7248 12216 7268
rect 12216 7248 12218 7268
rect 12162 6296 12218 6352
rect 12254 6196 12256 6216
rect 12256 6196 12308 6216
rect 12308 6196 12310 6216
rect 12254 6160 12310 6196
rect 12162 6024 12218 6080
rect 12990 15408 13046 15464
rect 12806 14864 12862 14920
rect 12898 11872 12954 11928
rect 19706 20324 19762 20360
rect 19706 20304 19708 20324
rect 19708 20304 19760 20324
rect 19760 20304 19762 20324
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 14646 17040 14702 17096
rect 13450 16632 13506 16688
rect 15842 18672 15898 18728
rect 16486 18536 16542 18592
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15658 17740 15714 17776
rect 15658 17720 15660 17740
rect 15660 17720 15712 17740
rect 15712 17720 15714 17740
rect 16670 18128 16726 18184
rect 16394 17448 16450 17504
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 16026 16632 16082 16688
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15382 15972 15438 16008
rect 15382 15952 15384 15972
rect 15384 15952 15436 15972
rect 15436 15952 15438 15972
rect 14830 12824 14886 12880
rect 13818 12144 13874 12200
rect 15014 12708 15070 12744
rect 15014 12688 15016 12708
rect 15016 12688 15068 12708
rect 15068 12688 15070 12708
rect 15474 13640 15530 13696
rect 15474 12552 15530 12608
rect 13358 9696 13414 9752
rect 13634 9696 13690 9752
rect 13174 7384 13230 7440
rect 13358 6976 13414 7032
rect 13174 5208 13230 5264
rect 11978 4120 12034 4176
rect 13266 3984 13322 4040
rect 15198 12008 15254 12064
rect 15198 11872 15254 11928
rect 15658 13776 15714 13832
rect 16670 17040 16726 17096
rect 18234 17584 18290 17640
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16302 14320 16358 14376
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 16486 13368 16542 13424
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 16026 11464 16082 11520
rect 16302 11328 16358 11384
rect 15750 10920 15806 10976
rect 15014 5888 15070 5944
rect 12254 3440 12310 3496
rect 12714 3440 12770 3496
rect 12070 3168 12126 3224
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 15750 10240 15806 10296
rect 16394 10240 16450 10296
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15566 9016 15622 9072
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 16486 8608 16542 8664
rect 16118 8372 16120 8392
rect 16120 8372 16172 8392
rect 16172 8372 16174 8392
rect 16118 8336 16174 8372
rect 15750 7792 15806 7848
rect 15566 6976 15622 7032
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 16394 7520 16450 7576
rect 17314 15272 17370 15328
rect 18602 15272 18658 15328
rect 18878 17484 18880 17504
rect 18880 17484 18932 17504
rect 18932 17484 18934 17504
rect 18878 17448 18934 17484
rect 18786 17176 18842 17232
rect 20074 18164 20076 18184
rect 20076 18164 20128 18184
rect 20128 18164 20130 18184
rect 20074 18128 20130 18164
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 20810 20440 20866 20496
rect 23202 20304 23258 20360
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 21270 18672 21326 18728
rect 21638 18300 21640 18320
rect 21640 18300 21692 18320
rect 21692 18300 21694 18320
rect 21638 18264 21694 18300
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 23662 18808 23718 18864
rect 23570 18536 23626 18592
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 19338 16224 19394 16280
rect 18786 15544 18842 15600
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 19246 15408 19302 15464
rect 18694 14456 18750 14512
rect 16854 11192 16910 11248
rect 17222 10784 17278 10840
rect 17222 10512 17278 10568
rect 17866 10104 17922 10160
rect 16762 7384 16818 7440
rect 17774 7112 17830 7168
rect 16486 6568 16542 6624
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 17682 6740 17684 6760
rect 17684 6740 17736 6760
rect 17736 6740 17738 6760
rect 17682 6704 17738 6740
rect 17958 6024 18014 6080
rect 19154 13640 19210 13696
rect 19338 13368 19394 13424
rect 19154 12960 19210 13016
rect 18970 12844 19026 12880
rect 18970 12824 18972 12844
rect 18972 12824 19024 12844
rect 19024 12824 19026 12844
rect 18878 12708 18934 12744
rect 18878 12688 18880 12708
rect 18880 12688 18932 12708
rect 18932 12688 18934 12708
rect 18970 9016 19026 9072
rect 18326 8900 18382 8936
rect 18326 8880 18328 8900
rect 18328 8880 18380 8900
rect 18380 8880 18382 8900
rect 19430 12552 19486 12608
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 19982 12824 20038 12880
rect 19706 12552 19762 12608
rect 18510 7812 18566 7848
rect 18510 7792 18512 7812
rect 18512 7792 18564 7812
rect 18564 7792 18566 7812
rect 18510 7384 18566 7440
rect 18510 6860 18566 6896
rect 18510 6840 18512 6860
rect 18512 6840 18564 6860
rect 18564 6840 18566 6860
rect 18234 6296 18290 6352
rect 18050 4528 18106 4584
rect 17958 3984 18014 4040
rect 18234 3984 18290 4040
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15014 2760 15070 2816
rect 16302 2760 16358 2816
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 18418 3848 18474 3904
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20258 12280 20314 12336
rect 19614 8336 19670 8392
rect 19614 6432 19670 6488
rect 19522 4528 19578 4584
rect 19982 4664 20038 4720
rect 20718 11872 20774 11928
rect 20718 11600 20774 11656
rect 20718 11464 20774 11520
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 20810 11328 20866 11384
rect 21362 10684 21364 10704
rect 21364 10684 21416 10704
rect 21416 10684 21418 10704
rect 21362 10648 21418 10684
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 21362 9016 21418 9072
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 20902 3984 20958 4040
rect 20810 3848 20866 3904
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 20442 3576 20498 3632
rect 19982 2488 20038 2544
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 22282 13368 22338 13424
rect 22006 12960 22062 13016
rect 22926 12860 22928 12880
rect 22928 12860 22980 12880
rect 22980 12860 22982 12880
rect 22926 12824 22982 12860
rect 22834 12688 22890 12744
rect 21822 11328 21878 11384
rect 22282 11328 22338 11384
rect 21638 9424 21694 9480
rect 22650 9580 22706 9616
rect 22650 9560 22652 9580
rect 22652 9560 22704 9580
rect 22704 9560 22706 9580
rect 21822 9016 21878 9072
rect 23938 17448 23994 17504
rect 24122 17176 24178 17232
rect 24306 15544 24362 15600
rect 24122 15272 24178 15328
rect 24398 14864 24454 14920
rect 24306 11756 24362 11792
rect 24306 11736 24308 11756
rect 24308 11736 24360 11756
rect 24360 11736 24362 11756
rect 24306 10532 24362 10568
rect 24306 10512 24308 10532
rect 24308 10512 24360 10532
rect 24360 10512 24362 10532
rect 23846 8628 23902 8664
rect 23846 8608 23848 8628
rect 23848 8608 23900 8628
rect 23900 8608 23902 8628
rect 24214 8472 24270 8528
rect 23570 7384 23626 7440
rect 24398 8084 24454 8120
rect 24398 8064 24400 8084
rect 24400 8064 24452 8084
rect 24452 8064 24454 8084
rect 24306 7520 24362 7576
rect 21730 5364 21786 5400
rect 21730 5344 21732 5364
rect 21732 5344 21784 5364
rect 21784 5344 21786 5364
rect 21638 4564 21640 4584
rect 21640 4564 21692 4584
rect 21692 4564 21694 4584
rect 21638 4528 21694 4564
rect 21822 4020 21824 4040
rect 21824 4020 21876 4040
rect 21876 4020 21878 4040
rect 21822 3984 21878 4020
rect 23570 4700 23572 4720
rect 23572 4700 23624 4720
rect 23624 4700 23626 4720
rect 23570 4664 23626 4700
rect 23662 3032 23718 3088
rect 24674 16496 24730 16552
rect 24766 16244 24822 16280
rect 24766 16224 24768 16244
rect 24768 16224 24820 16244
rect 24820 16224 24822 16244
rect 24582 15408 24638 15464
rect 24674 14592 24730 14648
rect 24766 13912 24822 13968
rect 25042 13776 25098 13832
rect 24766 12280 24822 12336
rect 24674 9460 24676 9480
rect 24676 9460 24728 9480
rect 24728 9460 24730 9480
rect 24674 9424 24730 9460
rect 24674 6296 24730 6352
rect 25410 23024 25466 23080
rect 26974 21800 27030 21856
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25226 21256 25282 21312
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25686 20440 25742 20496
rect 25410 19352 25466 19408
rect 25318 18808 25374 18864
rect 25502 18808 25558 18864
rect 25410 18536 25466 18592
rect 25226 15408 25282 15464
rect 25226 10784 25282 10840
rect 24858 9424 24914 9480
rect 25042 6976 25098 7032
rect 25594 18264 25650 18320
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25502 13368 25558 13424
rect 25410 12688 25466 12744
rect 25502 12280 25558 12336
rect 24858 6452 24914 6488
rect 25318 6568 25374 6624
rect 24858 6432 24860 6452
rect 24860 6432 24912 6452
rect 24912 6432 24914 6452
rect 24858 4548 24914 4584
rect 24858 4528 24860 4548
rect 24860 4528 24912 4548
rect 24912 4528 24914 4548
rect 25870 17584 25926 17640
rect 25778 16088 25834 16144
rect 25778 14456 25834 14512
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25686 13776 25742 13832
rect 25870 14320 25926 14376
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25778 13368 25834 13424
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 26514 18672 26570 18728
rect 26514 17176 26570 17232
rect 26698 11600 26754 11656
rect 26514 11212 26570 11248
rect 26514 11192 26516 11212
rect 26516 11192 26568 11212
rect 26568 11192 26570 11212
rect 26422 10648 26478 10704
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26054 9596 26056 9616
rect 26056 9596 26108 9616
rect 26108 9596 26110 9616
rect 26054 9560 26110 9596
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25962 7148 25964 7168
rect 25964 7148 26016 7168
rect 26016 7148 26018 7168
rect 25962 7112 26018 7148
rect 25594 6704 25650 6760
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26238 6180 26294 6216
rect 26238 6160 26240 6180
rect 26240 6160 26292 6180
rect 26292 6160 26294 6180
rect 25502 5636 25558 5672
rect 25502 5616 25504 5636
rect 25504 5616 25556 5636
rect 25556 5616 25558 5636
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26606 10412 26608 10432
rect 26608 10412 26660 10432
rect 26660 10412 26662 10432
rect 26606 10376 26662 10412
rect 26514 10124 26570 10160
rect 26514 10104 26516 10124
rect 26516 10104 26568 10124
rect 26568 10104 26570 10124
rect 26882 11056 26938 11112
rect 27434 13776 27490 13832
rect 27526 11736 27582 11792
rect 26974 10512 27030 10568
rect 26698 9288 26754 9344
rect 26698 8608 26754 8664
rect 26606 8472 26662 8528
rect 26790 8064 26846 8120
rect 26698 7384 26754 7440
rect 26790 6976 26846 7032
rect 26514 6296 26570 6352
rect 26606 5072 26662 5128
rect 27342 9596 27344 9616
rect 27344 9596 27396 9616
rect 27396 9596 27398 9616
rect 27342 9560 27398 9596
rect 26882 6296 26938 6352
rect 27710 6840 27766 6896
rect 26422 3712 26478 3768
rect 26514 3596 26570 3632
rect 26514 3576 26516 3596
rect 26516 3576 26568 3596
rect 26568 3576 26570 3596
rect 26698 3848 26754 3904
rect 26606 3304 26662 3360
rect 26330 2896 26386 2952
rect 25594 2760 25650 2816
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 26698 2080 26754 2136
rect 26606 1400 26662 1456
rect 2410 312 2466 368
rect 27710 4392 27766 4448
rect 27526 4020 27528 4040
rect 27528 4020 27580 4040
rect 27580 4020 27582 4040
rect 27526 3984 27582 4020
rect 27618 3712 27674 3768
rect 27526 3440 27582 3496
rect 26882 2508 26938 2544
rect 26882 2488 26884 2508
rect 26884 2488 26936 2508
rect 26936 2488 26938 2508
rect 29182 2760 29238 2816
rect 27710 2624 27766 2680
rect 27066 856 27122 912
rect 26790 312 26846 368
<< metal3 >>
rect 0 23626 480 23656
rect 3417 23626 3483 23629
rect 0 23624 3483 23626
rect 0 23568 3422 23624
rect 3478 23568 3483 23624
rect 0 23566 3483 23568
rect 0 23536 480 23566
rect 3417 23563 3483 23566
rect 25129 23626 25195 23629
rect 29520 23626 30000 23656
rect 25129 23624 30000 23626
rect 25129 23568 25134 23624
rect 25190 23568 30000 23624
rect 25129 23566 30000 23568
rect 25129 23563 25195 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 4153 23082 4219 23085
rect 0 23080 4219 23082
rect 0 23024 4158 23080
rect 4214 23024 4219 23080
rect 0 23022 4219 23024
rect 0 22992 480 23022
rect 4153 23019 4219 23022
rect 25405 23082 25471 23085
rect 29520 23082 30000 23112
rect 25405 23080 30000 23082
rect 25405 23024 25410 23080
rect 25466 23024 30000 23080
rect 25405 23022 30000 23024
rect 25405 23019 25471 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2957 22402 3023 22405
rect 0 22400 3023 22402
rect 0 22344 2962 22400
rect 3018 22344 3023 22400
rect 0 22342 3023 22344
rect 0 22312 480 22342
rect 2957 22339 3023 22342
rect 25446 22340 25452 22404
rect 25516 22402 25522 22404
rect 29520 22402 30000 22432
rect 25516 22342 30000 22402
rect 25516 22340 25522 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 4061 21858 4127 21861
rect 0 21856 4127 21858
rect 0 21800 4066 21856
rect 4122 21800 4127 21856
rect 0 21798 4127 21800
rect 0 21768 480 21798
rect 4061 21795 4127 21798
rect 26969 21858 27035 21861
rect 29520 21858 30000 21888
rect 26969 21856 30000 21858
rect 26969 21800 26974 21856
rect 27030 21800 30000 21856
rect 26969 21798 30000 21800
rect 26969 21795 27035 21798
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 29520 21768 30000 21798
rect 25944 21727 26264 21728
rect 0 21314 480 21344
rect 3693 21314 3759 21317
rect 0 21312 3759 21314
rect 0 21256 3698 21312
rect 3754 21256 3759 21312
rect 0 21254 3759 21256
rect 0 21224 480 21254
rect 3693 21251 3759 21254
rect 25221 21314 25287 21317
rect 29520 21314 30000 21344
rect 25221 21312 30000 21314
rect 25221 21256 25226 21312
rect 25282 21256 30000 21312
rect 25221 21254 30000 21256
rect 25221 21251 25287 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 1853 20634 1919 20637
rect 4981 20634 5047 20637
rect 29520 20634 30000 20664
rect 0 20574 1778 20634
rect 0 20544 480 20574
rect 1718 20498 1778 20574
rect 1853 20632 5047 20634
rect 1853 20576 1858 20632
rect 1914 20576 4986 20632
rect 5042 20576 5047 20632
rect 1853 20574 5047 20576
rect 1853 20571 1919 20574
rect 4981 20571 5047 20574
rect 26374 20574 30000 20634
rect 3417 20498 3483 20501
rect 1718 20496 3483 20498
rect 1718 20440 3422 20496
rect 3478 20440 3483 20496
rect 1718 20438 3483 20440
rect 3417 20435 3483 20438
rect 14917 20498 14983 20501
rect 20805 20498 20871 20501
rect 14917 20496 20871 20498
rect 14917 20440 14922 20496
rect 14978 20440 20810 20496
rect 20866 20440 20871 20496
rect 14917 20438 20871 20440
rect 14917 20435 14983 20438
rect 20805 20435 20871 20438
rect 25681 20498 25747 20501
rect 26374 20498 26434 20574
rect 29520 20544 30000 20574
rect 25681 20496 26434 20498
rect 25681 20440 25686 20496
rect 25742 20440 26434 20496
rect 25681 20438 26434 20440
rect 25681 20435 25747 20438
rect 6821 20362 6887 20365
rect 16665 20362 16731 20365
rect 6821 20360 16731 20362
rect 6821 20304 6826 20360
rect 6882 20304 16670 20360
rect 16726 20304 16731 20360
rect 6821 20302 16731 20304
rect 6821 20299 6887 20302
rect 16665 20299 16731 20302
rect 19701 20362 19767 20365
rect 23197 20362 23263 20365
rect 19701 20360 23263 20362
rect 19701 20304 19706 20360
rect 19762 20304 23202 20360
rect 23258 20304 23263 20360
rect 19701 20302 23263 20304
rect 19701 20299 19767 20302
rect 23197 20299 23263 20302
rect 10944 20160 11264 20161
rect 0 20090 480 20120
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 3877 20090 3943 20093
rect 0 20088 3943 20090
rect 0 20032 3882 20088
rect 3938 20032 3943 20088
rect 0 20030 3943 20032
rect 0 20000 480 20030
rect 3877 20027 3943 20030
rect 4061 20090 4127 20093
rect 5993 20090 6059 20093
rect 4061 20088 6059 20090
rect 4061 20032 4066 20088
rect 4122 20032 5998 20088
rect 6054 20032 6059 20088
rect 4061 20030 6059 20032
rect 4061 20027 4127 20030
rect 5993 20027 6059 20030
rect 24894 20028 24900 20092
rect 24964 20090 24970 20092
rect 29520 20090 30000 20120
rect 24964 20030 30000 20090
rect 24964 20028 24970 20030
rect 29520 20000 30000 20030
rect 7741 19954 7807 19957
rect 9857 19954 9923 19957
rect 7741 19952 9923 19954
rect 7741 19896 7746 19952
rect 7802 19896 9862 19952
rect 9918 19896 9923 19952
rect 7741 19894 9923 19896
rect 7741 19891 7807 19894
rect 9857 19891 9923 19894
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 0 19410 480 19440
rect 3141 19410 3207 19413
rect 0 19408 3207 19410
rect 0 19352 3146 19408
rect 3202 19352 3207 19408
rect 0 19350 3207 19352
rect 0 19320 480 19350
rect 3141 19347 3207 19350
rect 25405 19410 25471 19413
rect 29520 19410 30000 19440
rect 25405 19408 30000 19410
rect 25405 19352 25410 19408
rect 25466 19352 30000 19408
rect 25405 19350 30000 19352
rect 25405 19347 25471 19350
rect 29520 19320 30000 19350
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 0 18866 480 18896
rect 4521 18866 4587 18869
rect 0 18864 4587 18866
rect 0 18808 4526 18864
rect 4582 18808 4587 18864
rect 0 18806 4587 18808
rect 0 18776 480 18806
rect 4521 18803 4587 18806
rect 7649 18866 7715 18869
rect 23657 18866 23723 18869
rect 25313 18866 25379 18869
rect 7649 18864 25379 18866
rect 7649 18808 7654 18864
rect 7710 18808 23662 18864
rect 23718 18808 25318 18864
rect 25374 18808 25379 18864
rect 7649 18806 25379 18808
rect 7649 18803 7715 18806
rect 23657 18803 23723 18806
rect 25313 18803 25379 18806
rect 25497 18866 25563 18869
rect 29520 18866 30000 18896
rect 25497 18864 30000 18866
rect 25497 18808 25502 18864
rect 25558 18808 30000 18864
rect 25497 18806 30000 18808
rect 25497 18803 25563 18806
rect 29520 18776 30000 18806
rect 4153 18730 4219 18733
rect 4705 18730 4771 18733
rect 15837 18730 15903 18733
rect 21265 18730 21331 18733
rect 26509 18730 26575 18733
rect 4153 18728 26575 18730
rect 4153 18672 4158 18728
rect 4214 18672 4710 18728
rect 4766 18672 15842 18728
rect 15898 18672 21270 18728
rect 21326 18672 26514 18728
rect 26570 18672 26575 18728
rect 4153 18670 26575 18672
rect 4153 18667 4219 18670
rect 4705 18667 4771 18670
rect 15837 18667 15903 18670
rect 21265 18667 21331 18670
rect 26509 18667 26575 18670
rect 16481 18594 16547 18597
rect 23565 18594 23631 18597
rect 25405 18594 25471 18597
rect 16481 18592 25471 18594
rect 16481 18536 16486 18592
rect 16542 18536 23570 18592
rect 23626 18536 25410 18592
rect 25466 18536 25471 18592
rect 16481 18534 25471 18536
rect 16481 18531 16547 18534
rect 23565 18531 23631 18534
rect 25405 18531 25471 18534
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 7833 18458 7899 18461
rect 7833 18456 12266 18458
rect 7833 18400 7838 18456
rect 7894 18400 12266 18456
rect 7833 18398 12266 18400
rect 7833 18395 7899 18398
rect 0 18322 480 18352
rect 1577 18322 1643 18325
rect 0 18320 1643 18322
rect 0 18264 1582 18320
rect 1638 18264 1643 18320
rect 0 18262 1643 18264
rect 0 18232 480 18262
rect 1577 18259 1643 18262
rect 9305 18322 9371 18325
rect 12065 18322 12131 18325
rect 9305 18320 12131 18322
rect 9305 18264 9310 18320
rect 9366 18264 12070 18320
rect 12126 18264 12131 18320
rect 9305 18262 12131 18264
rect 12206 18322 12266 18398
rect 21633 18322 21699 18325
rect 25589 18322 25655 18325
rect 29520 18322 30000 18352
rect 12206 18320 30000 18322
rect 12206 18264 21638 18320
rect 21694 18264 25594 18320
rect 25650 18264 30000 18320
rect 12206 18262 30000 18264
rect 9305 18259 9371 18262
rect 12065 18259 12131 18262
rect 21633 18259 21699 18262
rect 25589 18259 25655 18262
rect 29520 18232 30000 18262
rect 2129 18186 2195 18189
rect 4797 18186 4863 18189
rect 16665 18186 16731 18189
rect 20069 18186 20135 18189
rect 2129 18184 20135 18186
rect 2129 18128 2134 18184
rect 2190 18128 4802 18184
rect 4858 18128 16670 18184
rect 16726 18128 20074 18184
rect 20130 18128 20135 18184
rect 2129 18126 20135 18128
rect 2129 18123 2195 18126
rect 4797 18123 4863 18126
rect 16665 18123 16731 18126
rect 20069 18123 20135 18126
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 3141 17778 3207 17781
rect 15653 17778 15719 17781
rect 3141 17776 15719 17778
rect 3141 17720 3146 17776
rect 3202 17720 15658 17776
rect 15714 17720 15719 17776
rect 3141 17718 15719 17720
rect 3141 17715 3207 17718
rect 15653 17715 15719 17718
rect 0 17642 480 17672
rect 3509 17642 3575 17645
rect 0 17640 3575 17642
rect 0 17584 3514 17640
rect 3570 17584 3575 17640
rect 0 17582 3575 17584
rect 0 17552 480 17582
rect 3509 17579 3575 17582
rect 8017 17642 8083 17645
rect 18229 17642 18295 17645
rect 8017 17640 18295 17642
rect 8017 17584 8022 17640
rect 8078 17584 18234 17640
rect 18290 17584 18295 17640
rect 8017 17582 18295 17584
rect 8017 17579 8083 17582
rect 18229 17579 18295 17582
rect 25865 17642 25931 17645
rect 29520 17642 30000 17672
rect 25865 17640 30000 17642
rect 25865 17584 25870 17640
rect 25926 17584 30000 17640
rect 25865 17582 30000 17584
rect 25865 17579 25931 17582
rect 29520 17552 30000 17582
rect 16389 17506 16455 17509
rect 18873 17506 18939 17509
rect 23933 17506 23999 17509
rect 16389 17504 23999 17506
rect 16389 17448 16394 17504
rect 16450 17448 18878 17504
rect 18934 17448 23938 17504
rect 23994 17448 23999 17504
rect 16389 17446 23999 17448
rect 16389 17443 16455 17446
rect 18873 17443 18939 17446
rect 23933 17443 23999 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 18781 17234 18847 17237
rect 24117 17234 24183 17237
rect 26509 17234 26575 17237
rect 18781 17232 26575 17234
rect 9308 17140 9874 17200
rect 18781 17176 18786 17232
rect 18842 17176 24122 17232
rect 24178 17176 26514 17232
rect 26570 17176 26575 17232
rect 18781 17174 26575 17176
rect 18781 17171 18847 17174
rect 24117 17171 24183 17174
rect 26509 17171 26575 17174
rect 0 17098 480 17128
rect 9308 17098 9368 17140
rect 0 17038 9368 17098
rect 9814 17098 9874 17140
rect 10225 17098 10291 17101
rect 9814 17096 10291 17098
rect 9814 17040 10230 17096
rect 10286 17040 10291 17096
rect 9814 17038 10291 17040
rect 0 17008 480 17038
rect 10225 17035 10291 17038
rect 10409 17098 10475 17101
rect 14641 17098 14707 17101
rect 10409 17096 14707 17098
rect 10409 17040 10414 17096
rect 10470 17040 14646 17096
rect 14702 17040 14707 17096
rect 10409 17038 14707 17040
rect 10409 17035 10475 17038
rect 14641 17035 14707 17038
rect 16665 17098 16731 17101
rect 29520 17098 30000 17128
rect 16665 17096 30000 17098
rect 16665 17040 16670 17096
rect 16726 17040 30000 17096
rect 16665 17038 30000 17040
rect 16665 17035 16731 17038
rect 29520 17008 30000 17038
rect 2681 16962 2747 16965
rect 8017 16962 8083 16965
rect 2681 16960 8083 16962
rect 2681 16904 2686 16960
rect 2742 16904 8022 16960
rect 8078 16904 8083 16960
rect 2681 16902 8083 16904
rect 2681 16899 2747 16902
rect 8017 16899 8083 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 2313 16826 2379 16829
rect 10409 16826 10475 16829
rect 2313 16824 10475 16826
rect 2313 16768 2318 16824
rect 2374 16768 10414 16824
rect 10470 16768 10475 16824
rect 2313 16766 10475 16768
rect 2313 16763 2379 16766
rect 10409 16763 10475 16766
rect 9121 16690 9187 16693
rect 13445 16690 13511 16693
rect 16021 16690 16087 16693
rect 9121 16688 12266 16690
rect 9121 16632 9126 16688
rect 9182 16632 12266 16688
rect 9121 16630 12266 16632
rect 9121 16627 9187 16630
rect 12206 16554 12266 16630
rect 13445 16688 16087 16690
rect 13445 16632 13450 16688
rect 13506 16632 16026 16688
rect 16082 16632 16087 16688
rect 13445 16630 16087 16632
rect 13445 16627 13511 16630
rect 16021 16627 16087 16630
rect 12709 16554 12775 16557
rect 24669 16554 24735 16557
rect 12206 16552 24735 16554
rect 12206 16496 12714 16552
rect 12770 16496 24674 16552
rect 24730 16496 24735 16552
rect 12206 16494 24735 16496
rect 12709 16491 12775 16494
rect 24669 16491 24735 16494
rect 0 16418 480 16448
rect 565 16418 631 16421
rect 29520 16418 30000 16448
rect 0 16416 631 16418
rect 0 16360 570 16416
rect 626 16360 631 16416
rect 0 16358 631 16360
rect 0 16328 480 16358
rect 565 16355 631 16358
rect 26374 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 19333 16282 19399 16285
rect 24761 16282 24827 16285
rect 19333 16280 24827 16282
rect 19333 16224 19338 16280
rect 19394 16224 24766 16280
rect 24822 16224 24827 16280
rect 19333 16222 24827 16224
rect 19333 16219 19399 16222
rect 24761 16219 24827 16222
rect 25773 16146 25839 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 25773 16144 26434 16146
rect 25773 16088 25778 16144
rect 25834 16088 26434 16144
rect 25773 16086 26434 16088
rect 25773 16083 25839 16086
rect 2129 16010 2195 16013
rect 10041 16010 10107 16013
rect 15377 16010 15443 16013
rect 2129 16008 15443 16010
rect 2129 15952 2134 16008
rect 2190 15952 10046 16008
rect 10102 15952 15382 16008
rect 15438 15952 15443 16008
rect 2129 15950 15443 15952
rect 2129 15947 2195 15950
rect 10041 15947 10107 15950
rect 15377 15947 15443 15950
rect 0 15874 480 15904
rect 3693 15874 3759 15877
rect 0 15872 3759 15874
rect 0 15816 3698 15872
rect 3754 15816 3759 15872
rect 0 15814 3759 15816
rect 0 15784 480 15814
rect 3693 15811 3759 15814
rect 25078 15812 25084 15876
rect 25148 15874 25154 15876
rect 29520 15874 30000 15904
rect 25148 15814 30000 15874
rect 25148 15812 25154 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 18781 15602 18847 15605
rect 24301 15602 24367 15605
rect 18781 15600 24367 15602
rect 18781 15544 18786 15600
rect 18842 15544 24306 15600
rect 24362 15544 24367 15600
rect 18781 15542 24367 15544
rect 18781 15539 18847 15542
rect 24301 15539 24367 15542
rect 8845 15466 8911 15469
rect 12985 15466 13051 15469
rect 19241 15466 19307 15469
rect 24577 15466 24643 15469
rect 8845 15464 18890 15466
rect 8845 15408 8850 15464
rect 8906 15408 12990 15464
rect 13046 15408 18890 15464
rect 8845 15406 18890 15408
rect 8845 15403 8911 15406
rect 12985 15403 13051 15406
rect 0 15330 480 15360
rect 4245 15330 4311 15333
rect 17309 15330 17375 15333
rect 18597 15330 18663 15333
rect 0 15328 4311 15330
rect 0 15272 4250 15328
rect 4306 15272 4311 15328
rect 0 15270 4311 15272
rect 0 15240 480 15270
rect 4245 15267 4311 15270
rect 16438 15328 18663 15330
rect 16438 15272 17314 15328
rect 17370 15272 18602 15328
rect 18658 15272 18663 15328
rect 16438 15270 18663 15272
rect 18830 15330 18890 15406
rect 19241 15464 24643 15466
rect 19241 15408 19246 15464
rect 19302 15408 24582 15464
rect 24638 15408 24643 15464
rect 19241 15406 24643 15408
rect 19241 15403 19307 15406
rect 24577 15403 24643 15406
rect 25221 15466 25287 15469
rect 25221 15464 26434 15466
rect 25221 15408 25226 15464
rect 25282 15408 26434 15464
rect 25221 15406 26434 15408
rect 25221 15403 25287 15406
rect 24117 15330 24183 15333
rect 18830 15328 24183 15330
rect 18830 15272 24122 15328
rect 24178 15272 24183 15328
rect 18830 15270 24183 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 10317 15058 10383 15061
rect 16438 15058 16498 15270
rect 17309 15267 17375 15270
rect 18597 15267 18663 15270
rect 24117 15267 24183 15270
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 10317 15056 16498 15058
rect 10317 15000 10322 15056
rect 10378 15000 16498 15056
rect 10317 14998 16498 15000
rect 10317 14995 10383 14998
rect 6269 14922 6335 14925
rect 12801 14922 12867 14925
rect 24393 14922 24459 14925
rect 6269 14920 24459 14922
rect 6269 14864 6274 14920
rect 6330 14864 12806 14920
rect 12862 14864 24398 14920
rect 24454 14864 24459 14920
rect 6269 14862 24459 14864
rect 6269 14859 6335 14862
rect 12801 14859 12867 14862
rect 24393 14859 24459 14862
rect 2865 14786 2931 14789
rect 5717 14786 5783 14789
rect 10317 14786 10383 14789
rect 2865 14784 10383 14786
rect 2865 14728 2870 14784
rect 2926 14728 5722 14784
rect 5778 14728 10322 14784
rect 10378 14728 10383 14784
rect 2865 14726 10383 14728
rect 2865 14723 2931 14726
rect 5717 14723 5783 14726
rect 10317 14723 10383 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 8845 14650 8911 14653
rect 0 14648 8911 14650
rect 0 14592 8850 14648
rect 8906 14592 8911 14648
rect 0 14590 8911 14592
rect 0 14560 480 14590
rect 8845 14587 8911 14590
rect 24669 14650 24735 14653
rect 29520 14650 30000 14680
rect 24669 14648 30000 14650
rect 24669 14592 24674 14648
rect 24730 14592 30000 14648
rect 24669 14590 30000 14592
rect 24669 14587 24735 14590
rect 29520 14560 30000 14590
rect 18689 14514 18755 14517
rect 25773 14514 25839 14517
rect 18689 14512 25839 14514
rect 18689 14456 18694 14512
rect 18750 14456 25778 14512
rect 25834 14456 25839 14512
rect 18689 14454 25839 14456
rect 18689 14451 18755 14454
rect 25773 14451 25839 14454
rect 16297 14378 16363 14381
rect 25865 14378 25931 14381
rect 16297 14376 25931 14378
rect 16297 14320 16302 14376
rect 16358 14320 25870 14376
rect 25926 14320 25931 14376
rect 16297 14318 25931 14320
rect 16297 14315 16363 14318
rect 25865 14315 25931 14318
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 2957 14106 3023 14109
rect 29520 14106 30000 14136
rect 0 14104 3023 14106
rect 0 14048 2962 14104
rect 3018 14048 3023 14104
rect 0 14046 3023 14048
rect 0 14016 480 14046
rect 2957 14043 3023 14046
rect 26374 14046 30000 14106
rect 24761 13970 24827 13973
rect 26374 13970 26434 14046
rect 29520 14016 30000 14046
rect 24761 13968 26434 13970
rect 24761 13912 24766 13968
rect 24822 13912 26434 13968
rect 24761 13910 26434 13912
rect 24761 13907 24827 13910
rect 5441 13834 5507 13837
rect 7649 13834 7715 13837
rect 5441 13832 7715 13834
rect 5441 13776 5446 13832
rect 5502 13776 7654 13832
rect 7710 13776 7715 13832
rect 5441 13774 7715 13776
rect 5441 13771 5507 13774
rect 7649 13771 7715 13774
rect 8201 13834 8267 13837
rect 10777 13834 10843 13837
rect 8201 13832 10843 13834
rect 8201 13776 8206 13832
rect 8262 13776 10782 13832
rect 10838 13776 10843 13832
rect 8201 13774 10843 13776
rect 8201 13771 8267 13774
rect 10777 13771 10843 13774
rect 15653 13834 15719 13837
rect 25037 13834 25103 13837
rect 25681 13834 25747 13837
rect 27429 13834 27495 13837
rect 15653 13832 15762 13834
rect 15653 13776 15658 13832
rect 15714 13776 15762 13832
rect 15653 13771 15762 13776
rect 25037 13832 27495 13834
rect 25037 13776 25042 13832
rect 25098 13776 25686 13832
rect 25742 13776 27434 13832
rect 27490 13776 27495 13832
rect 25037 13774 27495 13776
rect 25037 13771 25103 13774
rect 25681 13771 25747 13774
rect 27429 13771 27495 13774
rect 15469 13698 15535 13701
rect 15702 13698 15762 13771
rect 19149 13698 19215 13701
rect 15469 13696 19215 13698
rect 15469 13640 15474 13696
rect 15530 13640 19154 13696
rect 19210 13640 19215 13696
rect 15469 13638 19215 13640
rect 15469 13635 15535 13638
rect 19149 13635 19215 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 0 13426 480 13456
rect 2129 13426 2195 13429
rect 3601 13426 3667 13429
rect 0 13424 3667 13426
rect 0 13368 2134 13424
rect 2190 13368 3606 13424
rect 3662 13368 3667 13424
rect 0 13366 3667 13368
rect 0 13336 480 13366
rect 2129 13363 2195 13366
rect 3601 13363 3667 13366
rect 3877 13426 3943 13429
rect 7465 13426 7531 13429
rect 3877 13424 7531 13426
rect 3877 13368 3882 13424
rect 3938 13368 7470 13424
rect 7526 13368 7531 13424
rect 3877 13366 7531 13368
rect 3877 13363 3943 13366
rect 7465 13363 7531 13366
rect 7925 13426 7991 13429
rect 16481 13426 16547 13429
rect 19333 13426 19399 13429
rect 22277 13426 22343 13429
rect 7925 13424 22343 13426
rect 7925 13368 7930 13424
rect 7986 13368 16486 13424
rect 16542 13368 19338 13424
rect 19394 13368 22282 13424
rect 22338 13368 22343 13424
rect 7925 13366 22343 13368
rect 7925 13363 7991 13366
rect 16481 13363 16547 13366
rect 19333 13363 19399 13366
rect 22277 13363 22343 13366
rect 25497 13426 25563 13429
rect 25773 13426 25839 13429
rect 29520 13426 30000 13456
rect 25497 13424 30000 13426
rect 25497 13368 25502 13424
rect 25558 13368 25778 13424
rect 25834 13368 30000 13424
rect 25497 13366 30000 13368
rect 25497 13363 25563 13366
rect 25773 13363 25839 13366
rect 29520 13336 30000 13366
rect 2957 13290 3023 13293
rect 8201 13290 8267 13293
rect 2957 13288 8267 13290
rect 2957 13232 2962 13288
rect 3018 13232 8206 13288
rect 8262 13232 8267 13288
rect 2957 13230 8267 13232
rect 2957 13227 3023 13230
rect 8201 13227 8267 13230
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 7465 13018 7531 13021
rect 11421 13018 11487 13021
rect 7465 13016 11487 13018
rect 7465 12960 7470 13016
rect 7526 12960 11426 13016
rect 11482 12960 11487 13016
rect 7465 12958 11487 12960
rect 7465 12955 7531 12958
rect 11421 12955 11487 12958
rect 19149 13018 19215 13021
rect 22001 13018 22067 13021
rect 19149 13016 22067 13018
rect 19149 12960 19154 13016
rect 19210 12960 22006 13016
rect 22062 12960 22067 13016
rect 19149 12958 22067 12960
rect 19149 12955 19215 12958
rect 22001 12955 22067 12958
rect 0 12882 480 12912
rect 2313 12882 2379 12885
rect 7557 12882 7623 12885
rect 0 12880 7623 12882
rect 0 12824 2318 12880
rect 2374 12824 7562 12880
rect 7618 12824 7623 12880
rect 0 12822 7623 12824
rect 0 12792 480 12822
rect 2313 12819 2379 12822
rect 7557 12819 7623 12822
rect 8385 12882 8451 12885
rect 14825 12882 14891 12885
rect 18965 12882 19031 12885
rect 19977 12882 20043 12885
rect 8385 12880 20043 12882
rect 8385 12824 8390 12880
rect 8446 12824 14830 12880
rect 14886 12824 18970 12880
rect 19026 12824 19982 12880
rect 20038 12824 20043 12880
rect 8385 12822 20043 12824
rect 8385 12819 8451 12822
rect 14825 12819 14891 12822
rect 18965 12819 19031 12822
rect 19977 12819 20043 12822
rect 22921 12882 22987 12885
rect 29520 12882 30000 12912
rect 22921 12880 30000 12882
rect 22921 12824 22926 12880
rect 22982 12824 30000 12880
rect 22921 12822 30000 12824
rect 22921 12819 22987 12822
rect 29520 12792 30000 12822
rect 4521 12746 4587 12749
rect 11237 12746 11303 12749
rect 4521 12744 11303 12746
rect 4521 12688 4526 12744
rect 4582 12688 11242 12744
rect 11298 12688 11303 12744
rect 4521 12686 11303 12688
rect 4521 12683 4587 12686
rect 11237 12683 11303 12686
rect 11421 12746 11487 12749
rect 15009 12746 15075 12749
rect 11421 12744 15075 12746
rect 11421 12688 11426 12744
rect 11482 12688 15014 12744
rect 15070 12688 15075 12744
rect 11421 12686 15075 12688
rect 11421 12683 11487 12686
rect 15009 12683 15075 12686
rect 18873 12746 18939 12749
rect 22829 12746 22895 12749
rect 25405 12746 25471 12749
rect 18873 12744 22895 12746
rect 18873 12688 18878 12744
rect 18934 12688 22834 12744
rect 22890 12688 22895 12744
rect 18873 12686 22895 12688
rect 18873 12683 18939 12686
rect 22829 12683 22895 12686
rect 24902 12744 25471 12746
rect 24902 12688 25410 12744
rect 25466 12688 25471 12744
rect 24902 12686 25471 12688
rect 15469 12610 15535 12613
rect 11470 12608 15535 12610
rect 11470 12552 15474 12608
rect 15530 12552 15535 12608
rect 11470 12550 15535 12552
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 3325 12474 3391 12477
rect 7189 12474 7255 12477
rect 3325 12472 7255 12474
rect 3325 12416 3330 12472
rect 3386 12416 7194 12472
rect 7250 12416 7255 12472
rect 3325 12414 7255 12416
rect 3325 12411 3391 12414
rect 7189 12411 7255 12414
rect 0 12338 480 12368
rect 1945 12338 2011 12341
rect 0 12336 2011 12338
rect 0 12280 1950 12336
rect 2006 12280 2011 12336
rect 0 12278 2011 12280
rect 0 12248 480 12278
rect 1945 12275 2011 12278
rect 2313 12338 2379 12341
rect 2773 12338 2839 12341
rect 7925 12338 7991 12341
rect 9305 12338 9371 12341
rect 11470 12338 11530 12550
rect 15469 12547 15535 12550
rect 19425 12610 19491 12613
rect 19701 12610 19767 12613
rect 19425 12608 19767 12610
rect 19425 12552 19430 12608
rect 19486 12552 19706 12608
rect 19762 12552 19767 12608
rect 19425 12550 19767 12552
rect 19425 12547 19491 12550
rect 19701 12547 19767 12550
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 2313 12336 11530 12338
rect 2313 12280 2318 12336
rect 2374 12280 2778 12336
rect 2834 12280 7930 12336
rect 7986 12280 9310 12336
rect 9366 12280 11530 12336
rect 2313 12278 11530 12280
rect 12617 12338 12683 12341
rect 20253 12338 20319 12341
rect 24761 12338 24827 12341
rect 12617 12336 24827 12338
rect 12617 12280 12622 12336
rect 12678 12280 20258 12336
rect 20314 12280 24766 12336
rect 24822 12280 24827 12336
rect 12617 12278 24827 12280
rect 24902 12338 24962 12686
rect 25405 12683 25471 12686
rect 25497 12338 25563 12341
rect 29520 12338 30000 12368
rect 24902 12336 30000 12338
rect 24902 12280 25502 12336
rect 25558 12280 30000 12336
rect 24902 12278 30000 12280
rect 2313 12275 2379 12278
rect 2773 12275 2839 12278
rect 7925 12275 7991 12278
rect 9305 12275 9371 12278
rect 12617 12275 12683 12278
rect 20253 12275 20319 12278
rect 24761 12275 24827 12278
rect 25497 12275 25563 12278
rect 29520 12248 30000 12278
rect 2497 12202 2563 12205
rect 13813 12202 13879 12205
rect 2497 12200 13879 12202
rect 2497 12144 2502 12200
rect 2558 12144 13818 12200
rect 13874 12144 13879 12200
rect 2497 12142 13879 12144
rect 2497 12139 2563 12142
rect 13813 12139 13879 12142
rect 11605 12066 11671 12069
rect 15193 12066 15259 12069
rect 11605 12064 15259 12066
rect 11605 12008 11610 12064
rect 11666 12008 15198 12064
rect 15254 12008 15259 12064
rect 11605 12006 15259 12008
rect 11605 12003 11671 12006
rect 15193 12003 15259 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 10777 11930 10843 11933
rect 12617 11930 12683 11933
rect 10777 11928 12683 11930
rect 10777 11872 10782 11928
rect 10838 11872 12622 11928
rect 12678 11872 12683 11928
rect 10777 11870 12683 11872
rect 10777 11867 10843 11870
rect 12617 11867 12683 11870
rect 12893 11930 12959 11933
rect 15193 11930 15259 11933
rect 12893 11928 15259 11930
rect 12893 11872 12898 11928
rect 12954 11872 15198 11928
rect 15254 11872 15259 11928
rect 12893 11870 15259 11872
rect 12893 11867 12959 11870
rect 15193 11867 15259 11870
rect 20713 11930 20779 11933
rect 25630 11930 25636 11932
rect 20713 11928 25636 11930
rect 20713 11872 20718 11928
rect 20774 11872 25636 11928
rect 20713 11870 25636 11872
rect 20713 11867 20779 11870
rect 25630 11868 25636 11870
rect 25700 11868 25706 11932
rect 11329 11794 11395 11797
rect 24301 11794 24367 11797
rect 27521 11794 27587 11797
rect 11329 11792 27587 11794
rect 11329 11736 11334 11792
rect 11390 11736 24306 11792
rect 24362 11736 27526 11792
rect 27582 11736 27587 11792
rect 11329 11734 27587 11736
rect 11329 11731 11395 11734
rect 24301 11731 24367 11734
rect 27521 11731 27587 11734
rect 0 11658 480 11688
rect 2681 11658 2747 11661
rect 5257 11658 5323 11661
rect 20713 11658 20779 11661
rect 0 11656 2747 11658
rect 0 11600 2686 11656
rect 2742 11600 2747 11656
rect 0 11598 2747 11600
rect 0 11568 480 11598
rect 2681 11595 2747 11598
rect 5214 11656 20779 11658
rect 5214 11600 5262 11656
rect 5318 11600 20718 11656
rect 20774 11600 20779 11656
rect 5214 11598 20779 11600
rect 5214 11595 5323 11598
rect 20713 11595 20779 11598
rect 26693 11658 26759 11661
rect 29520 11658 30000 11688
rect 26693 11656 30000 11658
rect 26693 11600 26698 11656
rect 26754 11600 30000 11656
rect 26693 11598 30000 11600
rect 26693 11595 26759 11598
rect 1485 11522 1551 11525
rect 5214 11522 5274 11595
rect 29520 11568 30000 11598
rect 1485 11520 5274 11522
rect 1485 11464 1490 11520
rect 1546 11464 5274 11520
rect 1485 11462 5274 11464
rect 16021 11522 16087 11525
rect 20713 11522 20779 11525
rect 16021 11520 20779 11522
rect 16021 11464 16026 11520
rect 16082 11464 20718 11520
rect 20774 11464 20779 11520
rect 16021 11462 20779 11464
rect 1485 11459 1551 11462
rect 16021 11459 16087 11462
rect 20713 11459 20779 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 2405 11386 2471 11389
rect 4245 11386 4311 11389
rect 2405 11384 4311 11386
rect 2405 11328 2410 11384
rect 2466 11328 4250 11384
rect 4306 11328 4311 11384
rect 2405 11326 4311 11328
rect 2405 11323 2471 11326
rect 4245 11323 4311 11326
rect 16297 11386 16363 11389
rect 20805 11386 20871 11389
rect 16297 11384 20871 11386
rect 16297 11328 16302 11384
rect 16358 11328 20810 11384
rect 20866 11328 20871 11384
rect 16297 11326 20871 11328
rect 16297 11323 16363 11326
rect 20805 11323 20871 11326
rect 21817 11386 21883 11389
rect 22277 11386 22343 11389
rect 24894 11386 24900 11388
rect 21817 11384 24900 11386
rect 21817 11328 21822 11384
rect 21878 11328 22282 11384
rect 22338 11328 24900 11384
rect 21817 11326 24900 11328
rect 21817 11323 21883 11326
rect 22277 11323 22343 11326
rect 24894 11324 24900 11326
rect 24964 11324 24970 11388
rect 9581 11250 9647 11253
rect 12249 11250 12315 11253
rect 9581 11248 12315 11250
rect 9581 11192 9586 11248
rect 9642 11192 12254 11248
rect 12310 11192 12315 11248
rect 9581 11190 12315 11192
rect 9581 11187 9647 11190
rect 12249 11187 12315 11190
rect 16849 11250 16915 11253
rect 26509 11250 26575 11253
rect 16849 11248 26575 11250
rect 16849 11192 16854 11248
rect 16910 11192 26514 11248
rect 26570 11192 26575 11248
rect 16849 11190 26575 11192
rect 16849 11187 16915 11190
rect 26509 11187 26575 11190
rect 0 11114 480 11144
rect 1393 11114 1459 11117
rect 0 11112 1459 11114
rect 0 11056 1398 11112
rect 1454 11056 1459 11112
rect 0 11054 1459 11056
rect 0 11024 480 11054
rect 1393 11051 1459 11054
rect 1945 11114 2011 11117
rect 4613 11114 4679 11117
rect 9857 11114 9923 11117
rect 1945 11112 9923 11114
rect 1945 11056 1950 11112
rect 2006 11056 4618 11112
rect 4674 11056 9862 11112
rect 9918 11056 9923 11112
rect 1945 11054 9923 11056
rect 1945 11051 2011 11054
rect 4613 11051 4679 11054
rect 9857 11051 9923 11054
rect 26877 11114 26943 11117
rect 29520 11114 30000 11144
rect 26877 11112 30000 11114
rect 26877 11056 26882 11112
rect 26938 11056 30000 11112
rect 26877 11054 30000 11056
rect 26877 11051 26943 11054
rect 29520 11024 30000 11054
rect 8569 10978 8635 10981
rect 15745 10978 15811 10981
rect 8569 10976 15811 10978
rect 8569 10920 8574 10976
rect 8630 10920 15750 10976
rect 15806 10920 15811 10976
rect 8569 10918 15811 10920
rect 8569 10915 8635 10918
rect 15745 10915 15811 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 17217 10842 17283 10845
rect 25221 10842 25287 10845
rect 17217 10840 25287 10842
rect 17217 10784 17222 10840
rect 17278 10784 25226 10840
rect 25282 10784 25287 10840
rect 17217 10782 25287 10784
rect 17217 10779 17283 10782
rect 25221 10779 25287 10782
rect 5901 10706 5967 10709
rect 21357 10706 21423 10709
rect 26417 10706 26483 10709
rect 5901 10704 26483 10706
rect 5901 10648 5906 10704
rect 5962 10648 21362 10704
rect 21418 10648 26422 10704
rect 26478 10648 26483 10704
rect 5901 10646 26483 10648
rect 5901 10643 5967 10646
rect 21357 10643 21423 10646
rect 26417 10643 26483 10646
rect 3509 10570 3575 10573
rect 7649 10570 7715 10573
rect 8569 10570 8635 10573
rect 3509 10568 8635 10570
rect 3509 10512 3514 10568
rect 3570 10512 7654 10568
rect 7710 10512 8574 10568
rect 8630 10512 8635 10568
rect 3509 10510 8635 10512
rect 3509 10507 3575 10510
rect 7649 10507 7715 10510
rect 8569 10507 8635 10510
rect 10133 10570 10199 10573
rect 17217 10570 17283 10573
rect 24301 10570 24367 10573
rect 26969 10570 27035 10573
rect 10133 10568 17283 10570
rect 10133 10512 10138 10568
rect 10194 10512 17222 10568
rect 17278 10512 17283 10568
rect 10133 10510 17283 10512
rect 10133 10507 10199 10510
rect 17217 10507 17283 10510
rect 17358 10568 27035 10570
rect 17358 10512 24306 10568
rect 24362 10512 26974 10568
rect 27030 10512 27035 10568
rect 17358 10510 27035 10512
rect 0 10434 480 10464
rect 1577 10434 1643 10437
rect 0 10432 1643 10434
rect 0 10376 1582 10432
rect 1638 10376 1643 10432
rect 0 10374 1643 10376
rect 0 10344 480 10374
rect 1577 10371 1643 10374
rect 5625 10434 5691 10437
rect 10225 10434 10291 10437
rect 5625 10432 10291 10434
rect 5625 10376 5630 10432
rect 5686 10376 10230 10432
rect 10286 10376 10291 10432
rect 5625 10374 10291 10376
rect 5625 10371 5691 10374
rect 10225 10371 10291 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 5165 10298 5231 10301
rect 9213 10298 9279 10301
rect 5165 10296 9279 10298
rect 5165 10240 5170 10296
rect 5226 10240 9218 10296
rect 9274 10240 9279 10296
rect 5165 10238 9279 10240
rect 5165 10235 5231 10238
rect 9213 10235 9279 10238
rect 15745 10298 15811 10301
rect 16389 10298 16455 10301
rect 15745 10296 16455 10298
rect 15745 10240 15750 10296
rect 15806 10240 16394 10296
rect 16450 10240 16455 10296
rect 15745 10238 16455 10240
rect 15745 10235 15811 10238
rect 16389 10235 16455 10238
rect 7281 10162 7347 10165
rect 17358 10162 17418 10510
rect 24301 10507 24367 10510
rect 26969 10507 27035 10510
rect 26601 10434 26667 10437
rect 29520 10434 30000 10464
rect 26601 10432 30000 10434
rect 26601 10376 26606 10432
rect 26662 10376 30000 10432
rect 26601 10374 30000 10376
rect 26601 10371 26667 10374
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 7281 10160 17418 10162
rect 7281 10104 7286 10160
rect 7342 10104 17418 10160
rect 7281 10102 17418 10104
rect 17861 10162 17927 10165
rect 26509 10162 26575 10165
rect 17861 10160 26575 10162
rect 17861 10104 17866 10160
rect 17922 10104 26514 10160
rect 26570 10104 26575 10160
rect 17861 10102 26575 10104
rect 7281 10099 7347 10102
rect 17861 10099 17927 10102
rect 26509 10099 26575 10102
rect 1761 10026 1827 10029
rect 6177 10026 6243 10029
rect 1761 10024 6243 10026
rect 1761 9968 1766 10024
rect 1822 9968 6182 10024
rect 6238 9968 6243 10024
rect 1761 9966 6243 9968
rect 1761 9963 1827 9966
rect 6177 9963 6243 9966
rect 0 9890 480 9920
rect 1577 9890 1643 9893
rect 0 9888 1643 9890
rect 0 9832 1582 9888
rect 1638 9832 1643 9888
rect 0 9830 1643 9832
rect 0 9800 480 9830
rect 1577 9827 1643 9830
rect 4705 9890 4771 9893
rect 29520 9890 30000 9920
rect 4705 9888 5412 9890
rect 4705 9832 4710 9888
rect 4766 9832 5412 9888
rect 4705 9830 5412 9832
rect 4705 9827 4771 9830
rect 4705 9754 4771 9757
rect 5165 9754 5231 9757
rect 4705 9752 5231 9754
rect 4705 9696 4710 9752
rect 4766 9696 5170 9752
rect 5226 9696 5231 9752
rect 4705 9694 5231 9696
rect 4705 9691 4771 9694
rect 5165 9691 5231 9694
rect 5352 9618 5412 9830
rect 27478 9830 30000 9890
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 9759 26264 9760
rect 13353 9754 13419 9757
rect 13629 9754 13695 9757
rect 13353 9752 13695 9754
rect 13353 9696 13358 9752
rect 13414 9696 13634 9752
rect 13690 9696 13695 9752
rect 13353 9694 13695 9696
rect 13353 9691 13419 9694
rect 13629 9691 13695 9694
rect 7097 9618 7163 9621
rect 5352 9616 7163 9618
rect 5352 9560 7102 9616
rect 7158 9560 7163 9616
rect 5352 9558 7163 9560
rect 7097 9555 7163 9558
rect 22645 9618 22711 9621
rect 26049 9618 26115 9621
rect 22645 9616 26115 9618
rect 22645 9560 22650 9616
rect 22706 9560 26054 9616
rect 26110 9560 26115 9616
rect 22645 9558 26115 9560
rect 22645 9555 22711 9558
rect 26049 9555 26115 9558
rect 27337 9618 27403 9621
rect 27478 9618 27538 9830
rect 29520 9800 30000 9830
rect 27337 9616 27538 9618
rect 27337 9560 27342 9616
rect 27398 9560 27538 9616
rect 27337 9558 27538 9560
rect 27337 9555 27403 9558
rect 21633 9482 21699 9485
rect 24669 9482 24735 9485
rect 24853 9482 24919 9485
rect 21633 9480 24919 9482
rect 21633 9424 21638 9480
rect 21694 9424 24674 9480
rect 24730 9424 24858 9480
rect 24914 9424 24919 9480
rect 21633 9422 24919 9424
rect 21633 9419 21699 9422
rect 24669 9419 24735 9422
rect 24853 9419 24919 9422
rect 0 9346 480 9376
rect 1577 9346 1643 9349
rect 0 9344 1643 9346
rect 0 9288 1582 9344
rect 1638 9288 1643 9344
rect 0 9286 1643 9288
rect 0 9256 480 9286
rect 1577 9283 1643 9286
rect 26693 9346 26759 9349
rect 29520 9346 30000 9376
rect 26693 9344 30000 9346
rect 26693 9288 26698 9344
rect 26754 9288 30000 9344
rect 26693 9286 30000 9288
rect 26693 9283 26759 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 2405 9074 2471 9077
rect 15561 9074 15627 9077
rect 2405 9072 15627 9074
rect 2405 9016 2410 9072
rect 2466 9016 15566 9072
rect 15622 9016 15627 9072
rect 2405 9014 15627 9016
rect 2405 9011 2471 9014
rect 15561 9011 15627 9014
rect 18965 9074 19031 9077
rect 21357 9074 21423 9077
rect 21817 9074 21883 9077
rect 18965 9072 21883 9074
rect 18965 9016 18970 9072
rect 19026 9016 21362 9072
rect 21418 9016 21822 9072
rect 21878 9016 21883 9072
rect 18965 9014 21883 9016
rect 18965 9011 19031 9014
rect 21357 9011 21423 9014
rect 21817 9011 21883 9014
rect 7005 8938 7071 8941
rect 18321 8938 18387 8941
rect 7005 8936 18387 8938
rect 7005 8880 7010 8936
rect 7066 8880 18326 8936
rect 18382 8880 18387 8936
rect 7005 8878 18387 8880
rect 7005 8875 7071 8878
rect 18321 8875 18387 8878
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 1485 8666 1551 8669
rect 0 8664 1551 8666
rect 0 8608 1490 8664
rect 1546 8608 1551 8664
rect 0 8606 1551 8608
rect 0 8576 480 8606
rect 1485 8603 1551 8606
rect 16481 8666 16547 8669
rect 23841 8666 23907 8669
rect 26693 8666 26759 8669
rect 29520 8666 30000 8696
rect 16481 8664 25882 8666
rect 16481 8608 16486 8664
rect 16542 8608 23846 8664
rect 23902 8608 25882 8664
rect 16481 8606 25882 8608
rect 16481 8603 16547 8606
rect 23841 8603 23907 8606
rect 2037 8530 2103 8533
rect 24209 8530 24275 8533
rect 2037 8528 24275 8530
rect 2037 8472 2042 8528
rect 2098 8472 24214 8528
rect 24270 8472 24275 8528
rect 2037 8470 24275 8472
rect 25822 8530 25882 8606
rect 26693 8664 30000 8666
rect 26693 8608 26698 8664
rect 26754 8608 30000 8664
rect 26693 8606 30000 8608
rect 26693 8603 26759 8606
rect 29520 8576 30000 8606
rect 26601 8530 26667 8533
rect 25822 8528 26667 8530
rect 25822 8472 26606 8528
rect 26662 8472 26667 8528
rect 25822 8470 26667 8472
rect 2037 8467 2103 8470
rect 24209 8467 24275 8470
rect 26601 8467 26667 8470
rect 2129 8394 2195 8397
rect 7373 8394 7439 8397
rect 10777 8394 10843 8397
rect 2129 8392 10843 8394
rect 2129 8336 2134 8392
rect 2190 8336 7378 8392
rect 7434 8336 10782 8392
rect 10838 8336 10843 8392
rect 2129 8334 10843 8336
rect 2129 8331 2195 8334
rect 7373 8331 7439 8334
rect 10777 8331 10843 8334
rect 11789 8394 11855 8397
rect 16113 8394 16179 8397
rect 19609 8394 19675 8397
rect 11789 8392 19675 8394
rect 11789 8336 11794 8392
rect 11850 8336 16118 8392
rect 16174 8336 19614 8392
rect 19670 8336 19675 8392
rect 11789 8334 19675 8336
rect 11789 8331 11855 8334
rect 16113 8331 16179 8334
rect 19609 8331 19675 8334
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 1577 8122 1643 8125
rect 0 8120 1643 8122
rect 0 8064 1582 8120
rect 1638 8064 1643 8120
rect 0 8062 1643 8064
rect 0 8032 480 8062
rect 1577 8059 1643 8062
rect 24393 8122 24459 8125
rect 25078 8122 25084 8124
rect 24393 8120 25084 8122
rect 24393 8064 24398 8120
rect 24454 8064 25084 8120
rect 24393 8062 25084 8064
rect 24393 8059 24459 8062
rect 25078 8060 25084 8062
rect 25148 8060 25154 8124
rect 26785 8122 26851 8125
rect 29520 8122 30000 8152
rect 26785 8120 30000 8122
rect 26785 8064 26790 8120
rect 26846 8064 30000 8120
rect 26785 8062 30000 8064
rect 26785 8059 26851 8062
rect 29520 8032 30000 8062
rect 15745 7850 15811 7853
rect 18505 7850 18571 7853
rect 15745 7848 18571 7850
rect 15745 7792 15750 7848
rect 15806 7792 18510 7848
rect 18566 7792 18571 7848
rect 15745 7790 18571 7792
rect 15745 7787 15811 7790
rect 18505 7787 18571 7790
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 16389 7578 16455 7581
rect 24301 7578 24367 7581
rect 16389 7576 24367 7578
rect 16389 7520 16394 7576
rect 16450 7520 24306 7576
rect 24362 7520 24367 7576
rect 16389 7518 24367 7520
rect 16389 7515 16455 7518
rect 24301 7515 24367 7518
rect 0 7442 480 7472
rect 1393 7442 1459 7445
rect 0 7440 1459 7442
rect 0 7384 1398 7440
rect 1454 7384 1459 7440
rect 0 7382 1459 7384
rect 0 7352 480 7382
rect 1393 7379 1459 7382
rect 13169 7442 13235 7445
rect 16757 7442 16823 7445
rect 13169 7440 16823 7442
rect 13169 7384 13174 7440
rect 13230 7384 16762 7440
rect 16818 7384 16823 7440
rect 13169 7382 16823 7384
rect 13169 7379 13235 7382
rect 16757 7379 16823 7382
rect 18505 7442 18571 7445
rect 23565 7442 23631 7445
rect 18505 7440 23631 7442
rect 18505 7384 18510 7440
rect 18566 7384 23570 7440
rect 23626 7384 23631 7440
rect 18505 7382 23631 7384
rect 18505 7379 18571 7382
rect 23565 7379 23631 7382
rect 26693 7442 26759 7445
rect 29520 7442 30000 7472
rect 26693 7440 30000 7442
rect 26693 7384 26698 7440
rect 26754 7384 30000 7440
rect 26693 7382 30000 7384
rect 26693 7379 26759 7382
rect 29520 7352 30000 7382
rect 1945 7306 2011 7309
rect 5073 7306 5139 7309
rect 1945 7304 5139 7306
rect 1945 7248 1950 7304
rect 2006 7248 5078 7304
rect 5134 7248 5139 7304
rect 1945 7246 5139 7248
rect 1945 7243 2011 7246
rect 5073 7243 5139 7246
rect 6177 7306 6243 7309
rect 12157 7306 12223 7309
rect 6177 7304 17740 7306
rect 6177 7248 6182 7304
rect 6238 7248 12162 7304
rect 12218 7248 17740 7304
rect 6177 7246 17740 7248
rect 6177 7243 6243 7246
rect 12157 7243 12223 7246
rect 17680 7204 17740 7246
rect 20670 7212 21466 7272
rect 17680 7173 17786 7204
rect 17680 7170 17835 7173
rect 20670 7170 20730 7212
rect 17642 7168 20730 7170
rect 17642 7112 17774 7168
rect 17830 7112 20730 7168
rect 17642 7110 20730 7112
rect 21406 7170 21466 7212
rect 25957 7170 26023 7173
rect 21406 7168 26023 7170
rect 21406 7112 25962 7168
rect 26018 7112 26023 7168
rect 21406 7110 26023 7112
rect 17769 7107 17835 7110
rect 25957 7107 26023 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 13353 7034 13419 7037
rect 15561 7034 15627 7037
rect 13353 7032 15627 7034
rect 13353 6976 13358 7032
rect 13414 6976 15566 7032
rect 15622 6976 15627 7032
rect 13353 6974 15627 6976
rect 13353 6971 13419 6974
rect 15561 6971 15627 6974
rect 25037 7034 25103 7037
rect 26785 7034 26851 7037
rect 25037 7032 26851 7034
rect 25037 6976 25042 7032
rect 25098 6976 26790 7032
rect 26846 6976 26851 7032
rect 25037 6974 26851 6976
rect 25037 6971 25103 6974
rect 26785 6971 26851 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 6269 6898 6335 6901
rect 18505 6898 18571 6901
rect 6269 6896 18571 6898
rect 6269 6840 6274 6896
rect 6330 6840 18510 6896
rect 18566 6840 18571 6896
rect 6269 6838 18571 6840
rect 6269 6835 6335 6838
rect 18505 6835 18571 6838
rect 27705 6898 27771 6901
rect 29520 6898 30000 6928
rect 27705 6896 30000 6898
rect 27705 6840 27710 6896
rect 27766 6840 30000 6896
rect 27705 6838 30000 6840
rect 27705 6835 27771 6838
rect 29520 6808 30000 6838
rect 17677 6762 17743 6765
rect 25589 6762 25655 6765
rect 17677 6760 25655 6762
rect 17677 6704 17682 6760
rect 17738 6704 25594 6760
rect 25650 6704 25655 6760
rect 17677 6702 25655 6704
rect 17677 6699 17743 6702
rect 25589 6699 25655 6702
rect 16481 6626 16547 6629
rect 25313 6626 25379 6629
rect 16481 6624 25379 6626
rect 16481 6568 16486 6624
rect 16542 6568 25318 6624
rect 25374 6568 25379 6624
rect 16481 6566 25379 6568
rect 16481 6563 16547 6566
rect 25313 6563 25379 6566
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 19609 6490 19675 6493
rect 24853 6490 24919 6493
rect 19609 6488 25882 6490
rect 19609 6432 19614 6488
rect 19670 6432 24858 6488
rect 24914 6432 25882 6488
rect 19609 6430 25882 6432
rect 19609 6427 19675 6430
rect 24853 6427 24919 6430
rect 0 6354 480 6384
rect 1669 6354 1735 6357
rect 0 6352 1735 6354
rect 0 6296 1674 6352
rect 1730 6296 1735 6352
rect 0 6294 1735 6296
rect 0 6264 480 6294
rect 1669 6291 1735 6294
rect 2773 6354 2839 6357
rect 4797 6354 4863 6357
rect 2773 6352 4863 6354
rect 2773 6296 2778 6352
rect 2834 6296 4802 6352
rect 4858 6296 4863 6352
rect 2773 6294 4863 6296
rect 2773 6291 2839 6294
rect 4797 6291 4863 6294
rect 5073 6354 5139 6357
rect 12157 6354 12223 6357
rect 5073 6352 12223 6354
rect 5073 6296 5078 6352
rect 5134 6296 12162 6352
rect 12218 6296 12223 6352
rect 5073 6294 12223 6296
rect 5073 6291 5139 6294
rect 12157 6291 12223 6294
rect 18229 6354 18295 6357
rect 24669 6354 24735 6357
rect 18229 6352 24735 6354
rect 18229 6296 18234 6352
rect 18290 6296 24674 6352
rect 24730 6296 24735 6352
rect 18229 6294 24735 6296
rect 25822 6354 25882 6430
rect 26509 6354 26575 6357
rect 25822 6352 26575 6354
rect 25822 6296 26514 6352
rect 26570 6296 26575 6352
rect 25822 6294 26575 6296
rect 18229 6291 18295 6294
rect 24669 6291 24735 6294
rect 26509 6291 26575 6294
rect 26877 6354 26943 6357
rect 29520 6354 30000 6384
rect 26877 6352 30000 6354
rect 26877 6296 26882 6352
rect 26938 6296 30000 6352
rect 26877 6294 30000 6296
rect 26877 6291 26943 6294
rect 29520 6264 30000 6294
rect 5625 6218 5691 6221
rect 12249 6218 12315 6221
rect 26233 6218 26299 6221
rect 5625 6216 12315 6218
rect 5625 6160 5630 6216
rect 5686 6160 12254 6216
rect 12310 6160 12315 6216
rect 5625 6158 12315 6160
rect 5625 6155 5691 6158
rect 12249 6155 12315 6158
rect 12574 6158 17970 6218
rect 7925 6082 7991 6085
rect 9673 6082 9739 6085
rect 7925 6080 9739 6082
rect 7925 6024 7930 6080
rect 7986 6024 9678 6080
rect 9734 6024 9739 6080
rect 7925 6022 9739 6024
rect 7925 6019 7991 6022
rect 9673 6019 9739 6022
rect 12157 6082 12223 6085
rect 12574 6082 12634 6158
rect 12157 6080 12634 6082
rect 12157 6024 12162 6080
rect 12218 6024 12634 6080
rect 12157 6022 12634 6024
rect 17910 6085 17970 6158
rect 18830 6216 26299 6218
rect 18830 6160 26238 6216
rect 26294 6160 26299 6216
rect 18830 6158 26299 6160
rect 17910 6080 18019 6085
rect 17910 6024 17958 6080
rect 18014 6024 18019 6080
rect 17910 6022 18019 6024
rect 12157 6019 12223 6022
rect 17953 6019 18019 6022
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 15009 5946 15075 5949
rect 18830 5946 18890 6158
rect 26233 6155 26299 6158
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 15009 5944 18890 5946
rect 15009 5888 15014 5944
rect 15070 5888 18890 5944
rect 15009 5886 18890 5888
rect 15009 5883 15075 5886
rect 2405 5810 2471 5813
rect 11605 5810 11671 5813
rect 2405 5808 11671 5810
rect 2405 5752 2410 5808
rect 2466 5752 11610 5808
rect 11666 5752 11671 5808
rect 2405 5750 11671 5752
rect 2405 5747 2471 5750
rect 11605 5747 11671 5750
rect 0 5674 480 5704
rect 1577 5674 1643 5677
rect 0 5672 1643 5674
rect 0 5616 1582 5672
rect 1638 5616 1643 5672
rect 0 5614 1643 5616
rect 0 5584 480 5614
rect 1577 5611 1643 5614
rect 3141 5674 3207 5677
rect 4521 5674 4587 5677
rect 3141 5672 4587 5674
rect 3141 5616 3146 5672
rect 3202 5616 4526 5672
rect 4582 5616 4587 5672
rect 3141 5614 4587 5616
rect 3141 5611 3207 5614
rect 4521 5611 4587 5614
rect 7925 5674 7991 5677
rect 10961 5674 11027 5677
rect 17902 5674 17908 5676
rect 7925 5672 17908 5674
rect 7925 5616 7930 5672
rect 7986 5616 10966 5672
rect 11022 5616 17908 5672
rect 7925 5614 17908 5616
rect 7925 5611 7991 5614
rect 10961 5611 11027 5614
rect 17902 5612 17908 5614
rect 17972 5612 17978 5676
rect 25497 5674 25563 5677
rect 29520 5674 30000 5704
rect 25497 5672 30000 5674
rect 25497 5616 25502 5672
rect 25558 5616 30000 5672
rect 25497 5614 30000 5616
rect 25497 5611 25563 5614
rect 29520 5584 30000 5614
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 17902 5340 17908 5404
rect 17972 5402 17978 5404
rect 21725 5402 21791 5405
rect 17972 5400 21791 5402
rect 17972 5344 21730 5400
rect 21786 5344 21791 5400
rect 17972 5342 21791 5344
rect 17972 5340 17978 5342
rect 21725 5339 21791 5342
rect 2037 5266 2103 5269
rect 13169 5266 13235 5269
rect 2037 5264 13235 5266
rect 2037 5208 2042 5264
rect 2098 5208 13174 5264
rect 13230 5208 13235 5264
rect 2037 5206 13235 5208
rect 2037 5203 2103 5206
rect 13169 5203 13235 5206
rect 0 5130 480 5160
rect 1577 5130 1643 5133
rect 0 5128 1643 5130
rect 0 5072 1582 5128
rect 1638 5072 1643 5128
rect 0 5070 1643 5072
rect 0 5040 480 5070
rect 1577 5067 1643 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 19977 4722 20043 4725
rect 23565 4722 23631 4725
rect 19977 4720 23631 4722
rect 19977 4664 19982 4720
rect 20038 4664 23570 4720
rect 23626 4664 23631 4720
rect 19977 4662 23631 4664
rect 19977 4659 20043 4662
rect 23565 4659 23631 4662
rect 1393 4586 1459 4589
rect 1945 4586 2011 4589
rect 8017 4586 8083 4589
rect 8385 4586 8451 4589
rect 18045 4586 18111 4589
rect 19517 4586 19583 4589
rect 1393 4584 19583 4586
rect 1393 4528 1398 4584
rect 1454 4528 1950 4584
rect 2006 4528 8022 4584
rect 8078 4528 8390 4584
rect 8446 4528 18050 4584
rect 18106 4528 19522 4584
rect 19578 4528 19583 4584
rect 1393 4526 19583 4528
rect 1393 4523 1459 4526
rect 1945 4523 2011 4526
rect 8017 4523 8083 4526
rect 8385 4523 8451 4526
rect 18045 4523 18111 4526
rect 19517 4523 19583 4526
rect 21633 4586 21699 4589
rect 24853 4586 24919 4589
rect 21633 4584 24919 4586
rect 21633 4528 21638 4584
rect 21694 4528 24858 4584
rect 24914 4528 24919 4584
rect 21633 4526 24919 4528
rect 21633 4523 21699 4526
rect 24853 4523 24919 4526
rect 0 4450 480 4480
rect 1577 4450 1643 4453
rect 0 4448 1643 4450
rect 0 4392 1582 4448
rect 1638 4392 1643 4448
rect 0 4390 1643 4392
rect 0 4360 480 4390
rect 1577 4387 1643 4390
rect 27705 4450 27771 4453
rect 29520 4450 30000 4480
rect 27705 4448 30000 4450
rect 27705 4392 27710 4448
rect 27766 4392 30000 4448
rect 27705 4390 30000 4392
rect 27705 4387 27771 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 2497 4178 2563 4181
rect 11973 4178 12039 4181
rect 2497 4176 12039 4178
rect 2497 4120 2502 4176
rect 2558 4120 11978 4176
rect 12034 4120 12039 4176
rect 2497 4118 12039 4120
rect 2497 4115 2563 4118
rect 11973 4115 12039 4118
rect 2037 4042 2103 4045
rect 6269 4042 6335 4045
rect 2037 4040 6335 4042
rect 2037 3984 2042 4040
rect 2098 3984 6274 4040
rect 6330 3984 6335 4040
rect 2037 3982 6335 3984
rect 2037 3979 2103 3982
rect 6269 3979 6335 3982
rect 13261 4042 13327 4045
rect 17953 4042 18019 4045
rect 13261 4040 18019 4042
rect 13261 3984 13266 4040
rect 13322 3984 17958 4040
rect 18014 3984 18019 4040
rect 13261 3982 18019 3984
rect 13261 3979 13327 3982
rect 17953 3979 18019 3982
rect 18229 4042 18295 4045
rect 20897 4042 20963 4045
rect 18229 4040 20963 4042
rect 18229 3984 18234 4040
rect 18290 3984 20902 4040
rect 20958 3984 20963 4040
rect 18229 3982 20963 3984
rect 18229 3979 18295 3982
rect 20897 3979 20963 3982
rect 21817 4042 21883 4045
rect 27521 4042 27587 4045
rect 21817 4040 27587 4042
rect 21817 3984 21822 4040
rect 21878 3984 27526 4040
rect 27582 3984 27587 4040
rect 21817 3982 27587 3984
rect 21817 3979 21883 3982
rect 27521 3979 27587 3982
rect 0 3906 480 3936
rect 1577 3906 1643 3909
rect 0 3904 1643 3906
rect 0 3848 1582 3904
rect 1638 3848 1643 3904
rect 0 3846 1643 3848
rect 0 3816 480 3846
rect 1577 3843 1643 3846
rect 4797 3906 4863 3909
rect 8201 3906 8267 3909
rect 4797 3904 8267 3906
rect 4797 3848 4802 3904
rect 4858 3848 8206 3904
rect 8262 3848 8267 3904
rect 4797 3846 8267 3848
rect 4797 3843 4863 3846
rect 8201 3843 8267 3846
rect 18413 3906 18479 3909
rect 20805 3906 20871 3909
rect 18413 3904 20871 3906
rect 18413 3848 18418 3904
rect 18474 3848 20810 3904
rect 20866 3848 20871 3904
rect 18413 3846 20871 3848
rect 18413 3843 18479 3846
rect 20805 3843 20871 3846
rect 26693 3906 26759 3909
rect 29520 3906 30000 3936
rect 26693 3904 30000 3906
rect 26693 3848 26698 3904
rect 26754 3848 30000 3904
rect 26693 3846 30000 3848
rect 26693 3843 26759 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 4889 3770 4955 3773
rect 10777 3770 10843 3773
rect 4889 3768 10843 3770
rect 4889 3712 4894 3768
rect 4950 3712 10782 3768
rect 10838 3712 10843 3768
rect 4889 3710 10843 3712
rect 4889 3707 4955 3710
rect 10777 3707 10843 3710
rect 26417 3770 26483 3773
rect 27613 3770 27679 3773
rect 26417 3768 27679 3770
rect 26417 3712 26422 3768
rect 26478 3712 27618 3768
rect 27674 3712 27679 3768
rect 26417 3710 27679 3712
rect 26417 3707 26483 3710
rect 27613 3707 27679 3710
rect 2681 3634 2747 3637
rect 4705 3634 4771 3637
rect 2681 3632 4771 3634
rect 2681 3576 2686 3632
rect 2742 3576 4710 3632
rect 4766 3576 4771 3632
rect 2681 3574 4771 3576
rect 2681 3571 2747 3574
rect 4705 3571 4771 3574
rect 7097 3634 7163 3637
rect 9857 3634 9923 3637
rect 7097 3632 9923 3634
rect 7097 3576 7102 3632
rect 7158 3576 9862 3632
rect 9918 3576 9923 3632
rect 7097 3574 9923 3576
rect 7097 3571 7163 3574
rect 9857 3571 9923 3574
rect 20437 3634 20503 3637
rect 26509 3634 26575 3637
rect 20437 3632 26575 3634
rect 20437 3576 20442 3632
rect 20498 3576 26514 3632
rect 26570 3576 26575 3632
rect 20437 3574 26575 3576
rect 20437 3571 20503 3574
rect 26509 3571 26575 3574
rect 4337 3498 4403 3501
rect 12249 3498 12315 3501
rect 4337 3496 12315 3498
rect 4337 3440 4342 3496
rect 4398 3440 12254 3496
rect 12310 3440 12315 3496
rect 4337 3438 12315 3440
rect 4337 3435 4403 3438
rect 12249 3435 12315 3438
rect 12709 3498 12775 3501
rect 27521 3498 27587 3501
rect 12709 3496 27587 3498
rect 12709 3440 12714 3496
rect 12770 3440 27526 3496
rect 27582 3440 27587 3496
rect 12709 3438 27587 3440
rect 12709 3435 12775 3438
rect 27521 3435 27587 3438
rect 0 3362 480 3392
rect 2681 3362 2747 3365
rect 0 3360 2747 3362
rect 0 3304 2686 3360
rect 2742 3304 2747 3360
rect 0 3302 2747 3304
rect 0 3272 480 3302
rect 2681 3299 2747 3302
rect 26601 3362 26667 3365
rect 29520 3362 30000 3392
rect 26601 3360 30000 3362
rect 26601 3304 26606 3360
rect 26662 3304 30000 3360
rect 26601 3302 30000 3304
rect 26601 3299 26667 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 657 3226 723 3229
rect 10133 3226 10199 3229
rect 12065 3226 12131 3229
rect 657 3224 5826 3226
rect 657 3168 662 3224
rect 718 3168 5826 3224
rect 657 3166 5826 3168
rect 657 3163 723 3166
rect 2037 3090 2103 3093
rect 5533 3090 5599 3093
rect 2037 3088 5599 3090
rect 2037 3032 2042 3088
rect 2098 3032 5538 3088
rect 5594 3032 5599 3088
rect 2037 3030 5599 3032
rect 5766 3090 5826 3166
rect 10133 3224 12131 3226
rect 10133 3168 10138 3224
rect 10194 3168 12070 3224
rect 12126 3168 12131 3224
rect 10133 3166 12131 3168
rect 10133 3163 10199 3166
rect 12065 3163 12131 3166
rect 23657 3090 23723 3093
rect 5766 3088 23723 3090
rect 5766 3032 23662 3088
rect 23718 3032 23723 3088
rect 5766 3030 23723 3032
rect 2037 3027 2103 3030
rect 5533 3027 5599 3030
rect 23657 3027 23723 3030
rect 10225 2954 10291 2957
rect 26325 2954 26391 2957
rect 10225 2952 26391 2954
rect 10225 2896 10230 2952
rect 10286 2896 26330 2952
rect 26386 2896 26391 2952
rect 10225 2894 26391 2896
rect 10225 2891 10291 2894
rect 26325 2891 26391 2894
rect 2957 2818 3023 2821
rect 6361 2818 6427 2821
rect 2957 2816 6427 2818
rect 2957 2760 2962 2816
rect 3018 2760 6366 2816
rect 6422 2760 6427 2816
rect 2957 2758 6427 2760
rect 2957 2755 3023 2758
rect 6361 2755 6427 2758
rect 15009 2818 15075 2821
rect 16297 2818 16363 2821
rect 15009 2816 16363 2818
rect 15009 2760 15014 2816
rect 15070 2760 16302 2816
rect 16358 2760 16363 2816
rect 15009 2758 16363 2760
rect 15009 2755 15075 2758
rect 16297 2755 16363 2758
rect 25589 2818 25655 2821
rect 29177 2818 29243 2821
rect 25589 2816 29243 2818
rect 25589 2760 25594 2816
rect 25650 2760 29182 2816
rect 29238 2760 29243 2816
rect 25589 2758 29243 2760
rect 25589 2755 25655 2758
rect 29177 2755 29243 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 27705 2682 27771 2685
rect 29520 2682 30000 2712
rect 27705 2680 30000 2682
rect 27705 2624 27710 2680
rect 27766 2624 30000 2680
rect 27705 2622 30000 2624
rect 27705 2619 27771 2622
rect 29520 2592 30000 2622
rect 5533 2546 5599 2549
rect 9949 2546 10015 2549
rect 5533 2544 10015 2546
rect 5533 2488 5538 2544
rect 5594 2488 9954 2544
rect 10010 2488 10015 2544
rect 5533 2486 10015 2488
rect 5533 2483 5599 2486
rect 9949 2483 10015 2486
rect 19977 2546 20043 2549
rect 26877 2546 26943 2549
rect 19977 2544 26943 2546
rect 19977 2488 19982 2544
rect 20038 2488 26882 2544
rect 26938 2488 26943 2544
rect 19977 2486 26943 2488
rect 19977 2483 20043 2486
rect 26877 2483 26943 2486
rect 5944 2208 6264 2209
rect 0 2138 480 2168
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 1393 2138 1459 2141
rect 0 2136 1459 2138
rect 0 2080 1398 2136
rect 1454 2080 1459 2136
rect 0 2078 1459 2080
rect 0 2048 480 2078
rect 1393 2075 1459 2078
rect 26693 2138 26759 2141
rect 29520 2138 30000 2168
rect 26693 2136 30000 2138
rect 26693 2080 26698 2136
rect 26754 2080 30000 2136
rect 26693 2078 30000 2080
rect 26693 2075 26759 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1577 1458 1643 1461
rect 0 1456 1643 1458
rect 0 1400 1582 1456
rect 1638 1400 1643 1456
rect 0 1398 1643 1400
rect 0 1368 480 1398
rect 1577 1395 1643 1398
rect 26601 1458 26667 1461
rect 29520 1458 30000 1488
rect 26601 1456 30000 1458
rect 26601 1400 26606 1456
rect 26662 1400 30000 1456
rect 26601 1398 30000 1400
rect 26601 1395 26667 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 480 854
rect 1669 851 1735 854
rect 27061 914 27127 917
rect 29520 914 30000 944
rect 27061 912 30000 914
rect 27061 856 27066 912
rect 27122 856 30000 912
rect 27061 854 30000 856
rect 27061 851 27127 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 2405 370 2471 373
rect 0 368 2471 370
rect 0 312 2410 368
rect 2466 312 2471 368
rect 0 310 2471 312
rect 0 280 480 310
rect 2405 307 2471 310
rect 26785 370 26851 373
rect 29520 370 30000 400
rect 26785 368 30000 370
rect 26785 312 26790 368
rect 26846 312 30000 368
rect 26785 310 30000 312
rect 26785 307 26851 310
rect 29520 280 30000 310
<< via3 >>
rect 25452 22340 25516 22404
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 24900 20028 24964 20092
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 25084 15812 25148 15876
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 25636 11868 25700 11932
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 24900 11324 24964 11388
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 25084 8060 25148 8124
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 17908 5612 17972 5676
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 17908 5340 17972 5404
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 25451 22404 25517 22405
rect 25451 22340 25452 22404
rect 25516 22340 25517 22404
rect 25451 22339 25517 22340
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 24899 20092 24965 20093
rect 24899 20028 24900 20092
rect 24964 20028 24965 20092
rect 24899 20027 24965 20028
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 24902 11389 24962 20027
rect 25454 19410 25514 22339
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25454 19350 25882 19410
rect 25083 15876 25149 15877
rect 25083 15812 25084 15876
rect 25148 15812 25149 15876
rect 25083 15811 25149 15812
rect 24899 11388 24965 11389
rect 24899 11324 24900 11388
rect 24964 11324 24965 11388
rect 24899 11323 24965 11324
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 25086 8125 25146 15811
rect 25635 11932 25701 11933
rect 25635 11868 25636 11932
rect 25700 11930 25701 11932
rect 25822 11930 25882 19350
rect 25700 11870 25882 11930
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25700 11868 25701 11870
rect 25635 11867 25701 11868
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25083 8124 25149 8125
rect 25083 8060 25084 8124
rect 25148 8060 25149 8124
rect 25083 8059 25149 8060
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 17907 5676 17973 5677
rect 17907 5612 17908 5676
rect 17972 5612 17973 5676
rect 17907 5611 17973 5612
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 17910 5405 17970 5611
rect 17907 5404 17973 5405
rect 17907 5340 17908 5404
rect 17972 5340 17973 5404
rect 17907 5339 17973 5340
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604681595
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _56_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604681595
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1604681595
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2116 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 1604681595
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604681595
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604681595
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1604681595
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1604681595
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604681595
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 2668 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1604681595
transform 1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604681595
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 3772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 3036 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1604681595
transform 1 0 3956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1604681595
transform 1 0 4784 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1604681595
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 4324 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604681595
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_48
timestamp 1604681595
transform 1 0 5520 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1604681595
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4968 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1604681595
transform 1 0 5152 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1604681595
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_52
timestamp 1604681595
transform 1 0 5888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1604681595
transform 1 0 6348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1604681595
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604681595
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604681595
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604681595
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 6900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6992 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1604681595
transform 1 0 6992 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1604681595
transform 1 0 7820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1604681595
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1604681595
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1604681595
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 8372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1604681595
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 8556 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_85
timestamp 1604681595
transform 1 0 8924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1604681595
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 1604681595
transform 1 0 9292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 9200 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604681595
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_104
timestamp 1604681595
transform 1 0 10672 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1604681595
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9752 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9384 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1604681595
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_109
timestamp 1604681595
transform 1 0 11132 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 11316 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 11224 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1604681595
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_117
timestamp 1604681595
transform 1 0 11868 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1604681595
transform 1 0 12144 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_116
timestamp 1604681595
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604681595
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604681595
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604681595
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 13800 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_137
timestamp 1604681595
transform 1 0 13708 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_144
timestamp 1604681595
transform 1 0 14352 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604681595
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_154
timestamp 1604681595
transform 1 0 15272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_147
timestamp 1604681595
transform 1 0 14628 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1604681595
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_148
timestamp 1604681595
transform 1 0 14720 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 14720 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_158
timestamp 1604681595
transform 1 0 15640 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_156
timestamp 1604681595
transform 1 0 15456 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 15456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604681595
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_164
timestamp 1604681595
transform 1 0 16192 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_164
timestamp 1604681595
transform 1 0 16192 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 16284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16376 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_171
timestamp 1604681595
transform 1 0 16836 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_167
timestamp 1604681595
transform 1 0 16468 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_176
timestamp 1604681595
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1604681595
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1604681595
transform 1 0 18032 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1604681595
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1604681595
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604681595
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604681595
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 18216 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 18308 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1604681595
transform 1 0 19504 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_206
timestamp 1604681595
transform 1 0 20056 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_192
timestamp 1604681595
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_196
timestamp 1604681595
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_213
timestamp 1604681595
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1604681595
transform 1 0 20332 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1604681595
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_214
timestamp 1604681595
transform 1 0 20792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_210
timestamp 1604681595
transform 1 0 20424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604681595
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_222
timestamp 1604681595
transform 1 0 21528 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21344 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 21804 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21068 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_1_236
timestamp 1604681595
transform 1 0 22816 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 1604681595
transform 1 0 22356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 22540 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_245
timestamp 1604681595
transform 1 0 23644 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_249
timestamp 1604681595
transform 1 0 24012 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_247
timestamp 1604681595
transform 1 0 23828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604681595
transform 1 0 23828 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604681595
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604681595
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24104 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 24012 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_235
timestamp 1604681595
transform 1 0 22724 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604681595
transform 1 0 25392 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604681595
transform 1 0 25944 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 24840 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_256
timestamp 1604681595
transform 1 0 24656 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_260
timestamp 1604681595
transform 1 0 25024 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1604681595
transform 1 0 25760 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_255
timestamp 1604681595
transform 1 0 24564 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_259
timestamp 1604681595
transform 1 0 24932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604681595
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_271
timestamp 1604681595
transform 1 0 26036 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_278
timestamp 1604681595
transform 1 0 26680 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_272
timestamp 1604681595
transform 1 0 26128 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604681595
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1604681595
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_283
timestamp 1604681595
transform 1 0 27140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_288
timestamp 1604681595
transform 1 0 27600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_284
timestamp 1604681595
transform 1 0 27232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1604681595
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1604681595
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1604681595
transform 1 0 27416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1604681595
transform 1 0 26864 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1604681595
transform 1 0 27508 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_291
timestamp 1604681595
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604681595
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604681595
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1604681595
transform 1 0 28060 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_296
timestamp 1604681595
transform 1 0 28336 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604681595
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604681595
transform 1 0 2484 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604681595
transform 1 0 1380 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604681595
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604681595
transform 1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_7
timestamp 1604681595
transform 1 0 1748 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_11
timestamp 1604681595
transform 1 0 2116 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1604681595
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 4416 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604681595
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 3036 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_23
timestamp 1604681595
transform 1 0 3220 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_32
timestamp 1604681595
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_55
timestamp 1604681595
transform 1 0 6164 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1604681595
transform 1 0 7360 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_63
timestamp 1604681595
transform 1 0 6900 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_66
timestamp 1604681595
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_77
timestamp 1604681595
transform 1 0 8188 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 9844 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604681595
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_89
timestamp 1604681595
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1604681595
transform 1 0 9660 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1604681595
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 11132 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_2_105
timestamp 1604681595
transform 1 0 10764 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_128
timestamp 1604681595
transform 1 0 12880 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_140
timestamp 1604681595
transform 1 0 13984 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 16284 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604681595
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1604681595
transform 1 0 15088 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_154
timestamp 1604681595
transform 1 0 15272 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp 1604681595
transform 1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_184
timestamp 1604681595
transform 1 0 18032 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 19504 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_196
timestamp 1604681595
transform 1 0 19136 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_199
timestamp 1604681595
transform 1 0 19412 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1604681595
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 20884 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604681595
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21620 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1604681595
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1604681595
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_225
timestamp 1604681595
transform 1 0 21804 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604681595
transform 1 0 23460 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_237
timestamp 1604681595
transform 1 0 22908 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_247
timestamp 1604681595
transform 1 0 23828 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_259
timestamp 1604681595
transform 1 0 24932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1604681595
transform 1 0 26496 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604681595
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_271
timestamp 1604681595
transform 1 0 26036 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_280
timestamp 1604681595
transform 1 0 26864 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604681595
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_292
timestamp 1604681595
transform 1 0 27968 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_298
timestamp 1604681595
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604681595
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604681595
transform 1 0 2484 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604681595
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604681595
transform 1 0 2300 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604681595
transform 1 0 1932 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1604681595
transform 1 0 1748 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp 1604681595
transform 1 0 2116 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_19
timestamp 1604681595
transform 1 0 2852 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604681595
transform 1 0 3036 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4048 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 4784 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_23
timestamp 1604681595
transform 1 0 3220 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_31
timestamp 1604681595
transform 1 0 3956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1604681595
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_38
timestamp 1604681595
transform 1 0 4600 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 6808 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604681595
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_42
timestamp 1604681595
transform 1 0 4968 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_54
timestamp 1604681595
transform 1 0 6072 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_58
timestamp 1604681595
transform 1 0 6440 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 8648 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 7912 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1604681595
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1604681595
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_76
timestamp 1604681595
transform 1 0 8096 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 9384 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_88
timestamp 1604681595
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_92
timestamp 1604681595
transform 1 0 9568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_104
timestamp 1604681595
transform 1 0 10672 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604681595
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 12052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_110
timestamp 1604681595
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1604681595
transform 1 0 11500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1604681595
transform 1 0 11868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1604681595
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1604681595
transform 1 0 12420 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 12880 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1604681595
transform 1 0 12788 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1604681595
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_134
timestamp 1604681595
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_138
timestamp 1604681595
transform 1 0 13800 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1604681595
transform 1 0 16376 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15824 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_150
timestamp 1604681595
transform 1 0 14904 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1604681595
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1604681595
transform 1 0 16008 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604681595
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_175
timestamp 1604681595
transform 1 0 17204 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_184
timestamp 1604681595
transform 1 0 18032 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 18952 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1604681595
transform 1 0 18768 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1604681595
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_200
timestamp 1604681595
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1604681595
transform 1 0 21436 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 21252 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_213
timestamp 1604681595
transform 1 0 20700 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_217
timestamp 1604681595
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604681595
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 23828 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_230
timestamp 1604681595
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_234
timestamp 1604681595
transform 1 0 22632 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_242
timestamp 1604681595
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_245
timestamp 1604681595
transform 1 0 23644 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_249
timestamp 1604681595
transform 1 0 24012 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 24196 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_253
timestamp 1604681595
transform 1 0 24380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_265
timestamp 1604681595
transform 1 0 25484 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604681595
transform 1 0 27508 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604681595
transform 1 0 26404 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1604681595
transform 1 0 26956 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604681595
transform 1 0 26220 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_279
timestamp 1604681595
transform 1 0 26772 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_283
timestamp 1604681595
transform 1 0 27140 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_291
timestamp 1604681595
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604681595
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604681595
transform 1 0 28060 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_295
timestamp 1604681595
transform 1 0 28244 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604681595
transform 1 0 1380 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604681595
transform 1 0 2484 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604681595
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_7
timestamp 1604681595
transform 1 0 1748 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_19
timestamp 1604681595
transform 1 0 2852 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604681595
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3036 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_23
timestamp 1604681595
transform 1 0 3220 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1604681595
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 6808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_45
timestamp 1604681595
transform 1 0 5244 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1604681595
transform 1 0 6348 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_61
timestamp 1604681595
transform 1 0 6716 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7360 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 8372 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1604681595
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 1604681595
transform 1 0 8188 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1604681595
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604681595
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1604681595
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604681595
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1604681595
transform 1 0 11316 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 10764 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 11132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_107
timestamp 1604681595
transform 1 0 10948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1604681595
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_124
timestamp 1604681595
transform 1 0 12512 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1604681595
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_137
timestamp 1604681595
transform 1 0 13708 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604681595
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 15456 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1604681595
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1604681595
transform 1 0 15272 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_158
timestamp 1604681595
transform 1 0 15640 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_166
timestamp 1604681595
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_170
timestamp 1604681595
transform 1 0 16744 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1604681595
transform 1 0 17848 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1604681595
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_4_194
timestamp 1604681595
transform 1 0 18952 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_206
timestamp 1604681595
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604681595
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 21896 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_210
timestamp 1604681595
transform 1 0 20424 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_213
timestamp 1604681595
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_224
timestamp 1604681595
transform 1 0 21712 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_228
timestamp 1604681595
transform 1 0 22080 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 23460 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_4_240
timestamp 1604681595
transform 1 0 23184 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25392 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_262
timestamp 1604681595
transform 1 0 25208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_266
timestamp 1604681595
transform 1 0 25576 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1604681595
transform 1 0 26496 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604681595
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_274
timestamp 1604681595
transform 1 0 26312 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_280
timestamp 1604681595
transform 1 0 26864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604681595
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_292
timestamp 1604681595
transform 1 0 27968 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_298
timestamp 1604681595
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604681595
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604681595
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604681595
transform 1 0 1932 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604681595
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2852 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_7
timestamp 1604681595
transform 1 0 1748 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604681595
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1604681595
transform 1 0 2484 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 3036 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1604681595
transform 1 0 4784 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604681595
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 4968 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 5336 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1604681595
transform 1 0 5152 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_48
timestamp 1604681595
transform 1 0 5520 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_60
timestamp 1604681595
transform 1 0 6624 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1604681595
transform 1 0 6808 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 7176 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 6992 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 9660 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 9108 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_85
timestamp 1604681595
transform 1 0 8924 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp 1604681595
transform 1 0 9292 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_96
timestamp 1604681595
transform 1 0 9936 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604681595
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604681595
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 12604 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604681595
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604681595
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1604681595
transform 1 0 12420 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 13064 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_5_127
timestamp 1604681595
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1604681595
transform 1 0 16192 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1604681595
transform 1 0 14812 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1604681595
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1604681595
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1604681595
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604681595
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18216 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_173
timestamp 1604681595
transform 1 0 17020 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_184
timestamp 1604681595
transform 1 0 18032 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 19964 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1604681595
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_192
timestamp 1604681595
transform 1 0 18768 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1604681595
transform 1 0 19872 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1604681595
transform 1 0 20148 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20516 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21528 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21896 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1604681595
transform 1 0 21344 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_224
timestamp 1604681595
transform 1 0 21712 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_228
timestamp 1604681595
transform 1 0 22080 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604681595
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 22816 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_234
timestamp 1604681595
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_5_238
timestamp 1604681595
transform 1 0 23000 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1604681595
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25208 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604681595
transform 1 0 25024 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 24656 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_253
timestamp 1604681595
transform 1 0 24380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_258
timestamp 1604681595
transform 1 0 24840 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604681595
transform 1 0 27140 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1604681595
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_285
timestamp 1604681595
transform 1 0 27324 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604681595
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_297
timestamp 1604681595
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1604681595
transform 1 0 1380 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_7
timestamp 1604681595
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 1932 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604681595
transform 1 0 1564 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604681595
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604681595
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604681595
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_15
timestamp 1604681595
transform 1 0 2484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1604681595
transform 1 0 2116 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 1748 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1604681595
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_26
timestamp 1604681595
transform 1 0 3496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604681595
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604681595
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_36
timestamp 1604681595
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604681595
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604681595
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4600 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1604681595
transform 1 0 4232 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_7_47
timestamp 1604681595
transform 1 0 5428 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1604681595
transform 1 0 5060 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 5244 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604681595
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_57
timestamp 1604681595
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_53
timestamp 1604681595
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_59
timestamp 1604681595
transform 1 0 6532 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604681595
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_47
timestamp 1604681595
transform 1 0 5428 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_66
timestamp 1604681595
transform 1 0 7176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_68
timestamp 1604681595
transform 1 0 7360 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_65
timestamp 1604681595
transform 1 0 7084 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7544 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7544 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_7_79
timestamp 1604681595
transform 1 0 8372 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_79
timestamp 1604681595
transform 1 0 8372 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604681595
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604681595
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp 1604681595
transform 1 0 9660 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_87
timestamp 1604681595
transform 1 0 9108 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604681595
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_95
timestamp 1604681595
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_99
timestamp 1604681595
transform 1 0 10212 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10028 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_7_110
timestamp 1604681595
transform 1 0 11224 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_106
timestamp 1604681595
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_114
timestamp 1604681595
transform 1 0 11592 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 11040 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1604681595
transform 1 0 10764 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604681595
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1604681595
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_115
timestamp 1604681595
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604681595
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1604681595
transform 1 0 12328 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_133
timestamp 1604681595
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_127
timestamp 1604681595
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_135
timestamp 1604681595
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1604681595
transform 1 0 13156 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_140
timestamp 1604681595
transform 1 0 13984 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_136
timestamp 1604681595
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 13708 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13800 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_144
timestamp 1604681595
transform 1 0 14352 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1604681595
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 15272 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1604681595
transform 1 0 16376 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604681595
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 16192 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1604681595
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_156
timestamp 1604681595
transform 1 0 15456 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1604681595
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_175
timestamp 1604681595
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_173
timestamp 1604681595
transform 1 0 17020 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_179
timestamp 1604681595
transform 1 0 17572 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_180
timestamp 1604681595
transform 1 0 17664 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_177
timestamp 1604681595
transform 1 0 17388 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 17480 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604681595
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1604681595
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1604681595
transform 1 0 17756 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1604681595
transform 1 0 19228 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1604681595
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_194
timestamp 1604681595
transform 1 0 18952 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1604681595
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 19044 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1604681595
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_206
timestamp 1604681595
transform 1 0 20056 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_202
timestamp 1604681595
transform 1 0 19688 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1604681595
transform 1 0 19964 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604681595
transform 1 0 19780 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604681595
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_210
timestamp 1604681595
transform 1 0 20424 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1604681595
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_224
timestamp 1604681595
transform 1 0 21712 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_214
timestamp 1604681595
transform 1 0 20792 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_226
timestamp 1604681595
transform 1 0 21896 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 22448 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604681595
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 22632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23000 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_236
timestamp 1604681595
transform 1 0 22816 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_240
timestamp 1604681595
transform 1 0 23184 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604681595
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_260
timestamp 1604681595
transform 1 0 25024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_257
timestamp 1604681595
transform 1 0 24748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_268
timestamp 1604681595
transform 1 0 25760 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_264
timestamp 1604681595
transform 1 0 25392 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_267
timestamp 1604681595
transform 1 0 25668 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 25576 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 25208 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604681595
transform 1 0 25300 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604681595
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604681595
transform 1 0 26404 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604681595
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604681595
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604681595
transform 1 0 26956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604681595
transform 1 0 26220 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_280
timestamp 1604681595
transform 1 0 26864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_272
timestamp 1604681595
transform 1 0 26128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_279
timestamp 1604681595
transform 1 0 26772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_283
timestamp 1604681595
transform 1 0 27140 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604681595
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604681595
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_292
timestamp 1604681595
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_298
timestamp 1604681595
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_295
timestamp 1604681595
transform 1 0 28244 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604681595
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604681595
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604681595
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604681595
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604681595
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1604681595
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604681595
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1604681595
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_32
timestamp 1604681595
transform 1 0 4048 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5796 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_43
timestamp 1604681595
transform 1 0 5060 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_8_60
timestamp 1604681595
transform 1 0 6624 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 8280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_68
timestamp 1604681595
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_72
timestamp 1604681595
transform 1 0 7728 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604681595
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604681595
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_102
timestamp 1604681595
transform 1 0 10488 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1604681595
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_114
timestamp 1604681595
transform 1 0 11592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13432 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1604681595
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_130
timestamp 1604681595
transform 1 0 13064 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_143
timestamp 1604681595
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604681595
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 15640 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 16376 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16008 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1604681595
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_154
timestamp 1604681595
transform 1 0 15272 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_160
timestamp 1604681595
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_164
timestamp 1604681595
transform 1 0 16192 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1604681595
transform 1 0 17480 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_168
timestamp 1604681595
transform 1 0 16560 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_176
timestamp 1604681595
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_187
timestamp 1604681595
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 18492 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_191
timestamp 1604681595
transform 1 0 18676 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_199
timestamp 1604681595
transform 1 0 19412 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_202
timestamp 1604681595
transform 1 0 19688 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1604681595
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604681595
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21988 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604681595
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1604681595
transform 1 0 20884 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_219
timestamp 1604681595
transform 1 0 21252 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 1604681595
transform 1 0 22172 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1604681595
transform 1 0 22632 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_233
timestamp 1604681595
transform 1 0 22540 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_243
timestamp 1604681595
transform 1 0 23460 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24840 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 24564 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_257
timestamp 1604681595
transform 1 0 24748 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_267
timestamp 1604681595
transform 1 0 25668 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604681595
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604681595
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_271
timestamp 1604681595
transform 1 0 26036 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_274
timestamp 1604681595
transform 1 0 26312 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604681595
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604681595
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604681595
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604681595
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1564 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604681595
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604681595
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_24
timestamp 1604681595
transform 1 0 3312 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp 1604681595
transform 1 0 3680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604681595
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1604681595
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604681595
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1604681595
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604681595
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_53
timestamp 1604681595
transform 1 0 5980 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1604681595
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 8280 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 8096 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1604681595
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1604681595
transform 1 0 10028 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604681595
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 11776 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 11408 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1604681595
transform 1 0 11132 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_114
timestamp 1604681595
transform 1 0 11592 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1604681595
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1604681595
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604681595
transform 1 0 14168 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_134
timestamp 1604681595
transform 1 0 13432 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_145
timestamp 1604681595
transform 1 0 14444 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_151
timestamp 1604681595
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_154
timestamp 1604681595
transform 1 0 15272 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604681595
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604681595
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16652 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_167
timestamp 1604681595
transform 1 0 16468 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1604681595
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_187
timestamp 1604681595
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19504 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_prog_clk_A
timestamp 1604681595
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_191
timestamp 1604681595
transform 1 0 18676 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_197
timestamp 1604681595
transform 1 0 19228 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1604681595
transform 1 0 21988 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 21804 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_219
timestamp 1604681595
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_223
timestamp 1604681595
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604681595
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 24012 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_236
timestamp 1604681595
transform 1 0 22816 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_245
timestamp 1604681595
transform 1 0 23644 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24564 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604681595
transform 1 0 25944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_251
timestamp 1604681595
transform 1 0 24196 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_264
timestamp 1604681595
transform 1 0 25392 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_268
timestamp 1604681595
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26128 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_291
timestamp 1604681595
transform 1 0 27876 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604681595
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604681595
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604681595
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1604681595
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_11
timestamp 1604681595
transform 1 0 2116 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1604681595
transform 1 0 4140 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604681595
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_23
timestamp 1604681595
transform 1 0 3220 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 1604681595
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604681595
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_42
timestamp 1604681595
transform 1 0 4968 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_46
timestamp 1604681595
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_50
timestamp 1604681595
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_54
timestamp 1604681595
transform 1 0 6072 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_66
timestamp 1604681595
transform 1 0 7176 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_78
timestamp 1604681595
transform 1 0 8280 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604681595
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 9844 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10212 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_86
timestamp 1604681595
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604681595
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1604681595
transform 1 0 9660 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 1604681595
transform 1 0 10028 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_101
timestamp 1604681595
transform 1 0 10396 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 11684 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_10_113
timestamp 1604681595
transform 1 0 11500 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_134
timestamp 1604681595
transform 1 0 13432 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16008 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604681595
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_146
timestamp 1604681595
transform 1 0 14536 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1604681595
transform 1 0 15088 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_154
timestamp 1604681595
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_160
timestamp 1604681595
transform 1 0 15824 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_181
timestamp 1604681595
transform 1 0 17756 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 18492 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_192
timestamp 1604681595
transform 1 0 18768 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1604681595
transform 1 0 19872 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20976 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604681595
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_212
timestamp 1604681595
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_215
timestamp 1604681595
transform 1 0 20884 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 24012 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_235
timestamp 1604681595
transform 1 0 22724 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_247
timestamp 1604681595
transform 1 0 23828 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24288 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 25300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1604681595
transform 1 0 24196 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_261
timestamp 1604681595
transform 1 0 25116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_265
timestamp 1604681595
transform 1 0 25484 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604681595
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604681595
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_271
timestamp 1604681595
transform 1 0 26036 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_274
timestamp 1604681595
transform 1 0 26312 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604681595
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604681595
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604681595
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604681595
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604681595
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604681595
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604681595
transform 1 0 1932 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604681595
transform 1 0 2300 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1604681595
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1604681595
transform 1 0 2116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1604681595
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1604681595
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_27
timestamp 1604681595
transform 1 0 3588 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1604681595
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604681595
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 5704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1604681595
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_52
timestamp 1604681595
transform 1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_56
timestamp 1604681595
transform 1 0 6256 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1604681595
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1604681595
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 8188 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_74
timestamp 1604681595
transform 1 0 7912 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1604681595
transform 1 0 8372 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_83
timestamp 1604681595
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 9108 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604681595
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_106
timestamp 1604681595
transform 1 0 10856 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_118
timestamp 1604681595
transform 1 0 11960 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604681595
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_135
timestamp 1604681595
transform 1 0 13524 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_143
timestamp 1604681595
transform 1 0 14260 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_146
timestamp 1604681595
transform 1 0 14536 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1604681595
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_154
timestamp 1604681595
transform 1 0 15272 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604681595
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_167
timestamp 1604681595
transform 1 0 16468 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1604681595
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1604681595
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 18584 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18952 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 19320 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1604681595
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1604681595
transform 1 0 19136 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_200
timestamp 1604681595
transform 1 0 19504 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1604681595
transform 1 0 20884 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_prog_clk_A
timestamp 1604681595
transform 1 0 21344 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_212
timestamp 1604681595
transform 1 0 20608 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_218
timestamp 1604681595
transform 1 0 21160 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_222
timestamp 1604681595
transform 1 0 21528 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1604681595
transform 1 0 24012 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604681595
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23828 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23000 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_234
timestamp 1604681595
transform 1 0 22632 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_240
timestamp 1604681595
transform 1 0 23184 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_245
timestamp 1604681595
transform 1 0 23644 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_258
timestamp 1604681595
transform 1 0 24840 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_262
timestamp 1604681595
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_266
timestamp 1604681595
transform 1 0 25576 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604681595
transform 1 0 26496 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_274
timestamp 1604681595
transform 1 0 26312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_278
timestamp 1604681595
transform 1 0 26680 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_290
timestamp 1604681595
transform 1 0 27784 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604681595
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_298
timestamp 1604681595
transform 1 0 28520 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604681595
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604681595
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_7
timestamp 1604681595
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_19
timestamp 1604681595
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604681595
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_32
timestamp 1604681595
transform 1 0 4048 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_38
timestamp 1604681595
transform 1 0 4600 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_41
timestamp 1604681595
transform 1 0 4876 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 5428 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 7544 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_66
timestamp 1604681595
transform 1 0 7176 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_72
timestamp 1604681595
transform 1 0 7728 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_77
timestamp 1604681595
transform 1 0 8188 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604681595
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1604681595
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 8924 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_87
timestamp 1604681595
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_102
timestamp 1604681595
transform 1 0 10488 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1604681595
transform 1 0 11592 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_126
timestamp 1604681595
transform 1 0 12696 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_12_134
timestamp 1604681595
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604681595
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1604681595
transform 1 0 14536 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1604681595
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 18308 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_173
timestamp 1604681595
transform 1 0 17020 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_185
timestamp 1604681595
transform 1 0 18124 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1604681595
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_199
timestamp 1604681595
transform 1 0 19412 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604681595
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 21988 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21068 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1604681595
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_215
timestamp 1604681595
transform 1 0 20884 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_219
timestamp 1604681595
transform 1 0 21252 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_229
timestamp 1604681595
transform 1 0 22172 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23460 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_241
timestamp 1604681595
transform 1 0 23276 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 24656 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_252
timestamp 1604681595
transform 1 0 24288 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_258
timestamp 1604681595
transform 1 0 24840 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_270
timestamp 1604681595
transform 1 0 25944 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604681595
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604681595
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_274
timestamp 1604681595
transform 1 0 26312 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604681595
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604681595
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604681595
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604681595
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_7
timestamp 1604681595
transform 1 0 1748 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604681595
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604681595
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604681595
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604681595
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604681595
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_17
timestamp 1604681595
transform 1 0 2668 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_12
timestamp 1604681595
transform 1 0 2208 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 1604681595
transform 1 0 2484 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604681595
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 2024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604681595
transform 1 0 2484 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604681595
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604681595
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1604681595
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_21
timestamp 1604681595
transform 1 0 3036 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1604681595
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_23
timestamp 1604681595
transform 1 0 3220 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 3496 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604681595
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_40
timestamp 1604681595
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_36
timestamp 1604681595
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1604681595
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4048 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604681595
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1604681595
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1604681595
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1604681595
transform 1 0 6808 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1604681595
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1604681595
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1604681595
transform 1 0 7636 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_68
timestamp 1604681595
transform 1 0 7360 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_prog_clk_A
timestamp 1604681595
transform 1 0 7452 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1604681595
transform 1 0 7544 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1604681595
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1604681595
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp 1604681595
transform 1 0 7820 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 7820 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8004 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1604681595
transform 1 0 8924 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604681595
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1604681595
transform 1 0 9752 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1604681595
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_93
timestamp 1604681595
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_97
timestamp 1604681595
transform 1 0 10028 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 11040 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604681595
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 11040 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11408 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1604681595
transform 1 0 10856 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1604681595
transform 1 0 11224 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604681595
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_13_123
timestamp 1604681595
transform 1 0 12420 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_105
timestamp 1604681595
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13248 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_129
timestamp 1604681595
transform 1 0 12972 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_127
timestamp 1604681595
transform 1 0 12788 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_139
timestamp 1604681595
transform 1 0 13892 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604681595
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_147
timestamp 1604681595
transform 1 0 14628 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_156
timestamp 1604681595
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_151
timestamp 1604681595
transform 1 0 14996 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604681595
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1604681595
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_163
timestamp 1604681595
transform 1 0 16100 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_164
timestamp 1604681595
transform 1 0 16192 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_175
timestamp 1604681595
transform 1 0 17204 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_176
timestamp 1604681595
transform 1 0 17296 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_183
timestamp 1604681595
transform 1 0 17940 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1604681595
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604681595
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 18124 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604681595
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1604681595
transform 1 0 18308 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_196
timestamp 1604681595
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1604681595
transform 1 0 18584 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1604681595
transform 1 0 19780 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1604681595
transform 1 0 19412 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 19964 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 19320 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 19596 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1604681595
transform 1 0 20148 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_200
timestamp 1604681595
transform 1 0 19504 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1604681595
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_217
timestamp 1604681595
transform 1 0 21068 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_214
timestamp 1604681595
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_210
timestamp 1604681595
transform 1 0 20424 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604681595
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_223
timestamp 1604681595
transform 1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21804 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1604681595
transform 1 0 21988 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 20884 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1604681595
transform 1 0 23736 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604681595
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 23828 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_236
timestamp 1604681595
transform 1 0 22816 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_245
timestamp 1604681595
transform 1 0 23644 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_249
timestamp 1604681595
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_234
timestamp 1604681595
transform 1 0 22632 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604681595
transform 1 0 25300 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 24656 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 24196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_253
timestamp 1604681595
transform 1 0 24380 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_255
timestamp 1604681595
transform 1 0 24564 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_259
timestamp 1604681595
transform 1 0 24932 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_266
timestamp 1604681595
transform 1 0 25576 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604681595
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_279
timestamp 1604681595
transform 1 0 26772 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_275
timestamp 1604681595
transform 1 0 26404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604681595
transform 1 0 26588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604681595
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604681595
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_291
timestamp 1604681595
transform 1 0 27876 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_287
timestamp 1604681595
transform 1 0 27508 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604681595
transform 1 0 27692 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604681595
transform 1 0 27140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1604681595
transform 1 0 26864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604681595
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604681595
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_292
timestamp 1604681595
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_298
timestamp 1604681595
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 2024 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604681595
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604681595
transform 1 0 1564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1604681595
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_7
timestamp 1604681595
transform 1 0 1748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4508 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1604681595
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1604681595
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604681595
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1604681595
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_50
timestamp 1604681595
transform 1 0 5704 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604681595
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604681595
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1604681595
transform 1 0 6808 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8188 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1604681595
transform 1 0 7912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 6992 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1604681595
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1604681595
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9752 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_86
timestamp 1604681595
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 1604681595
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_103
timestamp 1604681595
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604681595
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 10764 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1604681595
transform 1 0 10948 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_111
timestamp 1604681595
transform 1 0 11316 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1604681595
transform 1 0 12052 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1604681595
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12880 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 14352 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 13984 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_127
timestamp 1604681595
transform 1 0 12788 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_130
timestamp 1604681595
transform 1 0 13064 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_134
timestamp 1604681595
transform 1 0 13432 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1604681595
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1604681595
transform 1 0 14904 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 14720 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_146
timestamp 1604681595
transform 1 0 14536 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1604681595
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1604681595
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604681595
transform 1 0 16468 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604681595
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_170
timestamp 1604681595
transform 1 0 16744 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_176
timestamp 1604681595
transform 1 0 17296 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 1604681595
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_184
timestamp 1604681595
transform 1 0 18032 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 19688 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1604681595
transform 1 0 19136 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1604681595
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_204
timestamp 1604681595
transform 1 0 19872 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604681595
transform 1 0 21712 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 22172 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 20976 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1604681595
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1604681595
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_227
timestamp 1604681595
transform 1 0 21988 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1604681595
transform 1 0 23828 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604681595
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 23000 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_231
timestamp 1604681595
transform 1 0 22356 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_237
timestamp 1604681595
transform 1 0 22908 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_240
timestamp 1604681595
transform 1 0 23184 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_245
timestamp 1604681595
transform 1 0 23644 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_256
timestamp 1604681595
transform 1 0 24656 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_268
timestamp 1604681595
transform 1 0 25760 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604681595
transform 1 0 26404 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604681595
transform 1 0 27508 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604681595
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604681595
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_274
timestamp 1604681595
transform 1 0 26312 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_279
timestamp 1604681595
transform 1 0 26772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_283
timestamp 1604681595
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_291
timestamp 1604681595
transform 1 0 27876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604681595
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604681595
transform 1 0 28060 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_295
timestamp 1604681595
transform 1 0 28244 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604681595
transform 1 0 2484 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604681595
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604681595
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 1932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 2300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1604681595
transform 1 0 1748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_11
timestamp 1604681595
transform 1 0 2116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_19
timestamp 1604681595
transform 1 0 2852 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604681595
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3036 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604681595
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604681595
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 5796 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 5244 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1604681595
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_47
timestamp 1604681595
transform 1 0 5428 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_60
timestamp 1604681595
transform 1 0 6624 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7820 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 7636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_68
timestamp 1604681595
transform 1 0 7360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1604681595
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1604681595
transform 1 0 10580 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604681595
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 9844 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1604681595
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_93
timestamp 1604681595
transform 1 0 9660 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_97
timestamp 1604681595
transform 1 0 10028 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_112
timestamp 1604681595
transform 1 0 11408 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_124
timestamp 1604681595
transform 1 0 12512 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 12880 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1604681595
transform 1 0 15548 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604681595
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_147
timestamp 1604681595
transform 1 0 14628 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1604681595
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1604681595
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18124 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16560 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 17940 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_170
timestamp 1604681595
transform 1 0 16744 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1604681595
transform 1 0 17848 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 19872 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 20240 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1604681595
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_198
timestamp 1604681595
transform 1 0 19320 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 1604681595
transform 1 0 20056 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1604681595
transform 1 0 21344 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604681595
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1604681595
transform 1 0 20424 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1604681595
transform 1 0 20884 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1604681595
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_229
timestamp 1604681595
transform 1 0 22172 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 23828 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 22724 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23092 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_237
timestamp 1604681595
transform 1 0 22908 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_241
timestamp 1604681595
transform 1 0 23276 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_249
timestamp 1604681595
transform 1 0 24012 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 24472 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 24840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 25208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_253
timestamp 1604681595
transform 1 0 24380 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_256
timestamp 1604681595
transform 1 0 24656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_260
timestamp 1604681595
transform 1 0 25024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_264
timestamp 1604681595
transform 1 0 25392 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604681595
transform 1 0 26496 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604681595
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604681595
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_280
timestamp 1604681595
transform 1 0 26864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604681595
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_292
timestamp 1604681595
transform 1 0 27968 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_298
timestamp 1604681595
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1656 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604681595
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1604681595
transform 1 0 1380 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4784 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 3588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1604681595
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1604681595
transform 1 0 3772 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_33
timestamp 1604681595
transform 1 0 4140 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604681595
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604681595
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 6256 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5888 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_49
timestamp 1604681595
transform 1 0 5612 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1604681595
transform 1 0 6072 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1604681595
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1604681595
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1604681595
transform 1 0 7820 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 7636 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 7268 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_66
timestamp 1604681595
transform 1 0 7176 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1604681595
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_82
timestamp 1604681595
transform 1 0 8648 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1604681595
transform 1 0 9660 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 1604681595
transform 1 0 9016 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_89
timestamp 1604681595
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1604681595
transform 1 0 10488 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1604681595
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604681595
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604681595
transform 1 0 11224 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1604681595
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_117
timestamp 1604681595
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 12052 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604681595
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604681595
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604681595
transform 1 0 13892 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1604681595
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1604681595
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1604681595
transform 1 0 15732 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_176
timestamp 1604681595
transform 1 0 17296 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_172
timestamp 1604681595
transform 1 0 16928 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_168
timestamp 1604681595
transform 1 0 16560 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_184
timestamp 1604681595
transform 1 0 18032 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604681595
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604681595
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18308 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1604681595
transform 1 0 19872 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 19688 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1604681595
transform 1 0 19136 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1604681595
transform 1 0 19504 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1604681595
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604681595
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604681595
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_234
timestamp 1604681595
transform 1 0 22632 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_230
timestamp 1604681595
transform 1 0 22264 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_237
timestamp 1604681595
transform 1 0 22908 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_241
timestamp 1604681595
transform 1 0 23276 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_245
timestamp 1604681595
transform 1 0 23644 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 23920 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604681595
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_250
timestamp 1604681595
transform 1 0 24104 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1604681595
transform 1 0 24472 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 24288 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25944 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 25576 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_263
timestamp 1604681595
transform 1 0 25300 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_268
timestamp 1604681595
transform 1 0 25760 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26128 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 27140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 27508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1604681595
transform 1 0 26956 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_285
timestamp 1604681595
transform 1 0 27324 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_289
timestamp 1604681595
transform 1 0 27692 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604681595
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_297
timestamp 1604681595
transform 1 0 28428 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1656 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604681595
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1604681595
transform 1 0 1380 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_15
timestamp 1604681595
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_19
timestamp 1604681595
transform 1 0 2852 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_23
timestamp 1604681595
transform 1 0 3220 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 3036 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1604681595
transform 1 0 3864 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1604681595
transform 1 0 3588 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 3680 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_32
timestamp 1604681595
transform 1 0 4048 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 4232 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604681595
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_36
timestamp 1604681595
transform 1 0 4416 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 4784 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604681595
transform 1 0 4968 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 6256 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_18_45
timestamp 1604681595
transform 1 0 5244 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_53
timestamp 1604681595
transform 1 0 5980 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 8188 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_75
timestamp 1604681595
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1604681595
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1604681595
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604681595
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604681595
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1604681595
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1604681595
transform 1 0 10856 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_18_105
timestamp 1604681595
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_115
timestamp 1604681595
transform 1 0 11684 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_127
timestamp 1604681595
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_139
timestamp 1604681595
transform 1 0 13892 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604681595
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16284 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_149
timestamp 1604681595
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1604681595
transform 1 0 16100 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18308 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 18124 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 16652 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 1604681595
transform 1 0 16468 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_171
timestamp 1604681595
transform 1 0 16836 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1604681595
transform 1 0 17940 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_206
timestamp 1604681595
transform 1 0 20056 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604681595
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 21896 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_224
timestamp 1604681595
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_228
timestamp 1604681595
transform 1 0 22080 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1604681595
transform 1 0 22724 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 24104 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_234
timestamp 1604681595
transform 1 0 22632 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_244
timestamp 1604681595
transform 1 0 23552 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1604681595
transform 1 0 24288 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 25668 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_261
timestamp 1604681595
transform 1 0 25116 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_269
timestamp 1604681595
transform 1 0 25852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1604681595
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604681595
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604681595
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_285
timestamp 1604681595
transform 1 0 27324 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604681595
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1604681595
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1604681595
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604681595
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 1656 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1656 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604681595
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604681595
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 1840 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_17
timestamp 1604681595
transform 1 0 2668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1604681595
transform 1 0 2668 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 2852 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604681595
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1604681595
transform 1 0 3588 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 1604681595
transform 1 0 3036 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_25
timestamp 1604681595
transform 1 0 3404 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_21
timestamp 1604681595
transform 1 0 3036 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 3680 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 3220 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 3680 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_32
timestamp 1604681595
transform 1 0 4048 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_37
timestamp 1604681595
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604681595
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 4232 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_41
timestamp 1604681595
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604681595
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 5060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1604681595
transform 1 0 5244 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_49
timestamp 1604681595
transform 1 0 5612 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_62
timestamp 1604681595
transform 1 0 6808 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_43
timestamp 1604681595
transform 1 0 5060 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_55
timestamp 1604681595
transform 1 0 6164 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1604681595
transform 1 0 7268 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604681595
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_67
timestamp 1604681595
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1604681595
transform 1 0 7452 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1604681595
transform 1 0 8004 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_78
timestamp 1604681595
transform 1 0 8280 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8556 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604681595
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_100
timestamp 1604681595
transform 1 0 10304 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1604681595
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1604681595
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_107
timestamp 1604681595
transform 1 0 10948 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604681595
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_108
timestamp 1604681595
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 10764 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1604681595
transform 1 0 11224 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604681595
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_119
timestamp 1604681595
transform 1 0 12052 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1604681595
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1604681595
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604681595
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1604681595
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604681595
transform 1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 13248 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_135
timestamp 1604681595
transform 1 0 13524 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_145
timestamp 1604681595
transform 1 0 14444 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1604681595
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_134
timestamp 1604681595
transform 1 0 13432 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_150
timestamp 1604681595
transform 1 0 14904 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1604681595
transform 1 0 14536 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_149
timestamp 1604681595
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14628 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604681595
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15180 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1604681595
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604681595
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 16284 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_166
timestamp 1604681595
transform 1 0 16376 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_167
timestamp 1604681595
transform 1 0 16468 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_177
timestamp 1604681595
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1604681595
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_170
timestamp 1604681595
transform 1 0 16744 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1604681595
transform 1 0 16836 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_184
timestamp 1604681595
transform 1 0 18032 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1604681595
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604681595
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_180
timestamp 1604681595
transform 1 0 17664 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 19504 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1604681595
transform 1 0 19688 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 19320 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 18952 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 19504 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_192
timestamp 1604681595
transform 1 0 18768 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_196
timestamp 1604681595
transform 1 0 19136 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_192
timestamp 1604681595
transform 1 0 18768 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_205
timestamp 1604681595
transform 1 0 19964 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604681595
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_prog_clk_A
timestamp 1604681595
transform 1 0 20516 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_219
timestamp 1604681595
transform 1 0 21252 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_213
timestamp 1604681595
transform 1 0 20700 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1604681595
transform 1 0 20884 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_227
timestamp 1604681595
transform 1 0 21988 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_237
timestamp 1604681595
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_233
timestamp 1604681595
transform 1 0 22540 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 23092 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1604681595
transform 1 0 22356 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_248
timestamp 1604681595
transform 1 0 23920 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_240
timestamp 1604681595
transform 1 0 23184 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1604681595
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_241
timestamp 1604681595
transform 1 0 23276 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23920 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604681595
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 24104 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1604681595
transform 1 0 24104 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1604681595
transform 1 0 25668 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_259
timestamp 1604681595
transform 1 0 24932 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_252
timestamp 1604681595
transform 1 0 24288 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_264
timestamp 1604681595
transform 1 0 25392 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_269
timestamp 1604681595
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604681595
transform 1 0 27232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604681595
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_276
timestamp 1604681595
transform 1 0 26496 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_287
timestamp 1604681595
transform 1 0 27508 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_273
timestamp 1604681595
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1604681595
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1604681595
transform 1 0 27600 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604681595
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604681595
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1604681595
transform 1 0 28336 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 1840 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604681595
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 1656 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1604681595
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 4324 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 3772 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_27
timestamp 1604681595
transform 1 0 3588 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1604681595
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604681595
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 5336 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_44
timestamp 1604681595
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1604681595
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_52
timestamp 1604681595
transform 1 0 5888 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1604681595
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_62
timestamp 1604681595
transform 1 0 6808 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8188 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_70
timestamp 1604681595
transform 1 0 7544 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1604681595
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_prog_clk_A
timestamp 1604681595
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1604681595
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_90
timestamp 1604681595
transform 1 0 9384 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_102
timestamp 1604681595
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1604681595
transform 1 0 10764 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1604681595
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604681595
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604681595
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604681595
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 13800 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604681595
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1604681595
transform 1 0 13616 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_140
timestamp 1604681595
transform 1 0 13984 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15732 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 15548 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 15180 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 14812 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_148
timestamp 1604681595
transform 1 0 14720 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_151
timestamp 1604681595
transform 1 0 14996 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_155
timestamp 1604681595
transform 1 0 15364 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604681595
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_168
timestamp 1604681595
transform 1 0 16560 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_172
timestamp 1604681595
transform 1 0 16928 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604681595
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_184
timestamp 1604681595
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19228 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19044 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 18676 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_190
timestamp 1604681595
transform 1 0 18584 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1604681595
transform 1 0 18860 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 21804 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_216
timestamp 1604681595
transform 1 0 20976 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_220
timestamp 1604681595
transform 1 0 21344 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_223
timestamp 1604681595
transform 1 0 21620 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_227
timestamp 1604681595
transform 1 0 21988 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604681595
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23920 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_239
timestamp 1604681595
transform 1 0 23092 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1604681595
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_245
timestamp 1604681595
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_250
timestamp 1604681595
transform 1 0 24104 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 25852 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 24288 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_254
timestamp 1604681595
transform 1 0 24472 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_266
timestamp 1604681595
transform 1 0 25576 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 26036 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_21_290
timestamp 1604681595
transform 1 0 27784 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604681595
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_298
timestamp 1604681595
transform 1 0 28520 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604681595
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 1748 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 2116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 2484 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1604681595
transform 1 0 1380 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_9
timestamp 1604681595
transform 1 0 1932 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 1604681595
transform 1 0 2300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1604681595
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604681595
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 4324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_21
timestamp 1604681595
transform 1 0 3036 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604681595
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 1604681595
transform 1 0 4048 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_37
timestamp 1604681595
transform 1 0 4508 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1604681595
transform 1 0 4876 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 4968 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_61
timestamp 1604681595
transform 1 0 6716 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1604681595
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_73
timestamp 1604681595
transform 1 0 7820 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1604681595
transform 1 0 8372 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1604681595
transform 1 0 8740 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604681595
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1604681595
transform 1 0 8832 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_87
timestamp 1604681595
transform 1 0 9108 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1604681595
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1604681595
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1604681595
transform 1 0 11500 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 12512 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 11316 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1604681595
transform 1 0 10948 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_122
timestamp 1604681595
transform 1 0 12328 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1604681595
transform 1 0 13064 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_126
timestamp 1604681595
transform 1 0 12696 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_139
timestamp 1604681595
transform 1 0 13892 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 16100 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604681595
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1604681595
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1604681595
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_160
timestamp 1604681595
transform 1 0 15824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_182
timestamp 1604681595
transform 1 0 17848 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_190
timestamp 1604681595
transform 1 0 18584 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_195
timestamp 1604681595
transform 1 0 19044 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_199
timestamp 1604681595
transform 1 0 19412 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_202
timestamp 1604681595
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_206
timestamp 1604681595
transform 1 0 20056 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 21436 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604681595
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1604681595
transform 1 0 20516 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 1604681595
transform 1 0 20424 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_215
timestamp 1604681595
transform 1 0 20884 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23920 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_22_240
timestamp 1604681595
transform 1 0 23184 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604681595
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604681595
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1604681595
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1604681595
transform 1 0 27600 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604681595
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1604681595
transform 1 0 28336 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1604681595
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604681595
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604681595
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1604681595
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604681595
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604681595
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1604681595
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1604681595
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604681595
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1604681595
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1604681595
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1604681595
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 7636 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_prog_clk_A
timestamp 1604681595
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_67
timestamp 1604681595
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 9660 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_90
timestamp 1604681595
transform 1 0 9384 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_95
timestamp 1604681595
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_99
timestamp 1604681595
transform 1 0 10212 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1604681595
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604681595
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 11500 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_111
timestamp 1604681595
transform 1 0 11316 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_115
timestamp 1604681595
transform 1 0 11684 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_119
timestamp 1604681595
transform 1 0 12052 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_132
timestamp 1604681595
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1604681595
transform 1 0 15640 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 15088 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_146
timestamp 1604681595
transform 1 0 14536 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1604681595
transform 1 0 14904 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1604681595
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604681595
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_prog_clk_A
timestamp 1604681595
transform 1 0 18216 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_167
timestamp 1604681595
transform 1 0 16468 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1604681595
transform 1 0 17572 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_184
timestamp 1604681595
transform 1 0 18032 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 19504 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1604681595
transform 1 0 18768 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_188
timestamp 1604681595
transform 1 0 18400 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1604681595
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_199
timestamp 1604681595
transform 1 0 19412 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_219
timestamp 1604681595
transform 1 0 21252 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_229
timestamp 1604681595
transform 1 0 22172 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604681595
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_233
timestamp 1604681595
transform 1 0 22540 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1604681595
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1604681595
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1604681595
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_269
timestamp 1604681595
transform 1 0 25852 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604681595
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_275
timestamp 1604681595
transform 1 0 26404 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_278
timestamp 1604681595
transform 1 0 26680 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_290
timestamp 1604681595
transform 1 0 27784 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604681595
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_298
timestamp 1604681595
transform 1 0 28520 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1604681595
transform 1 0 1748 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604681595
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 2760 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604681595
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_16
timestamp 1604681595
transform 1 0 2576 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1604681595
transform 1 0 2944 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604681595
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_28
timestamp 1604681595
transform 1 0 3680 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1604681595
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1604681595
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_56
timestamp 1604681595
transform 1 0 6256 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1604681595
transform 1 0 7084 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_64
timestamp 1604681595
transform 1 0 6992 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1604681595
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1604681595
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 9660 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604681595
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_112
timestamp 1604681595
transform 1 0 11408 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_120
timestamp 1604681595
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1604681595
transform 1 0 12604 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 12788 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1604681595
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1604681595
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604681595
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_173
timestamp 1604681595
transform 1 0 17020 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_185
timestamp 1604681595
transform 1 0 18124 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1604681595
transform 1 0 18860 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_190
timestamp 1604681595
transform 1 0 18584 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1604681595
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 21988 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604681595
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1604681595
transform 1 0 20884 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_246
timestamp 1604681595
transform 1 0 23736 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 24472 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 24840 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 25852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_256
timestamp 1604681595
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_260
timestamp 1604681595
transform 1 0 25024 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_268
timestamp 1604681595
transform 1 0 25760 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604681595
transform 1 0 26496 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604681595
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1604681595
transform 1 0 26036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_280
timestamp 1604681595
transform 1 0 26864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604681595
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_292
timestamp 1604681595
transform 1 0 27968 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_298
timestamp 1604681595
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 2208 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604681595
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 1840 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1604681595
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1604681595
transform 1 0 1748 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_10
timestamp 1604681595
transform 1 0 2024 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_31
timestamp 1604681595
transform 1 0 3956 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_39
timestamp 1604681595
transform 1 0 4692 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 6808 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604681595
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1604681595
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_46
timestamp 1604681595
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_58
timestamp 1604681595
transform 1 0 6440 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_81
timestamp 1604681595
transform 1 0 8556 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1604681595
transform 1 0 9844 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 9660 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 9292 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_prog_clk_A
timestamp 1604681595
transform 1 0 10672 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_91
timestamp 1604681595
transform 1 0 9476 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_98
timestamp 1604681595
transform 1 0 10120 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_102
timestamp 1604681595
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 12420 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604681595
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_106
timestamp 1604681595
transform 1 0 10856 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604681595
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604681595
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_142
timestamp 1604681595
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1604681595
transform 1 0 15456 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 15272 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1604681595
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_152
timestamp 1604681595
transform 1 0 15088 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_165
timestamp 1604681595
transform 1 0 16284 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1604681595
transform 1 0 16652 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 16836 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 16468 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_173
timestamp 1604681595
transform 1 0 17020 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 17204 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1604681595
transform 1 0 17388 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 1604681595
transform 1 0 18032 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 18216 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604681595
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1604681595
transform 1 0 18400 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 19412 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 20148 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1604681595
transform 1 0 19228 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_201
timestamp 1604681595
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1604681595
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 21252 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 21620 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_209
timestamp 1604681595
transform 1 0 20332 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_217
timestamp 1604681595
transform 1 0 21068 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1604681595
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1604681595
transform 1 0 21804 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604681595
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 24104 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_237
timestamp 1604681595
transform 1 0 22908 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_241
timestamp 1604681595
transform 1 0 23276 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1604681595
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_249
timestamp 1604681595
transform 1 0 24012 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 25852 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1604681595
transform 1 0 24288 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 25300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 25668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_261
timestamp 1604681595
transform 1 0 25116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_265
timestamp 1604681595
transform 1 0 25484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_288
timestamp 1604681595
transform 1 0 27600 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604681595
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_296
timestamp 1604681595
transform 1 0 28336 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1604681595
transform 1 0 1748 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604681595
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_3
timestamp 1604681595
transform 1 0 1380 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 1656 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604681595
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604681595
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604681595
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1604681595
transform 1 0 1840 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1604681595
transform 1 0 1840 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1604681595
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_17
timestamp 1604681595
transform 1 0 2668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 2852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 2852 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604681595
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_21
timestamp 1604681595
transform 1 0 3036 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1604681595
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_21
timestamp 1604681595
transform 1 0 3036 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604681595
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_37
timestamp 1604681595
transform 1 0 4508 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1604681595
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_37
timestamp 1604681595
transform 1 0 4508 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 1604681595
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1604681595
transform 1 0 4784 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4784 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604681595
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_59
timestamp 1604681595
transform 1 0 6532 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_49
timestamp 1604681595
transform 1 0 5612 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604681595
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp 1604681595
transform 1 0 6348 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1604681595
transform 1 0 6808 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 8004 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_71
timestamp 1604681595
transform 1 0 7636 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_83
timestamp 1604681595
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1604681595
transform 1 0 7544 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1604681595
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_77
timestamp 1604681595
transform 1 0 8188 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1604681595
transform 1 0 8556 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_88
timestamp 1604681595
transform 1 0 9200 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 9016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604681595
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604681595
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604681595
transform 1 0 9016 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1604681595
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1604681595
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1604681595
transform 1 0 10212 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1604681595
transform 1 0 9844 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 10396 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 10028 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_102
timestamp 1604681595
transform 1 0 10488 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 12328 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604681595
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_114
timestamp 1604681595
transform 1 0 11592 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_27_107
timestamp 1604681595
transform 1 0 10948 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_119
timestamp 1604681595
transform 1 0 12052 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604681595
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_141
timestamp 1604681595
transform 1 0 14076 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1604681595
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1604681595
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1604681595
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1604681595
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_154
timestamp 1604681595
transform 1 0 15272 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1604681595
transform 1 0 14812 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604681595
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1604681595
transform 1 0 15088 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1604681595
transform 1 0 15456 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_165
timestamp 1604681595
transform 1 0 16284 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1604681595
transform 1 0 15916 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 16100 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1604681595
transform 1 0 16284 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_173
timestamp 1604681595
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1604681595
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__S
timestamp 1604681595
transform 1 0 16468 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1604681595
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1604681595
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604681595
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_177
timestamp 1604681595
transform 1 0 17388 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_177
timestamp 1604681595
transform 1 0 17388 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604681595
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_185
timestamp 1604681595
transform 1 0 18124 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1604681595
transform 1 0 18400 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1604681595
transform 1 0 18400 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 20056 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1604681595
transform 1 0 19228 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_197
timestamp 1604681595
transform 1 0 19228 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_205
timestamp 1604681595
transform 1 0 19964 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 1604681595
transform 1 0 20240 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 20608 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1604681595
transform 1 0 20884 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604681595
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 20424 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_209
timestamp 1604681595
transform 1 0 20332 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_224
timestamp 1604681595
transform 1 0 21712 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_235
timestamp 1604681595
transform 1 0 22724 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_231
timestamp 1604681595
transform 1 0 22356 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 22540 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1604681595
transform 1 0 24104 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_245
timestamp 1604681595
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604681595
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1604681595
transform 1 0 24104 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 23920 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1604681595
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604681595
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_236
timestamp 1604681595
transform 1 0 22816 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1604681595
transform 1 0 24472 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1604681595
transform 1 0 24472 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1604681595
transform 1 0 24288 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1604681595
transform 1 0 24288 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1604681595
transform 1 0 25300 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_263
timestamp 1604681595
transform 1 0 25300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604681595
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604681595
transform 1 0 26496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1604681595
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1604681595
transform 1 0 27600 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_275
timestamp 1604681595
transform 1 0 26404 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_278
timestamp 1604681595
transform 1 0 26680 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_290
timestamp 1604681595
transform 1 0 27784 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604681595
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604681595
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1604681595
transform 1 0 28336 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1604681595
transform 1 0 28520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604681595
transform 1 0 1380 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604681595
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604681595
transform 1 0 1932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 2300 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1604681595
transform 1 0 1748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1604681595
transform 1 0 2116 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1604681595
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1604681595
transform 1 0 2852 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1604681595
transform 1 0 4324 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604681595
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 3772 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1604681595
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1604681595
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 5336 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1604681595
transform 1 0 5152 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_48
timestamp 1604681595
transform 1 0 5520 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1604681595
transform 1 0 6624 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604681595
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 7728 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_66
timestamp 1604681595
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1604681595
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_74
timestamp 1604681595
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604681595
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604681595
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604681595
transform 1 0 9016 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1604681595
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1604681595
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_102
timestamp 1604681595
transform 1 0 10488 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_114
timestamp 1604681595
transform 1 0 11592 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_122
timestamp 1604681595
transform 1 0 12328 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_125
timestamp 1604681595
transform 1 0 12604 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 13616 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 13984 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_133
timestamp 1604681595
transform 1 0 13340 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1604681595
transform 1 0 13800 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_142
timestamp 1604681595
transform 1 0 14168 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1604681595
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604681595
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 14996 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_146
timestamp 1604681595
transform 1 0 14536 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1604681595
transform 1 0 14812 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_163
timestamp 1604681595
transform 1 0 16100 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1604681595
transform 1 0 16836 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_28_180
timestamp 1604681595
transform 1 0 17664 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 18400 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 20240 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1604681595
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_202
timestamp 1604681595
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1604681595
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604681595
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1604681595
transform 1 0 20424 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_224
timestamp 1604681595
transform 1 0 21712 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1604681595
transform 1 0 23920 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__S
timestamp 1604681595
transform 1 0 23736 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 23368 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_236
timestamp 1604681595
transform 1 0 22816 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_244
timestamp 1604681595
transform 1 0 23552 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__S
timestamp 1604681595
transform 1 0 24932 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_257
timestamp 1604681595
transform 1 0 24748 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_261
timestamp 1604681595
transform 1 0 25116 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_269
timestamp 1604681595
transform 1 0 25852 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604681595
transform 1 0 26496 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604681595
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 26128 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_274
timestamp 1604681595
transform 1 0 26312 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_280
timestamp 1604681595
transform 1 0 26864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604681595
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_292
timestamp 1604681595
transform 1 0 27968 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_298
timestamp 1604681595
transform 1 0 28520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 1656 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604681595
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1604681595
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1604681595
transform 1 0 4232 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 3680 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_25
timestamp 1604681595
transform 1 0 3404 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_30
timestamp 1604681595
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1604681595
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 5244 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1604681595
transform 1 0 5796 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_47
timestamp 1604681595
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1604681595
transform 1 0 6348 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604681595
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604681595
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1604681595
transform 1 0 8648 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604681595
transform 1 0 7084 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 8096 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604681595
transform 1 0 8464 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1604681595
transform 1 0 7912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1604681595
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 10672 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_91
timestamp 1604681595
transform 1 0 9476 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_103
timestamp 1604681595
transform 1 0 10580 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604681595
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604681595
transform 1 0 11040 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1604681595
transform 1 0 10856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_110
timestamp 1604681595
transform 1 0 11224 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604681595
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1604681595
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1604681595
transform 1 0 14904 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1604681595
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_159
timestamp 1604681595
transform 1 0 15732 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_164
timestamp 1604681595
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604681595
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 18216 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_168
timestamp 1604681595
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_172
timestamp 1604681595
transform 1 0 16928 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_180
timestamp 1604681595
transform 1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_184
timestamp 1604681595
transform 1 0 18032 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1604681595
transform 1 0 20240 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1604681595
transform 1 0 18400 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_192
timestamp 1604681595
transform 1 0 18768 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_204
timestamp 1604681595
transform 1 0 19872 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 21252 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 21620 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 21988 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_217
timestamp 1604681595
transform 1 0 21068 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1604681595
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1604681595
transform 1 0 21804 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1604681595
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1604681595
transform 1 0 23736 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604681595
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1604681595
transform 1 0 23368 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__S
timestamp 1604681595
transform 1 0 23000 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_0__A0
timestamp 1604681595
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_233
timestamp 1604681595
transform 1 0 22540 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_236
timestamp 1604681595
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_240
timestamp 1604681595
transform 1 0 23184 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_245
timestamp 1604681595
transform 1 0 23644 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604681595
transform 1 0 25944 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A1
timestamp 1604681595
transform 1 0 24748 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_255
timestamp 1604681595
transform 1 0 24564 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_259
timestamp 1604681595
transform 1 0 24932 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_267
timestamp 1604681595
transform 1 0 25668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 26128 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_291
timestamp 1604681595
transform 1 0 27876 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604681595
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604681595
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604681595
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1604681595
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1604681595
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1604681595
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1604681595
transform 1 0 4324 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604681595
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1604681595
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_32
timestamp 1604681595
transform 1 0 4048 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1604681595
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_56
timestamp 1604681595
transform 1 0 6256 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604681595
transform 1 0 7360 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604681595
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1604681595
transform 1 0 6992 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_67
timestamp 1604681595
transform 1 0 7268 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_77
timestamp 1604681595
transform 1 0 8188 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_81
timestamp 1604681595
transform 1 0 8556 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604681595
transform 1 0 10672 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604681595
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604681595
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1604681595
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1604681595
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_93
timestamp 1604681595
transform 1 0 9660 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_101
timestamp 1604681595
transform 1 0 10396 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_30_123
timestamp 1604681595
transform 1 0 12420 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1604681595
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 13064 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_129
timestamp 1604681595
transform 1 0 12972 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_132
timestamp 1604681595
transform 1 0 13248 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_145
timestamp 1604681595
transform 1 0 14444 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1604681595
transform 1 0 16008 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604681595
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 15548 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_0__A1
timestamp 1604681595
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_149
timestamp 1604681595
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1604681595
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_154
timestamp 1604681595
transform 1 0 15272 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_159
timestamp 1604681595
transform 1 0 15732 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 18216 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_30_171
timestamp 1604681595
transform 1 0 16836 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_183
timestamp 1604681595
transform 1 0 17940 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 20240 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_205
timestamp 1604681595
transform 1 0 19964 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1604681595
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604681595
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1604681595
transform 1 0 20424 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_224
timestamp 1604681595
transform 1 0 21712 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1604681595
transform 1 0 23368 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_30_236
timestamp 1604681595
transform 1 0 22816 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1604681595
transform 1 0 25484 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__S
timestamp 1604681595
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 24932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_251
timestamp 1604681595
transform 1 0 24196 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_257
timestamp 1604681595
transform 1 0 24748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_261
timestamp 1604681595
transform 1 0 25116 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_267
timestamp 1604681595
transform 1 0 25668 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604681595
transform 1 0 26496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604681595
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_279
timestamp 1604681595
transform 1 0 26772 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_291
timestamp 1604681595
transform 1 0 27876 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604681595
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604681595
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604681595
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1604681595
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604681595
transform 1 0 4416 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 4876 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1604681595
transform 1 0 3588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_35
timestamp 1604681595
transform 1 0 4324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1604681595
transform 1 0 4692 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604681595
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 5244 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_43
timestamp 1604681595
transform 1 0 5060 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1604681595
transform 1 0 5428 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1604681595
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1604681595
transform 1 0 6808 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604681595
transform 1 0 7360 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 7176 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 8740 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_77
timestamp 1604681595
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1604681595
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604681595
transform 1 0 8924 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_88
timestamp 1604681595
transform 1 0 9200 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_100
timestamp 1604681595
transform 1 0 10304 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604681595
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 10948 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1604681595
transform 1 0 10764 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_109
timestamp 1604681595
transform 1 0 11132 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_121
timestamp 1604681595
transform 1 0 12236 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1604681595
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 13064 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 12880 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 1604681595
transform 1 0 12788 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1604681595
transform 1 0 15548 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 15364 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1604681595
transform 1 0 14812 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_153
timestamp 1604681595
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1604681595
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604681595
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_170
timestamp 1604681595
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_174
timestamp 1604681595
transform 1 0 17112 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1604681595
transform 1 0 17848 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1604681595
transform 1 0 18032 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1604681595
transform 1 0 19136 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_208
timestamp 1604681595
transform 1 0 20240 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604681595
transform 1 0 20332 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 21804 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 22172 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_212
timestamp 1604681595
transform 1 0 20608 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_224
timestamp 1604681595
transform 1 0 21712 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_227
timestamp 1604681595
transform 1 0 21988 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1604681595
transform 1 0 23644 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604681595
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 23000 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_231
timestamp 1604681595
transform 1 0 22356 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1604681595
transform 1 0 22908 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_240
timestamp 1604681595
transform 1 0 23184 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1604681595
transform 1 0 25484 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1604681595
transform 1 0 25300 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__S
timestamp 1604681595
transform 1 0 24932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_254
timestamp 1604681595
transform 1 0 24472 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_258
timestamp 1604681595
transform 1 0 24840 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_261
timestamp 1604681595
transform 1 0 25116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1604681595
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A0
timestamp 1604681595
transform 1 0 26864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__S
timestamp 1604681595
transform 1 0 27232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_274
timestamp 1604681595
transform 1 0 26312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1604681595
transform 1 0 26680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_282
timestamp 1604681595
transform 1 0 27048 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_286
timestamp 1604681595
transform 1 0 27416 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604681595
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_298
timestamp 1604681595
transform 1 0 28520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604681595
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 2944 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604681595
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_15
timestamp 1604681595
transform 1 0 2484 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_19
timestamp 1604681595
transform 1 0 2852 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 4600 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604681595
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_22
timestamp 1604681595
transform 1 0 3128 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604681595
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_32
timestamp 1604681595
transform 1 0 4048 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_57
timestamp 1604681595
transform 1 0 6348 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_61
timestamp 1604681595
transform 1 0 6716 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604681595
transform 1 0 7084 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 8464 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_64
timestamp 1604681595
transform 1 0 6992 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_74
timestamp 1604681595
transform 1 0 7912 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_82
timestamp 1604681595
transform 1 0 8648 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 10580 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604681595
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604681595
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_93
timestamp 1604681595
transform 1 0 9660 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1604681595
transform 1 0 10396 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_122
timestamp 1604681595
transform 1 0 12328 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604681595
transform 1 0 13892 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_134
timestamp 1604681595
transform 1 0 13432 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_138
timestamp 1604681595
transform 1 0 13800 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1604681595
transform 1 0 14076 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1604681595
transform 1 0 16100 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604681595
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l3_in_1__A1
timestamp 1604681595
transform 1 0 15548 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_154
timestamp 1604681595
transform 1 0 15272 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_159
timestamp 1604681595
transform 1 0 15732 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604681595
transform 1 0 17664 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_172
timestamp 1604681595
transform 1 0 16928 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_183
timestamp 1604681595
transform 1 0 17940 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604681595
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_195
timestamp 1604681595
transform 1 0 19044 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1604681595
transform 1 0 19596 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 21804 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604681595
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604681595
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_215
timestamp 1604681595
transform 1 0 20884 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_223
timestamp 1604681595
transform 1 0 21620 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__A1
timestamp 1604681595
transform 1 0 23736 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_244
timestamp 1604681595
transform 1 0 23552 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_248
timestamp 1604681595
transform 1 0 23920 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1604681595
transform 1 0 24564 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l3_in_1__A0
timestamp 1604681595
transform 1 0 24380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_252
timestamp 1604681595
transform 1 0 24288 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_264
timestamp 1604681595
transform 1 0 25392 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1604681595
transform 1 0 26496 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604681595
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_272
timestamp 1604681595
transform 1 0 26128 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_285
timestamp 1604681595
transform 1 0 27324 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604681595
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_297
timestamp 1604681595
transform 1 0 28428 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_10
timestamp 1604681595
transform 1 0 2024 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1604681595
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604681595
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604681595
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604681595
transform 1 0 1656 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_14
timestamp 1604681595
transform 1 0 2392 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 2760 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604681595
transform 1 0 2208 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604681595
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604681595
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 2944 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604681595
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1604681595
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604681595
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1604681595
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604681595
transform 1 0 6808 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604681595
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604681595
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604681595
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604681595
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1604681595
transform 1 0 5796 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604681595
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1604681595
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_56
timestamp 1604681595
transform 1 0 6256 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 8464 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_71
timestamp 1604681595
transform 1 0 7636 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_77
timestamp 1604681595
transform 1 0 8188 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1604681595
transform 1 0 7176 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_78
timestamp 1604681595
transform 1 0 8280 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604681595
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_99
timestamp 1604681595
transform 1 0 10212 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1604681595
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604681595
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604681595
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_111
timestamp 1604681595
transform 1 0 11316 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_119
timestamp 1604681595
transform 1 0 12052 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604681595
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604681595
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1604681595
transform 1 0 11868 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604681595
transform 1 0 13892 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604681595
transform 1 0 13708 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1604681595
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1604681595
transform 1 0 12972 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1604681595
transform 1 0 14076 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604681595
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_158
timestamp 1604681595
transform 1 0 15640 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_166
timestamp 1604681595
transform 1 0 16376 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604681595
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1604681595
transform 1 0 16376 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604681595
transform 1 0 16652 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604681595
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604681595
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1604681595
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_179
timestamp 1604681595
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1604681595
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1604681595
transform 1 0 17480 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604681595
transform 1 0 19412 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_mode_io__0.ltile_physical_iopad_0.EMBEDDED_IO_mem.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604681595
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1604681595
transform 1 0 19136 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1604681595
transform 1 0 18584 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1604681595
transform 1 0 19688 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1604681595
transform 1 0 20884 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604681595
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1604681595
transform 1 0 21344 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_218
timestamp 1604681595
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_222
timestamp 1604681595
transform 1 0 21528 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_219
timestamp 1604681595
transform 1 0 21252 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604681595
transform 1 0 23644 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604681595
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604681595
transform 1 0 23368 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604681595
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_234
timestamp 1604681595
transform 1 0 22632 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_231
timestamp 1604681595
transform 1 0 22356 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_243
timestamp 1604681595
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_247
timestamp 1604681595
transform 1 0 23828 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_264
timestamp 1604681595
transform 1 0 25392 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_259
timestamp 1604681595
transform 1 0 24932 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1604681595
transform 1 0 26404 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604681595
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1604681595
transform 1 0 26956 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_272
timestamp 1604681595
transform 1 0 26128 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_279
timestamp 1604681595
transform 1 0 26772 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_283
timestamp 1604681595
transform 1 0 27140 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1604681595
transform 1 0 26036 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604681595
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604681595
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604681595
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604681595
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_295
timestamp 1604681595
transform 1 0 28244 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604681595
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604681595
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604681595
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604681595
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604681595
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604681595
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604681595
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604681595
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604681595
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604681595
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604681595
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604681595
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604681595
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604681595
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604681595
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604681595
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604681595
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604681595
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604681595
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604681595
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604681595
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604681595
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604681595
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604681595
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604681595
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604681595
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604681595
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604681595
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604681595
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604681595
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604681595
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604681595
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604681595
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604681595
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604681595
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604681595
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604681595
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604681595
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604681595
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604681595
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604681595
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604681595
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 2042 0 2098 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 4986 23520 5042 24000 6 SC_IN_TOP
port 1 nsew default input
rlabel metal2 s 3514 0 3570 480 6 SC_OUT_BOT
port 2 nsew default tristate
rlabel metal2 s 8298 23520 8354 24000 6 SC_OUT_TOP
port 3 nsew default tristate
rlabel metal2 s 4894 0 4950 480 6 bottom_grid_pin_0_
port 4 nsew default tristate
rlabel metal2 s 19154 0 19210 480 6 bottom_grid_pin_10_
port 5 nsew default tristate
rlabel metal2 s 20626 0 20682 480 6 bottom_grid_pin_11_
port 6 nsew default tristate
rlabel metal2 s 22006 0 22062 480 6 bottom_grid_pin_12_
port 7 nsew default tristate
rlabel metal2 s 23478 0 23534 480 6 bottom_grid_pin_13_
port 8 nsew default tristate
rlabel metal2 s 24858 0 24914 480 6 bottom_grid_pin_14_
port 9 nsew default tristate
rlabel metal2 s 26330 0 26386 480 6 bottom_grid_pin_15_
port 10 nsew default tristate
rlabel metal2 s 6366 0 6422 480 6 bottom_grid_pin_1_
port 11 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 bottom_grid_pin_2_
port 12 nsew default tristate
rlabel metal2 s 9218 0 9274 480 6 bottom_grid_pin_3_
port 13 nsew default tristate
rlabel metal2 s 10598 0 10654 480 6 bottom_grid_pin_4_
port 14 nsew default tristate
rlabel metal2 s 12070 0 12126 480 6 bottom_grid_pin_5_
port 15 nsew default tristate
rlabel metal2 s 13450 0 13506 480 6 bottom_grid_pin_6_
port 16 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 bottom_grid_pin_7_
port 17 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 bottom_grid_pin_8_
port 18 nsew default tristate
rlabel metal2 s 17774 0 17830 480 6 bottom_grid_pin_9_
port 19 nsew default tristate
rlabel metal2 s 27710 0 27766 480 6 bottom_width_0_height_0__pin_0_
port 20 nsew default input
rlabel metal2 s 29182 0 29238 480 6 bottom_width_0_height_0__pin_1_lower
port 21 nsew default tristate
rlabel metal2 s 662 0 718 480 6 bottom_width_0_height_0__pin_1_upper
port 22 nsew default tristate
rlabel metal2 s 11610 23520 11666 24000 6 ccff_head
port 23 nsew default input
rlabel metal2 s 14922 23520 14978 24000 6 ccff_tail
port 24 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 25 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 26 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 27 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 28 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 29 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 30 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 31 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 32 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 33 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 34 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 35 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 36 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 37 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 38 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 39 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 40 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 41 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 42 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 43 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 44 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 45 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 46 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 47 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 48 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 49 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 50 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 51 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 52 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 53 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 54 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 55 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 56 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 57 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 58 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 59 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 60 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 61 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 62 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 63 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 64 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 65 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 66 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 67 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 68 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 69 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 70 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 71 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 72 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 73 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 74 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 75 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 76 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 77 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 78 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 79 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 80 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 81 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 82 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 83 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 84 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 85 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 86 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 87 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 88 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 89 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 90 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 91 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 92 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 93 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 94 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 95 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 96 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 97 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 98 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 99 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 100 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 101 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 102 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 103 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 104 nsew default tristate
rlabel metal2 s 21638 23520 21694 24000 6 gfpga_pad_EMBEDDED_IO_SOC_DIR
port 105 nsew default tristate
rlabel metal2 s 24950 23520 25006 24000 6 gfpga_pad_EMBEDDED_IO_SOC_IN
port 106 nsew default input
rlabel metal2 s 28262 23520 28318 24000 6 gfpga_pad_EMBEDDED_IO_SOC_OUT
port 107 nsew default tristate
rlabel metal2 s 1674 23520 1730 24000 6 prog_clk
port 108 nsew default input
rlabel metal2 s 18326 23520 18382 24000 6 top_grid_pin_0_
port 109 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 110 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 111 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
