magic
tech sky130A
magscale 1 2
timestamp 1604668008
<< locali >>
rect 12081 2839 12115 3145
<< viali >>
rect 5641 36873 5675 36907
rect 5457 36669 5491 36703
rect 6009 36669 6043 36703
rect 4905 36329 4939 36363
rect 6009 36329 6043 36363
rect 4721 36193 4755 36227
rect 5825 36193 5859 36227
rect 2973 35785 3007 35819
rect 4077 35785 4111 35819
rect 5181 35785 5215 35819
rect 7481 35785 7515 35819
rect 9873 35717 9907 35751
rect 4813 35649 4847 35683
rect 2789 35581 2823 35615
rect 3801 35581 3835 35615
rect 3893 35581 3927 35615
rect 4997 35581 5031 35615
rect 7297 35581 7331 35615
rect 9689 35581 9723 35615
rect 3433 35445 3467 35479
rect 5641 35445 5675 35479
rect 6009 35445 6043 35479
rect 7941 35445 7975 35479
rect 10333 35445 10367 35479
rect 1593 35241 1627 35275
rect 2697 35241 2731 35275
rect 5089 35241 5123 35275
rect 6469 35241 6503 35275
rect 7573 35241 7607 35275
rect 1409 35105 1443 35139
rect 2513 35105 2547 35139
rect 4905 35105 4939 35139
rect 6285 35105 6319 35139
rect 7389 35105 7423 35139
rect 8493 35105 8527 35139
rect 9945 35105 9979 35139
rect 9689 35037 9723 35071
rect 12357 35037 12391 35071
rect 8677 34969 8711 35003
rect 7941 34901 7975 34935
rect 9505 34901 9539 34935
rect 11069 34901 11103 34935
rect 12909 34901 12943 34935
rect 1593 34697 1627 34731
rect 2697 34697 2731 34731
rect 7297 34697 7331 34731
rect 9689 34697 9723 34731
rect 11897 34697 11931 34731
rect 12265 34629 12299 34663
rect 3341 34561 3375 34595
rect 9873 34561 9907 34595
rect 13001 34561 13035 34595
rect 1409 34493 1443 34527
rect 1961 34493 1995 34527
rect 2421 34493 2455 34527
rect 2513 34493 2547 34527
rect 3065 34493 3099 34527
rect 3525 34493 3559 34527
rect 5549 34493 5583 34527
rect 6377 34493 6411 34527
rect 7389 34493 7423 34527
rect 7656 34493 7690 34527
rect 9321 34493 9355 34527
rect 3792 34425 3826 34459
rect 10140 34425 10174 34459
rect 12817 34425 12851 34459
rect 12909 34425 12943 34459
rect 4905 34357 4939 34391
rect 8769 34357 8803 34391
rect 11253 34357 11287 34391
rect 12449 34357 12483 34391
rect 2421 34153 2455 34187
rect 9505 34153 9539 34187
rect 9873 34153 9907 34187
rect 1685 34085 1719 34119
rect 11253 34085 11287 34119
rect 12072 34085 12106 34119
rect 2237 34017 2271 34051
rect 4977 34017 5011 34051
rect 7941 34017 7975 34051
rect 10517 34017 10551 34051
rect 11805 34017 11839 34051
rect 4721 33949 4755 33983
rect 8033 33949 8067 33983
rect 8217 33949 8251 33983
rect 10609 33949 10643 33983
rect 10793 33949 10827 33983
rect 7481 33881 7515 33915
rect 3617 33813 3651 33847
rect 6101 33813 6135 33847
rect 7021 33813 7055 33847
rect 7573 33813 7607 33847
rect 10149 33813 10183 33847
rect 13185 33813 13219 33847
rect 1593 33609 1627 33643
rect 3065 33609 3099 33643
rect 4169 33609 4203 33643
rect 5273 33609 5307 33643
rect 6285 33609 6319 33643
rect 8861 33609 8895 33643
rect 9413 33609 9447 33643
rect 11989 33609 12023 33643
rect 9689 33541 9723 33575
rect 10425 33541 10459 33575
rect 4997 33473 5031 33507
rect 6653 33473 6687 33507
rect 11253 33473 11287 33507
rect 13001 33473 13035 33507
rect 13461 33473 13495 33507
rect 1409 33405 1443 33439
rect 2881 33405 2915 33439
rect 3985 33405 4019 33439
rect 5089 33405 5123 33439
rect 5733 33405 5767 33439
rect 6837 33405 6871 33439
rect 9505 33405 9539 33439
rect 10057 33405 10091 33439
rect 12817 33405 12851 33439
rect 13829 33405 13863 33439
rect 1961 33337 1995 33371
rect 7082 33337 7116 33371
rect 11069 33337 11103 33371
rect 2329 33269 2363 33303
rect 3525 33269 3559 33303
rect 4629 33269 4663 33303
rect 8217 33269 8251 33303
rect 10609 33269 10643 33303
rect 10977 33269 11011 33303
rect 11621 33269 11655 33303
rect 12449 33269 12483 33303
rect 12909 33269 12943 33303
rect 1593 33065 1627 33099
rect 6101 33065 6135 33099
rect 7297 33065 7331 33099
rect 7665 33065 7699 33099
rect 10241 33065 10275 33099
rect 10517 33065 10551 33099
rect 11161 33065 11195 33099
rect 12265 33065 12299 33099
rect 12725 33065 12759 33099
rect 6929 32997 6963 33031
rect 11069 32997 11103 33031
rect 1409 32929 1443 32963
rect 12633 32929 12667 32963
rect 6193 32861 6227 32895
rect 6377 32861 6411 32895
rect 7757 32861 7791 32895
rect 7849 32861 7883 32895
rect 9689 32861 9723 32895
rect 11345 32861 11379 32895
rect 12817 32861 12851 32895
rect 10701 32793 10735 32827
rect 3341 32725 3375 32759
rect 4721 32725 4755 32759
rect 5733 32725 5767 32759
rect 8309 32725 8343 32759
rect 11805 32725 11839 32759
rect 13277 32725 13311 32759
rect 1593 32521 1627 32555
rect 5457 32521 5491 32555
rect 6193 32521 6227 32555
rect 6653 32521 6687 32555
rect 9137 32521 9171 32555
rect 9965 32521 9999 32555
rect 10793 32521 10827 32555
rect 11805 32521 11839 32555
rect 12173 32521 12207 32555
rect 12449 32521 12483 32555
rect 13829 32521 13863 32555
rect 5825 32453 5859 32487
rect 10333 32453 10367 32487
rect 13461 32453 13495 32487
rect 3801 32385 3835 32419
rect 11253 32385 11287 32419
rect 11437 32385 11471 32419
rect 13001 32385 13035 32419
rect 3709 32317 3743 32351
rect 7297 32317 7331 32351
rect 7757 32317 7791 32351
rect 8024 32317 8058 32351
rect 12909 32317 12943 32351
rect 3157 32249 3191 32283
rect 3249 32181 3283 32215
rect 3617 32181 3651 32215
rect 4629 32181 4663 32215
rect 10701 32181 10735 32215
rect 11161 32181 11195 32215
rect 12817 32181 12851 32215
rect 3341 31977 3375 32011
rect 6561 31977 6595 32011
rect 7021 31977 7055 32011
rect 8585 31977 8619 32011
rect 9689 31977 9723 32011
rect 10057 31977 10091 32011
rect 10149 31977 10183 32011
rect 10793 31977 10827 32011
rect 11253 31977 11287 32011
rect 11529 31977 11563 32011
rect 12541 31977 12575 32011
rect 4322 31909 4356 31943
rect 6929 31909 6963 31943
rect 4077 31773 4111 31807
rect 6469 31773 6503 31807
rect 7113 31773 7147 31807
rect 8125 31773 8159 31807
rect 10333 31773 10367 31807
rect 12817 31773 12851 31807
rect 5457 31637 5491 31671
rect 7849 31637 7883 31671
rect 4169 31433 4203 31467
rect 6929 31433 6963 31467
rect 7941 31433 7975 31467
rect 8493 31433 8527 31467
rect 9873 31433 9907 31467
rect 13553 31433 13587 31467
rect 2513 31365 2547 31399
rect 6285 31365 6319 31399
rect 10057 31365 10091 31399
rect 3617 31297 3651 31331
rect 5089 31297 5123 31331
rect 7573 31297 7607 31331
rect 8309 31297 8343 31331
rect 8953 31297 8987 31331
rect 9045 31297 9079 31331
rect 10609 31297 10643 31331
rect 11069 31297 11103 31331
rect 2881 31229 2915 31263
rect 8861 31229 8895 31263
rect 10425 31229 10459 31263
rect 13369 31229 13403 31263
rect 13829 31229 13863 31263
rect 2145 31161 2179 31195
rect 5549 31161 5583 31195
rect 2973 31093 3007 31127
rect 3341 31093 3375 31127
rect 3433 31093 3467 31127
rect 4537 31093 4571 31127
rect 4905 31093 4939 31127
rect 4997 31093 5031 31127
rect 6653 31093 6687 31127
rect 7297 31093 7331 31127
rect 7389 31093 7423 31127
rect 9505 31093 9539 31127
rect 10517 31093 10551 31127
rect 4077 30889 4111 30923
rect 6837 30889 6871 30923
rect 7573 30889 7607 30923
rect 8585 30889 8619 30923
rect 10425 30889 10459 30923
rect 10793 30889 10827 30923
rect 13001 30889 13035 30923
rect 3801 30821 3835 30855
rect 11888 30821 11922 30855
rect 4445 30753 4479 30787
rect 6929 30753 6963 30787
rect 11621 30753 11655 30787
rect 2973 30685 3007 30719
rect 4537 30685 4571 30719
rect 4721 30685 4755 30719
rect 5089 30685 5123 30719
rect 7021 30685 7055 30719
rect 6377 30617 6411 30651
rect 6469 30549 6503 30583
rect 10057 30549 10091 30583
rect 3801 30345 3835 30379
rect 5917 30345 5951 30379
rect 11621 30345 11655 30379
rect 12081 30345 12115 30379
rect 3433 30277 3467 30311
rect 4629 30277 4663 30311
rect 4169 30209 4203 30243
rect 5181 30209 5215 30243
rect 7297 30209 7331 30243
rect 7481 30209 7515 30243
rect 10241 30209 10275 30243
rect 7849 30141 7883 30175
rect 9229 30141 9263 30175
rect 10057 30141 10091 30175
rect 4997 30073 5031 30107
rect 6193 30073 6227 30107
rect 6653 30073 6687 30107
rect 9505 30073 9539 30107
rect 10149 30073 10183 30107
rect 4537 30005 4571 30039
rect 5089 30005 5123 30039
rect 6837 30005 6871 30039
rect 7205 30005 7239 30039
rect 9689 30005 9723 30039
rect 1593 29801 1627 29835
rect 4353 29801 4387 29835
rect 5733 29801 5767 29835
rect 6561 29801 6595 29835
rect 7665 29801 7699 29835
rect 9965 29801 9999 29835
rect 4629 29733 4663 29767
rect 6929 29733 6963 29767
rect 7573 29733 7607 29767
rect 1409 29665 1443 29699
rect 5641 29665 5675 29699
rect 8033 29665 8067 29699
rect 10600 29665 10634 29699
rect 5825 29597 5859 29631
rect 8125 29597 8159 29631
rect 8217 29597 8251 29631
rect 10333 29597 10367 29631
rect 5273 29461 5307 29495
rect 8769 29461 8803 29495
rect 11713 29461 11747 29495
rect 1593 29257 1627 29291
rect 1961 29257 1995 29291
rect 4077 29257 4111 29291
rect 4629 29257 4663 29291
rect 6009 29257 6043 29291
rect 6469 29257 6503 29291
rect 10701 29257 10735 29291
rect 8033 29189 8067 29223
rect 5181 29121 5215 29155
rect 5733 29121 5767 29155
rect 8677 29121 8711 29155
rect 10057 29121 10091 29155
rect 10241 29121 10275 29155
rect 1409 29053 1443 29087
rect 7297 29053 7331 29087
rect 8493 29053 8527 29087
rect 9413 29053 9447 29087
rect 9965 29053 9999 29087
rect 2329 28985 2363 29019
rect 4537 28985 4571 29019
rect 4997 28985 5031 29019
rect 7665 28985 7699 29019
rect 8401 28985 8435 29019
rect 5089 28917 5123 28951
rect 9045 28917 9079 28951
rect 9597 28917 9631 28951
rect 11069 28917 11103 28951
rect 2421 28713 2455 28747
rect 4905 28713 4939 28747
rect 10241 28713 10275 28747
rect 2789 28645 2823 28679
rect 11428 28645 11462 28679
rect 5273 28577 5307 28611
rect 6817 28577 6851 28611
rect 9965 28577 9999 28611
rect 2881 28509 2915 28543
rect 3065 28509 3099 28543
rect 5365 28509 5399 28543
rect 5549 28509 5583 28543
rect 6561 28509 6595 28543
rect 11161 28509 11195 28543
rect 7941 28441 7975 28475
rect 8953 28441 8987 28475
rect 12541 28441 12575 28475
rect 4629 28373 4663 28407
rect 8585 28373 8619 28407
rect 10701 28373 10735 28407
rect 2513 28169 2547 28203
rect 3157 28169 3191 28203
rect 5089 28169 5123 28203
rect 5641 28169 5675 28203
rect 7297 28169 7331 28203
rect 10609 28169 10643 28203
rect 12081 28169 12115 28203
rect 2881 28033 2915 28067
rect 11161 28033 11195 28067
rect 3709 27965 3743 27999
rect 8125 27965 8159 27999
rect 8392 27965 8426 27999
rect 11621 27965 11655 27999
rect 3954 27897 3988 27931
rect 6561 27897 6595 27931
rect 7941 27897 7975 27931
rect 10425 27897 10459 27931
rect 11069 27897 11103 27931
rect 3617 27829 3651 27863
rect 6101 27829 6135 27863
rect 6837 27829 6871 27863
rect 9505 27829 9539 27863
rect 10977 27829 11011 27863
rect 3801 27625 3835 27659
rect 4997 27625 5031 27659
rect 6653 27625 6687 27659
rect 7941 27625 7975 27659
rect 10057 27625 10091 27659
rect 10609 27625 10643 27659
rect 2881 27557 2915 27591
rect 5540 27557 5574 27591
rect 9045 27557 9079 27591
rect 11244 27557 11278 27591
rect 2789 27489 2823 27523
rect 8401 27489 8435 27523
rect 3065 27421 3099 27455
rect 5273 27421 5307 27455
rect 8493 27421 8527 27455
rect 8585 27421 8619 27455
rect 10977 27421 11011 27455
rect 2421 27353 2455 27387
rect 8033 27285 8067 27319
rect 12357 27285 12391 27319
rect 12909 27285 12943 27319
rect 1777 27081 1811 27115
rect 3985 27081 4019 27115
rect 5733 27081 5767 27115
rect 6837 27081 6871 27115
rect 9505 27081 9539 27115
rect 9873 27081 9907 27115
rect 11345 27081 11379 27115
rect 2145 27013 2179 27047
rect 2421 27013 2455 27047
rect 6561 27013 6595 27047
rect 7389 26945 7423 26979
rect 8861 26945 8895 26979
rect 8953 26945 8987 26979
rect 10609 26945 10643 26979
rect 13001 26945 13035 26979
rect 2605 26877 2639 26911
rect 6285 26877 6319 26911
rect 7297 26877 7331 26911
rect 8033 26877 8067 26911
rect 8769 26877 8803 26911
rect 2872 26809 2906 26843
rect 7205 26809 7239 26843
rect 10333 26809 10367 26843
rect 12817 26809 12851 26843
rect 5273 26741 5307 26775
rect 8401 26741 8435 26775
rect 9965 26741 9999 26775
rect 10425 26741 10459 26775
rect 10977 26741 11011 26775
rect 11805 26741 11839 26775
rect 12173 26741 12207 26775
rect 12449 26741 12483 26775
rect 12909 26741 12943 26775
rect 2973 26537 3007 26571
rect 6561 26537 6595 26571
rect 7205 26537 7239 26571
rect 7757 26537 7791 26571
rect 8217 26537 8251 26571
rect 9137 26537 9171 26571
rect 10333 26537 10367 26571
rect 10793 26537 10827 26571
rect 8125 26469 8159 26503
rect 5448 26401 5482 26435
rect 10701 26401 10735 26435
rect 12164 26401 12198 26435
rect 5181 26333 5215 26367
rect 8309 26333 8343 26367
rect 9965 26333 9999 26367
rect 10885 26333 10919 26367
rect 11897 26333 11931 26367
rect 2605 26265 2639 26299
rect 8861 26265 8895 26299
rect 13277 26265 13311 26299
rect 6837 25993 6871 26027
rect 7941 25993 7975 26027
rect 8309 25993 8343 26027
rect 10609 25993 10643 26027
rect 10885 25993 10919 26027
rect 5641 25857 5675 25891
rect 6285 25857 6319 25891
rect 7481 25857 7515 25891
rect 8585 25857 8619 25891
rect 9413 25857 9447 25891
rect 10057 25857 10091 25891
rect 11069 25857 11103 25891
rect 12633 25857 12667 25891
rect 6653 25789 6687 25823
rect 7205 25789 7239 25823
rect 9873 25789 9907 25823
rect 11897 25789 11931 25823
rect 9045 25721 9079 25755
rect 5181 25653 5215 25687
rect 7297 25653 7331 25687
rect 9505 25653 9539 25687
rect 9965 25653 9999 25687
rect 1593 25449 1627 25483
rect 6929 25449 6963 25483
rect 9505 25449 9539 25483
rect 10793 25449 10827 25483
rect 1409 25313 1443 25347
rect 10057 25313 10091 25347
rect 4537 25245 4571 25279
rect 10149 25245 10183 25279
rect 10333 25245 10367 25279
rect 9689 25177 9723 25211
rect 8033 25109 8067 25143
rect 9045 24905 9079 24939
rect 9781 24905 9815 24939
rect 10057 24837 10091 24871
rect 4353 24769 4387 24803
rect 4905 24769 4939 24803
rect 5089 24769 5123 24803
rect 5457 24769 5491 24803
rect 7481 24769 7515 24803
rect 8493 24769 8527 24803
rect 9321 24769 9355 24803
rect 10701 24769 10735 24803
rect 11437 24769 11471 24803
rect 1961 24701 1995 24735
rect 3985 24701 4019 24735
rect 4813 24701 4847 24735
rect 7757 24701 7791 24735
rect 8401 24701 8435 24735
rect 10425 24701 10459 24735
rect 2228 24633 2262 24667
rect 1869 24565 1903 24599
rect 3341 24565 3375 24599
rect 4445 24565 4479 24599
rect 7941 24565 7975 24599
rect 8309 24565 8343 24599
rect 10517 24565 10551 24599
rect 11069 24565 11103 24599
rect 1593 24361 1627 24395
rect 2329 24361 2363 24395
rect 2697 24361 2731 24395
rect 4077 24361 4111 24395
rect 7113 24361 7147 24395
rect 7665 24361 7699 24395
rect 10149 24361 10183 24395
rect 10793 24361 10827 24395
rect 7573 24293 7607 24327
rect 4445 24225 4479 24259
rect 10057 24225 10091 24259
rect 11520 24225 11554 24259
rect 2789 24157 2823 24191
rect 2973 24157 3007 24191
rect 4537 24157 4571 24191
rect 4721 24157 4755 24191
rect 7849 24157 7883 24191
rect 10241 24157 10275 24191
rect 11253 24157 11287 24191
rect 2053 24021 2087 24055
rect 3433 24021 3467 24055
rect 5273 24021 5307 24055
rect 7205 24021 7239 24055
rect 9689 24021 9723 24055
rect 12633 24021 12667 24055
rect 2329 23817 2363 23851
rect 5365 23817 5399 23851
rect 6653 23817 6687 23851
rect 9137 23817 9171 23851
rect 9781 23817 9815 23851
rect 10425 23817 10459 23851
rect 4353 23749 4387 23783
rect 5733 23749 5767 23783
rect 7297 23749 7331 23783
rect 1961 23681 1995 23715
rect 3433 23681 3467 23715
rect 3893 23681 3927 23715
rect 4997 23681 5031 23715
rect 4261 23613 4295 23647
rect 4721 23613 4755 23647
rect 7757 23613 7791 23647
rect 8024 23613 8058 23647
rect 2697 23545 2731 23579
rect 4813 23545 4847 23579
rect 2789 23477 2823 23511
rect 3157 23477 3191 23511
rect 3249 23477 3283 23511
rect 7573 23477 7607 23511
rect 10149 23477 10183 23511
rect 11253 23477 11287 23511
rect 11713 23477 11747 23511
rect 1593 23273 1627 23307
rect 2329 23273 2363 23307
rect 2421 23273 2455 23307
rect 3893 23273 3927 23307
rect 4445 23273 4479 23307
rect 5917 23273 5951 23307
rect 7021 23273 7055 23307
rect 7389 23273 7423 23307
rect 8401 23273 8435 23307
rect 11069 23273 11103 23307
rect 12633 23273 12667 23307
rect 1961 23205 1995 23239
rect 2789 23205 2823 23239
rect 8033 23205 8067 23239
rect 12541 23205 12575 23239
rect 1409 23137 1443 23171
rect 4804 23137 4838 23171
rect 9689 23137 9723 23171
rect 9956 23137 9990 23171
rect 2881 23069 2915 23103
rect 3065 23069 3099 23103
rect 4537 23069 4571 23103
rect 6561 23069 6595 23103
rect 7481 23069 7515 23103
rect 7573 23069 7607 23103
rect 12817 23069 12851 23103
rect 6929 23001 6963 23035
rect 12173 22933 12207 22967
rect 13277 22933 13311 22967
rect 1869 22729 1903 22763
rect 4077 22729 4111 22763
rect 8217 22729 8251 22763
rect 8953 22729 8987 22763
rect 9321 22729 9355 22763
rect 10885 22729 10919 22763
rect 11437 22729 11471 22763
rect 2237 22661 2271 22695
rect 2513 22661 2547 22695
rect 5089 22661 5123 22695
rect 11805 22661 11839 22695
rect 2697 22593 2731 22627
rect 5641 22593 5675 22627
rect 5825 22593 5859 22627
rect 9505 22593 9539 22627
rect 13093 22593 13127 22627
rect 13829 22593 13863 22627
rect 2964 22525 2998 22559
rect 5549 22525 5583 22559
rect 6837 22525 6871 22559
rect 7093 22525 7127 22559
rect 12265 22525 12299 22559
rect 12909 22525 12943 22559
rect 6193 22457 6227 22491
rect 9772 22457 9806 22491
rect 12817 22457 12851 22491
rect 13461 22457 13495 22491
rect 4721 22389 4755 22423
rect 5181 22389 5215 22423
rect 6561 22389 6595 22423
rect 12449 22389 12483 22423
rect 1685 22185 1719 22219
rect 2789 22185 2823 22219
rect 3249 22185 3283 22219
rect 4813 22185 4847 22219
rect 6377 22185 6411 22219
rect 7573 22185 7607 22219
rect 10057 22185 10091 22219
rect 11253 22185 11287 22219
rect 12817 22185 12851 22219
rect 5264 22117 5298 22151
rect 11713 22117 11747 22151
rect 2421 22049 2455 22083
rect 4997 22049 5031 22083
rect 7941 22049 7975 22083
rect 9137 22049 9171 22083
rect 11161 22049 11195 22083
rect 11621 22049 11655 22083
rect 7481 21981 7515 22015
rect 8033 21981 8067 22015
rect 8125 21981 8159 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 11897 21981 11931 22015
rect 9505 21913 9539 21947
rect 4445 21845 4479 21879
rect 7113 21845 7147 21879
rect 9689 21845 9723 21879
rect 10793 21845 10827 21879
rect 12541 21845 12575 21879
rect 1593 21641 1627 21675
rect 3157 21641 3191 21675
rect 4721 21641 4755 21675
rect 7389 21641 7423 21675
rect 9781 21641 9815 21675
rect 11345 21641 11379 21675
rect 12449 21641 12483 21675
rect 6653 21573 6687 21607
rect 8217 21573 8251 21607
rect 3709 21505 3743 21539
rect 5273 21505 5307 21539
rect 7757 21505 7791 21539
rect 8769 21505 8803 21539
rect 10701 21505 10735 21539
rect 13001 21505 13035 21539
rect 1409 21437 1443 21471
rect 3065 21437 3099 21471
rect 3525 21437 3559 21471
rect 10425 21437 10459 21471
rect 12173 21437 12207 21471
rect 12817 21437 12851 21471
rect 1961 21369 1995 21403
rect 4629 21369 4663 21403
rect 8677 21369 8711 21403
rect 9413 21369 9447 21403
rect 10517 21369 10551 21403
rect 12909 21369 12943 21403
rect 3617 21301 3651 21335
rect 5089 21301 5123 21335
rect 5181 21301 5215 21335
rect 5825 21301 5859 21335
rect 8033 21301 8067 21335
rect 8585 21301 8619 21335
rect 10057 21301 10091 21335
rect 11805 21301 11839 21335
rect 5181 21097 5215 21131
rect 9505 21097 9539 21131
rect 10609 21097 10643 21131
rect 11069 21097 11103 21131
rect 12173 21097 12207 21131
rect 6929 21029 6963 21063
rect 11437 21029 11471 21063
rect 7481 20961 7515 20995
rect 10057 20961 10091 20995
rect 11529 20961 11563 20995
rect 7573 20893 7607 20927
rect 7757 20893 7791 20927
rect 11621 20893 11655 20927
rect 6561 20825 6595 20859
rect 3249 20757 3283 20791
rect 3801 20757 3835 20791
rect 4813 20757 4847 20791
rect 7113 20757 7147 20791
rect 8309 20757 8343 20791
rect 9137 20757 9171 20791
rect 12541 20757 12575 20791
rect 6837 20553 6871 20587
rect 9045 20553 9079 20587
rect 6285 20485 6319 20519
rect 10609 20485 10643 20519
rect 4261 20417 4295 20451
rect 7297 20417 7331 20451
rect 7481 20417 7515 20451
rect 8953 20417 8987 20451
rect 9597 20417 9631 20451
rect 11161 20417 11195 20451
rect 11989 20417 12023 20451
rect 3617 20349 3651 20383
rect 7205 20349 7239 20383
rect 8217 20349 8251 20383
rect 9413 20349 9447 20383
rect 10977 20349 11011 20383
rect 5733 20281 5767 20315
rect 10149 20281 10183 20315
rect 11069 20281 11103 20315
rect 3709 20213 3743 20247
rect 4077 20213 4111 20247
rect 4169 20213 4203 20247
rect 6561 20213 6595 20247
rect 7849 20213 7883 20247
rect 9505 20213 9539 20247
rect 10425 20213 10459 20247
rect 11621 20213 11655 20247
rect 3801 20009 3835 20043
rect 4537 20009 4571 20043
rect 4905 20009 4939 20043
rect 7757 20009 7791 20043
rect 9137 20009 9171 20043
rect 9965 20009 9999 20043
rect 11161 20009 11195 20043
rect 12909 20009 12943 20043
rect 6644 19941 6678 19975
rect 6377 19873 6411 19907
rect 10333 19873 10367 19907
rect 11796 19873 11830 19907
rect 4997 19805 5031 19839
rect 5089 19805 5123 19839
rect 10425 19805 10459 19839
rect 10517 19805 10551 19839
rect 11529 19805 11563 19839
rect 6101 19465 6135 19499
rect 7205 19465 7239 19499
rect 10517 19465 10551 19499
rect 11069 19465 11103 19499
rect 11897 19465 11931 19499
rect 7849 19329 7883 19363
rect 11529 19329 11563 19363
rect 2789 19261 2823 19295
rect 2881 19261 2915 19295
rect 7573 19261 7607 19295
rect 9045 19261 9079 19295
rect 9137 19261 9171 19295
rect 3126 19193 3160 19227
rect 5181 19193 5215 19227
rect 6469 19193 6503 19227
rect 9382 19193 9416 19227
rect 4261 19125 4295 19159
rect 4905 19125 4939 19159
rect 5365 19125 5399 19159
rect 7113 19125 7147 19159
rect 7665 19125 7699 19159
rect 8309 19125 8343 19159
rect 7205 18921 7239 18955
rect 7665 18921 7699 18955
rect 4905 18785 4939 18819
rect 5172 18785 5206 18819
rect 8401 18785 8435 18819
rect 8493 18717 8527 18751
rect 8585 18717 8619 18751
rect 10333 18717 10367 18751
rect 2973 18581 3007 18615
rect 4537 18581 4571 18615
rect 6285 18581 6319 18615
rect 8033 18581 8067 18615
rect 9229 18581 9263 18615
rect 10057 18581 10091 18615
rect 1593 18377 1627 18411
rect 4813 18377 4847 18411
rect 4353 18309 4387 18343
rect 5365 18241 5399 18275
rect 6193 18241 6227 18275
rect 1409 18173 1443 18207
rect 3985 18173 4019 18207
rect 5181 18173 5215 18207
rect 7941 18173 7975 18207
rect 8033 18173 8067 18207
rect 7205 18105 7239 18139
rect 7573 18105 7607 18139
rect 8300 18105 8334 18139
rect 1961 18037 1995 18071
rect 4721 18037 4755 18071
rect 5273 18037 5307 18071
rect 5825 18037 5859 18071
rect 9413 18037 9447 18071
rect 5273 17833 5307 17867
rect 7757 17833 7791 17867
rect 8217 17833 8251 17867
rect 8125 17697 8159 17731
rect 10057 17697 10091 17731
rect 11621 17697 11655 17731
rect 11888 17697 11922 17731
rect 5365 17629 5399 17663
rect 5549 17629 5583 17663
rect 8309 17629 8343 17663
rect 10149 17629 10183 17663
rect 10241 17629 10275 17663
rect 4905 17561 4939 17595
rect 7665 17561 7699 17595
rect 9689 17561 9723 17595
rect 3065 17493 3099 17527
rect 6929 17493 6963 17527
rect 7297 17493 7331 17527
rect 8769 17493 8803 17527
rect 10701 17493 10735 17527
rect 13001 17493 13035 17527
rect 4077 17289 4111 17323
rect 4353 17289 4387 17323
rect 7941 17289 7975 17323
rect 8585 17289 8619 17323
rect 10149 17289 10183 17323
rect 11621 17289 11655 17323
rect 2973 17221 3007 17255
rect 10057 17221 10091 17255
rect 3433 17153 3467 17187
rect 3525 17153 3559 17187
rect 5549 17153 5583 17187
rect 7297 17153 7331 17187
rect 7481 17153 7515 17187
rect 9137 17153 9171 17187
rect 10701 17153 10735 17187
rect 2881 17085 2915 17119
rect 4813 17085 4847 17119
rect 5365 17085 5399 17119
rect 5917 17085 5951 17119
rect 6653 17085 6687 17119
rect 10609 17085 10643 17119
rect 2513 17017 2547 17051
rect 3341 17017 3375 17051
rect 5273 17017 5307 17051
rect 10517 17017 10551 17051
rect 11161 17017 11195 17051
rect 4905 16949 4939 16983
rect 6837 16949 6871 16983
rect 7205 16949 7239 16983
rect 8493 16949 8527 16983
rect 8953 16949 8987 16983
rect 9045 16949 9079 16983
rect 9689 16949 9723 16983
rect 12081 16949 12115 16983
rect 2421 16745 2455 16779
rect 2789 16745 2823 16779
rect 4077 16745 4111 16779
rect 4537 16745 4571 16779
rect 5089 16745 5123 16779
rect 7665 16745 7699 16779
rect 8217 16745 8251 16779
rect 9505 16745 9539 16779
rect 11621 16745 11655 16779
rect 2881 16677 2915 16711
rect 4445 16609 4479 16643
rect 5457 16609 5491 16643
rect 6541 16609 6575 16643
rect 8585 16609 8619 16643
rect 9873 16609 9907 16643
rect 10241 16609 10275 16643
rect 10508 16609 10542 16643
rect 3065 16541 3099 16575
rect 4629 16541 4663 16575
rect 6285 16541 6319 16575
rect 1593 16201 1627 16235
rect 2053 16201 2087 16235
rect 4261 16201 4295 16235
rect 6837 16201 6871 16235
rect 9229 16201 9263 16235
rect 10701 16201 10735 16235
rect 11345 16201 11379 16235
rect 6653 16065 6687 16099
rect 7297 16065 7331 16099
rect 7481 16065 7515 16099
rect 9321 16065 9355 16099
rect 1409 15997 1443 16031
rect 2789 15997 2823 16031
rect 2881 15997 2915 16031
rect 5917 15997 5951 16031
rect 6285 15997 6319 16031
rect 7205 15997 7239 16031
rect 2421 15929 2455 15963
rect 3126 15929 3160 15963
rect 4813 15929 4847 15963
rect 9566 15929 9600 15963
rect 7941 15861 7975 15895
rect 1593 15657 1627 15691
rect 2513 15657 2547 15691
rect 2973 15657 3007 15691
rect 4629 15657 4663 15691
rect 6929 15657 6963 15691
rect 7389 15657 7423 15691
rect 9413 15657 9447 15691
rect 9873 15657 9907 15691
rect 10885 15657 10919 15691
rect 12541 15657 12575 15691
rect 4353 15589 4387 15623
rect 11897 15589 11931 15623
rect 5161 15521 5195 15555
rect 7757 15521 7791 15555
rect 10241 15521 10275 15555
rect 11805 15521 11839 15555
rect 4905 15453 4939 15487
rect 7849 15453 7883 15487
rect 7941 15453 7975 15487
rect 10333 15453 10367 15487
rect 10517 15453 10551 15487
rect 11989 15453 12023 15487
rect 7205 15385 7239 15419
rect 11437 15385 11471 15419
rect 6285 15317 6319 15351
rect 1961 15113 1995 15147
rect 4077 15113 4111 15147
rect 5181 15113 5215 15147
rect 5549 15113 5583 15147
rect 10333 15113 10367 15147
rect 10885 15113 10919 15147
rect 9965 15045 9999 15079
rect 3617 14977 3651 15011
rect 4629 14977 4663 15011
rect 13001 14977 13035 15011
rect 1409 14909 1443 14943
rect 3985 14909 4019 14943
rect 4445 14909 4479 14943
rect 7849 14909 7883 14943
rect 12909 14909 12943 14943
rect 8116 14841 8150 14875
rect 12265 14841 12299 14875
rect 12817 14841 12851 14875
rect 1593 14773 1627 14807
rect 4537 14773 4571 14807
rect 6561 14773 6595 14807
rect 7113 14773 7147 14807
rect 7481 14773 7515 14807
rect 9229 14773 9263 14807
rect 11161 14773 11195 14807
rect 11345 14773 11379 14807
rect 11897 14773 11931 14807
rect 12449 14773 12483 14807
rect 4353 14569 4387 14603
rect 4721 14569 4755 14603
rect 5181 14569 5215 14603
rect 8033 14569 8067 14603
rect 9505 14569 9539 14603
rect 10241 14569 10275 14603
rect 11529 14569 11563 14603
rect 7481 14501 7515 14535
rect 5089 14433 5123 14467
rect 7389 14433 7423 14467
rect 10609 14433 10643 14467
rect 11805 14433 11839 14467
rect 12061 14433 12095 14467
rect 5365 14365 5399 14399
rect 7573 14365 7607 14399
rect 10149 14365 10183 14399
rect 10701 14365 10735 14399
rect 10793 14365 10827 14399
rect 6561 14297 6595 14331
rect 7021 14297 7055 14331
rect 6929 14229 6963 14263
rect 8401 14229 8435 14263
rect 8861 14229 8895 14263
rect 13185 14229 13219 14263
rect 4813 14025 4847 14059
rect 6193 14025 6227 14059
rect 6653 14025 6687 14059
rect 7849 14025 7883 14059
rect 8401 14025 8435 14059
rect 10241 14025 10275 14059
rect 10425 14025 10459 14059
rect 11805 14025 11839 14059
rect 12173 14025 12207 14059
rect 12449 14025 12483 14059
rect 8309 13957 8343 13991
rect 9597 13957 9631 13991
rect 5089 13889 5123 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 8861 13889 8895 13923
rect 8953 13889 8987 13923
rect 9965 13889 9999 13923
rect 10977 13889 11011 13923
rect 11437 13889 11471 13923
rect 13093 13889 13127 13923
rect 13461 13889 13495 13923
rect 5457 13821 5491 13855
rect 10793 13821 10827 13855
rect 12909 13821 12943 13855
rect 7205 13753 7239 13787
rect 6837 13685 6871 13719
rect 8769 13685 8803 13719
rect 10885 13685 10919 13719
rect 12817 13685 12851 13719
rect 1593 13481 1627 13515
rect 6285 13481 6319 13515
rect 8033 13481 8067 13515
rect 8493 13481 8527 13515
rect 9965 13481 9999 13515
rect 11621 13481 11655 13515
rect 11989 13481 12023 13515
rect 12633 13481 12667 13515
rect 6377 13413 6411 13447
rect 7941 13413 7975 13447
rect 1409 13345 1443 13379
rect 8401 13345 8435 13379
rect 10425 13345 10459 13379
rect 12081 13345 12115 13379
rect 6469 13277 6503 13311
rect 8585 13277 8619 13311
rect 10517 13277 10551 13311
rect 10701 13277 10735 13311
rect 12173 13277 12207 13311
rect 10057 13209 10091 13243
rect 11069 13209 11103 13243
rect 2697 13141 2731 13175
rect 5917 13141 5951 13175
rect 7021 13141 7055 13175
rect 7481 13141 7515 13175
rect 9137 13141 9171 13175
rect 6009 12937 6043 12971
rect 7389 12937 7423 12971
rect 8769 12937 8803 12971
rect 10333 12937 10367 12971
rect 11253 12937 11287 12971
rect 11713 12937 11747 12971
rect 12633 12937 12667 12971
rect 5641 12869 5675 12903
rect 11989 12869 12023 12903
rect 6653 12801 6687 12835
rect 7941 12801 7975 12835
rect 8493 12801 8527 12835
rect 2605 12733 2639 12767
rect 2861 12733 2895 12767
rect 7757 12733 7791 12767
rect 8953 12733 8987 12767
rect 1685 12665 1719 12699
rect 7297 12665 7331 12699
rect 7849 12665 7883 12699
rect 9220 12665 9254 12699
rect 2513 12597 2547 12631
rect 3985 12597 4019 12631
rect 10885 12597 10919 12631
rect 5457 12393 5491 12427
rect 6101 12393 6135 12427
rect 6561 12393 6595 12427
rect 7573 12393 7607 12427
rect 8125 12393 8159 12427
rect 8585 12393 8619 12427
rect 10057 12393 10091 12427
rect 11713 12393 11747 12427
rect 4344 12257 4378 12291
rect 6929 12257 6963 12291
rect 10600 12257 10634 12291
rect 4077 12189 4111 12223
rect 7021 12189 7055 12223
rect 7205 12189 7239 12223
rect 10333 12189 10367 12223
rect 2605 12053 2639 12087
rect 6377 12053 6411 12087
rect 9045 12053 9079 12087
rect 2421 11849 2455 11883
rect 3893 11849 3927 11883
rect 4537 11849 4571 11883
rect 6653 11849 6687 11883
rect 8769 11849 8803 11883
rect 10333 11849 10367 11883
rect 10701 11849 10735 11883
rect 2513 11713 2547 11747
rect 5641 11713 5675 11747
rect 6009 11713 6043 11747
rect 2780 11645 2814 11679
rect 7389 11645 7423 11679
rect 7656 11645 7690 11679
rect 4905 11577 4939 11611
rect 5457 11577 5491 11611
rect 4997 11509 5031 11543
rect 5365 11509 5399 11543
rect 7205 11509 7239 11543
rect 4169 11305 4203 11339
rect 5089 11305 5123 11339
rect 5181 11305 5215 11339
rect 6653 11305 6687 11339
rect 8125 11305 8159 11339
rect 2789 11237 2823 11271
rect 4629 11237 4663 11271
rect 7012 11237 7046 11271
rect 5549 11169 5583 11203
rect 2881 11101 2915 11135
rect 3065 11101 3099 11135
rect 5641 11101 5675 11135
rect 5733 11101 5767 11135
rect 6745 11101 6779 11135
rect 2421 10965 2455 10999
rect 2513 10761 2547 10795
rect 2789 10761 2823 10795
rect 2973 10761 3007 10795
rect 2145 10693 2179 10727
rect 4537 10693 4571 10727
rect 6837 10693 6871 10727
rect 3617 10625 3651 10659
rect 5181 10625 5215 10659
rect 5917 10625 5951 10659
rect 7481 10625 7515 10659
rect 7849 10625 7883 10659
rect 3341 10557 3375 10591
rect 3433 10557 3467 10591
rect 4997 10489 5031 10523
rect 6653 10489 6687 10523
rect 7205 10489 7239 10523
rect 1777 10421 1811 10455
rect 3985 10421 4019 10455
rect 4445 10421 4479 10455
rect 4905 10421 4939 10455
rect 6285 10421 6319 10455
rect 7297 10421 7331 10455
rect 8401 10421 8435 10455
rect 12449 10421 12483 10455
rect 1593 10217 1627 10251
rect 2421 10217 2455 10251
rect 3433 10217 3467 10251
rect 5273 10217 5307 10251
rect 5917 10217 5951 10251
rect 6561 10217 6595 10251
rect 6929 10217 6963 10251
rect 13369 10217 13403 10251
rect 2329 10149 2363 10183
rect 4905 10149 4939 10183
rect 5641 10149 5675 10183
rect 7573 10149 7607 10183
rect 10762 10149 10796 10183
rect 1409 10081 1443 10115
rect 2789 10081 2823 10115
rect 7021 10081 7055 10115
rect 10517 10081 10551 10115
rect 13461 10081 13495 10115
rect 2881 10013 2915 10047
rect 3065 10013 3099 10047
rect 7205 10013 7239 10047
rect 13553 10013 13587 10047
rect 4537 9877 4571 9911
rect 9321 9877 9355 9911
rect 10425 9877 10459 9911
rect 11897 9877 11931 9911
rect 12449 9877 12483 9911
rect 12909 9877 12943 9911
rect 13001 9877 13035 9911
rect 2881 9673 2915 9707
rect 7113 9673 7147 9707
rect 7481 9673 7515 9707
rect 10517 9673 10551 9707
rect 4445 9605 4479 9639
rect 12265 9605 12299 9639
rect 12449 9605 12483 9639
rect 13461 9605 13495 9639
rect 13829 9605 13863 9639
rect 2421 9537 2455 9571
rect 3525 9537 3559 9571
rect 3985 9537 4019 9571
rect 5089 9537 5123 9571
rect 9689 9537 9723 9571
rect 9873 9537 9907 9571
rect 11345 9537 11379 9571
rect 13001 9537 13035 9571
rect 1685 9469 1719 9503
rect 2789 9469 2823 9503
rect 3249 9469 3283 9503
rect 6561 9469 6595 9503
rect 9137 9469 9171 9503
rect 11161 9469 11195 9503
rect 12817 9469 12851 9503
rect 2053 9401 2087 9435
rect 4905 9401 4939 9435
rect 9597 9401 9631 9435
rect 11253 9401 11287 9435
rect 3341 9333 3375 9367
rect 4353 9333 4387 9367
rect 4813 9333 4847 9367
rect 8677 9333 8711 9367
rect 9229 9333 9263 9367
rect 10793 9333 10827 9367
rect 11897 9333 11931 9367
rect 12909 9333 12943 9367
rect 1593 9129 1627 9163
rect 2513 9129 2547 9163
rect 2973 9129 3007 9163
rect 5457 9129 5491 9163
rect 8401 9129 8435 9163
rect 9689 9129 9723 9163
rect 10149 9129 10183 9163
rect 3433 9061 3467 9095
rect 4322 9061 4356 9095
rect 11980 9061 12014 9095
rect 10057 8993 10091 9027
rect 11713 8993 11747 9027
rect 4077 8925 4111 8959
rect 8493 8925 8527 8959
rect 8585 8925 8619 8959
rect 10333 8925 10367 8959
rect 9045 8857 9079 8891
rect 11529 8857 11563 8891
rect 7389 8789 7423 8823
rect 7849 8789 7883 8823
rect 8033 8789 8067 8823
rect 10885 8789 10919 8823
rect 11253 8789 11287 8823
rect 13093 8789 13127 8823
rect 3341 8585 3375 8619
rect 7297 8585 7331 8619
rect 8769 8585 8803 8619
rect 10241 8585 10275 8619
rect 11437 8585 11471 8619
rect 12449 8585 12483 8619
rect 10793 8517 10827 8551
rect 11713 8517 11747 8551
rect 3249 8449 3283 8483
rect 3801 8449 3835 8483
rect 3985 8449 4019 8483
rect 7849 8449 7883 8483
rect 8401 8449 8435 8483
rect 13001 8449 13035 8483
rect 6561 8381 6595 8415
rect 8861 8381 8895 8415
rect 12265 8381 12299 8415
rect 6285 8313 6319 8347
rect 7205 8313 7239 8347
rect 7665 8313 7699 8347
rect 7757 8313 7791 8347
rect 9106 8313 9140 8347
rect 12817 8313 12851 8347
rect 3709 8245 3743 8279
rect 4445 8245 4479 8279
rect 4721 8245 4755 8279
rect 12909 8245 12943 8279
rect 1869 8041 1903 8075
rect 3433 8041 3467 8075
rect 10149 8041 10183 8075
rect 10517 8041 10551 8075
rect 10701 8041 10735 8075
rect 11161 8041 11195 8075
rect 12541 8041 12575 8075
rect 8953 7973 8987 8007
rect 12817 7973 12851 8007
rect 4804 7905 4838 7939
rect 7288 7905 7322 7939
rect 11069 7905 11103 7939
rect 4537 7837 4571 7871
rect 7021 7837 7055 7871
rect 9689 7837 9723 7871
rect 11345 7837 11379 7871
rect 5917 7701 5951 7735
rect 6561 7701 6595 7735
rect 6929 7701 6963 7735
rect 8401 7701 8435 7735
rect 3157 7497 3191 7531
rect 8033 7497 8067 7531
rect 10333 7497 10367 7531
rect 11713 7497 11747 7531
rect 8585 7429 8619 7463
rect 11345 7429 11379 7463
rect 1777 7361 1811 7395
rect 4261 7361 4295 7395
rect 5641 7361 5675 7395
rect 7481 7361 7515 7395
rect 7665 7361 7699 7395
rect 9137 7361 9171 7395
rect 9597 7361 9631 7395
rect 10793 7361 10827 7395
rect 10885 7361 10919 7395
rect 7389 7293 7423 7327
rect 9045 7293 9079 7327
rect 2022 7225 2056 7259
rect 4905 7225 4939 7259
rect 5549 7225 5583 7259
rect 6285 7225 6319 7259
rect 1593 7157 1627 7191
rect 4537 7157 4571 7191
rect 5089 7157 5123 7191
rect 5457 7157 5491 7191
rect 6561 7157 6595 7191
rect 7021 7157 7055 7191
rect 8493 7157 8527 7191
rect 8953 7157 8987 7191
rect 10241 7157 10275 7191
rect 10701 7157 10735 7191
rect 5181 6953 5215 6987
rect 7389 6953 7423 6987
rect 7941 6953 7975 6987
rect 8309 6953 8343 6987
rect 8401 6953 8435 6987
rect 10793 6953 10827 6987
rect 11161 6953 11195 6987
rect 10425 6885 10459 6919
rect 1409 6817 1443 6851
rect 2421 6817 2455 6851
rect 2881 6817 2915 6851
rect 5724 6817 5758 6851
rect 7849 6817 7883 6851
rect 9689 6817 9723 6851
rect 12081 6817 12115 6851
rect 12348 6817 12382 6851
rect 5457 6749 5491 6783
rect 8493 6749 8527 6783
rect 2605 6681 2639 6715
rect 4629 6681 4663 6715
rect 1593 6613 1627 6647
rect 6837 6613 6871 6647
rect 8953 6613 8987 6647
rect 9873 6613 9907 6647
rect 13461 6613 13495 6647
rect 2053 6409 2087 6443
rect 5917 6409 5951 6443
rect 7113 6409 7147 6443
rect 7849 6409 7883 6443
rect 9321 6409 9355 6443
rect 12173 6409 12207 6443
rect 12633 6409 12667 6443
rect 5549 6341 5583 6375
rect 3709 6273 3743 6307
rect 4997 6273 5031 6307
rect 5181 6273 5215 6307
rect 8861 6273 8895 6307
rect 10425 6273 10459 6307
rect 10885 6273 10919 6307
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 4077 6205 4111 6239
rect 7205 6205 7239 6239
rect 9781 6205 9815 6239
rect 4445 6137 4479 6171
rect 4905 6137 4939 6171
rect 8217 6137 8251 6171
rect 10241 6137 10275 6171
rect 10333 6137 10367 6171
rect 1593 6069 1627 6103
rect 2421 6069 2455 6103
rect 2697 6069 2731 6103
rect 3065 6069 3099 6103
rect 4537 6069 4571 6103
rect 6653 6069 6687 6103
rect 7389 6069 7423 6103
rect 8309 6069 8343 6103
rect 8677 6069 8711 6103
rect 8769 6069 8803 6103
rect 9873 6069 9907 6103
rect 4353 5865 4387 5899
rect 7389 5865 7423 5899
rect 4813 5797 4847 5831
rect 6276 5797 6310 5831
rect 9873 5797 9907 5831
rect 12072 5797 12106 5831
rect 1409 5729 1443 5763
rect 2881 5729 2915 5763
rect 7941 5729 7975 5763
rect 8493 5729 8527 5763
rect 9505 5729 9539 5763
rect 10609 5729 10643 5763
rect 11345 5729 11379 5763
rect 4905 5661 4939 5695
rect 5089 5661 5123 5695
rect 6009 5661 6043 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 11805 5661 11839 5695
rect 8677 5593 8711 5627
rect 10241 5593 10275 5627
rect 1593 5525 1627 5559
rect 2513 5525 2547 5559
rect 3065 5525 3099 5559
rect 3433 5525 3467 5559
rect 3893 5525 3927 5559
rect 4445 5525 4479 5559
rect 5549 5525 5583 5559
rect 5917 5525 5951 5559
rect 8309 5525 8343 5559
rect 13185 5525 13219 5559
rect 1593 5321 1627 5355
rect 2881 5321 2915 5355
rect 4353 5321 4387 5355
rect 6561 5321 6595 5355
rect 7389 5321 7423 5355
rect 8033 5321 8067 5355
rect 9505 5321 9539 5355
rect 10793 5321 10827 5355
rect 11805 5321 11839 5355
rect 12265 5321 12299 5355
rect 10701 5253 10735 5287
rect 8125 5185 8159 5219
rect 11345 5185 11379 5219
rect 1777 5117 1811 5151
rect 2973 5117 3007 5151
rect 5641 5117 5675 5151
rect 6193 5117 6227 5151
rect 6837 5117 6871 5151
rect 10333 5117 10367 5151
rect 11161 5117 11195 5151
rect 2421 5049 2455 5083
rect 3218 5049 3252 5083
rect 8392 5049 8426 5083
rect 11253 5049 11287 5083
rect 1961 4981 1995 5015
rect 4905 4981 4939 5015
rect 5365 4981 5399 5015
rect 5825 4981 5859 5015
rect 7021 4981 7055 5015
rect 12449 4981 12483 5015
rect 2421 4777 2455 4811
rect 2881 4777 2915 4811
rect 4077 4777 4111 4811
rect 4537 4777 4571 4811
rect 5181 4777 5215 4811
rect 6561 4777 6595 4811
rect 7205 4777 7239 4811
rect 8401 4777 8435 4811
rect 9505 4777 9539 4811
rect 10609 4777 10643 4811
rect 12541 4777 12575 4811
rect 2329 4709 2363 4743
rect 4445 4709 4479 4743
rect 6009 4709 6043 4743
rect 6469 4709 6503 4743
rect 9137 4709 9171 4743
rect 10517 4709 10551 4743
rect 2789 4641 2823 4675
rect 8493 4641 8527 4675
rect 10977 4641 11011 4675
rect 1409 4573 1443 4607
rect 1961 4573 1995 4607
rect 2973 4573 3007 4607
rect 3893 4573 3927 4607
rect 4721 4573 4755 4607
rect 6653 4573 6687 4607
rect 8677 4573 8711 4607
rect 11069 4573 11103 4607
rect 11161 4573 11195 4607
rect 12633 4573 12667 4607
rect 12725 4573 12759 4607
rect 6101 4505 6135 4539
rect 7573 4505 7607 4539
rect 7941 4505 7975 4539
rect 3433 4437 3467 4471
rect 5549 4437 5583 4471
rect 8033 4437 8067 4471
rect 10149 4437 10183 4471
rect 12173 4437 12207 4471
rect 13185 4437 13219 4471
rect 2145 4233 2179 4267
rect 3985 4233 4019 4267
rect 4813 4233 4847 4267
rect 6193 4233 6227 4267
rect 6837 4233 6871 4267
rect 8033 4233 8067 4267
rect 11069 4233 11103 4267
rect 12265 4233 12299 4267
rect 13829 4233 13863 4267
rect 6561 4165 6595 4199
rect 5641 4097 5675 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 9137 4097 9171 4131
rect 9505 4097 9539 4131
rect 10701 4097 10735 4131
rect 13093 4097 13127 4131
rect 13461 4097 13495 4131
rect 1501 4029 1535 4063
rect 2513 4029 2547 4063
rect 2605 4029 2639 4063
rect 2872 4029 2906 4063
rect 5457 4029 5491 4063
rect 7205 4029 7239 4063
rect 8953 4029 8987 4063
rect 9965 4029 9999 4063
rect 10517 4029 10551 4063
rect 11437 4029 11471 4063
rect 12817 4029 12851 4063
rect 5549 3961 5583 3995
rect 1685 3893 1719 3927
rect 5089 3893 5123 3927
rect 8493 3893 8527 3927
rect 8861 3893 8895 3927
rect 10057 3893 10091 3927
rect 10425 3893 10459 3927
rect 11805 3893 11839 3927
rect 12449 3893 12483 3927
rect 12909 3893 12943 3927
rect 1685 3689 1719 3723
rect 3525 3689 3559 3723
rect 3893 3689 3927 3723
rect 4721 3689 4755 3723
rect 7665 3689 7699 3723
rect 8033 3689 8067 3723
rect 8769 3689 8803 3723
rect 9505 3689 9539 3723
rect 10333 3689 10367 3723
rect 10609 3689 10643 3723
rect 10977 3689 11011 3723
rect 2513 3621 2547 3655
rect 4629 3621 4663 3655
rect 5181 3621 5215 3655
rect 6193 3621 6227 3655
rect 8125 3621 8159 3655
rect 9137 3621 9171 3655
rect 1777 3553 1811 3587
rect 2881 3553 2915 3587
rect 5089 3553 5123 3587
rect 6285 3553 6319 3587
rect 6929 3553 6963 3587
rect 7297 3553 7331 3587
rect 9689 3553 9723 3587
rect 11161 3553 11195 3587
rect 11417 3553 11451 3587
rect 5273 3485 5307 3519
rect 5825 3485 5859 3519
rect 8217 3485 8251 3519
rect 3065 3417 3099 3451
rect 6469 3417 6503 3451
rect 12541 3417 12575 3451
rect 1961 3349 1995 3383
rect 9873 3349 9907 3383
rect 13093 3349 13127 3383
rect 1777 3145 1811 3179
rect 2973 3145 3007 3179
rect 5641 3145 5675 3179
rect 6377 3145 6411 3179
rect 7205 3145 7239 3179
rect 10149 3145 10183 3179
rect 10793 3145 10827 3179
rect 11437 3145 11471 3179
rect 12081 3145 12115 3179
rect 12173 3145 12207 3179
rect 12449 3145 12483 3179
rect 2237 3077 2271 3111
rect 4261 3009 4295 3043
rect 7665 3009 7699 3043
rect 7849 3009 7883 3043
rect 2053 2941 2087 2975
rect 2605 2941 2639 2975
rect 3157 2941 3191 2975
rect 3709 2941 3743 2975
rect 4528 2941 4562 2975
rect 7113 2941 7147 2975
rect 7573 2941 7607 2975
rect 8769 2941 8803 2975
rect 11161 2941 11195 2975
rect 11253 2941 11287 2975
rect 4169 2873 4203 2907
rect 8309 2873 8343 2907
rect 9014 2873 9048 2907
rect 11897 2873 11931 2907
rect 13093 3009 13127 3043
rect 13461 3009 13495 3043
rect 12909 2873 12943 2907
rect 3341 2805 3375 2839
rect 8677 2805 8711 2839
rect 12081 2805 12115 2839
rect 12817 2805 12851 2839
rect 1961 2601 1995 2635
rect 4261 2601 4295 2635
rect 4721 2601 4755 2635
rect 5273 2601 5307 2635
rect 7113 2601 7147 2635
rect 7481 2601 7515 2635
rect 8125 2601 8159 2635
rect 8493 2601 8527 2635
rect 11713 2601 11747 2635
rect 12449 2601 12483 2635
rect 12633 2601 12667 2635
rect 3525 2533 3559 2567
rect 9229 2533 9263 2567
rect 10026 2533 10060 2567
rect 13093 2533 13127 2567
rect 1777 2465 1811 2499
rect 2881 2465 2915 2499
rect 5181 2465 5215 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 8033 2465 8067 2499
rect 9597 2465 9631 2499
rect 9781 2465 9815 2499
rect 13001 2465 13035 2499
rect 13645 2465 13679 2499
rect 3893 2397 3927 2431
rect 5365 2397 5399 2431
rect 6193 2397 6227 2431
rect 6745 2397 6779 2431
rect 8585 2397 8619 2431
rect 8769 2397 8803 2431
rect 13277 2397 13311 2431
rect 14013 2397 14047 2431
rect 2421 2329 2455 2363
rect 4813 2329 4847 2363
rect 3065 2261 3099 2295
rect 11161 2261 11195 2295
<< metal1 >>
rect 1104 37562 14812 37584
rect 1104 37510 6315 37562
rect 6367 37510 6379 37562
rect 6431 37510 6443 37562
rect 6495 37510 6507 37562
rect 6559 37510 11648 37562
rect 11700 37510 11712 37562
rect 11764 37510 11776 37562
rect 11828 37510 11840 37562
rect 11892 37510 14812 37562
rect 1104 37488 14812 37510
rect 1104 37018 14812 37040
rect 1104 36966 3648 37018
rect 3700 36966 3712 37018
rect 3764 36966 3776 37018
rect 3828 36966 3840 37018
rect 3892 36966 8982 37018
rect 9034 36966 9046 37018
rect 9098 36966 9110 37018
rect 9162 36966 9174 37018
rect 9226 36966 14315 37018
rect 14367 36966 14379 37018
rect 14431 36966 14443 37018
rect 14495 36966 14507 37018
rect 14559 36966 14812 37018
rect 1104 36944 14812 36966
rect 5629 36907 5687 36913
rect 5629 36873 5641 36907
rect 5675 36904 5687 36907
rect 6178 36904 6184 36916
rect 5675 36876 6184 36904
rect 5675 36873 5687 36876
rect 5629 36867 5687 36873
rect 6178 36864 6184 36876
rect 6236 36864 6242 36916
rect 5258 36660 5264 36712
rect 5316 36700 5322 36712
rect 5445 36703 5503 36709
rect 5445 36700 5457 36703
rect 5316 36672 5457 36700
rect 5316 36660 5322 36672
rect 5445 36669 5457 36672
rect 5491 36700 5503 36703
rect 5997 36703 6055 36709
rect 5997 36700 6009 36703
rect 5491 36672 6009 36700
rect 5491 36669 5503 36672
rect 5445 36663 5503 36669
rect 5997 36669 6009 36672
rect 6043 36669 6055 36703
rect 5997 36663 6055 36669
rect 1104 36474 14812 36496
rect 1104 36422 6315 36474
rect 6367 36422 6379 36474
rect 6431 36422 6443 36474
rect 6495 36422 6507 36474
rect 6559 36422 11648 36474
rect 11700 36422 11712 36474
rect 11764 36422 11776 36474
rect 11828 36422 11840 36474
rect 11892 36422 14812 36474
rect 1104 36400 14812 36422
rect 4893 36363 4951 36369
rect 4893 36329 4905 36363
rect 4939 36360 4951 36363
rect 5350 36360 5356 36372
rect 4939 36332 5356 36360
rect 4939 36329 4951 36332
rect 4893 36323 4951 36329
rect 5350 36320 5356 36332
rect 5408 36320 5414 36372
rect 5997 36363 6055 36369
rect 5997 36329 6009 36363
rect 6043 36360 6055 36363
rect 6638 36360 6644 36372
rect 6043 36332 6644 36360
rect 6043 36329 6055 36332
rect 5997 36323 6055 36329
rect 6638 36320 6644 36332
rect 6696 36320 6702 36372
rect 4706 36224 4712 36236
rect 4667 36196 4712 36224
rect 4706 36184 4712 36196
rect 4764 36184 4770 36236
rect 5813 36227 5871 36233
rect 5813 36193 5825 36227
rect 5859 36224 5871 36227
rect 5994 36224 6000 36236
rect 5859 36196 6000 36224
rect 5859 36193 5871 36196
rect 5813 36187 5871 36193
rect 5994 36184 6000 36196
rect 6052 36184 6058 36236
rect 1104 35930 14812 35952
rect 1104 35878 3648 35930
rect 3700 35878 3712 35930
rect 3764 35878 3776 35930
rect 3828 35878 3840 35930
rect 3892 35878 8982 35930
rect 9034 35878 9046 35930
rect 9098 35878 9110 35930
rect 9162 35878 9174 35930
rect 9226 35878 14315 35930
rect 14367 35878 14379 35930
rect 14431 35878 14443 35930
rect 14495 35878 14507 35930
rect 14559 35878 14812 35930
rect 1104 35856 14812 35878
rect 2961 35819 3019 35825
rect 2961 35785 2973 35819
rect 3007 35816 3019 35819
rect 3326 35816 3332 35828
rect 3007 35788 3332 35816
rect 3007 35785 3019 35788
rect 2961 35779 3019 35785
rect 3326 35776 3332 35788
rect 3384 35776 3390 35828
rect 3418 35776 3424 35828
rect 3476 35816 3482 35828
rect 4065 35819 4123 35825
rect 4065 35816 4077 35819
rect 3476 35788 4077 35816
rect 3476 35776 3482 35788
rect 4065 35785 4077 35788
rect 4111 35785 4123 35819
rect 4065 35779 4123 35785
rect 4246 35776 4252 35828
rect 4304 35816 4310 35828
rect 5169 35819 5227 35825
rect 5169 35816 5181 35819
rect 4304 35788 5181 35816
rect 4304 35776 4310 35788
rect 5169 35785 5181 35788
rect 5215 35785 5227 35819
rect 5169 35779 5227 35785
rect 7374 35776 7380 35828
rect 7432 35816 7438 35828
rect 7469 35819 7527 35825
rect 7469 35816 7481 35819
rect 7432 35788 7481 35816
rect 7432 35776 7438 35788
rect 7469 35785 7481 35788
rect 7515 35785 7527 35819
rect 7469 35779 7527 35785
rect 9858 35748 9864 35760
rect 9819 35720 9864 35748
rect 9858 35708 9864 35720
rect 9916 35708 9922 35760
rect 4706 35640 4712 35692
rect 4764 35680 4770 35692
rect 4801 35683 4859 35689
rect 4801 35680 4813 35683
rect 4764 35652 4813 35680
rect 4764 35640 4770 35652
rect 4801 35649 4813 35652
rect 4847 35680 4859 35683
rect 5810 35680 5816 35692
rect 4847 35652 5816 35680
rect 4847 35649 4859 35652
rect 4801 35643 4859 35649
rect 5810 35640 5816 35652
rect 5868 35640 5874 35692
rect 2777 35615 2835 35621
rect 2777 35581 2789 35615
rect 2823 35612 2835 35615
rect 3789 35615 3847 35621
rect 2823 35584 3464 35612
rect 2823 35581 2835 35584
rect 2777 35575 2835 35581
rect 3436 35485 3464 35584
rect 3789 35581 3801 35615
rect 3835 35612 3847 35615
rect 3881 35615 3939 35621
rect 3881 35612 3893 35615
rect 3835 35584 3893 35612
rect 3835 35581 3847 35584
rect 3789 35575 3847 35581
rect 3881 35581 3893 35584
rect 3927 35612 3939 35615
rect 4062 35612 4068 35624
rect 3927 35584 4068 35612
rect 3927 35581 3939 35584
rect 3881 35575 3939 35581
rect 4062 35572 4068 35584
rect 4120 35572 4126 35624
rect 4985 35615 5043 35621
rect 4985 35581 4997 35615
rect 5031 35612 5043 35615
rect 7285 35615 7343 35621
rect 5031 35584 5672 35612
rect 5031 35581 5043 35584
rect 4985 35575 5043 35581
rect 5644 35488 5672 35584
rect 7285 35581 7297 35615
rect 7331 35612 7343 35615
rect 9677 35615 9735 35621
rect 7331 35584 7972 35612
rect 7331 35581 7343 35584
rect 7285 35575 7343 35581
rect 3421 35479 3479 35485
rect 3421 35445 3433 35479
rect 3467 35476 3479 35479
rect 3510 35476 3516 35488
rect 3467 35448 3516 35476
rect 3467 35445 3479 35448
rect 3421 35439 3479 35445
rect 3510 35436 3516 35448
rect 3568 35436 3574 35488
rect 5626 35476 5632 35488
rect 5587 35448 5632 35476
rect 5626 35436 5632 35448
rect 5684 35436 5690 35488
rect 5994 35476 6000 35488
rect 5955 35448 6000 35476
rect 5994 35436 6000 35448
rect 6052 35436 6058 35488
rect 7944 35485 7972 35584
rect 9677 35581 9689 35615
rect 9723 35612 9735 35615
rect 9723 35584 10364 35612
rect 9723 35581 9735 35584
rect 9677 35575 9735 35581
rect 7929 35479 7987 35485
rect 7929 35445 7941 35479
rect 7975 35476 7987 35479
rect 9582 35476 9588 35488
rect 7975 35448 9588 35476
rect 7975 35445 7987 35448
rect 7929 35439 7987 35445
rect 9582 35436 9588 35448
rect 9640 35436 9646 35488
rect 10336 35485 10364 35584
rect 10321 35479 10379 35485
rect 10321 35445 10333 35479
rect 10367 35476 10379 35479
rect 10686 35476 10692 35488
rect 10367 35448 10692 35476
rect 10367 35445 10379 35448
rect 10321 35439 10379 35445
rect 10686 35436 10692 35448
rect 10744 35436 10750 35488
rect 1104 35386 14812 35408
rect 1104 35334 6315 35386
rect 6367 35334 6379 35386
rect 6431 35334 6443 35386
rect 6495 35334 6507 35386
rect 6559 35334 11648 35386
rect 11700 35334 11712 35386
rect 11764 35334 11776 35386
rect 11828 35334 11840 35386
rect 11892 35334 14812 35386
rect 1104 35312 14812 35334
rect 934 35232 940 35284
rect 992 35272 998 35284
rect 1581 35275 1639 35281
rect 1581 35272 1593 35275
rect 992 35244 1593 35272
rect 992 35232 998 35244
rect 1581 35241 1593 35244
rect 1627 35241 1639 35275
rect 1581 35235 1639 35241
rect 2130 35232 2136 35284
rect 2188 35272 2194 35284
rect 2685 35275 2743 35281
rect 2685 35272 2697 35275
rect 2188 35244 2697 35272
rect 2188 35232 2194 35244
rect 2685 35241 2697 35244
rect 2731 35241 2743 35275
rect 5074 35272 5080 35284
rect 5035 35244 5080 35272
rect 2685 35235 2743 35241
rect 5074 35232 5080 35244
rect 5132 35232 5138 35284
rect 5718 35232 5724 35284
rect 5776 35272 5782 35284
rect 6457 35275 6515 35281
rect 6457 35272 6469 35275
rect 5776 35244 6469 35272
rect 5776 35232 5782 35244
rect 6457 35241 6469 35244
rect 6503 35241 6515 35275
rect 7558 35272 7564 35284
rect 7519 35244 7564 35272
rect 6457 35235 6515 35241
rect 7558 35232 7564 35244
rect 7616 35232 7622 35284
rect 1397 35139 1455 35145
rect 1397 35105 1409 35139
rect 1443 35136 1455 35139
rect 1670 35136 1676 35148
rect 1443 35108 1676 35136
rect 1443 35105 1455 35108
rect 1397 35099 1455 35105
rect 1670 35096 1676 35108
rect 1728 35096 1734 35148
rect 2501 35139 2559 35145
rect 2501 35105 2513 35139
rect 2547 35136 2559 35139
rect 3418 35136 3424 35148
rect 2547 35108 3424 35136
rect 2547 35105 2559 35108
rect 2501 35099 2559 35105
rect 3418 35096 3424 35108
rect 3476 35096 3482 35148
rect 4890 35136 4896 35148
rect 4851 35108 4896 35136
rect 4890 35096 4896 35108
rect 4948 35096 4954 35148
rect 6270 35136 6276 35148
rect 6231 35108 6276 35136
rect 6270 35096 6276 35108
rect 6328 35096 6334 35148
rect 7377 35139 7435 35145
rect 7377 35105 7389 35139
rect 7423 35136 7435 35139
rect 7650 35136 7656 35148
rect 7423 35108 7656 35136
rect 7423 35105 7435 35108
rect 7377 35099 7435 35105
rect 7650 35096 7656 35108
rect 7708 35096 7714 35148
rect 8481 35139 8539 35145
rect 8481 35105 8493 35139
rect 8527 35136 8539 35139
rect 8754 35136 8760 35148
rect 8527 35108 8760 35136
rect 8527 35105 8539 35108
rect 8481 35099 8539 35105
rect 8754 35096 8760 35108
rect 8812 35096 8818 35148
rect 9490 35096 9496 35148
rect 9548 35136 9554 35148
rect 9933 35139 9991 35145
rect 9933 35136 9945 35139
rect 9548 35108 9945 35136
rect 9548 35096 9554 35108
rect 9933 35105 9945 35108
rect 9979 35105 9991 35139
rect 9933 35099 9991 35105
rect 9674 35028 9680 35080
rect 9732 35068 9738 35080
rect 12342 35068 12348 35080
rect 9732 35040 9777 35068
rect 12303 35040 12348 35068
rect 9732 35028 9738 35040
rect 12342 35028 12348 35040
rect 12400 35028 12406 35080
rect 6914 34960 6920 35012
rect 6972 35000 6978 35012
rect 8665 35003 8723 35009
rect 8665 35000 8677 35003
rect 6972 34972 8677 35000
rect 6972 34960 6978 34972
rect 8665 34969 8677 34972
rect 8711 34969 8723 35003
rect 8665 34963 8723 34969
rect 7926 34932 7932 34944
rect 7887 34904 7932 34932
rect 7926 34892 7932 34904
rect 7984 34892 7990 34944
rect 9493 34935 9551 34941
rect 9493 34901 9505 34935
rect 9539 34932 9551 34935
rect 10778 34932 10784 34944
rect 9539 34904 10784 34932
rect 9539 34901 9551 34904
rect 9493 34895 9551 34901
rect 10778 34892 10784 34904
rect 10836 34932 10842 34944
rect 11057 34935 11115 34941
rect 11057 34932 11069 34935
rect 10836 34904 11069 34932
rect 10836 34892 10842 34904
rect 11057 34901 11069 34904
rect 11103 34901 11115 34935
rect 12894 34932 12900 34944
rect 12855 34904 12900 34932
rect 11057 34895 11115 34901
rect 12894 34892 12900 34904
rect 12952 34892 12958 34944
rect 1104 34842 14812 34864
rect 1104 34790 3648 34842
rect 3700 34790 3712 34842
rect 3764 34790 3776 34842
rect 3828 34790 3840 34842
rect 3892 34790 8982 34842
rect 9034 34790 9046 34842
rect 9098 34790 9110 34842
rect 9162 34790 9174 34842
rect 9226 34790 14315 34842
rect 14367 34790 14379 34842
rect 14431 34790 14443 34842
rect 14495 34790 14507 34842
rect 14559 34790 14812 34842
rect 1104 34768 14812 34790
rect 198 34688 204 34740
rect 256 34728 262 34740
rect 1581 34731 1639 34737
rect 1581 34728 1593 34731
rect 256 34700 1593 34728
rect 256 34688 262 34700
rect 1581 34697 1593 34700
rect 1627 34697 1639 34731
rect 2682 34728 2688 34740
rect 2643 34700 2688 34728
rect 1581 34691 1639 34697
rect 2682 34688 2688 34700
rect 2740 34688 2746 34740
rect 7285 34731 7343 34737
rect 7285 34697 7297 34731
rect 7331 34728 7343 34731
rect 7650 34728 7656 34740
rect 7331 34700 7656 34728
rect 7331 34697 7343 34700
rect 7285 34691 7343 34697
rect 7650 34688 7656 34700
rect 7708 34688 7714 34740
rect 9674 34688 9680 34740
rect 9732 34728 9738 34740
rect 11885 34731 11943 34737
rect 9732 34700 9777 34728
rect 9732 34688 9738 34700
rect 11885 34697 11897 34731
rect 11931 34728 11943 34731
rect 12342 34728 12348 34740
rect 11931 34700 12348 34728
rect 11931 34697 11943 34700
rect 11885 34691 11943 34697
rect 12342 34688 12348 34700
rect 12400 34688 12406 34740
rect 3329 34595 3387 34601
rect 3329 34561 3341 34595
rect 3375 34592 3387 34595
rect 9692 34592 9720 34688
rect 12253 34663 12311 34669
rect 12253 34629 12265 34663
rect 12299 34660 12311 34663
rect 12299 34632 13124 34660
rect 12299 34629 12311 34632
rect 12253 34623 12311 34629
rect 9858 34592 9864 34604
rect 3375 34564 3556 34592
rect 9692 34564 9864 34592
rect 3375 34561 3387 34564
rect 3329 34555 3387 34561
rect 1397 34527 1455 34533
rect 1397 34493 1409 34527
rect 1443 34524 1455 34527
rect 1949 34527 2007 34533
rect 1949 34524 1961 34527
rect 1443 34496 1961 34524
rect 1443 34493 1455 34496
rect 1397 34487 1455 34493
rect 1949 34493 1961 34496
rect 1995 34524 2007 34527
rect 2222 34524 2228 34536
rect 1995 34496 2228 34524
rect 1995 34493 2007 34496
rect 1949 34487 2007 34493
rect 2222 34484 2228 34496
rect 2280 34484 2286 34536
rect 2409 34527 2467 34533
rect 2409 34493 2421 34527
rect 2455 34524 2467 34527
rect 2498 34524 2504 34536
rect 2455 34496 2504 34524
rect 2455 34493 2467 34496
rect 2409 34487 2467 34493
rect 2498 34484 2504 34496
rect 2556 34484 2562 34536
rect 3053 34527 3111 34533
rect 3053 34493 3065 34527
rect 3099 34524 3111 34527
rect 3418 34524 3424 34536
rect 3099 34496 3424 34524
rect 3099 34493 3111 34496
rect 3053 34487 3111 34493
rect 3418 34484 3424 34496
rect 3476 34484 3482 34536
rect 3528 34533 3556 34564
rect 9858 34552 9864 34564
rect 9916 34552 9922 34604
rect 12066 34552 12072 34604
rect 12124 34592 12130 34604
rect 12894 34592 12900 34604
rect 12124 34564 12900 34592
rect 12124 34552 12130 34564
rect 12894 34552 12900 34564
rect 12952 34592 12958 34604
rect 12989 34595 13047 34601
rect 12989 34592 13001 34595
rect 12952 34564 13001 34592
rect 12952 34552 12958 34564
rect 12989 34561 13001 34564
rect 13035 34561 13047 34595
rect 12989 34555 13047 34561
rect 3513 34527 3571 34533
rect 3513 34493 3525 34527
rect 3559 34524 3571 34527
rect 3559 34496 4200 34524
rect 3559 34493 3571 34496
rect 3513 34487 3571 34493
rect 3780 34459 3838 34465
rect 3780 34425 3792 34459
rect 3826 34456 3838 34459
rect 3970 34456 3976 34468
rect 3826 34428 3976 34456
rect 3826 34425 3838 34428
rect 3780 34419 3838 34425
rect 3970 34416 3976 34428
rect 4028 34416 4034 34468
rect 4172 34456 4200 34496
rect 4890 34484 4896 34536
rect 4948 34524 4954 34536
rect 5537 34527 5595 34533
rect 5537 34524 5549 34527
rect 4948 34496 5549 34524
rect 4948 34484 4954 34496
rect 5537 34493 5549 34496
rect 5583 34524 5595 34527
rect 5902 34524 5908 34536
rect 5583 34496 5908 34524
rect 5583 34493 5595 34496
rect 5537 34487 5595 34493
rect 5902 34484 5908 34496
rect 5960 34484 5966 34536
rect 6270 34484 6276 34536
rect 6328 34524 6334 34536
rect 6365 34527 6423 34533
rect 6365 34524 6377 34527
rect 6328 34496 6377 34524
rect 6328 34484 6334 34496
rect 6365 34493 6377 34496
rect 6411 34524 6423 34527
rect 6822 34524 6828 34536
rect 6411 34496 6828 34524
rect 6411 34493 6423 34496
rect 6365 34487 6423 34493
rect 6822 34484 6828 34496
rect 6880 34484 6886 34536
rect 7374 34524 7380 34536
rect 7335 34496 7380 34524
rect 7374 34484 7380 34496
rect 7432 34484 7438 34536
rect 7644 34527 7702 34533
rect 7644 34493 7656 34527
rect 7690 34524 7702 34527
rect 7926 34524 7932 34536
rect 7690 34496 7932 34524
rect 7690 34493 7702 34496
rect 7644 34487 7702 34493
rect 7926 34484 7932 34496
rect 7984 34484 7990 34536
rect 8754 34484 8760 34536
rect 8812 34524 8818 34536
rect 9309 34527 9367 34533
rect 9309 34524 9321 34527
rect 8812 34496 9321 34524
rect 8812 34484 8818 34496
rect 9309 34493 9321 34496
rect 9355 34493 9367 34527
rect 9309 34487 9367 34493
rect 12342 34484 12348 34536
rect 12400 34484 12406 34536
rect 13096 34524 13124 34632
rect 13170 34524 13176 34536
rect 12912 34496 13176 34524
rect 4706 34456 4712 34468
rect 4172 34428 4712 34456
rect 4706 34416 4712 34428
rect 4764 34416 4770 34468
rect 10128 34459 10186 34465
rect 10128 34425 10140 34459
rect 10174 34456 10186 34459
rect 10778 34456 10784 34468
rect 10174 34428 10784 34456
rect 10174 34425 10186 34428
rect 10128 34419 10186 34425
rect 10778 34416 10784 34428
rect 10836 34416 10842 34468
rect 12360 34456 12388 34484
rect 12912 34465 12940 34496
rect 13170 34484 13176 34496
rect 13228 34484 13234 34536
rect 12805 34459 12863 34465
rect 12805 34456 12817 34459
rect 12360 34428 12817 34456
rect 12805 34425 12817 34428
rect 12851 34425 12863 34459
rect 12805 34419 12863 34425
rect 12897 34459 12955 34465
rect 12897 34425 12909 34459
rect 12943 34425 12955 34459
rect 12897 34419 12955 34425
rect 4798 34348 4804 34400
rect 4856 34388 4862 34400
rect 4893 34391 4951 34397
rect 4893 34388 4905 34391
rect 4856 34360 4905 34388
rect 4856 34348 4862 34360
rect 4893 34357 4905 34360
rect 4939 34357 4951 34391
rect 4893 34351 4951 34357
rect 8757 34391 8815 34397
rect 8757 34357 8769 34391
rect 8803 34388 8815 34391
rect 8846 34388 8852 34400
rect 8803 34360 8852 34388
rect 8803 34357 8815 34360
rect 8757 34351 8815 34357
rect 8846 34348 8852 34360
rect 8904 34388 8910 34400
rect 9490 34388 9496 34400
rect 8904 34360 9496 34388
rect 8904 34348 8910 34360
rect 9490 34348 9496 34360
rect 9548 34348 9554 34400
rect 11238 34388 11244 34400
rect 11199 34360 11244 34388
rect 11238 34348 11244 34360
rect 11296 34348 11302 34400
rect 12434 34348 12440 34400
rect 12492 34388 12498 34400
rect 12492 34360 12537 34388
rect 12492 34348 12498 34360
rect 1104 34298 14812 34320
rect 1104 34246 6315 34298
rect 6367 34246 6379 34298
rect 6431 34246 6443 34298
rect 6495 34246 6507 34298
rect 6559 34246 11648 34298
rect 11700 34246 11712 34298
rect 11764 34246 11776 34298
rect 11828 34246 11840 34298
rect 11892 34246 14812 34298
rect 1104 34224 14812 34246
rect 1394 34144 1400 34196
rect 1452 34184 1458 34196
rect 2409 34187 2467 34193
rect 2409 34184 2421 34187
rect 1452 34156 2421 34184
rect 1452 34144 1458 34156
rect 2409 34153 2421 34156
rect 2455 34153 2467 34187
rect 9490 34184 9496 34196
rect 9451 34156 9496 34184
rect 2409 34147 2467 34153
rect 9490 34144 9496 34156
rect 9548 34144 9554 34196
rect 9858 34184 9864 34196
rect 9819 34156 9864 34184
rect 9858 34144 9864 34156
rect 9916 34184 9922 34196
rect 9916 34156 11100 34184
rect 9916 34144 9922 34156
rect 1670 34116 1676 34128
rect 1631 34088 1676 34116
rect 1670 34076 1676 34088
rect 1728 34076 1734 34128
rect 11072 34060 11100 34156
rect 11238 34116 11244 34128
rect 11151 34088 11244 34116
rect 11238 34076 11244 34088
rect 11296 34116 11302 34128
rect 12066 34125 12072 34128
rect 12060 34116 12072 34125
rect 11296 34088 12072 34116
rect 11296 34076 11302 34088
rect 12060 34079 12072 34088
rect 12066 34076 12072 34079
rect 12124 34076 12130 34128
rect 2225 34051 2283 34057
rect 2225 34017 2237 34051
rect 2271 34048 2283 34051
rect 2590 34048 2596 34060
rect 2271 34020 2596 34048
rect 2271 34017 2283 34020
rect 2225 34011 2283 34017
rect 2590 34008 2596 34020
rect 2648 34008 2654 34060
rect 4798 34008 4804 34060
rect 4856 34048 4862 34060
rect 4965 34051 5023 34057
rect 4965 34048 4977 34051
rect 4856 34020 4977 34048
rect 4856 34008 4862 34020
rect 4965 34017 4977 34020
rect 5011 34017 5023 34051
rect 4965 34011 5023 34017
rect 6270 34008 6276 34060
rect 6328 34048 6334 34060
rect 7929 34051 7987 34057
rect 7929 34048 7941 34051
rect 6328 34020 7941 34048
rect 6328 34008 6334 34020
rect 7929 34017 7941 34020
rect 7975 34048 7987 34051
rect 8478 34048 8484 34060
rect 7975 34020 8484 34048
rect 7975 34017 7987 34020
rect 7929 34011 7987 34017
rect 8478 34008 8484 34020
rect 8536 34008 8542 34060
rect 8570 34008 8576 34060
rect 8628 34048 8634 34060
rect 10226 34048 10232 34060
rect 8628 34020 10232 34048
rect 8628 34008 8634 34020
rect 10226 34008 10232 34020
rect 10284 34048 10290 34060
rect 10505 34051 10563 34057
rect 10505 34048 10517 34051
rect 10284 34020 10517 34048
rect 10284 34008 10290 34020
rect 10505 34017 10517 34020
rect 10551 34017 10563 34051
rect 11054 34048 11060 34060
rect 10967 34020 11060 34048
rect 10505 34011 10563 34017
rect 11054 34008 11060 34020
rect 11112 34048 11118 34060
rect 11790 34048 11796 34060
rect 11112 34020 11796 34048
rect 11112 34008 11118 34020
rect 11790 34008 11796 34020
rect 11848 34008 11854 34060
rect 4706 33980 4712 33992
rect 4667 33952 4712 33980
rect 4706 33940 4712 33952
rect 4764 33940 4770 33992
rect 8021 33983 8079 33989
rect 8021 33980 8033 33983
rect 7024 33952 8033 33980
rect 3605 33847 3663 33853
rect 3605 33813 3617 33847
rect 3651 33844 3663 33847
rect 3970 33844 3976 33856
rect 3651 33816 3976 33844
rect 3651 33813 3663 33816
rect 3605 33807 3663 33813
rect 3970 33804 3976 33816
rect 4028 33804 4034 33856
rect 6086 33844 6092 33856
rect 6047 33816 6092 33844
rect 6086 33804 6092 33816
rect 6144 33804 6150 33856
rect 6914 33804 6920 33856
rect 6972 33844 6978 33856
rect 7024 33853 7052 33952
rect 8021 33949 8033 33952
rect 8067 33949 8079 33983
rect 8021 33943 8079 33949
rect 8205 33983 8263 33989
rect 8205 33949 8217 33983
rect 8251 33980 8263 33983
rect 8846 33980 8852 33992
rect 8251 33952 8852 33980
rect 8251 33949 8263 33952
rect 8205 33943 8263 33949
rect 8846 33940 8852 33952
rect 8904 33940 8910 33992
rect 10318 33940 10324 33992
rect 10376 33980 10382 33992
rect 10597 33983 10655 33989
rect 10597 33980 10609 33983
rect 10376 33952 10609 33980
rect 10376 33940 10382 33952
rect 10597 33949 10609 33952
rect 10643 33949 10655 33983
rect 10778 33980 10784 33992
rect 10739 33952 10784 33980
rect 10597 33943 10655 33949
rect 10778 33940 10784 33952
rect 10836 33940 10842 33992
rect 7374 33872 7380 33924
rect 7432 33912 7438 33924
rect 7469 33915 7527 33921
rect 7469 33912 7481 33915
rect 7432 33884 7481 33912
rect 7432 33872 7438 33884
rect 7469 33881 7481 33884
rect 7515 33912 7527 33915
rect 7834 33912 7840 33924
rect 7515 33884 7840 33912
rect 7515 33881 7527 33884
rect 7469 33875 7527 33881
rect 7834 33872 7840 33884
rect 7892 33872 7898 33924
rect 7009 33847 7067 33853
rect 7009 33844 7021 33847
rect 6972 33816 7021 33844
rect 6972 33804 6978 33816
rect 7009 33813 7021 33816
rect 7055 33813 7067 33847
rect 7558 33844 7564 33856
rect 7519 33816 7564 33844
rect 7009 33807 7067 33813
rect 7558 33804 7564 33816
rect 7616 33804 7622 33856
rect 10137 33847 10195 33853
rect 10137 33813 10149 33847
rect 10183 33844 10195 33847
rect 10502 33844 10508 33856
rect 10183 33816 10508 33844
rect 10183 33813 10195 33816
rect 10137 33807 10195 33813
rect 10502 33804 10508 33816
rect 10560 33804 10566 33856
rect 12894 33804 12900 33856
rect 12952 33844 12958 33856
rect 13173 33847 13231 33853
rect 13173 33844 13185 33847
rect 12952 33816 13185 33844
rect 12952 33804 12958 33816
rect 13173 33813 13185 33816
rect 13219 33813 13231 33847
rect 13173 33807 13231 33813
rect 1104 33754 14812 33776
rect 1104 33702 3648 33754
rect 3700 33702 3712 33754
rect 3764 33702 3776 33754
rect 3828 33702 3840 33754
rect 3892 33702 8982 33754
rect 9034 33702 9046 33754
rect 9098 33702 9110 33754
rect 9162 33702 9174 33754
rect 9226 33702 14315 33754
rect 14367 33702 14379 33754
rect 14431 33702 14443 33754
rect 14495 33702 14507 33754
rect 14559 33702 14812 33754
rect 1104 33680 14812 33702
rect 1486 33600 1492 33652
rect 1544 33640 1550 33652
rect 1581 33643 1639 33649
rect 1581 33640 1593 33643
rect 1544 33612 1593 33640
rect 1544 33600 1550 33612
rect 1581 33609 1593 33612
rect 1627 33609 1639 33643
rect 1581 33603 1639 33609
rect 2958 33600 2964 33652
rect 3016 33640 3022 33652
rect 3053 33643 3111 33649
rect 3053 33640 3065 33643
rect 3016 33612 3065 33640
rect 3016 33600 3022 33612
rect 3053 33609 3065 33612
rect 3099 33609 3111 33643
rect 4154 33640 4160 33652
rect 4115 33612 4160 33640
rect 3053 33603 3111 33609
rect 4154 33600 4160 33612
rect 4212 33600 4218 33652
rect 4982 33600 4988 33652
rect 5040 33640 5046 33652
rect 5261 33643 5319 33649
rect 5261 33640 5273 33643
rect 5040 33612 5273 33640
rect 5040 33600 5046 33612
rect 5261 33609 5273 33612
rect 5307 33609 5319 33643
rect 6270 33640 6276 33652
rect 6231 33612 6276 33640
rect 5261 33603 5319 33609
rect 6270 33600 6276 33612
rect 6328 33600 6334 33652
rect 8846 33640 8852 33652
rect 8807 33612 8852 33640
rect 8846 33600 8852 33612
rect 8904 33600 8910 33652
rect 9401 33643 9459 33649
rect 9401 33609 9413 33643
rect 9447 33640 9459 33643
rect 10778 33640 10784 33652
rect 9447 33612 10784 33640
rect 9447 33609 9459 33612
rect 9401 33603 9459 33609
rect 10778 33600 10784 33612
rect 10836 33600 10842 33652
rect 11790 33600 11796 33652
rect 11848 33640 11854 33652
rect 11977 33643 12035 33649
rect 11977 33640 11989 33643
rect 11848 33612 11989 33640
rect 11848 33600 11854 33612
rect 11977 33609 11989 33612
rect 12023 33609 12035 33643
rect 11977 33603 12035 33609
rect 9674 33572 9680 33584
rect 9635 33544 9680 33572
rect 9674 33532 9680 33544
rect 9732 33532 9738 33584
rect 10318 33532 10324 33584
rect 10376 33572 10382 33584
rect 10413 33575 10471 33581
rect 10413 33572 10425 33575
rect 10376 33544 10425 33572
rect 10376 33532 10382 33544
rect 10413 33541 10425 33544
rect 10459 33541 10471 33575
rect 10413 33535 10471 33541
rect 4706 33464 4712 33516
rect 4764 33504 4770 33516
rect 4985 33507 5043 33513
rect 4985 33504 4997 33507
rect 4764 33476 4997 33504
rect 4764 33464 4770 33476
rect 4985 33473 4997 33476
rect 5031 33504 5043 33507
rect 6641 33507 6699 33513
rect 6641 33504 6653 33507
rect 5031 33476 6653 33504
rect 5031 33473 5043 33476
rect 4985 33467 5043 33473
rect 6641 33473 6653 33476
rect 6687 33504 6699 33507
rect 11238 33504 11244 33516
rect 6687 33476 6868 33504
rect 11199 33476 11244 33504
rect 6687 33473 6699 33476
rect 6641 33467 6699 33473
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33405 1455 33439
rect 1397 33399 1455 33405
rect 2869 33439 2927 33445
rect 2869 33405 2881 33439
rect 2915 33436 2927 33439
rect 3973 33439 4031 33445
rect 2915 33408 3556 33436
rect 2915 33405 2927 33408
rect 2869 33399 2927 33405
rect 1412 33368 1440 33399
rect 1946 33368 1952 33380
rect 1412 33340 1952 33368
rect 1946 33328 1952 33340
rect 2004 33328 2010 33380
rect 2317 33303 2375 33309
rect 2317 33269 2329 33303
rect 2363 33300 2375 33303
rect 2590 33300 2596 33312
rect 2363 33272 2596 33300
rect 2363 33269 2375 33272
rect 2317 33263 2375 33269
rect 2590 33260 2596 33272
rect 2648 33260 2654 33312
rect 3528 33309 3556 33408
rect 3973 33405 3985 33439
rect 4019 33436 4031 33439
rect 5077 33439 5135 33445
rect 4019 33408 4660 33436
rect 4019 33405 4031 33408
rect 3973 33399 4031 33405
rect 4632 33312 4660 33408
rect 5077 33405 5089 33439
rect 5123 33436 5135 33439
rect 5721 33439 5779 33445
rect 5721 33436 5733 33439
rect 5123 33408 5733 33436
rect 5123 33405 5135 33408
rect 5077 33399 5135 33405
rect 5721 33405 5733 33408
rect 5767 33436 5779 33439
rect 6730 33436 6736 33448
rect 5767 33408 6736 33436
rect 5767 33405 5779 33408
rect 5721 33399 5779 33405
rect 6730 33396 6736 33408
rect 6788 33396 6794 33448
rect 6840 33445 6868 33476
rect 11238 33464 11244 33476
rect 11296 33464 11302 33516
rect 12894 33464 12900 33516
rect 12952 33504 12958 33516
rect 12989 33507 13047 33513
rect 12989 33504 13001 33507
rect 12952 33476 13001 33504
rect 12952 33464 12958 33476
rect 12989 33473 13001 33476
rect 13035 33504 13047 33507
rect 13449 33507 13507 33513
rect 13449 33504 13461 33507
rect 13035 33476 13461 33504
rect 13035 33473 13047 33476
rect 12989 33467 13047 33473
rect 13449 33473 13461 33476
rect 13495 33473 13507 33507
rect 13449 33467 13507 33473
rect 6825 33439 6883 33445
rect 6825 33405 6837 33439
rect 6871 33436 6883 33439
rect 7834 33436 7840 33448
rect 6871 33408 7840 33436
rect 6871 33405 6883 33408
rect 6825 33399 6883 33405
rect 7834 33396 7840 33408
rect 7892 33396 7898 33448
rect 9493 33439 9551 33445
rect 9493 33405 9505 33439
rect 9539 33436 9551 33439
rect 10045 33439 10103 33445
rect 10045 33436 10057 33439
rect 9539 33408 10057 33436
rect 9539 33405 9551 33408
rect 9493 33399 9551 33405
rect 10045 33405 10057 33408
rect 10091 33436 10103 33439
rect 11146 33436 11152 33448
rect 10091 33408 11152 33436
rect 10091 33405 10103 33408
rect 10045 33399 10103 33405
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 12434 33396 12440 33448
rect 12492 33436 12498 33448
rect 12805 33439 12863 33445
rect 12805 33436 12817 33439
rect 12492 33408 12817 33436
rect 12492 33396 12498 33408
rect 12805 33405 12817 33408
rect 12851 33436 12863 33439
rect 13817 33439 13875 33445
rect 13817 33436 13829 33439
rect 12851 33408 13829 33436
rect 12851 33405 12863 33408
rect 12805 33399 12863 33405
rect 13817 33405 13829 33408
rect 13863 33405 13875 33439
rect 13817 33399 13875 33405
rect 6086 33328 6092 33380
rect 6144 33368 6150 33380
rect 7098 33377 7104 33380
rect 7070 33371 7104 33377
rect 7070 33368 7082 33371
rect 6144 33340 7082 33368
rect 6144 33328 6150 33340
rect 7070 33337 7082 33340
rect 7156 33368 7162 33380
rect 7156 33340 7218 33368
rect 7070 33331 7104 33337
rect 7098 33328 7104 33331
rect 7156 33328 7162 33340
rect 10502 33328 10508 33380
rect 10560 33368 10566 33380
rect 11057 33371 11115 33377
rect 11057 33368 11069 33371
rect 10560 33340 11069 33368
rect 10560 33328 10566 33340
rect 11057 33337 11069 33340
rect 11103 33337 11115 33371
rect 11057 33331 11115 33337
rect 3513 33303 3571 33309
rect 3513 33269 3525 33303
rect 3559 33300 3571 33303
rect 4062 33300 4068 33312
rect 3559 33272 4068 33300
rect 3559 33269 3571 33272
rect 3513 33263 3571 33269
rect 4062 33260 4068 33272
rect 4120 33260 4126 33312
rect 4614 33300 4620 33312
rect 4575 33272 4620 33300
rect 4614 33260 4620 33272
rect 4672 33260 4678 33312
rect 6822 33260 6828 33312
rect 6880 33300 6886 33312
rect 7466 33300 7472 33312
rect 6880 33272 7472 33300
rect 6880 33260 6886 33272
rect 7466 33260 7472 33272
rect 7524 33300 7530 33312
rect 8205 33303 8263 33309
rect 8205 33300 8217 33303
rect 7524 33272 8217 33300
rect 7524 33260 7530 33272
rect 8205 33269 8217 33272
rect 8251 33269 8263 33303
rect 10594 33300 10600 33312
rect 10555 33272 10600 33300
rect 8205 33263 8263 33269
rect 10594 33260 10600 33272
rect 10652 33260 10658 33312
rect 10778 33260 10784 33312
rect 10836 33300 10842 33312
rect 10965 33303 11023 33309
rect 10965 33300 10977 33303
rect 10836 33272 10977 33300
rect 10836 33260 10842 33272
rect 10965 33269 10977 33272
rect 11011 33300 11023 33303
rect 11609 33303 11667 33309
rect 11609 33300 11621 33303
rect 11011 33272 11621 33300
rect 11011 33269 11023 33272
rect 10965 33263 11023 33269
rect 11609 33269 11621 33272
rect 11655 33269 11667 33303
rect 11609 33263 11667 33269
rect 12342 33260 12348 33312
rect 12400 33300 12406 33312
rect 12437 33303 12495 33309
rect 12437 33300 12449 33303
rect 12400 33272 12449 33300
rect 12400 33260 12406 33272
rect 12437 33269 12449 33272
rect 12483 33269 12495 33303
rect 12894 33300 12900 33312
rect 12855 33272 12900 33300
rect 12437 33263 12495 33269
rect 12894 33260 12900 33272
rect 12952 33260 12958 33312
rect 1104 33210 14812 33232
rect 1104 33158 6315 33210
rect 6367 33158 6379 33210
rect 6431 33158 6443 33210
rect 6495 33158 6507 33210
rect 6559 33158 11648 33210
rect 11700 33158 11712 33210
rect 11764 33158 11776 33210
rect 11828 33158 11840 33210
rect 11892 33158 14812 33210
rect 1104 33136 14812 33158
rect 1578 33096 1584 33108
rect 1539 33068 1584 33096
rect 1578 33056 1584 33068
rect 1636 33056 1642 33108
rect 5442 33056 5448 33108
rect 5500 33096 5506 33108
rect 6089 33099 6147 33105
rect 6089 33096 6101 33099
rect 5500 33068 6101 33096
rect 5500 33056 5506 33068
rect 6089 33065 6101 33068
rect 6135 33096 6147 33099
rect 7285 33099 7343 33105
rect 7285 33096 7297 33099
rect 6135 33068 7297 33096
rect 6135 33065 6147 33068
rect 6089 33059 6147 33065
rect 7285 33065 7297 33068
rect 7331 33065 7343 33099
rect 7285 33059 7343 33065
rect 7374 33056 7380 33108
rect 7432 33096 7438 33108
rect 7653 33099 7711 33105
rect 7653 33096 7665 33099
rect 7432 33068 7665 33096
rect 7432 33056 7438 33068
rect 7653 33065 7665 33068
rect 7699 33096 7711 33099
rect 8018 33096 8024 33108
rect 7699 33068 8024 33096
rect 7699 33065 7711 33068
rect 7653 33059 7711 33065
rect 8018 33056 8024 33068
rect 8076 33056 8082 33108
rect 9950 33056 9956 33108
rect 10008 33096 10014 33108
rect 10226 33096 10232 33108
rect 10008 33068 10232 33096
rect 10008 33056 10014 33068
rect 10226 33056 10232 33068
rect 10284 33056 10290 33108
rect 10502 33096 10508 33108
rect 10463 33068 10508 33096
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 10594 33056 10600 33108
rect 10652 33096 10658 33108
rect 11149 33099 11207 33105
rect 11149 33096 11161 33099
rect 10652 33068 11161 33096
rect 10652 33056 10658 33068
rect 11149 33065 11161 33068
rect 11195 33096 11207 33099
rect 12253 33099 12311 33105
rect 12253 33096 12265 33099
rect 11195 33068 12265 33096
rect 11195 33065 11207 33068
rect 11149 33059 11207 33065
rect 12253 33065 12265 33068
rect 12299 33065 12311 33099
rect 12710 33096 12716 33108
rect 12671 33068 12716 33096
rect 12253 33059 12311 33065
rect 12710 33056 12716 33068
rect 12768 33056 12774 33108
rect 6917 33031 6975 33037
rect 6917 32997 6929 33031
rect 6963 33028 6975 33031
rect 7098 33028 7104 33040
rect 6963 33000 7104 33028
rect 6963 32997 6975 33000
rect 6917 32991 6975 32997
rect 7098 32988 7104 33000
rect 7156 33028 7162 33040
rect 11057 33031 11115 33037
rect 7156 33000 7788 33028
rect 7156 32988 7162 33000
rect 1394 32960 1400 32972
rect 1355 32932 1400 32960
rect 1394 32920 1400 32932
rect 1452 32920 1458 32972
rect 7760 32960 7788 33000
rect 11057 32997 11069 33031
rect 11103 33028 11115 33031
rect 11514 33028 11520 33040
rect 11103 33000 11520 33028
rect 11103 32997 11115 33000
rect 11057 32991 11115 32997
rect 11514 32988 11520 33000
rect 11572 33028 11578 33040
rect 12342 33028 12348 33040
rect 11572 33000 12348 33028
rect 11572 32988 11578 33000
rect 12342 32988 12348 33000
rect 12400 32988 12406 33040
rect 12618 32960 12624 32972
rect 7760 32932 7880 32960
rect 12579 32932 12624 32960
rect 6178 32892 6184 32904
rect 6139 32864 6184 32892
rect 6178 32852 6184 32864
rect 6236 32852 6242 32904
rect 6362 32892 6368 32904
rect 6275 32864 6368 32892
rect 6362 32852 6368 32864
rect 6420 32892 6426 32904
rect 6822 32892 6828 32904
rect 6420 32864 6828 32892
rect 6420 32852 6426 32864
rect 6822 32852 6828 32864
rect 6880 32852 6886 32904
rect 7282 32852 7288 32904
rect 7340 32892 7346 32904
rect 7742 32892 7748 32904
rect 7340 32864 7748 32892
rect 7340 32852 7346 32864
rect 7742 32852 7748 32864
rect 7800 32852 7806 32904
rect 7852 32901 7880 32932
rect 12618 32920 12624 32932
rect 12676 32920 12682 32972
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 10042 32892 10048 32904
rect 9723 32864 10048 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 10042 32852 10048 32864
rect 10100 32852 10106 32904
rect 10318 32852 10324 32904
rect 10376 32892 10382 32904
rect 11333 32895 11391 32901
rect 11333 32892 11345 32895
rect 10376 32864 11345 32892
rect 10376 32852 10382 32864
rect 11333 32861 11345 32864
rect 11379 32892 11391 32895
rect 12342 32892 12348 32904
rect 11379 32864 12348 32892
rect 11379 32861 11391 32864
rect 11333 32855 11391 32861
rect 12342 32852 12348 32864
rect 12400 32852 12406 32904
rect 12802 32892 12808 32904
rect 12763 32864 12808 32892
rect 12802 32852 12808 32864
rect 12860 32852 12866 32904
rect 9858 32784 9864 32836
rect 9916 32824 9922 32836
rect 10689 32827 10747 32833
rect 10689 32824 10701 32827
rect 9916 32796 10701 32824
rect 9916 32784 9922 32796
rect 10689 32793 10701 32796
rect 10735 32793 10747 32827
rect 10689 32787 10747 32793
rect 11146 32784 11152 32836
rect 11204 32824 11210 32836
rect 12066 32824 12072 32836
rect 11204 32796 12072 32824
rect 11204 32784 11210 32796
rect 12066 32784 12072 32796
rect 12124 32784 12130 32836
rect 3326 32756 3332 32768
rect 3287 32728 3332 32756
rect 3326 32716 3332 32728
rect 3384 32716 3390 32768
rect 4154 32716 4160 32768
rect 4212 32756 4218 32768
rect 4709 32759 4767 32765
rect 4709 32756 4721 32759
rect 4212 32728 4721 32756
rect 4212 32716 4218 32728
rect 4709 32725 4721 32728
rect 4755 32756 4767 32759
rect 4798 32756 4804 32768
rect 4755 32728 4804 32756
rect 4755 32725 4767 32728
rect 4709 32719 4767 32725
rect 4798 32716 4804 32728
rect 4856 32716 4862 32768
rect 5718 32756 5724 32768
rect 5679 32728 5724 32756
rect 5718 32716 5724 32728
rect 5776 32716 5782 32768
rect 8294 32756 8300 32768
rect 8255 32728 8300 32756
rect 8294 32716 8300 32728
rect 8352 32716 8358 32768
rect 11238 32716 11244 32768
rect 11296 32756 11302 32768
rect 11790 32756 11796 32768
rect 11296 32728 11796 32756
rect 11296 32716 11302 32728
rect 11790 32716 11796 32728
rect 11848 32716 11854 32768
rect 12434 32716 12440 32768
rect 12492 32756 12498 32768
rect 12894 32756 12900 32768
rect 12492 32728 12900 32756
rect 12492 32716 12498 32728
rect 12894 32716 12900 32728
rect 12952 32756 12958 32768
rect 13265 32759 13323 32765
rect 13265 32756 13277 32759
rect 12952 32728 13277 32756
rect 12952 32716 12958 32728
rect 13265 32725 13277 32728
rect 13311 32725 13323 32759
rect 13265 32719 13323 32725
rect 1104 32666 14812 32688
rect 1104 32614 3648 32666
rect 3700 32614 3712 32666
rect 3764 32614 3776 32666
rect 3828 32614 3840 32666
rect 3892 32614 8982 32666
rect 9034 32614 9046 32666
rect 9098 32614 9110 32666
rect 9162 32614 9174 32666
rect 9226 32614 14315 32666
rect 14367 32614 14379 32666
rect 14431 32614 14443 32666
rect 14495 32614 14507 32666
rect 14559 32614 14812 32666
rect 1104 32592 14812 32614
rect 1394 32512 1400 32564
rect 1452 32552 1458 32564
rect 1581 32555 1639 32561
rect 1581 32552 1593 32555
rect 1452 32524 1593 32552
rect 1452 32512 1458 32524
rect 1581 32521 1593 32524
rect 1627 32521 1639 32555
rect 5442 32552 5448 32564
rect 5403 32524 5448 32552
rect 1581 32515 1639 32521
rect 5442 32512 5448 32524
rect 5500 32512 5506 32564
rect 6178 32552 6184 32564
rect 6139 32524 6184 32552
rect 6178 32512 6184 32524
rect 6236 32512 6242 32564
rect 6641 32555 6699 32561
rect 6641 32521 6653 32555
rect 6687 32552 6699 32555
rect 7374 32552 7380 32564
rect 6687 32524 7380 32552
rect 6687 32521 6699 32524
rect 6641 32515 6699 32521
rect 7374 32512 7380 32524
rect 7432 32512 7438 32564
rect 7926 32512 7932 32564
rect 7984 32552 7990 32564
rect 8386 32552 8392 32564
rect 7984 32524 8392 32552
rect 7984 32512 7990 32524
rect 8386 32512 8392 32524
rect 8444 32552 8450 32564
rect 9125 32555 9183 32561
rect 9125 32552 9137 32555
rect 8444 32524 9137 32552
rect 8444 32512 8450 32524
rect 9125 32521 9137 32524
rect 9171 32521 9183 32555
rect 9125 32515 9183 32521
rect 9953 32555 10011 32561
rect 9953 32521 9965 32555
rect 9999 32552 10011 32555
rect 10594 32552 10600 32564
rect 9999 32524 10600 32552
rect 9999 32521 10011 32524
rect 9953 32515 10011 32521
rect 10594 32512 10600 32524
rect 10652 32512 10658 32564
rect 10778 32552 10784 32564
rect 10739 32524 10784 32552
rect 10778 32512 10784 32524
rect 10836 32512 10842 32564
rect 11790 32552 11796 32564
rect 11751 32524 11796 32552
rect 11790 32512 11796 32524
rect 11848 32512 11854 32564
rect 12066 32512 12072 32564
rect 12124 32552 12130 32564
rect 12161 32555 12219 32561
rect 12161 32552 12173 32555
rect 12124 32524 12173 32552
rect 12124 32512 12130 32524
rect 12161 32521 12173 32524
rect 12207 32552 12219 32555
rect 12250 32552 12256 32564
rect 12207 32524 12256 32552
rect 12207 32521 12219 32524
rect 12161 32515 12219 32521
rect 12250 32512 12256 32524
rect 12308 32512 12314 32564
rect 12434 32512 12440 32564
rect 12492 32552 12498 32564
rect 12492 32524 12537 32552
rect 12492 32512 12498 32524
rect 12618 32512 12624 32564
rect 12676 32552 12682 32564
rect 13817 32555 13875 32561
rect 13817 32552 13829 32555
rect 12676 32524 13829 32552
rect 12676 32512 12682 32524
rect 13817 32521 13829 32524
rect 13863 32521 13875 32555
rect 13817 32515 13875 32521
rect 5813 32487 5871 32493
rect 5813 32453 5825 32487
rect 5859 32484 5871 32487
rect 6362 32484 6368 32496
rect 5859 32456 6368 32484
rect 5859 32453 5871 32456
rect 5813 32447 5871 32453
rect 6362 32444 6368 32456
rect 6420 32444 6426 32496
rect 10318 32484 10324 32496
rect 10279 32456 10324 32484
rect 10318 32444 10324 32456
rect 10376 32444 10382 32496
rect 3326 32376 3332 32428
rect 3384 32416 3390 32428
rect 3786 32416 3792 32428
rect 3384 32388 3792 32416
rect 3384 32376 3390 32388
rect 3786 32376 3792 32388
rect 3844 32376 3850 32428
rect 10778 32376 10784 32428
rect 10836 32416 10842 32428
rect 11241 32419 11299 32425
rect 11241 32416 11253 32419
rect 10836 32388 11253 32416
rect 10836 32376 10842 32388
rect 11241 32385 11253 32388
rect 11287 32385 11299 32419
rect 11241 32379 11299 32385
rect 11425 32419 11483 32425
rect 11425 32385 11437 32419
rect 11471 32416 11483 32419
rect 11808 32416 11836 32512
rect 12710 32444 12716 32496
rect 12768 32484 12774 32496
rect 13449 32487 13507 32493
rect 13449 32484 13461 32487
rect 12768 32456 13461 32484
rect 12768 32444 12774 32456
rect 13449 32453 13461 32456
rect 13495 32453 13507 32487
rect 13449 32447 13507 32453
rect 12989 32419 13047 32425
rect 12989 32416 13001 32419
rect 11471 32388 13001 32416
rect 11471 32385 11483 32388
rect 11425 32379 11483 32385
rect 12989 32385 13001 32388
rect 13035 32385 13047 32419
rect 12989 32379 13047 32385
rect 3694 32348 3700 32360
rect 3655 32320 3700 32348
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 7282 32348 7288 32360
rect 7243 32320 7288 32348
rect 7282 32308 7288 32320
rect 7340 32308 7346 32360
rect 7745 32351 7803 32357
rect 7745 32317 7757 32351
rect 7791 32348 7803 32351
rect 7834 32348 7840 32360
rect 7791 32320 7840 32348
rect 7791 32317 7803 32320
rect 7745 32311 7803 32317
rect 7834 32308 7840 32320
rect 7892 32308 7898 32360
rect 8018 32357 8024 32360
rect 8012 32348 8024 32357
rect 7931 32320 8024 32348
rect 8012 32311 8024 32320
rect 8076 32348 8082 32360
rect 8294 32348 8300 32360
rect 8076 32320 8300 32348
rect 8018 32308 8024 32311
rect 8076 32308 8082 32320
rect 8294 32308 8300 32320
rect 8352 32308 8358 32360
rect 12526 32308 12532 32360
rect 12584 32348 12590 32360
rect 12897 32351 12955 32357
rect 12897 32348 12909 32351
rect 12584 32320 12909 32348
rect 12584 32308 12590 32320
rect 12897 32317 12909 32320
rect 12943 32348 12955 32351
rect 13170 32348 13176 32360
rect 12943 32320 13176 32348
rect 12943 32317 12955 32320
rect 12897 32311 12955 32317
rect 13170 32308 13176 32320
rect 13228 32308 13234 32360
rect 3145 32283 3203 32289
rect 3145 32249 3157 32283
rect 3191 32280 3203 32283
rect 3191 32252 3648 32280
rect 3191 32249 3203 32252
rect 3145 32243 3203 32249
rect 3620 32224 3648 32252
rect 3234 32212 3240 32224
rect 3195 32184 3240 32212
rect 3234 32172 3240 32184
rect 3292 32172 3298 32224
rect 3602 32212 3608 32224
rect 3563 32184 3608 32212
rect 3602 32172 3608 32184
rect 3660 32172 3666 32224
rect 4617 32215 4675 32221
rect 4617 32181 4629 32215
rect 4663 32212 4675 32215
rect 4982 32212 4988 32224
rect 4663 32184 4988 32212
rect 4663 32181 4675 32184
rect 4617 32175 4675 32181
rect 4982 32172 4988 32184
rect 5040 32172 5046 32224
rect 10686 32212 10692 32224
rect 10599 32184 10692 32212
rect 10686 32172 10692 32184
rect 10744 32212 10750 32224
rect 11146 32212 11152 32224
rect 10744 32184 11152 32212
rect 10744 32172 10750 32184
rect 11146 32172 11152 32184
rect 11204 32172 11210 32224
rect 12250 32172 12256 32224
rect 12308 32212 12314 32224
rect 12805 32215 12863 32221
rect 12805 32212 12817 32215
rect 12308 32184 12817 32212
rect 12308 32172 12314 32184
rect 12805 32181 12817 32184
rect 12851 32181 12863 32215
rect 12805 32175 12863 32181
rect 1104 32122 14812 32144
rect 1104 32070 6315 32122
rect 6367 32070 6379 32122
rect 6431 32070 6443 32122
rect 6495 32070 6507 32122
rect 6559 32070 11648 32122
rect 11700 32070 11712 32122
rect 11764 32070 11776 32122
rect 11828 32070 11840 32122
rect 11892 32070 14812 32122
rect 1104 32048 14812 32070
rect 3329 32011 3387 32017
rect 3329 31977 3341 32011
rect 3375 32008 3387 32011
rect 3694 32008 3700 32020
rect 3375 31980 3700 32008
rect 3375 31977 3387 31980
rect 3329 31971 3387 31977
rect 3694 31968 3700 31980
rect 3752 31968 3758 32020
rect 6178 31968 6184 32020
rect 6236 32008 6242 32020
rect 6549 32011 6607 32017
rect 6549 32008 6561 32011
rect 6236 31980 6561 32008
rect 6236 31968 6242 31980
rect 6549 31977 6561 31980
rect 6595 31977 6607 32011
rect 6549 31971 6607 31977
rect 6638 31968 6644 32020
rect 6696 32008 6702 32020
rect 7009 32011 7067 32017
rect 7009 32008 7021 32011
rect 6696 31980 7021 32008
rect 6696 31968 6702 31980
rect 7009 31977 7021 31980
rect 7055 31977 7067 32011
rect 7009 31971 7067 31977
rect 8573 32011 8631 32017
rect 8573 31977 8585 32011
rect 8619 32008 8631 32011
rect 8846 32008 8852 32020
rect 8619 31980 8852 32008
rect 8619 31977 8631 31980
rect 8573 31971 8631 31977
rect 8846 31968 8852 31980
rect 8904 32008 8910 32020
rect 9677 32011 9735 32017
rect 9677 32008 9689 32011
rect 8904 31980 9689 32008
rect 8904 31968 8910 31980
rect 9677 31977 9689 31980
rect 9723 31977 9735 32011
rect 10042 32008 10048 32020
rect 10003 31980 10048 32008
rect 9677 31971 9735 31977
rect 10042 31968 10048 31980
rect 10100 31968 10106 32020
rect 10137 32011 10195 32017
rect 10137 31977 10149 32011
rect 10183 32008 10195 32011
rect 10226 32008 10232 32020
rect 10183 31980 10232 32008
rect 10183 31977 10195 31980
rect 10137 31971 10195 31977
rect 3786 31900 3792 31952
rect 3844 31940 3850 31952
rect 4310 31943 4368 31949
rect 4310 31940 4322 31943
rect 3844 31912 4322 31940
rect 3844 31900 3850 31912
rect 4310 31909 4322 31912
rect 4356 31940 4368 31943
rect 4798 31940 4804 31952
rect 4356 31912 4804 31940
rect 4356 31909 4368 31912
rect 4310 31903 4368 31909
rect 4798 31900 4804 31912
rect 4856 31900 4862 31952
rect 6822 31900 6828 31952
rect 6880 31940 6886 31952
rect 6917 31943 6975 31949
rect 6917 31940 6929 31943
rect 6880 31912 6929 31940
rect 6880 31900 6886 31912
rect 6917 31909 6929 31912
rect 6963 31940 6975 31943
rect 7190 31940 7196 31952
rect 6963 31912 7196 31940
rect 6963 31909 6975 31912
rect 6917 31903 6975 31909
rect 7190 31900 7196 31912
rect 7248 31900 7254 31952
rect 9674 31832 9680 31884
rect 9732 31872 9738 31884
rect 10152 31872 10180 31971
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 10318 31968 10324 32020
rect 10376 32008 10382 32020
rect 10778 32008 10784 32020
rect 10376 31980 10784 32008
rect 10376 31968 10382 31980
rect 10778 31968 10784 31980
rect 10836 31968 10842 32020
rect 11238 32008 11244 32020
rect 11199 31980 11244 32008
rect 11238 31968 11244 31980
rect 11296 31968 11302 32020
rect 11514 32008 11520 32020
rect 11475 31980 11520 32008
rect 11514 31968 11520 31980
rect 11572 31968 11578 32020
rect 12526 32008 12532 32020
rect 12487 31980 12532 32008
rect 12526 31968 12532 31980
rect 12584 31968 12590 32020
rect 9732 31844 10180 31872
rect 9732 31832 9738 31844
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31773 4123 31807
rect 4065 31767 4123 31773
rect 6457 31807 6515 31813
rect 6457 31773 6469 31807
rect 6503 31804 6515 31807
rect 6503 31776 6868 31804
rect 6503 31773 6515 31776
rect 6457 31767 6515 31773
rect 4080 31668 4108 31767
rect 6840 31736 6868 31776
rect 7098 31764 7104 31816
rect 7156 31804 7162 31816
rect 7926 31804 7932 31816
rect 7156 31776 7932 31804
rect 7156 31764 7162 31776
rect 7926 31764 7932 31776
rect 7984 31804 7990 31816
rect 8113 31807 8171 31813
rect 8113 31804 8125 31807
rect 7984 31776 8125 31804
rect 7984 31764 7990 31776
rect 8113 31773 8125 31776
rect 8159 31773 8171 31807
rect 8113 31767 8171 31773
rect 9582 31764 9588 31816
rect 9640 31764 9646 31816
rect 10321 31807 10379 31813
rect 10321 31773 10333 31807
rect 10367 31804 10379 31807
rect 12802 31804 12808 31816
rect 10367 31776 10401 31804
rect 12360 31776 12808 31804
rect 10367 31773 10379 31776
rect 10321 31767 10379 31773
rect 7374 31736 7380 31748
rect 6840 31708 7380 31736
rect 7374 31696 7380 31708
rect 7432 31696 7438 31748
rect 9600 31680 9628 31764
rect 9766 31696 9772 31748
rect 9824 31696 9830 31748
rect 9950 31696 9956 31748
rect 10008 31736 10014 31748
rect 10336 31736 10364 31767
rect 10594 31736 10600 31748
rect 10008 31708 10600 31736
rect 10008 31696 10014 31708
rect 10594 31696 10600 31708
rect 10652 31696 10658 31748
rect 4246 31668 4252 31680
rect 4080 31640 4252 31668
rect 4246 31628 4252 31640
rect 4304 31668 4310 31680
rect 4706 31668 4712 31680
rect 4304 31640 4712 31668
rect 4304 31628 4310 31640
rect 4706 31628 4712 31640
rect 4764 31628 4770 31680
rect 5074 31628 5080 31680
rect 5132 31668 5138 31680
rect 5445 31671 5503 31677
rect 5445 31668 5457 31671
rect 5132 31640 5457 31668
rect 5132 31628 5138 31640
rect 5445 31637 5457 31640
rect 5491 31637 5503 31671
rect 7834 31668 7840 31680
rect 7795 31640 7840 31668
rect 5445 31631 5503 31637
rect 7834 31628 7840 31640
rect 7892 31628 7898 31680
rect 9582 31628 9588 31680
rect 9640 31628 9646 31680
rect 9784 31668 9812 31696
rect 10686 31668 10692 31680
rect 9784 31640 10692 31668
rect 10686 31628 10692 31640
rect 10744 31628 10750 31680
rect 12066 31628 12072 31680
rect 12124 31668 12130 31680
rect 12360 31668 12388 31776
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 12124 31640 12388 31668
rect 12124 31628 12130 31640
rect 1104 31578 14812 31600
rect 1104 31526 3648 31578
rect 3700 31526 3712 31578
rect 3764 31526 3776 31578
rect 3828 31526 3840 31578
rect 3892 31526 8982 31578
rect 9034 31526 9046 31578
rect 9098 31526 9110 31578
rect 9162 31526 9174 31578
rect 9226 31526 14315 31578
rect 14367 31526 14379 31578
rect 14431 31526 14443 31578
rect 14495 31526 14507 31578
rect 14559 31526 14812 31578
rect 1104 31504 14812 31526
rect 4157 31467 4215 31473
rect 4157 31433 4169 31467
rect 4203 31464 4215 31467
rect 4246 31464 4252 31476
rect 4203 31436 4252 31464
rect 4203 31433 4215 31436
rect 4157 31427 4215 31433
rect 4246 31424 4252 31436
rect 4304 31424 4310 31476
rect 6914 31464 6920 31476
rect 6875 31436 6920 31464
rect 6914 31424 6920 31436
rect 6972 31424 6978 31476
rect 7926 31464 7932 31476
rect 7887 31436 7932 31464
rect 7926 31424 7932 31436
rect 7984 31424 7990 31476
rect 8294 31424 8300 31476
rect 8352 31464 8358 31476
rect 8481 31467 8539 31473
rect 8481 31464 8493 31467
rect 8352 31436 8493 31464
rect 8352 31424 8358 31436
rect 8481 31433 8493 31436
rect 8527 31433 8539 31467
rect 8481 31427 8539 31433
rect 9674 31424 9680 31476
rect 9732 31464 9738 31476
rect 9861 31467 9919 31473
rect 9861 31464 9873 31467
rect 9732 31436 9873 31464
rect 9732 31424 9738 31436
rect 9861 31433 9873 31436
rect 9907 31464 9919 31467
rect 13538 31464 13544 31476
rect 9907 31436 10456 31464
rect 13499 31436 13544 31464
rect 9907 31433 9919 31436
rect 9861 31427 9919 31433
rect 2501 31399 2559 31405
rect 2501 31365 2513 31399
rect 2547 31396 2559 31399
rect 3510 31396 3516 31408
rect 2547 31368 3516 31396
rect 2547 31365 2559 31368
rect 2501 31359 2559 31365
rect 3510 31356 3516 31368
rect 3568 31356 3574 31408
rect 6273 31399 6331 31405
rect 6273 31365 6285 31399
rect 6319 31396 6331 31399
rect 6822 31396 6828 31408
rect 6319 31368 6828 31396
rect 6319 31365 6331 31368
rect 6273 31359 6331 31365
rect 6822 31356 6828 31368
rect 6880 31356 6886 31408
rect 10045 31399 10103 31405
rect 10045 31396 10057 31399
rect 8956 31368 10057 31396
rect 3605 31331 3663 31337
rect 3605 31297 3617 31331
rect 3651 31328 3663 31331
rect 4062 31328 4068 31340
rect 3651 31300 4068 31328
rect 3651 31297 3663 31300
rect 3605 31291 3663 31297
rect 2869 31263 2927 31269
rect 2869 31229 2881 31263
rect 2915 31260 2927 31263
rect 3620 31260 3648 31291
rect 4062 31288 4068 31300
rect 4120 31288 4126 31340
rect 5074 31328 5080 31340
rect 5035 31300 5080 31328
rect 5074 31288 5080 31300
rect 5132 31288 5138 31340
rect 7558 31328 7564 31340
rect 7471 31300 7564 31328
rect 7558 31288 7564 31300
rect 7616 31328 7622 31340
rect 8202 31328 8208 31340
rect 7616 31300 8208 31328
rect 7616 31288 7622 31300
rect 8202 31288 8208 31300
rect 8260 31328 8266 31340
rect 8297 31331 8355 31337
rect 8297 31328 8309 31331
rect 8260 31300 8309 31328
rect 8260 31288 8266 31300
rect 8297 31297 8309 31300
rect 8343 31297 8355 31331
rect 8297 31291 8355 31297
rect 2915 31232 3648 31260
rect 2915 31229 2927 31232
rect 2869 31223 2927 31229
rect 2133 31195 2191 31201
rect 2133 31161 2145 31195
rect 2179 31192 2191 31195
rect 2179 31164 3372 31192
rect 2179 31161 2191 31164
rect 2133 31155 2191 31161
rect 3344 31136 3372 31164
rect 4798 31152 4804 31204
rect 4856 31192 4862 31204
rect 5537 31195 5595 31201
rect 5537 31192 5549 31195
rect 4856 31164 5549 31192
rect 4856 31152 4862 31164
rect 5537 31161 5549 31164
rect 5583 31161 5595 31195
rect 8312 31192 8340 31291
rect 8570 31288 8576 31340
rect 8628 31328 8634 31340
rect 8956 31337 8984 31368
rect 10045 31365 10057 31368
rect 10091 31365 10103 31399
rect 10045 31359 10103 31365
rect 8941 31331 8999 31337
rect 8941 31328 8953 31331
rect 8628 31300 8953 31328
rect 8628 31288 8634 31300
rect 8941 31297 8953 31300
rect 8987 31297 8999 31331
rect 8941 31291 8999 31297
rect 9033 31331 9091 31337
rect 9033 31297 9045 31331
rect 9079 31297 9091 31331
rect 9033 31291 9091 31297
rect 8846 31260 8852 31272
rect 8807 31232 8852 31260
rect 8846 31220 8852 31232
rect 8904 31220 8910 31272
rect 9048 31260 9076 31291
rect 10428 31269 10456 31436
rect 13538 31424 13544 31436
rect 13596 31424 13602 31476
rect 10594 31328 10600 31340
rect 10555 31300 10600 31328
rect 10594 31288 10600 31300
rect 10652 31328 10658 31340
rect 11057 31331 11115 31337
rect 11057 31328 11069 31331
rect 10652 31300 11069 31328
rect 10652 31288 10658 31300
rect 11057 31297 11069 31300
rect 11103 31297 11115 31331
rect 11057 31291 11115 31297
rect 8956 31232 9076 31260
rect 10413 31263 10471 31269
rect 8956 31192 8984 31232
rect 10413 31229 10425 31263
rect 10459 31229 10471 31263
rect 10413 31223 10471 31229
rect 13357 31263 13415 31269
rect 13357 31229 13369 31263
rect 13403 31260 13415 31263
rect 13446 31260 13452 31272
rect 13403 31232 13452 31260
rect 13403 31229 13415 31232
rect 13357 31223 13415 31229
rect 13446 31220 13452 31232
rect 13504 31260 13510 31272
rect 13817 31263 13875 31269
rect 13817 31260 13829 31263
rect 13504 31232 13829 31260
rect 13504 31220 13510 31232
rect 13817 31229 13829 31232
rect 13863 31229 13875 31263
rect 13817 31223 13875 31229
rect 8312 31164 8984 31192
rect 5537 31155 5595 31161
rect 2866 31084 2872 31136
rect 2924 31124 2930 31136
rect 2961 31127 3019 31133
rect 2961 31124 2973 31127
rect 2924 31096 2973 31124
rect 2924 31084 2930 31096
rect 2961 31093 2973 31096
rect 3007 31093 3019 31127
rect 3326 31124 3332 31136
rect 3287 31096 3332 31124
rect 2961 31087 3019 31093
rect 3326 31084 3332 31096
rect 3384 31084 3390 31136
rect 3421 31127 3479 31133
rect 3421 31093 3433 31127
rect 3467 31124 3479 31127
rect 3510 31124 3516 31136
rect 3467 31096 3516 31124
rect 3467 31093 3479 31096
rect 3421 31087 3479 31093
rect 3510 31084 3516 31096
rect 3568 31124 3574 31136
rect 4525 31127 4583 31133
rect 4525 31124 4537 31127
rect 3568 31096 4537 31124
rect 3568 31084 3574 31096
rect 4525 31093 4537 31096
rect 4571 31093 4583 31127
rect 4890 31124 4896 31136
rect 4851 31096 4896 31124
rect 4525 31087 4583 31093
rect 4890 31084 4896 31096
rect 4948 31084 4954 31136
rect 4982 31084 4988 31136
rect 5040 31124 5046 31136
rect 6638 31124 6644 31136
rect 5040 31096 5085 31124
rect 6599 31096 6644 31124
rect 5040 31084 5046 31096
rect 6638 31084 6644 31096
rect 6696 31084 6702 31136
rect 7282 31124 7288 31136
rect 7243 31096 7288 31124
rect 7282 31084 7288 31096
rect 7340 31084 7346 31136
rect 7374 31084 7380 31136
rect 7432 31124 7438 31136
rect 7742 31124 7748 31136
rect 7432 31096 7748 31124
rect 7432 31084 7438 31096
rect 7742 31084 7748 31096
rect 7800 31084 7806 31136
rect 8478 31084 8484 31136
rect 8536 31124 8542 31136
rect 9493 31127 9551 31133
rect 9493 31124 9505 31127
rect 8536 31096 9505 31124
rect 8536 31084 8542 31096
rect 9493 31093 9505 31096
rect 9539 31124 9551 31127
rect 9766 31124 9772 31136
rect 9539 31096 9772 31124
rect 9539 31093 9551 31096
rect 9493 31087 9551 31093
rect 9766 31084 9772 31096
rect 9824 31084 9830 31136
rect 10502 31124 10508 31136
rect 10463 31096 10508 31124
rect 10502 31084 10508 31096
rect 10560 31084 10566 31136
rect 1104 31034 14812 31056
rect 1104 30982 6315 31034
rect 6367 30982 6379 31034
rect 6431 30982 6443 31034
rect 6495 30982 6507 31034
rect 6559 30982 11648 31034
rect 11700 30982 11712 31034
rect 11764 30982 11776 31034
rect 11828 30982 11840 31034
rect 11892 30982 14812 31034
rect 1104 30960 14812 30982
rect 3326 30880 3332 30932
rect 3384 30920 3390 30932
rect 4065 30923 4123 30929
rect 4065 30920 4077 30923
rect 3384 30892 4077 30920
rect 3384 30880 3390 30892
rect 4065 30889 4077 30892
rect 4111 30889 4123 30923
rect 6822 30920 6828 30932
rect 6783 30892 6828 30920
rect 4065 30883 4123 30889
rect 6822 30880 6828 30892
rect 6880 30880 6886 30932
rect 7558 30920 7564 30932
rect 7519 30892 7564 30920
rect 7558 30880 7564 30892
rect 7616 30880 7622 30932
rect 8570 30920 8576 30932
rect 8531 30892 8576 30920
rect 8570 30880 8576 30892
rect 8628 30880 8634 30932
rect 10042 30880 10048 30932
rect 10100 30920 10106 30932
rect 10413 30923 10471 30929
rect 10413 30920 10425 30923
rect 10100 30892 10425 30920
rect 10100 30880 10106 30892
rect 10413 30889 10425 30892
rect 10459 30889 10471 30923
rect 10413 30883 10471 30889
rect 10594 30880 10600 30932
rect 10652 30920 10658 30932
rect 10781 30923 10839 30929
rect 10781 30920 10793 30923
rect 10652 30892 10793 30920
rect 10652 30880 10658 30892
rect 10781 30889 10793 30892
rect 10827 30889 10839 30923
rect 10781 30883 10839 30889
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 12989 30923 13047 30929
rect 12989 30920 13001 30923
rect 12492 30892 13001 30920
rect 12492 30880 12498 30892
rect 12989 30889 13001 30892
rect 13035 30889 13047 30923
rect 12989 30883 13047 30889
rect 3234 30812 3240 30864
rect 3292 30852 3298 30864
rect 3789 30855 3847 30861
rect 3789 30852 3801 30855
rect 3292 30824 3801 30852
rect 3292 30812 3298 30824
rect 3789 30821 3801 30824
rect 3835 30852 3847 30855
rect 4890 30852 4896 30864
rect 3835 30824 4896 30852
rect 3835 30821 3847 30824
rect 3789 30815 3847 30821
rect 4890 30812 4896 30824
rect 4948 30812 4954 30864
rect 11876 30855 11934 30861
rect 11876 30821 11888 30855
rect 11922 30852 11934 30855
rect 12066 30852 12072 30864
rect 11922 30824 12072 30852
rect 11922 30821 11934 30824
rect 11876 30815 11934 30821
rect 12066 30812 12072 30824
rect 12124 30812 12130 30864
rect 4430 30784 4436 30796
rect 4391 30756 4436 30784
rect 4430 30744 4436 30756
rect 4488 30744 4494 30796
rect 6178 30744 6184 30796
rect 6236 30784 6242 30796
rect 6917 30787 6975 30793
rect 6917 30784 6929 30787
rect 6236 30756 6929 30784
rect 6236 30744 6242 30756
rect 6917 30753 6929 30756
rect 6963 30753 6975 30787
rect 6917 30747 6975 30753
rect 7098 30744 7104 30796
rect 7156 30744 7162 30796
rect 11054 30744 11060 30796
rect 11112 30784 11118 30796
rect 11606 30784 11612 30796
rect 11112 30756 11612 30784
rect 11112 30744 11118 30756
rect 11606 30744 11612 30756
rect 11664 30744 11670 30796
rect 2961 30719 3019 30725
rect 2961 30685 2973 30719
rect 3007 30716 3019 30719
rect 4154 30716 4160 30728
rect 3007 30688 4160 30716
rect 3007 30685 3019 30688
rect 2961 30679 3019 30685
rect 4154 30676 4160 30688
rect 4212 30676 4218 30728
rect 4522 30716 4528 30728
rect 4483 30688 4528 30716
rect 4522 30676 4528 30688
rect 4580 30676 4586 30728
rect 4706 30716 4712 30728
rect 4667 30688 4712 30716
rect 4706 30676 4712 30688
rect 4764 30716 4770 30728
rect 5074 30716 5080 30728
rect 4764 30688 5080 30716
rect 4764 30676 4770 30688
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 6822 30676 6828 30728
rect 6880 30716 6886 30728
rect 7009 30719 7067 30725
rect 7009 30716 7021 30719
rect 6880 30688 7021 30716
rect 6880 30676 6886 30688
rect 7009 30685 7021 30688
rect 7055 30716 7067 30719
rect 7116 30716 7144 30744
rect 7055 30688 7144 30716
rect 7055 30685 7067 30688
rect 7009 30679 7067 30685
rect 6365 30651 6423 30657
rect 6365 30617 6377 30651
rect 6411 30648 6423 30651
rect 7282 30648 7288 30660
rect 6411 30620 7288 30648
rect 6411 30617 6423 30620
rect 6365 30611 6423 30617
rect 7282 30608 7288 30620
rect 7340 30608 7346 30660
rect 6457 30583 6515 30589
rect 6457 30549 6469 30583
rect 6503 30580 6515 30583
rect 6914 30580 6920 30592
rect 6503 30552 6920 30580
rect 6503 30549 6515 30552
rect 6457 30543 6515 30549
rect 6914 30540 6920 30552
rect 6972 30540 6978 30592
rect 9766 30540 9772 30592
rect 9824 30580 9830 30592
rect 10045 30583 10103 30589
rect 10045 30580 10057 30583
rect 9824 30552 10057 30580
rect 9824 30540 9830 30552
rect 10045 30549 10057 30552
rect 10091 30580 10103 30583
rect 10502 30580 10508 30592
rect 10091 30552 10508 30580
rect 10091 30549 10103 30552
rect 10045 30543 10103 30549
rect 10502 30540 10508 30552
rect 10560 30540 10566 30592
rect 1104 30490 14812 30512
rect 1104 30438 3648 30490
rect 3700 30438 3712 30490
rect 3764 30438 3776 30490
rect 3828 30438 3840 30490
rect 3892 30438 8982 30490
rect 9034 30438 9046 30490
rect 9098 30438 9110 30490
rect 9162 30438 9174 30490
rect 9226 30438 14315 30490
rect 14367 30438 14379 30490
rect 14431 30438 14443 30490
rect 14495 30438 14507 30490
rect 14559 30438 14812 30490
rect 1104 30416 14812 30438
rect 3789 30379 3847 30385
rect 3789 30345 3801 30379
rect 3835 30376 3847 30379
rect 3970 30376 3976 30388
rect 3835 30348 3976 30376
rect 3835 30345 3847 30348
rect 3789 30339 3847 30345
rect 3970 30336 3976 30348
rect 4028 30376 4034 30388
rect 4706 30376 4712 30388
rect 4028 30348 4712 30376
rect 4028 30336 4034 30348
rect 4706 30336 4712 30348
rect 4764 30336 4770 30388
rect 5905 30379 5963 30385
rect 5905 30345 5917 30379
rect 5951 30376 5963 30379
rect 6822 30376 6828 30388
rect 5951 30348 6828 30376
rect 5951 30345 5963 30348
rect 5905 30339 5963 30345
rect 6822 30336 6828 30348
rect 6880 30336 6886 30388
rect 11606 30376 11612 30388
rect 11567 30348 11612 30376
rect 11606 30336 11612 30348
rect 11664 30336 11670 30388
rect 12066 30376 12072 30388
rect 12027 30348 12072 30376
rect 12066 30336 12072 30348
rect 12124 30336 12130 30388
rect 3421 30311 3479 30317
rect 3421 30277 3433 30311
rect 3467 30308 3479 30311
rect 4430 30308 4436 30320
rect 3467 30280 4436 30308
rect 3467 30277 3479 30280
rect 3421 30271 3479 30277
rect 4430 30268 4436 30280
rect 4488 30308 4494 30320
rect 4617 30311 4675 30317
rect 4617 30308 4629 30311
rect 4488 30280 4629 30308
rect 4488 30268 4494 30280
rect 4617 30277 4629 30280
rect 4663 30277 4675 30311
rect 4617 30271 4675 30277
rect 4062 30200 4068 30252
rect 4120 30240 4126 30252
rect 4157 30243 4215 30249
rect 4157 30240 4169 30243
rect 4120 30212 4169 30240
rect 4120 30200 4126 30212
rect 4157 30209 4169 30212
rect 4203 30240 4215 30243
rect 4798 30240 4804 30252
rect 4203 30212 4804 30240
rect 4203 30209 4215 30212
rect 4157 30203 4215 30209
rect 4798 30200 4804 30212
rect 4856 30240 4862 30252
rect 5169 30243 5227 30249
rect 5169 30240 5181 30243
rect 4856 30212 5181 30240
rect 4856 30200 4862 30212
rect 5169 30209 5181 30212
rect 5215 30209 5227 30243
rect 5169 30203 5227 30209
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7285 30243 7343 30249
rect 7285 30240 7297 30243
rect 6972 30212 7297 30240
rect 6972 30200 6978 30212
rect 7285 30209 7297 30212
rect 7331 30209 7343 30243
rect 7466 30240 7472 30252
rect 7427 30212 7472 30240
rect 7285 30203 7343 30209
rect 5810 30132 5816 30184
rect 5868 30172 5874 30184
rect 7300 30172 7328 30203
rect 7466 30200 7472 30212
rect 7524 30200 7530 30252
rect 10226 30240 10232 30252
rect 10187 30212 10232 30240
rect 10226 30200 10232 30212
rect 10284 30200 10290 30252
rect 7837 30175 7895 30181
rect 7837 30172 7849 30175
rect 5868 30144 6684 30172
rect 7300 30144 7849 30172
rect 5868 30132 5874 30144
rect 4154 30064 4160 30116
rect 4212 30104 4218 30116
rect 4985 30107 5043 30113
rect 4985 30104 4997 30107
rect 4212 30076 4997 30104
rect 4212 30064 4218 30076
rect 4985 30073 4997 30076
rect 5031 30073 5043 30107
rect 6178 30104 6184 30116
rect 6139 30076 6184 30104
rect 4985 30067 5043 30073
rect 6178 30064 6184 30076
rect 6236 30064 6242 30116
rect 6656 30113 6684 30144
rect 7837 30141 7849 30144
rect 7883 30141 7895 30175
rect 7837 30135 7895 30141
rect 8110 30132 8116 30184
rect 8168 30172 8174 30184
rect 9217 30175 9275 30181
rect 9217 30172 9229 30175
rect 8168 30144 9229 30172
rect 8168 30132 8174 30144
rect 9217 30141 9229 30144
rect 9263 30172 9275 30175
rect 9950 30172 9956 30184
rect 9263 30144 9956 30172
rect 9263 30141 9275 30144
rect 9217 30135 9275 30141
rect 9950 30132 9956 30144
rect 10008 30172 10014 30184
rect 10045 30175 10103 30181
rect 10045 30172 10057 30175
rect 10008 30144 10057 30172
rect 10008 30132 10014 30144
rect 10045 30141 10057 30144
rect 10091 30141 10103 30175
rect 10045 30135 10103 30141
rect 6641 30107 6699 30113
rect 6641 30073 6653 30107
rect 6687 30104 6699 30107
rect 6687 30076 7236 30104
rect 6687 30073 6699 30076
rect 6641 30067 6699 30073
rect 7208 30048 7236 30076
rect 8846 30064 8852 30116
rect 8904 30104 8910 30116
rect 9493 30107 9551 30113
rect 9493 30104 9505 30107
rect 8904 30076 9505 30104
rect 8904 30064 8910 30076
rect 9493 30073 9505 30076
rect 9539 30104 9551 30107
rect 10137 30107 10195 30113
rect 10137 30104 10149 30107
rect 9539 30076 10149 30104
rect 9539 30073 9551 30076
rect 9493 30067 9551 30073
rect 10137 30073 10149 30076
rect 10183 30073 10195 30107
rect 10137 30067 10195 30073
rect 4525 30039 4583 30045
rect 4525 30005 4537 30039
rect 4571 30036 4583 30039
rect 5074 30036 5080 30048
rect 4571 30008 5080 30036
rect 4571 30005 4583 30008
rect 4525 29999 4583 30005
rect 5074 29996 5080 30008
rect 5132 29996 5138 30048
rect 6822 30036 6828 30048
rect 6783 30008 6828 30036
rect 6822 29996 6828 30008
rect 6880 29996 6886 30048
rect 7190 30036 7196 30048
rect 7151 30008 7196 30036
rect 7190 29996 7196 30008
rect 7248 29996 7254 30048
rect 9674 30036 9680 30048
rect 9635 30008 9680 30036
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 1104 29946 14812 29968
rect 1104 29894 6315 29946
rect 6367 29894 6379 29946
rect 6431 29894 6443 29946
rect 6495 29894 6507 29946
rect 6559 29894 11648 29946
rect 11700 29894 11712 29946
rect 11764 29894 11776 29946
rect 11828 29894 11840 29946
rect 11892 29894 14812 29946
rect 1104 29872 14812 29894
rect 1578 29832 1584 29844
rect 1539 29804 1584 29832
rect 1578 29792 1584 29804
rect 1636 29792 1642 29844
rect 4341 29835 4399 29841
rect 4341 29801 4353 29835
rect 4387 29832 4399 29835
rect 4522 29832 4528 29844
rect 4387 29804 4528 29832
rect 4387 29801 4399 29804
rect 4341 29795 4399 29801
rect 4522 29792 4528 29804
rect 4580 29792 4586 29844
rect 5718 29832 5724 29844
rect 5679 29804 5724 29832
rect 5718 29792 5724 29804
rect 5776 29792 5782 29844
rect 6549 29835 6607 29841
rect 6549 29801 6561 29835
rect 6595 29832 6607 29835
rect 6730 29832 6736 29844
rect 6595 29804 6736 29832
rect 6595 29801 6607 29804
rect 6549 29795 6607 29801
rect 6730 29792 6736 29804
rect 6788 29792 6794 29844
rect 7282 29792 7288 29844
rect 7340 29832 7346 29844
rect 7653 29835 7711 29841
rect 7653 29832 7665 29835
rect 7340 29804 7665 29832
rect 7340 29792 7346 29804
rect 7653 29801 7665 29804
rect 7699 29801 7711 29835
rect 7653 29795 7711 29801
rect 8018 29792 8024 29844
rect 8076 29792 8082 29844
rect 9953 29835 10011 29841
rect 9953 29801 9965 29835
rect 9999 29832 10011 29835
rect 10226 29832 10232 29844
rect 9999 29804 10232 29832
rect 9999 29801 10011 29804
rect 9953 29795 10011 29801
rect 10226 29792 10232 29804
rect 10284 29832 10290 29844
rect 10284 29804 11100 29832
rect 10284 29792 10290 29804
rect 4154 29724 4160 29776
rect 4212 29764 4218 29776
rect 4617 29767 4675 29773
rect 4617 29764 4629 29767
rect 4212 29736 4629 29764
rect 4212 29724 4218 29736
rect 4617 29733 4629 29736
rect 4663 29733 4675 29767
rect 4617 29727 4675 29733
rect 6917 29767 6975 29773
rect 6917 29733 6929 29767
rect 6963 29764 6975 29767
rect 7466 29764 7472 29776
rect 6963 29736 7472 29764
rect 6963 29733 6975 29736
rect 6917 29727 6975 29733
rect 7466 29724 7472 29736
rect 7524 29724 7530 29776
rect 7561 29767 7619 29773
rect 7561 29733 7573 29767
rect 7607 29764 7619 29767
rect 8036 29764 8064 29792
rect 10962 29764 10968 29776
rect 7607 29736 8248 29764
rect 7607 29733 7619 29736
rect 7561 29727 7619 29733
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29696 1455 29699
rect 2314 29696 2320 29708
rect 1443 29668 2320 29696
rect 1443 29665 1455 29668
rect 1397 29659 1455 29665
rect 2314 29656 2320 29668
rect 2372 29656 2378 29708
rect 5629 29699 5687 29705
rect 5629 29665 5641 29699
rect 5675 29696 5687 29699
rect 6822 29696 6828 29708
rect 5675 29668 6828 29696
rect 5675 29665 5687 29668
rect 5629 29659 5687 29665
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 8018 29696 8024 29708
rect 7979 29668 8024 29696
rect 8018 29656 8024 29668
rect 8076 29656 8082 29708
rect 8220 29640 8248 29736
rect 10336 29736 10968 29764
rect 5810 29628 5816 29640
rect 5771 29600 5816 29628
rect 5810 29588 5816 29600
rect 5868 29588 5874 29640
rect 8113 29631 8171 29637
rect 8113 29597 8125 29631
rect 8159 29597 8171 29631
rect 8113 29591 8171 29597
rect 5258 29492 5264 29504
rect 5219 29464 5264 29492
rect 5258 29452 5264 29464
rect 5316 29452 5322 29504
rect 8128 29492 8156 29591
rect 8202 29588 8208 29640
rect 8260 29628 8266 29640
rect 10336 29637 10364 29736
rect 10962 29724 10968 29736
rect 11020 29724 11026 29776
rect 11072 29708 11100 29804
rect 10588 29699 10646 29705
rect 10588 29665 10600 29699
rect 10634 29696 10646 29699
rect 11054 29696 11060 29708
rect 10634 29668 11060 29696
rect 10634 29665 10646 29668
rect 10588 29659 10646 29665
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 10321 29631 10379 29637
rect 8260 29600 8305 29628
rect 8260 29588 8266 29600
rect 10321 29597 10333 29631
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 8757 29495 8815 29501
rect 8757 29492 8769 29495
rect 8128 29464 8769 29492
rect 8757 29461 8769 29464
rect 8803 29492 8815 29495
rect 9582 29492 9588 29504
rect 8803 29464 9588 29492
rect 8803 29461 8815 29464
rect 8757 29455 8815 29461
rect 9582 29452 9588 29464
rect 9640 29452 9646 29504
rect 10226 29452 10232 29504
rect 10284 29492 10290 29504
rect 11701 29495 11759 29501
rect 11701 29492 11713 29495
rect 10284 29464 11713 29492
rect 10284 29452 10290 29464
rect 11701 29461 11713 29464
rect 11747 29461 11759 29495
rect 11701 29455 11759 29461
rect 1104 29402 14812 29424
rect 1104 29350 3648 29402
rect 3700 29350 3712 29402
rect 3764 29350 3776 29402
rect 3828 29350 3840 29402
rect 3892 29350 8982 29402
rect 9034 29350 9046 29402
rect 9098 29350 9110 29402
rect 9162 29350 9174 29402
rect 9226 29350 14315 29402
rect 14367 29350 14379 29402
rect 14431 29350 14443 29402
rect 14495 29350 14507 29402
rect 14559 29350 14812 29402
rect 1104 29328 14812 29350
rect 1578 29288 1584 29300
rect 1539 29260 1584 29288
rect 1578 29248 1584 29260
rect 1636 29248 1642 29300
rect 1949 29291 2007 29297
rect 1949 29257 1961 29291
rect 1995 29288 2007 29291
rect 2682 29288 2688 29300
rect 1995 29260 2688 29288
rect 1995 29257 2007 29260
rect 1949 29251 2007 29257
rect 1397 29087 1455 29093
rect 1397 29053 1409 29087
rect 1443 29084 1455 29087
rect 1964 29084 1992 29251
rect 2682 29248 2688 29260
rect 2740 29248 2746 29300
rect 4062 29288 4068 29300
rect 4023 29260 4068 29288
rect 4062 29248 4068 29260
rect 4120 29248 4126 29300
rect 4522 29248 4528 29300
rect 4580 29288 4586 29300
rect 4617 29291 4675 29297
rect 4617 29288 4629 29291
rect 4580 29260 4629 29288
rect 4580 29248 4586 29260
rect 4617 29257 4629 29260
rect 4663 29257 4675 29291
rect 4617 29251 4675 29257
rect 5718 29248 5724 29300
rect 5776 29288 5782 29300
rect 5997 29291 6055 29297
rect 5997 29288 6009 29291
rect 5776 29260 6009 29288
rect 5776 29248 5782 29260
rect 5997 29257 6009 29260
rect 6043 29257 6055 29291
rect 5997 29251 6055 29257
rect 6457 29291 6515 29297
rect 6457 29257 6469 29291
rect 6503 29288 6515 29291
rect 6822 29288 6828 29300
rect 6503 29260 6828 29288
rect 6503 29257 6515 29260
rect 6457 29251 6515 29257
rect 6822 29248 6828 29260
rect 6880 29248 6886 29300
rect 10689 29291 10747 29297
rect 10689 29257 10701 29291
rect 10735 29288 10747 29291
rect 10962 29288 10968 29300
rect 10735 29260 10968 29288
rect 10735 29257 10747 29260
rect 10689 29251 10747 29257
rect 10962 29248 10968 29260
rect 11020 29248 11026 29300
rect 4080 29152 4108 29248
rect 8021 29223 8079 29229
rect 8021 29189 8033 29223
rect 8067 29220 8079 29223
rect 8110 29220 8116 29232
rect 8067 29192 8116 29220
rect 8067 29189 8079 29192
rect 8021 29183 8079 29189
rect 8110 29180 8116 29192
rect 8168 29180 8174 29232
rect 5074 29152 5080 29164
rect 4080 29124 5080 29152
rect 5074 29112 5080 29124
rect 5132 29152 5138 29164
rect 5169 29155 5227 29161
rect 5169 29152 5181 29155
rect 5132 29124 5181 29152
rect 5132 29112 5138 29124
rect 5169 29121 5181 29124
rect 5215 29121 5227 29155
rect 5169 29115 5227 29121
rect 5721 29155 5779 29161
rect 5721 29121 5733 29155
rect 5767 29152 5779 29155
rect 5810 29152 5816 29164
rect 5767 29124 5816 29152
rect 5767 29121 5779 29124
rect 5721 29115 5779 29121
rect 5810 29112 5816 29124
rect 5868 29112 5874 29164
rect 8665 29155 8723 29161
rect 8665 29121 8677 29155
rect 8711 29152 8723 29155
rect 9030 29152 9036 29164
rect 8711 29124 9036 29152
rect 8711 29121 8723 29124
rect 8665 29115 8723 29121
rect 9030 29112 9036 29124
rect 9088 29112 9094 29164
rect 9674 29112 9680 29164
rect 9732 29152 9738 29164
rect 10042 29152 10048 29164
rect 9732 29124 10048 29152
rect 9732 29112 9738 29124
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 10226 29152 10232 29164
rect 10187 29124 10232 29152
rect 10226 29112 10232 29124
rect 10284 29112 10290 29164
rect 7282 29084 7288 29096
rect 1443 29056 1992 29084
rect 7243 29056 7288 29084
rect 1443 29053 1455 29056
rect 1397 29047 1455 29053
rect 7282 29044 7288 29056
rect 7340 29084 7346 29096
rect 7834 29084 7840 29096
rect 7340 29056 7840 29084
rect 7340 29044 7346 29056
rect 7834 29044 7840 29056
rect 7892 29084 7898 29096
rect 8481 29087 8539 29093
rect 8481 29084 8493 29087
rect 7892 29056 8493 29084
rect 7892 29044 7898 29056
rect 8481 29053 8493 29056
rect 8527 29084 8539 29087
rect 9401 29087 9459 29093
rect 9401 29084 9413 29087
rect 8527 29056 9413 29084
rect 8527 29053 8539 29056
rect 8481 29047 8539 29053
rect 9401 29053 9413 29056
rect 9447 29084 9459 29087
rect 9953 29087 10011 29093
rect 9953 29084 9965 29087
rect 9447 29056 9965 29084
rect 9447 29053 9459 29056
rect 9401 29047 9459 29053
rect 9953 29053 9965 29056
rect 9999 29053 10011 29087
rect 9953 29047 10011 29053
rect 11146 29044 11152 29096
rect 11204 29084 11210 29096
rect 11204 29056 12020 29084
rect 11204 29044 11210 29056
rect 11992 29028 12020 29056
rect 2314 29016 2320 29028
rect 2275 28988 2320 29016
rect 2314 28976 2320 28988
rect 2372 28976 2378 29028
rect 4525 29019 4583 29025
rect 4525 28985 4537 29019
rect 4571 29016 4583 29019
rect 4985 29019 5043 29025
rect 4985 29016 4997 29019
rect 4571 28988 4997 29016
rect 4571 28985 4583 28988
rect 4525 28979 4583 28985
rect 4985 28985 4997 28988
rect 5031 29016 5043 29019
rect 5994 29016 6000 29028
rect 5031 28988 6000 29016
rect 5031 28985 5043 28988
rect 4985 28979 5043 28985
rect 5994 28976 6000 28988
rect 6052 28976 6058 29028
rect 7006 28976 7012 29028
rect 7064 29016 7070 29028
rect 7653 29019 7711 29025
rect 7653 29016 7665 29019
rect 7064 28988 7665 29016
rect 7064 28976 7070 28988
rect 7653 28985 7665 28988
rect 7699 29016 7711 29019
rect 8018 29016 8024 29028
rect 7699 28988 8024 29016
rect 7699 28985 7711 28988
rect 7653 28979 7711 28985
rect 8018 28976 8024 28988
rect 8076 28976 8082 29028
rect 8389 29019 8447 29025
rect 8389 28985 8401 29019
rect 8435 29016 8447 29019
rect 8570 29016 8576 29028
rect 8435 28988 8576 29016
rect 8435 28985 8447 28988
rect 8389 28979 8447 28985
rect 8570 28976 8576 28988
rect 8628 28976 8634 29028
rect 11974 28976 11980 29028
rect 12032 28976 12038 29028
rect 4246 28908 4252 28960
rect 4304 28948 4310 28960
rect 5077 28951 5135 28957
rect 5077 28948 5089 28951
rect 4304 28920 5089 28948
rect 4304 28908 4310 28920
rect 5077 28917 5089 28920
rect 5123 28917 5135 28951
rect 5077 28911 5135 28917
rect 5166 28908 5172 28960
rect 5224 28948 5230 28960
rect 5350 28948 5356 28960
rect 5224 28920 5356 28948
rect 5224 28908 5230 28920
rect 5350 28908 5356 28920
rect 5408 28908 5414 28960
rect 9030 28948 9036 28960
rect 8991 28920 9036 28948
rect 9030 28908 9036 28920
rect 9088 28908 9094 28960
rect 9582 28948 9588 28960
rect 9543 28920 9588 28948
rect 9582 28908 9588 28920
rect 9640 28908 9646 28960
rect 11054 28948 11060 28960
rect 10967 28920 11060 28948
rect 11054 28908 11060 28920
rect 11112 28948 11118 28960
rect 12526 28948 12532 28960
rect 11112 28920 12532 28948
rect 11112 28908 11118 28920
rect 12526 28908 12532 28920
rect 12584 28908 12590 28960
rect 1104 28858 14812 28880
rect 1104 28806 6315 28858
rect 6367 28806 6379 28858
rect 6431 28806 6443 28858
rect 6495 28806 6507 28858
rect 6559 28806 11648 28858
rect 11700 28806 11712 28858
rect 11764 28806 11776 28858
rect 11828 28806 11840 28858
rect 11892 28806 14812 28858
rect 1104 28784 14812 28806
rect 2406 28744 2412 28756
rect 2367 28716 2412 28744
rect 2406 28704 2412 28716
rect 2464 28704 2470 28756
rect 4890 28744 4896 28756
rect 4851 28716 4896 28744
rect 4890 28704 4896 28716
rect 4948 28704 4954 28756
rect 10042 28704 10048 28756
rect 10100 28744 10106 28756
rect 10229 28747 10287 28753
rect 10229 28744 10241 28747
rect 10100 28716 10241 28744
rect 10100 28704 10106 28716
rect 10229 28713 10241 28716
rect 10275 28713 10287 28747
rect 10229 28707 10287 28713
rect 1670 28636 1676 28688
rect 1728 28676 1734 28688
rect 2590 28676 2596 28688
rect 1728 28648 2596 28676
rect 1728 28636 1734 28648
rect 2590 28636 2596 28648
rect 2648 28676 2654 28688
rect 2777 28679 2835 28685
rect 2777 28676 2789 28679
rect 2648 28648 2789 28676
rect 2648 28636 2654 28648
rect 2777 28645 2789 28648
rect 2823 28645 2835 28679
rect 6086 28676 6092 28688
rect 2777 28639 2835 28645
rect 5276 28648 6092 28676
rect 5276 28617 5304 28648
rect 6086 28636 6092 28648
rect 6144 28636 6150 28688
rect 11416 28679 11474 28685
rect 11416 28645 11428 28679
rect 11462 28676 11474 28679
rect 12342 28676 12348 28688
rect 11462 28648 12348 28676
rect 11462 28645 11474 28648
rect 11416 28639 11474 28645
rect 12342 28636 12348 28648
rect 12400 28636 12406 28688
rect 5261 28611 5319 28617
rect 5261 28577 5273 28611
rect 5307 28577 5319 28611
rect 6805 28611 6863 28617
rect 6805 28608 6817 28611
rect 5261 28571 5319 28577
rect 5552 28580 6817 28608
rect 5552 28552 5580 28580
rect 6805 28577 6817 28580
rect 6851 28608 6863 28611
rect 7282 28608 7288 28620
rect 6851 28580 7288 28608
rect 6851 28577 6863 28580
rect 6805 28571 6863 28577
rect 7282 28568 7288 28580
rect 7340 28568 7346 28620
rect 9953 28611 10011 28617
rect 9953 28577 9965 28611
rect 9999 28608 10011 28611
rect 10226 28608 10232 28620
rect 9999 28580 10232 28608
rect 9999 28577 10011 28580
rect 9953 28571 10011 28577
rect 10226 28568 10232 28580
rect 10284 28568 10290 28620
rect 2866 28540 2872 28552
rect 2827 28512 2872 28540
rect 2866 28500 2872 28512
rect 2924 28500 2930 28552
rect 2958 28500 2964 28552
rect 3016 28540 3022 28552
rect 3053 28543 3111 28549
rect 3053 28540 3065 28543
rect 3016 28512 3065 28540
rect 3016 28500 3022 28512
rect 3053 28509 3065 28512
rect 3099 28540 3111 28543
rect 5074 28540 5080 28552
rect 3099 28512 5080 28540
rect 3099 28509 3111 28512
rect 3053 28503 3111 28509
rect 5074 28500 5080 28512
rect 5132 28500 5138 28552
rect 5350 28540 5356 28552
rect 5311 28512 5356 28540
rect 5350 28500 5356 28512
rect 5408 28500 5414 28552
rect 5534 28540 5540 28552
rect 5495 28512 5540 28540
rect 5534 28500 5540 28512
rect 5592 28500 5598 28552
rect 6546 28540 6552 28552
rect 6507 28512 6552 28540
rect 6546 28500 6552 28512
rect 6604 28500 6610 28552
rect 10962 28500 10968 28552
rect 11020 28540 11026 28552
rect 11149 28543 11207 28549
rect 11149 28540 11161 28543
rect 11020 28512 11161 28540
rect 11020 28500 11026 28512
rect 11149 28509 11161 28512
rect 11195 28509 11207 28543
rect 11149 28503 11207 28509
rect 7929 28475 7987 28481
rect 7929 28441 7941 28475
rect 7975 28472 7987 28475
rect 8386 28472 8392 28484
rect 7975 28444 8392 28472
rect 7975 28441 7987 28444
rect 7929 28435 7987 28441
rect 8386 28432 8392 28444
rect 8444 28472 8450 28484
rect 8941 28475 8999 28481
rect 8941 28472 8953 28475
rect 8444 28444 8953 28472
rect 8444 28432 8450 28444
rect 8941 28441 8953 28444
rect 8987 28472 8999 28475
rect 9030 28472 9036 28484
rect 8987 28444 9036 28472
rect 8987 28441 8999 28444
rect 8941 28435 8999 28441
rect 9030 28432 9036 28444
rect 9088 28472 9094 28484
rect 12526 28472 12532 28484
rect 9088 28444 10732 28472
rect 12487 28444 12532 28472
rect 9088 28432 9094 28444
rect 10704 28416 10732 28444
rect 12526 28432 12532 28444
rect 12584 28432 12590 28484
rect 4246 28364 4252 28416
rect 4304 28404 4310 28416
rect 4617 28407 4675 28413
rect 4617 28404 4629 28407
rect 4304 28376 4629 28404
rect 4304 28364 4310 28376
rect 4617 28373 4629 28376
rect 4663 28373 4675 28407
rect 8570 28404 8576 28416
rect 8531 28376 8576 28404
rect 4617 28367 4675 28373
rect 8570 28364 8576 28376
rect 8628 28364 8634 28416
rect 10686 28404 10692 28416
rect 10647 28376 10692 28404
rect 10686 28364 10692 28376
rect 10744 28364 10750 28416
rect 1104 28314 14812 28336
rect 1104 28262 3648 28314
rect 3700 28262 3712 28314
rect 3764 28262 3776 28314
rect 3828 28262 3840 28314
rect 3892 28262 8982 28314
rect 9034 28262 9046 28314
rect 9098 28262 9110 28314
rect 9162 28262 9174 28314
rect 9226 28262 14315 28314
rect 14367 28262 14379 28314
rect 14431 28262 14443 28314
rect 14495 28262 14507 28314
rect 14559 28262 14812 28314
rect 1104 28240 14812 28262
rect 2501 28203 2559 28209
rect 2501 28169 2513 28203
rect 2547 28200 2559 28203
rect 2590 28200 2596 28212
rect 2547 28172 2596 28200
rect 2547 28169 2559 28172
rect 2501 28163 2559 28169
rect 2590 28160 2596 28172
rect 2648 28160 2654 28212
rect 2866 28160 2872 28212
rect 2924 28200 2930 28212
rect 3145 28203 3203 28209
rect 3145 28200 3157 28203
rect 2924 28172 3157 28200
rect 2924 28160 2930 28172
rect 3145 28169 3157 28172
rect 3191 28169 3203 28203
rect 5074 28200 5080 28212
rect 5035 28172 5080 28200
rect 3145 28163 3203 28169
rect 5074 28160 5080 28172
rect 5132 28160 5138 28212
rect 5534 28160 5540 28212
rect 5592 28200 5598 28212
rect 5629 28203 5687 28209
rect 5629 28200 5641 28203
rect 5592 28172 5641 28200
rect 5592 28160 5598 28172
rect 5629 28169 5641 28172
rect 5675 28169 5687 28203
rect 7282 28200 7288 28212
rect 7243 28172 7288 28200
rect 5629 28163 5687 28169
rect 7282 28160 7288 28172
rect 7340 28160 7346 28212
rect 9674 28160 9680 28212
rect 9732 28200 9738 28212
rect 10597 28203 10655 28209
rect 10597 28200 10609 28203
rect 9732 28172 10609 28200
rect 9732 28160 9738 28172
rect 10597 28169 10609 28172
rect 10643 28169 10655 28203
rect 10597 28163 10655 28169
rect 12069 28203 12127 28209
rect 12069 28169 12081 28203
rect 12115 28200 12127 28203
rect 12342 28200 12348 28212
rect 12115 28172 12348 28200
rect 12115 28169 12127 28172
rect 12069 28163 12127 28169
rect 12342 28160 12348 28172
rect 12400 28160 12406 28212
rect 2869 28067 2927 28073
rect 2869 28033 2881 28067
rect 2915 28064 2927 28067
rect 2958 28064 2964 28076
rect 2915 28036 2964 28064
rect 2915 28033 2927 28036
rect 2869 28027 2927 28033
rect 2958 28024 2964 28036
rect 3016 28024 3022 28076
rect 10686 28024 10692 28076
rect 10744 28064 10750 28076
rect 11149 28067 11207 28073
rect 11149 28064 11161 28067
rect 10744 28036 11161 28064
rect 10744 28024 10750 28036
rect 11149 28033 11161 28036
rect 11195 28033 11207 28067
rect 11149 28027 11207 28033
rect 8386 28005 8392 28008
rect 3697 27999 3755 28005
rect 3697 27965 3709 27999
rect 3743 27965 3755 27999
rect 3697 27959 3755 27965
rect 8113 27999 8171 28005
rect 8113 27965 8125 27999
rect 8159 27965 8171 27999
rect 8380 27996 8392 28005
rect 8347 27968 8392 27996
rect 8113 27959 8171 27965
rect 8380 27959 8392 27968
rect 2682 27820 2688 27872
rect 2740 27860 2746 27872
rect 3605 27863 3663 27869
rect 3605 27860 3617 27863
rect 2740 27832 3617 27860
rect 2740 27820 2746 27832
rect 3605 27829 3617 27832
rect 3651 27860 3663 27863
rect 3712 27860 3740 27959
rect 3786 27888 3792 27940
rect 3844 27928 3850 27940
rect 3942 27931 4000 27937
rect 3942 27928 3954 27931
rect 3844 27900 3954 27928
rect 3844 27888 3850 27900
rect 3942 27897 3954 27900
rect 3988 27897 4000 27931
rect 3942 27891 4000 27897
rect 5166 27888 5172 27940
rect 5224 27928 5230 27940
rect 6546 27928 6552 27940
rect 5224 27900 6552 27928
rect 5224 27888 5230 27900
rect 6546 27888 6552 27900
rect 6604 27928 6610 27940
rect 7926 27928 7932 27940
rect 6604 27900 7932 27928
rect 6604 27888 6610 27900
rect 7926 27888 7932 27900
rect 7984 27928 7990 27940
rect 8128 27928 8156 27959
rect 8386 27956 8392 27959
rect 8444 27956 8450 28008
rect 10962 27956 10968 28008
rect 11020 27996 11026 28008
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11020 27968 11621 27996
rect 11020 27956 11026 27968
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 7984 27900 8156 27928
rect 7984 27888 7990 27900
rect 10042 27888 10048 27940
rect 10100 27928 10106 27940
rect 10413 27931 10471 27937
rect 10413 27928 10425 27931
rect 10100 27900 10425 27928
rect 10100 27888 10106 27900
rect 10413 27897 10425 27900
rect 10459 27928 10471 27931
rect 11057 27931 11115 27937
rect 11057 27928 11069 27931
rect 10459 27900 11069 27928
rect 10459 27897 10471 27900
rect 10413 27891 10471 27897
rect 11057 27897 11069 27900
rect 11103 27897 11115 27931
rect 11057 27891 11115 27897
rect 4062 27860 4068 27872
rect 3651 27832 4068 27860
rect 3651 27829 3663 27832
rect 3605 27823 3663 27829
rect 4062 27820 4068 27832
rect 4120 27820 4126 27872
rect 6086 27860 6092 27872
rect 6047 27832 6092 27860
rect 6086 27820 6092 27832
rect 6144 27820 6150 27872
rect 6822 27860 6828 27872
rect 6783 27832 6828 27860
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 8294 27820 8300 27872
rect 8352 27860 8358 27872
rect 9493 27863 9551 27869
rect 9493 27860 9505 27863
rect 8352 27832 9505 27860
rect 8352 27820 8358 27832
rect 9493 27829 9505 27832
rect 9539 27829 9551 27863
rect 9493 27823 9551 27829
rect 10502 27820 10508 27872
rect 10560 27860 10566 27872
rect 10965 27863 11023 27869
rect 10965 27860 10977 27863
rect 10560 27832 10977 27860
rect 10560 27820 10566 27832
rect 10965 27829 10977 27832
rect 11011 27860 11023 27863
rect 11330 27860 11336 27872
rect 11011 27832 11336 27860
rect 11011 27829 11023 27832
rect 10965 27823 11023 27829
rect 11330 27820 11336 27832
rect 11388 27820 11394 27872
rect 1104 27770 14812 27792
rect 1104 27718 6315 27770
rect 6367 27718 6379 27770
rect 6431 27718 6443 27770
rect 6495 27718 6507 27770
rect 6559 27718 11648 27770
rect 11700 27718 11712 27770
rect 11764 27718 11776 27770
rect 11828 27718 11840 27770
rect 11892 27718 14812 27770
rect 1104 27696 14812 27718
rect 3786 27656 3792 27668
rect 3747 27628 3792 27656
rect 3786 27616 3792 27628
rect 3844 27616 3850 27668
rect 4985 27659 5043 27665
rect 4985 27625 4997 27659
rect 5031 27656 5043 27659
rect 5350 27656 5356 27668
rect 5031 27628 5356 27656
rect 5031 27625 5043 27628
rect 4985 27619 5043 27625
rect 5350 27616 5356 27628
rect 5408 27616 5414 27668
rect 6641 27659 6699 27665
rect 6641 27625 6653 27659
rect 6687 27656 6699 27659
rect 7282 27656 7288 27668
rect 6687 27628 7288 27656
rect 6687 27625 6699 27628
rect 6641 27619 6699 27625
rect 7282 27616 7288 27628
rect 7340 27616 7346 27668
rect 7929 27659 7987 27665
rect 7929 27625 7941 27659
rect 7975 27656 7987 27659
rect 8386 27656 8392 27668
rect 7975 27628 8392 27656
rect 7975 27625 7987 27628
rect 7929 27619 7987 27625
rect 8386 27616 8392 27628
rect 8444 27616 8450 27668
rect 10045 27659 10103 27665
rect 10045 27625 10057 27659
rect 10091 27656 10103 27659
rect 10226 27656 10232 27668
rect 10091 27628 10232 27656
rect 10091 27625 10103 27628
rect 10045 27619 10103 27625
rect 10226 27616 10232 27628
rect 10284 27616 10290 27668
rect 10502 27616 10508 27668
rect 10560 27656 10566 27668
rect 10597 27659 10655 27665
rect 10597 27656 10609 27659
rect 10560 27628 10609 27656
rect 10560 27616 10566 27628
rect 10597 27625 10609 27628
rect 10643 27625 10655 27659
rect 10597 27619 10655 27625
rect 11146 27616 11152 27668
rect 11204 27656 11210 27668
rect 12158 27656 12164 27668
rect 11204 27628 12164 27656
rect 11204 27616 11210 27628
rect 12158 27616 12164 27628
rect 12216 27616 12222 27668
rect 2222 27548 2228 27600
rect 2280 27588 2286 27600
rect 2869 27591 2927 27597
rect 2869 27588 2881 27591
rect 2280 27560 2881 27588
rect 2280 27548 2286 27560
rect 2869 27557 2881 27560
rect 2915 27557 2927 27591
rect 2869 27551 2927 27557
rect 5528 27591 5586 27597
rect 5528 27557 5540 27591
rect 5574 27588 5586 27591
rect 5810 27588 5816 27600
rect 5574 27560 5816 27588
rect 5574 27557 5586 27560
rect 5528 27551 5586 27557
rect 5810 27548 5816 27560
rect 5868 27548 5874 27600
rect 8404 27588 8432 27616
rect 8404 27560 8524 27588
rect 2130 27480 2136 27532
rect 2188 27520 2194 27532
rect 2774 27520 2780 27532
rect 2188 27492 2780 27520
rect 2188 27480 2194 27492
rect 2774 27480 2780 27492
rect 2832 27520 2838 27532
rect 2832 27492 2877 27520
rect 2832 27480 2838 27492
rect 8294 27480 8300 27532
rect 8352 27520 8358 27532
rect 8389 27523 8447 27529
rect 8389 27520 8401 27523
rect 8352 27492 8401 27520
rect 8352 27480 8358 27492
rect 8389 27489 8401 27492
rect 8435 27489 8447 27523
rect 8496 27520 8524 27560
rect 8754 27548 8760 27600
rect 8812 27588 8818 27600
rect 9030 27588 9036 27600
rect 8812 27560 9036 27588
rect 8812 27548 8818 27560
rect 9030 27548 9036 27560
rect 9088 27548 9094 27600
rect 10244 27588 10272 27616
rect 11232 27591 11290 27597
rect 11232 27588 11244 27591
rect 10244 27560 11244 27588
rect 11232 27557 11244 27560
rect 11278 27588 11290 27591
rect 11330 27588 11336 27600
rect 11278 27560 11336 27588
rect 11278 27557 11290 27560
rect 11232 27551 11290 27557
rect 11330 27548 11336 27560
rect 11388 27548 11394 27600
rect 9950 27520 9956 27532
rect 8496 27492 8616 27520
rect 8389 27483 8447 27489
rect 3053 27455 3111 27461
rect 3053 27421 3065 27455
rect 3099 27452 3111 27455
rect 3786 27452 3792 27464
rect 3099 27424 3792 27452
rect 3099 27421 3111 27424
rect 3053 27415 3111 27421
rect 3786 27412 3792 27424
rect 3844 27412 3850 27464
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 5166 27452 5172 27464
rect 4212 27424 5172 27452
rect 4212 27412 4218 27424
rect 5166 27412 5172 27424
rect 5224 27452 5230 27464
rect 5261 27455 5319 27461
rect 5261 27452 5273 27455
rect 5224 27424 5273 27452
rect 5224 27412 5230 27424
rect 5261 27421 5273 27424
rect 5307 27421 5319 27455
rect 5261 27415 5319 27421
rect 7926 27412 7932 27464
rect 7984 27452 7990 27464
rect 8588 27461 8616 27492
rect 9600 27492 9956 27520
rect 8481 27455 8539 27461
rect 8481 27452 8493 27455
rect 7984 27424 8493 27452
rect 7984 27412 7990 27424
rect 8481 27421 8493 27424
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 8573 27455 8631 27461
rect 8573 27421 8585 27455
rect 8619 27421 8631 27455
rect 8573 27415 8631 27421
rect 2409 27387 2467 27393
rect 2409 27353 2421 27387
rect 2455 27384 2467 27387
rect 2866 27384 2872 27396
rect 2455 27356 2872 27384
rect 2455 27353 2467 27356
rect 2409 27347 2467 27353
rect 2866 27344 2872 27356
rect 2924 27344 2930 27396
rect 8496 27384 8524 27415
rect 8846 27384 8852 27396
rect 8496 27356 8852 27384
rect 8846 27344 8852 27356
rect 8904 27344 8910 27396
rect 8018 27316 8024 27328
rect 7979 27288 8024 27316
rect 8018 27276 8024 27288
rect 8076 27276 8082 27328
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 8478 27316 8484 27328
rect 8352 27288 8484 27316
rect 8352 27276 8358 27288
rect 8478 27276 8484 27288
rect 8536 27316 8542 27328
rect 9600 27316 9628 27492
rect 9950 27480 9956 27492
rect 10008 27480 10014 27532
rect 10962 27452 10968 27464
rect 10923 27424 10968 27452
rect 10962 27412 10968 27424
rect 11020 27412 11026 27464
rect 8536 27288 9628 27316
rect 8536 27276 8542 27288
rect 9766 27276 9772 27328
rect 9824 27316 9830 27328
rect 10042 27316 10048 27328
rect 9824 27288 10048 27316
rect 9824 27276 9830 27288
rect 10042 27276 10048 27288
rect 10100 27276 10106 27328
rect 12158 27276 12164 27328
rect 12216 27316 12222 27328
rect 12345 27319 12403 27325
rect 12345 27316 12357 27319
rect 12216 27288 12357 27316
rect 12216 27276 12222 27288
rect 12345 27285 12357 27288
rect 12391 27285 12403 27319
rect 12345 27279 12403 27285
rect 12802 27276 12808 27328
rect 12860 27316 12866 27328
rect 12897 27319 12955 27325
rect 12897 27316 12909 27319
rect 12860 27288 12909 27316
rect 12860 27276 12866 27288
rect 12897 27285 12909 27288
rect 12943 27285 12955 27319
rect 12897 27279 12955 27285
rect 1104 27226 14812 27248
rect 1104 27174 3648 27226
rect 3700 27174 3712 27226
rect 3764 27174 3776 27226
rect 3828 27174 3840 27226
rect 3892 27174 8982 27226
rect 9034 27174 9046 27226
rect 9098 27174 9110 27226
rect 9162 27174 9174 27226
rect 9226 27174 14315 27226
rect 14367 27174 14379 27226
rect 14431 27174 14443 27226
rect 14495 27174 14507 27226
rect 14559 27174 14812 27226
rect 1104 27152 14812 27174
rect 1765 27115 1823 27121
rect 1765 27081 1777 27115
rect 1811 27112 1823 27115
rect 3970 27112 3976 27124
rect 1811 27084 3976 27112
rect 1811 27081 1823 27084
rect 1765 27075 1823 27081
rect 3970 27072 3976 27084
rect 4028 27072 4034 27124
rect 5721 27115 5779 27121
rect 5721 27081 5733 27115
rect 5767 27112 5779 27115
rect 5810 27112 5816 27124
rect 5767 27084 5816 27112
rect 5767 27081 5779 27084
rect 5721 27075 5779 27081
rect 5810 27072 5816 27084
rect 5868 27072 5874 27124
rect 6086 27072 6092 27124
rect 6144 27112 6150 27124
rect 6825 27115 6883 27121
rect 6825 27112 6837 27115
rect 6144 27084 6837 27112
rect 6144 27072 6150 27084
rect 6825 27081 6837 27084
rect 6871 27081 6883 27115
rect 9490 27112 9496 27124
rect 6825 27075 6883 27081
rect 8864 27084 9496 27112
rect 2130 27044 2136 27056
rect 2091 27016 2136 27044
rect 2130 27004 2136 27016
rect 2188 27004 2194 27056
rect 2222 27004 2228 27056
rect 2280 27044 2286 27056
rect 2409 27047 2467 27053
rect 2409 27044 2421 27047
rect 2280 27016 2421 27044
rect 2280 27004 2286 27016
rect 2409 27013 2421 27016
rect 2455 27013 2467 27047
rect 5828 27044 5856 27072
rect 6178 27044 6184 27056
rect 5828 27016 6184 27044
rect 2409 27007 2467 27013
rect 6178 27004 6184 27016
rect 6236 27044 6242 27056
rect 6549 27047 6607 27053
rect 6549 27044 6561 27047
rect 6236 27016 6561 27044
rect 6236 27004 6242 27016
rect 6549 27013 6561 27016
rect 6595 27044 6607 27047
rect 6595 27016 7420 27044
rect 6595 27013 6607 27016
rect 6549 27007 6607 27013
rect 7392 26985 7420 27016
rect 8864 26985 8892 27084
rect 9490 27072 9496 27084
rect 9548 27072 9554 27124
rect 9861 27115 9919 27121
rect 9861 27112 9873 27115
rect 9692 27084 9873 27112
rect 7377 26979 7435 26985
rect 7377 26945 7389 26979
rect 7423 26945 7435 26979
rect 7377 26939 7435 26945
rect 8849 26979 8907 26985
rect 8849 26945 8861 26979
rect 8895 26945 8907 26979
rect 8849 26939 8907 26945
rect 8938 26936 8944 26988
rect 8996 26976 9002 26988
rect 8996 26948 9041 26976
rect 8996 26936 9002 26948
rect 2406 26868 2412 26920
rect 2464 26908 2470 26920
rect 2593 26911 2651 26917
rect 2593 26908 2605 26911
rect 2464 26880 2605 26908
rect 2464 26868 2470 26880
rect 2593 26877 2605 26880
rect 2639 26908 2651 26911
rect 2682 26908 2688 26920
rect 2639 26880 2688 26908
rect 2639 26877 2651 26880
rect 2593 26871 2651 26877
rect 2682 26868 2688 26880
rect 2740 26868 2746 26920
rect 6273 26911 6331 26917
rect 6273 26877 6285 26911
rect 6319 26908 6331 26911
rect 6822 26908 6828 26920
rect 6319 26880 6828 26908
rect 6319 26877 6331 26880
rect 6273 26871 6331 26877
rect 6822 26868 6828 26880
rect 6880 26908 6886 26920
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 6880 26880 7297 26908
rect 6880 26868 6886 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 7926 26868 7932 26920
rect 7984 26908 7990 26920
rect 8021 26911 8079 26917
rect 8021 26908 8033 26911
rect 7984 26880 8033 26908
rect 7984 26868 7990 26880
rect 8021 26877 8033 26880
rect 8067 26877 8079 26911
rect 8754 26908 8760 26920
rect 8715 26880 8760 26908
rect 8021 26871 8079 26877
rect 8754 26868 8760 26880
rect 8812 26868 8818 26920
rect 2860 26843 2918 26849
rect 2860 26809 2872 26843
rect 2906 26840 2918 26843
rect 2958 26840 2964 26852
rect 2906 26812 2964 26840
rect 2906 26809 2918 26812
rect 2860 26803 2918 26809
rect 2958 26800 2964 26812
rect 3016 26800 3022 26852
rect 5994 26800 6000 26852
rect 6052 26840 6058 26852
rect 6362 26840 6368 26852
rect 6052 26812 6368 26840
rect 6052 26800 6058 26812
rect 6362 26800 6368 26812
rect 6420 26800 6426 26852
rect 7190 26840 7196 26852
rect 7103 26812 7196 26840
rect 7190 26800 7196 26812
rect 7248 26840 7254 26852
rect 9692 26840 9720 27084
rect 9861 27081 9873 27084
rect 9907 27112 9919 27115
rect 9950 27112 9956 27124
rect 9907 27084 9956 27112
rect 9907 27081 9919 27084
rect 9861 27075 9919 27081
rect 9950 27072 9956 27084
rect 10008 27072 10014 27124
rect 10134 27072 10140 27124
rect 10192 27112 10198 27124
rect 10778 27112 10784 27124
rect 10192 27084 10784 27112
rect 10192 27072 10198 27084
rect 10778 27072 10784 27084
rect 10836 27072 10842 27124
rect 11330 27112 11336 27124
rect 11291 27084 11336 27112
rect 11330 27072 11336 27084
rect 11388 27072 11394 27124
rect 9766 27004 9772 27056
rect 9824 27044 9830 27056
rect 10410 27044 10416 27056
rect 9824 27016 10416 27044
rect 9824 27004 9830 27016
rect 10410 27004 10416 27016
rect 10468 27004 10474 27056
rect 10597 26979 10655 26985
rect 10597 26945 10609 26979
rect 10643 26976 10655 26979
rect 10870 26976 10876 26988
rect 10643 26948 10876 26976
rect 10643 26945 10655 26948
rect 10597 26939 10655 26945
rect 10870 26936 10876 26948
rect 10928 26976 10934 26988
rect 11348 26976 11376 27072
rect 10928 26948 11376 26976
rect 10928 26936 10934 26948
rect 12158 26936 12164 26988
rect 12216 26976 12222 26988
rect 12989 26979 13047 26985
rect 12989 26976 13001 26979
rect 12216 26948 13001 26976
rect 12216 26936 12222 26948
rect 12989 26945 13001 26948
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 9858 26868 9864 26920
rect 9916 26908 9922 26920
rect 10410 26908 10416 26920
rect 9916 26880 10416 26908
rect 9916 26868 9922 26880
rect 10410 26868 10416 26880
rect 10468 26868 10474 26920
rect 10321 26843 10379 26849
rect 10321 26840 10333 26843
rect 7248 26812 8432 26840
rect 9692 26812 10333 26840
rect 7248 26800 7254 26812
rect 5166 26732 5172 26784
rect 5224 26772 5230 26784
rect 8404 26781 8432 26812
rect 10321 26809 10333 26812
rect 10367 26809 10379 26843
rect 12802 26840 12808 26852
rect 12763 26812 12808 26840
rect 10321 26803 10379 26809
rect 12802 26800 12808 26812
rect 12860 26800 12866 26852
rect 5261 26775 5319 26781
rect 5261 26772 5273 26775
rect 5224 26744 5273 26772
rect 5224 26732 5230 26744
rect 5261 26741 5273 26744
rect 5307 26741 5319 26775
rect 5261 26735 5319 26741
rect 8389 26775 8447 26781
rect 8389 26741 8401 26775
rect 8435 26741 8447 26775
rect 9950 26772 9956 26784
rect 9911 26744 9956 26772
rect 8389 26735 8447 26741
rect 9950 26732 9956 26744
rect 10008 26732 10014 26784
rect 10413 26775 10471 26781
rect 10413 26741 10425 26775
rect 10459 26772 10471 26775
rect 10502 26772 10508 26784
rect 10459 26744 10508 26772
rect 10459 26741 10471 26744
rect 10413 26735 10471 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10962 26772 10968 26784
rect 10923 26744 10968 26772
rect 10962 26732 10968 26744
rect 11020 26732 11026 26784
rect 11514 26732 11520 26784
rect 11572 26772 11578 26784
rect 11793 26775 11851 26781
rect 11793 26772 11805 26775
rect 11572 26744 11805 26772
rect 11572 26732 11578 26744
rect 11793 26741 11805 26744
rect 11839 26741 11851 26775
rect 12158 26772 12164 26784
rect 12119 26744 12164 26772
rect 11793 26735 11851 26741
rect 12158 26732 12164 26744
rect 12216 26732 12222 26784
rect 12434 26732 12440 26784
rect 12492 26772 12498 26784
rect 12894 26772 12900 26784
rect 12492 26744 12537 26772
rect 12855 26744 12900 26772
rect 12492 26732 12498 26744
rect 12894 26732 12900 26744
rect 12952 26732 12958 26784
rect 1104 26682 14812 26704
rect 1104 26630 6315 26682
rect 6367 26630 6379 26682
rect 6431 26630 6443 26682
rect 6495 26630 6507 26682
rect 6559 26630 11648 26682
rect 11700 26630 11712 26682
rect 11764 26630 11776 26682
rect 11828 26630 11840 26682
rect 11892 26630 14812 26682
rect 1104 26608 14812 26630
rect 2958 26568 2964 26580
rect 2919 26540 2964 26568
rect 2958 26528 2964 26540
rect 3016 26528 3022 26580
rect 6178 26528 6184 26580
rect 6236 26568 6242 26580
rect 6549 26571 6607 26577
rect 6549 26568 6561 26571
rect 6236 26540 6561 26568
rect 6236 26528 6242 26540
rect 6549 26537 6561 26540
rect 6595 26537 6607 26571
rect 7190 26568 7196 26580
rect 7151 26540 7196 26568
rect 6549 26531 6607 26537
rect 7190 26528 7196 26540
rect 7248 26528 7254 26580
rect 7742 26568 7748 26580
rect 7703 26540 7748 26568
rect 7742 26528 7748 26540
rect 7800 26528 7806 26580
rect 8018 26528 8024 26580
rect 8076 26568 8082 26580
rect 8205 26571 8263 26577
rect 8205 26568 8217 26571
rect 8076 26540 8217 26568
rect 8076 26528 8082 26540
rect 8205 26537 8217 26540
rect 8251 26568 8263 26571
rect 8294 26568 8300 26580
rect 8251 26540 8300 26568
rect 8251 26537 8263 26540
rect 8205 26531 8263 26537
rect 8294 26528 8300 26540
rect 8352 26528 8358 26580
rect 8938 26528 8944 26580
rect 8996 26568 9002 26580
rect 9125 26571 9183 26577
rect 9125 26568 9137 26571
rect 8996 26540 9137 26568
rect 8996 26528 9002 26540
rect 9125 26537 9137 26540
rect 9171 26537 9183 26571
rect 10318 26568 10324 26580
rect 10279 26540 10324 26568
rect 9125 26531 9183 26537
rect 10318 26528 10324 26540
rect 10376 26528 10382 26580
rect 10686 26528 10692 26580
rect 10744 26568 10750 26580
rect 10781 26571 10839 26577
rect 10781 26568 10793 26571
rect 10744 26540 10793 26568
rect 10744 26528 10750 26540
rect 10781 26537 10793 26540
rect 10827 26537 10839 26571
rect 10781 26531 10839 26537
rect 11514 26528 11520 26580
rect 11572 26568 11578 26580
rect 12894 26568 12900 26580
rect 11572 26540 12900 26568
rect 11572 26528 11578 26540
rect 12894 26528 12900 26540
rect 12952 26528 12958 26580
rect 8110 26500 8116 26512
rect 8071 26472 8116 26500
rect 8110 26460 8116 26472
rect 8168 26460 8174 26512
rect 5442 26441 5448 26444
rect 5436 26432 5448 26441
rect 5403 26404 5448 26432
rect 5436 26395 5448 26404
rect 5442 26392 5448 26395
rect 5500 26392 5506 26444
rect 10686 26432 10692 26444
rect 10647 26404 10692 26432
rect 10686 26392 10692 26404
rect 10744 26392 10750 26444
rect 12158 26441 12164 26444
rect 12152 26432 12164 26441
rect 12119 26404 12164 26432
rect 12152 26395 12164 26404
rect 12158 26392 12164 26395
rect 12216 26392 12222 26444
rect 5166 26364 5172 26376
rect 5127 26336 5172 26364
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 7926 26324 7932 26376
rect 7984 26364 7990 26376
rect 8202 26364 8208 26376
rect 7984 26336 8208 26364
rect 7984 26324 7990 26336
rect 8202 26324 8208 26336
rect 8260 26364 8266 26376
rect 8297 26367 8355 26373
rect 8297 26364 8309 26367
rect 8260 26336 8309 26364
rect 8260 26324 8266 26336
rect 8297 26333 8309 26336
rect 8343 26333 8355 26367
rect 8297 26327 8355 26333
rect 9858 26324 9864 26376
rect 9916 26364 9922 26376
rect 9953 26367 10011 26373
rect 9953 26364 9965 26367
rect 9916 26336 9965 26364
rect 9916 26324 9922 26336
rect 9953 26333 9965 26336
rect 9999 26364 10011 26367
rect 10502 26364 10508 26376
rect 9999 26336 10508 26364
rect 9999 26333 10011 26336
rect 9953 26327 10011 26333
rect 10502 26324 10508 26336
rect 10560 26324 10566 26376
rect 10870 26364 10876 26376
rect 10831 26336 10876 26364
rect 10870 26324 10876 26336
rect 10928 26324 10934 26376
rect 11882 26364 11888 26376
rect 11843 26336 11888 26364
rect 11882 26324 11888 26336
rect 11940 26324 11946 26376
rect 2406 26256 2412 26308
rect 2464 26296 2470 26308
rect 2593 26299 2651 26305
rect 2593 26296 2605 26299
rect 2464 26268 2605 26296
rect 2464 26256 2470 26268
rect 2593 26265 2605 26268
rect 2639 26265 2651 26299
rect 2593 26259 2651 26265
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 8849 26299 8907 26305
rect 8849 26296 8861 26299
rect 8536 26268 8861 26296
rect 8536 26256 8542 26268
rect 8849 26265 8861 26268
rect 8895 26296 8907 26299
rect 9490 26296 9496 26308
rect 8895 26268 9496 26296
rect 8895 26265 8907 26268
rect 8849 26259 8907 26265
rect 9490 26256 9496 26268
rect 9548 26256 9554 26308
rect 13262 26296 13268 26308
rect 13223 26268 13268 26296
rect 13262 26256 13268 26268
rect 13320 26256 13326 26308
rect 1104 26138 14812 26160
rect 1104 26086 3648 26138
rect 3700 26086 3712 26138
rect 3764 26086 3776 26138
rect 3828 26086 3840 26138
rect 3892 26086 8982 26138
rect 9034 26086 9046 26138
rect 9098 26086 9110 26138
rect 9162 26086 9174 26138
rect 9226 26086 14315 26138
rect 14367 26086 14379 26138
rect 14431 26086 14443 26138
rect 14495 26086 14507 26138
rect 14559 26086 14812 26138
rect 1104 26064 14812 26086
rect 6822 26024 6828 26036
rect 6783 25996 6828 26024
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 7926 26024 7932 26036
rect 7887 25996 7932 26024
rect 7926 25984 7932 25996
rect 7984 25984 7990 26036
rect 8294 26024 8300 26036
rect 8255 25996 8300 26024
rect 8294 25984 8300 25996
rect 8352 25984 8358 26036
rect 10594 26024 10600 26036
rect 10555 25996 10600 26024
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 10873 26027 10931 26033
rect 10873 26024 10885 26027
rect 10744 25996 10885 26024
rect 10744 25984 10750 25996
rect 10873 25993 10885 25996
rect 10919 26024 10931 26027
rect 10919 25996 11100 26024
rect 10919 25993 10931 25996
rect 10873 25987 10931 25993
rect 5534 25848 5540 25900
rect 5592 25888 5598 25900
rect 5629 25891 5687 25897
rect 5629 25888 5641 25891
rect 5592 25860 5641 25888
rect 5592 25848 5598 25860
rect 5629 25857 5641 25860
rect 5675 25888 5687 25891
rect 6273 25891 6331 25897
rect 6273 25888 6285 25891
rect 5675 25860 6285 25888
rect 5675 25857 5687 25860
rect 5629 25851 5687 25857
rect 6273 25857 6285 25860
rect 6319 25888 6331 25891
rect 7466 25888 7472 25900
rect 6319 25860 7472 25888
rect 6319 25857 6331 25860
rect 6273 25851 6331 25857
rect 7466 25848 7472 25860
rect 7524 25848 7530 25900
rect 8294 25848 8300 25900
rect 8352 25888 8358 25900
rect 11072 25897 11100 25996
rect 12158 25916 12164 25968
rect 12216 25916 12222 25968
rect 8573 25891 8631 25897
rect 8573 25888 8585 25891
rect 8352 25860 8585 25888
rect 8352 25848 8358 25860
rect 8573 25857 8585 25860
rect 8619 25857 8631 25891
rect 8573 25851 8631 25857
rect 9401 25891 9459 25897
rect 9401 25857 9413 25891
rect 9447 25888 9459 25891
rect 10045 25891 10103 25897
rect 10045 25888 10057 25891
rect 9447 25860 10057 25888
rect 9447 25857 9459 25860
rect 9401 25851 9459 25857
rect 10045 25857 10057 25860
rect 10091 25857 10103 25891
rect 10045 25851 10103 25857
rect 11057 25891 11115 25897
rect 11057 25857 11069 25891
rect 11103 25857 11115 25891
rect 12176 25888 12204 25916
rect 12621 25891 12679 25897
rect 12621 25888 12633 25891
rect 11057 25851 11115 25857
rect 11716 25860 12633 25888
rect 6641 25823 6699 25829
rect 6641 25789 6653 25823
rect 6687 25820 6699 25823
rect 7193 25823 7251 25829
rect 7193 25820 7205 25823
rect 6687 25792 7205 25820
rect 6687 25789 6699 25792
rect 6641 25783 6699 25789
rect 7193 25789 7205 25792
rect 7239 25820 7251 25823
rect 8662 25820 8668 25832
rect 7239 25792 8668 25820
rect 7239 25789 7251 25792
rect 7193 25783 7251 25789
rect 8662 25780 8668 25792
rect 8720 25780 8726 25832
rect 9861 25823 9919 25829
rect 9861 25789 9873 25823
rect 9907 25820 9919 25823
rect 9950 25820 9956 25832
rect 9907 25792 9956 25820
rect 9907 25789 9919 25792
rect 9861 25783 9919 25789
rect 9950 25780 9956 25792
rect 10008 25780 10014 25832
rect 10060 25820 10088 25851
rect 11716 25820 11744 25860
rect 12621 25857 12633 25860
rect 12667 25857 12679 25891
rect 12621 25851 12679 25857
rect 11882 25820 11888 25832
rect 10060 25792 11744 25820
rect 11795 25792 11888 25820
rect 9033 25755 9091 25761
rect 9033 25721 9045 25755
rect 9079 25752 9091 25755
rect 9079 25724 9628 25752
rect 9079 25721 9091 25724
rect 9033 25715 9091 25721
rect 9600 25696 9628 25724
rect 10962 25712 10968 25764
rect 11020 25752 11026 25764
rect 11799 25752 11827 25792
rect 11882 25780 11888 25792
rect 11940 25780 11946 25832
rect 11020 25724 11827 25752
rect 11020 25712 11026 25724
rect 5166 25684 5172 25696
rect 5127 25656 5172 25684
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 7282 25644 7288 25696
rect 7340 25684 7346 25696
rect 9490 25684 9496 25696
rect 7340 25656 7385 25684
rect 9451 25656 9496 25684
rect 7340 25644 7346 25656
rect 9490 25644 9496 25656
rect 9548 25644 9554 25696
rect 9582 25644 9588 25696
rect 9640 25684 9646 25696
rect 9953 25687 10011 25693
rect 9953 25684 9965 25687
rect 9640 25656 9965 25684
rect 9640 25644 9646 25656
rect 9953 25653 9965 25656
rect 9999 25653 10011 25687
rect 9953 25647 10011 25653
rect 1104 25594 14812 25616
rect 1104 25542 6315 25594
rect 6367 25542 6379 25594
rect 6431 25542 6443 25594
rect 6495 25542 6507 25594
rect 6559 25542 11648 25594
rect 11700 25542 11712 25594
rect 11764 25542 11776 25594
rect 11828 25542 11840 25594
rect 11892 25542 14812 25594
rect 1104 25520 14812 25542
rect 1578 25480 1584 25492
rect 1539 25452 1584 25480
rect 1578 25440 1584 25452
rect 1636 25440 1642 25492
rect 6917 25483 6975 25489
rect 6917 25449 6929 25483
rect 6963 25480 6975 25483
rect 7282 25480 7288 25492
rect 6963 25452 7288 25480
rect 6963 25449 6975 25452
rect 6917 25443 6975 25449
rect 7282 25440 7288 25452
rect 7340 25440 7346 25492
rect 9493 25483 9551 25489
rect 9493 25449 9505 25483
rect 9539 25480 9551 25483
rect 9950 25480 9956 25492
rect 9539 25452 9956 25480
rect 9539 25449 9551 25452
rect 9493 25443 9551 25449
rect 9950 25440 9956 25452
rect 10008 25440 10014 25492
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25480 10839 25483
rect 10870 25480 10876 25492
rect 10827 25452 10876 25480
rect 10827 25449 10839 25452
rect 10781 25443 10839 25449
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 10045 25347 10103 25353
rect 10045 25313 10057 25347
rect 10091 25344 10103 25347
rect 11054 25344 11060 25356
rect 10091 25316 11060 25344
rect 10091 25313 10103 25316
rect 10045 25307 10103 25313
rect 11054 25304 11060 25316
rect 11112 25304 11118 25356
rect 4522 25276 4528 25288
rect 4483 25248 4528 25276
rect 4522 25236 4528 25248
rect 4580 25236 4586 25288
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 10137 25279 10195 25285
rect 10137 25276 10149 25279
rect 9548 25248 10149 25276
rect 9548 25236 9554 25248
rect 10137 25245 10149 25248
rect 10183 25245 10195 25279
rect 10318 25276 10324 25288
rect 10279 25248 10324 25276
rect 10137 25239 10195 25245
rect 10318 25236 10324 25248
rect 10376 25236 10382 25288
rect 10594 25236 10600 25288
rect 10652 25276 10658 25288
rect 10778 25276 10784 25288
rect 10652 25248 10784 25276
rect 10652 25236 10658 25248
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 9674 25208 9680 25220
rect 9635 25180 9680 25208
rect 9674 25168 9680 25180
rect 9732 25168 9738 25220
rect 8021 25143 8079 25149
rect 8021 25109 8033 25143
rect 8067 25140 8079 25143
rect 8202 25140 8208 25152
rect 8067 25112 8208 25140
rect 8067 25109 8079 25112
rect 8021 25103 8079 25109
rect 8202 25100 8208 25112
rect 8260 25100 8266 25152
rect 10226 25100 10232 25152
rect 10284 25140 10290 25152
rect 10502 25140 10508 25152
rect 10284 25112 10508 25140
rect 10284 25100 10290 25112
rect 10502 25100 10508 25112
rect 10560 25100 10566 25152
rect 1104 25050 14812 25072
rect 1104 24998 3648 25050
rect 3700 24998 3712 25050
rect 3764 24998 3776 25050
rect 3828 24998 3840 25050
rect 3892 24998 8982 25050
rect 9034 24998 9046 25050
rect 9098 24998 9110 25050
rect 9162 24998 9174 25050
rect 9226 24998 14315 25050
rect 14367 24998 14379 25050
rect 14431 24998 14443 25050
rect 14495 24998 14507 25050
rect 14559 24998 14812 25050
rect 1104 24976 14812 24998
rect 9033 24939 9091 24945
rect 9033 24905 9045 24939
rect 9079 24936 9091 24939
rect 9490 24936 9496 24948
rect 9079 24908 9496 24936
rect 9079 24905 9091 24908
rect 9033 24899 9091 24905
rect 9490 24896 9496 24908
rect 9548 24896 9554 24948
rect 9769 24939 9827 24945
rect 9769 24905 9781 24939
rect 9815 24936 9827 24939
rect 10318 24936 10324 24948
rect 9815 24908 10324 24936
rect 9815 24905 9827 24908
rect 9769 24899 9827 24905
rect 10318 24896 10324 24908
rect 10376 24896 10382 24948
rect 10045 24871 10103 24877
rect 8496 24840 9628 24868
rect 4341 24803 4399 24809
rect 4341 24769 4353 24803
rect 4387 24800 4399 24803
rect 4890 24800 4896 24812
rect 4387 24772 4896 24800
rect 4387 24769 4399 24772
rect 4341 24763 4399 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 4982 24760 4988 24812
rect 5040 24800 5046 24812
rect 5077 24803 5135 24809
rect 5077 24800 5089 24803
rect 5040 24772 5089 24800
rect 5040 24760 5046 24772
rect 5077 24769 5089 24772
rect 5123 24800 5135 24803
rect 5445 24803 5503 24809
rect 5445 24800 5457 24803
rect 5123 24772 5457 24800
rect 5123 24769 5135 24772
rect 5077 24763 5135 24769
rect 5445 24769 5457 24772
rect 5491 24769 5503 24803
rect 5445 24763 5503 24769
rect 7469 24803 7527 24809
rect 7469 24769 7481 24803
rect 7515 24800 7527 24803
rect 8018 24800 8024 24812
rect 7515 24772 8024 24800
rect 7515 24769 7527 24772
rect 7469 24763 7527 24769
rect 8018 24760 8024 24772
rect 8076 24800 8082 24812
rect 8496 24809 8524 24840
rect 8481 24803 8539 24809
rect 8481 24800 8493 24803
rect 8076 24772 8493 24800
rect 8076 24760 8082 24772
rect 8481 24769 8493 24772
rect 8527 24769 8539 24803
rect 9306 24800 9312 24812
rect 9267 24772 9312 24800
rect 8481 24763 8539 24769
rect 9306 24760 9312 24772
rect 9364 24760 9370 24812
rect 9600 24800 9628 24840
rect 10045 24837 10057 24871
rect 10091 24868 10103 24871
rect 11514 24868 11520 24880
rect 10091 24840 11520 24868
rect 10091 24837 10103 24840
rect 10045 24831 10103 24837
rect 11514 24828 11520 24840
rect 11572 24828 11578 24880
rect 10226 24800 10232 24812
rect 9600 24772 10232 24800
rect 10226 24760 10232 24772
rect 10284 24760 10290 24812
rect 10689 24803 10747 24809
rect 10689 24769 10701 24803
rect 10735 24800 10747 24803
rect 10870 24800 10876 24812
rect 10735 24772 10876 24800
rect 10735 24769 10747 24772
rect 10689 24763 10747 24769
rect 10870 24760 10876 24772
rect 10928 24760 10934 24812
rect 11054 24760 11060 24812
rect 11112 24800 11118 24812
rect 11425 24803 11483 24809
rect 11425 24800 11437 24803
rect 11112 24772 11437 24800
rect 11112 24760 11118 24772
rect 11425 24769 11437 24772
rect 11471 24800 11483 24803
rect 12342 24800 12348 24812
rect 11471 24772 12348 24800
rect 11471 24769 11483 24772
rect 11425 24763 11483 24769
rect 12342 24760 12348 24772
rect 12400 24760 12406 24812
rect 1949 24735 2007 24741
rect 1949 24701 1961 24735
rect 1995 24701 2007 24735
rect 1949 24695 2007 24701
rect 3973 24735 4031 24741
rect 3973 24701 3985 24735
rect 4019 24732 4031 24735
rect 4522 24732 4528 24744
rect 4019 24704 4528 24732
rect 4019 24701 4031 24704
rect 3973 24695 4031 24701
rect 1857 24599 1915 24605
rect 1857 24565 1869 24599
rect 1903 24596 1915 24599
rect 1964 24596 1992 24695
rect 4522 24692 4528 24704
rect 4580 24732 4586 24744
rect 4801 24735 4859 24741
rect 4801 24732 4813 24735
rect 4580 24704 4813 24732
rect 4580 24692 4586 24704
rect 4801 24701 4813 24704
rect 4847 24701 4859 24735
rect 4801 24695 4859 24701
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 7745 24735 7803 24741
rect 7745 24732 7757 24735
rect 7708 24704 7757 24732
rect 7708 24692 7714 24704
rect 7745 24701 7757 24704
rect 7791 24732 7803 24735
rect 8389 24735 8447 24741
rect 8389 24732 8401 24735
rect 7791 24704 8401 24732
rect 7791 24701 7803 24704
rect 7745 24695 7803 24701
rect 8389 24701 8401 24704
rect 8435 24732 8447 24735
rect 8754 24732 8760 24744
rect 8435 24704 8760 24732
rect 8435 24701 8447 24704
rect 8389 24695 8447 24701
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 8846 24692 8852 24744
rect 8904 24732 8910 24744
rect 9324 24732 9352 24760
rect 10413 24735 10471 24741
rect 10413 24732 10425 24735
rect 8904 24704 10425 24732
rect 8904 24692 8910 24704
rect 10413 24701 10425 24704
rect 10459 24701 10471 24735
rect 10413 24695 10471 24701
rect 2222 24673 2228 24676
rect 2216 24664 2228 24673
rect 2183 24636 2228 24664
rect 2216 24627 2228 24636
rect 2222 24624 2228 24627
rect 2280 24624 2286 24676
rect 2406 24596 2412 24608
rect 1903 24568 2412 24596
rect 1903 24565 1915 24568
rect 1857 24559 1915 24565
rect 2406 24556 2412 24568
rect 2464 24556 2470 24608
rect 2958 24556 2964 24608
rect 3016 24596 3022 24608
rect 3329 24599 3387 24605
rect 3329 24596 3341 24599
rect 3016 24568 3341 24596
rect 3016 24556 3022 24568
rect 3329 24565 3341 24568
rect 3375 24565 3387 24599
rect 4430 24596 4436 24608
rect 4391 24568 4436 24596
rect 3329 24559 3387 24565
rect 4430 24556 4436 24568
rect 4488 24556 4494 24608
rect 7926 24596 7932 24608
rect 7887 24568 7932 24596
rect 7926 24556 7932 24568
rect 7984 24556 7990 24608
rect 8202 24556 8208 24608
rect 8260 24596 8266 24608
rect 8297 24599 8355 24605
rect 8297 24596 8309 24599
rect 8260 24568 8309 24596
rect 8260 24556 8266 24568
rect 8297 24565 8309 24568
rect 8343 24596 8355 24599
rect 8478 24596 8484 24608
rect 8343 24568 8484 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 8478 24556 8484 24568
rect 8536 24596 8542 24608
rect 10134 24596 10140 24608
rect 8536 24568 10140 24596
rect 8536 24556 8542 24568
rect 10134 24556 10140 24568
rect 10192 24596 10198 24608
rect 10505 24599 10563 24605
rect 10505 24596 10517 24599
rect 10192 24568 10517 24596
rect 10192 24556 10198 24568
rect 10505 24565 10517 24568
rect 10551 24596 10563 24599
rect 11057 24599 11115 24605
rect 11057 24596 11069 24599
rect 10551 24568 11069 24596
rect 10551 24565 10563 24568
rect 10505 24559 10563 24565
rect 11057 24565 11069 24568
rect 11103 24565 11115 24599
rect 11057 24559 11115 24565
rect 1104 24506 14812 24528
rect 1104 24454 6315 24506
rect 6367 24454 6379 24506
rect 6431 24454 6443 24506
rect 6495 24454 6507 24506
rect 6559 24454 11648 24506
rect 11700 24454 11712 24506
rect 11764 24454 11776 24506
rect 11828 24454 11840 24506
rect 11892 24454 14812 24506
rect 1104 24432 14812 24454
rect 1394 24352 1400 24404
rect 1452 24392 1458 24404
rect 1581 24395 1639 24401
rect 1581 24392 1593 24395
rect 1452 24364 1593 24392
rect 1452 24352 1458 24364
rect 1581 24361 1593 24364
rect 1627 24392 1639 24395
rect 2317 24395 2375 24401
rect 2317 24392 2329 24395
rect 1627 24364 2329 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 2317 24361 2329 24364
rect 2363 24361 2375 24395
rect 2682 24392 2688 24404
rect 2595 24364 2688 24392
rect 2317 24355 2375 24361
rect 2682 24352 2688 24364
rect 2740 24392 2746 24404
rect 4065 24395 4123 24401
rect 4065 24392 4077 24395
rect 2740 24364 4077 24392
rect 2740 24352 2746 24364
rect 4065 24361 4077 24364
rect 4111 24361 4123 24395
rect 4065 24355 4123 24361
rect 7101 24395 7159 24401
rect 7101 24361 7113 24395
rect 7147 24392 7159 24395
rect 7653 24395 7711 24401
rect 7653 24392 7665 24395
rect 7147 24364 7665 24392
rect 7147 24361 7159 24364
rect 7101 24355 7159 24361
rect 7653 24361 7665 24364
rect 7699 24392 7711 24395
rect 7926 24392 7932 24404
rect 7699 24364 7932 24392
rect 7699 24361 7711 24364
rect 7653 24355 7711 24361
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 9858 24352 9864 24404
rect 9916 24392 9922 24404
rect 10137 24395 10195 24401
rect 10137 24392 10149 24395
rect 9916 24364 10149 24392
rect 9916 24352 9922 24364
rect 10137 24361 10149 24364
rect 10183 24361 10195 24395
rect 10137 24355 10195 24361
rect 10781 24395 10839 24401
rect 10781 24361 10793 24395
rect 10827 24392 10839 24395
rect 10870 24392 10876 24404
rect 10827 24364 10876 24392
rect 10827 24361 10839 24364
rect 10781 24355 10839 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 7558 24324 7564 24336
rect 7519 24296 7564 24324
rect 7558 24284 7564 24296
rect 7616 24284 7622 24336
rect 4062 24216 4068 24268
rect 4120 24256 4126 24268
rect 4430 24256 4436 24268
rect 4120 24228 4436 24256
rect 4120 24216 4126 24228
rect 4430 24216 4436 24228
rect 4488 24216 4494 24268
rect 9674 24216 9680 24268
rect 9732 24256 9738 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9732 24228 10057 24256
rect 9732 24216 9738 24228
rect 10045 24225 10057 24228
rect 10091 24256 10103 24259
rect 10318 24256 10324 24268
rect 10091 24228 10324 24256
rect 10091 24225 10103 24228
rect 10045 24219 10103 24225
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 11514 24265 11520 24268
rect 11508 24256 11520 24265
rect 11475 24228 11520 24256
rect 11508 24219 11520 24228
rect 11514 24216 11520 24219
rect 11572 24216 11578 24268
rect 2406 24148 2412 24200
rect 2464 24188 2470 24200
rect 2777 24191 2835 24197
rect 2777 24188 2789 24191
rect 2464 24160 2789 24188
rect 2464 24148 2470 24160
rect 2777 24157 2789 24160
rect 2823 24157 2835 24191
rect 2958 24188 2964 24200
rect 2919 24160 2964 24188
rect 2777 24151 2835 24157
rect 2958 24148 2964 24160
rect 3016 24148 3022 24200
rect 4522 24188 4528 24200
rect 4483 24160 4528 24188
rect 4522 24148 4528 24160
rect 4580 24148 4586 24200
rect 4706 24188 4712 24200
rect 4667 24160 4712 24188
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 7837 24191 7895 24197
rect 7837 24157 7849 24191
rect 7883 24188 7895 24191
rect 7926 24188 7932 24200
rect 7883 24160 7932 24188
rect 7883 24157 7895 24160
rect 7837 24151 7895 24157
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 10226 24148 10232 24200
rect 10284 24188 10290 24200
rect 10284 24160 10329 24188
rect 10284 24148 10290 24160
rect 10962 24148 10968 24200
rect 11020 24188 11026 24200
rect 11241 24191 11299 24197
rect 11241 24188 11253 24191
rect 11020 24160 11253 24188
rect 11020 24148 11026 24160
rect 11241 24157 11253 24160
rect 11287 24157 11299 24191
rect 11241 24151 11299 24157
rect 2041 24055 2099 24061
rect 2041 24021 2053 24055
rect 2087 24052 2099 24055
rect 2222 24052 2228 24064
rect 2087 24024 2228 24052
rect 2087 24021 2099 24024
rect 2041 24015 2099 24021
rect 2222 24012 2228 24024
rect 2280 24012 2286 24064
rect 3421 24055 3479 24061
rect 3421 24021 3433 24055
rect 3467 24052 3479 24055
rect 3510 24052 3516 24064
rect 3467 24024 3516 24052
rect 3467 24021 3479 24024
rect 3421 24015 3479 24021
rect 3510 24012 3516 24024
rect 3568 24012 3574 24064
rect 4430 24012 4436 24064
rect 4488 24052 4494 24064
rect 4890 24052 4896 24064
rect 4488 24024 4896 24052
rect 4488 24012 4494 24024
rect 4890 24012 4896 24024
rect 4948 24012 4954 24064
rect 5261 24055 5319 24061
rect 5261 24021 5273 24055
rect 5307 24052 5319 24055
rect 5534 24052 5540 24064
rect 5307 24024 5540 24052
rect 5307 24021 5319 24024
rect 5261 24015 5319 24021
rect 5534 24012 5540 24024
rect 5592 24012 5598 24064
rect 7190 24052 7196 24064
rect 7151 24024 7196 24052
rect 7190 24012 7196 24024
rect 7248 24012 7254 24064
rect 9674 24052 9680 24064
rect 9635 24024 9680 24052
rect 9674 24012 9680 24024
rect 9732 24012 9738 24064
rect 12434 24012 12440 24064
rect 12492 24052 12498 24064
rect 12621 24055 12679 24061
rect 12621 24052 12633 24055
rect 12492 24024 12633 24052
rect 12492 24012 12498 24024
rect 12621 24021 12633 24024
rect 12667 24021 12679 24055
rect 12621 24015 12679 24021
rect 1104 23962 14812 23984
rect 1104 23910 3648 23962
rect 3700 23910 3712 23962
rect 3764 23910 3776 23962
rect 3828 23910 3840 23962
rect 3892 23910 8982 23962
rect 9034 23910 9046 23962
rect 9098 23910 9110 23962
rect 9162 23910 9174 23962
rect 9226 23910 14315 23962
rect 14367 23910 14379 23962
rect 14431 23910 14443 23962
rect 14495 23910 14507 23962
rect 14559 23910 14812 23962
rect 1104 23888 14812 23910
rect 2317 23851 2375 23857
rect 2317 23817 2329 23851
rect 2363 23848 2375 23851
rect 2958 23848 2964 23860
rect 2363 23820 2964 23848
rect 2363 23817 2375 23820
rect 2317 23811 2375 23817
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 4706 23848 4712 23860
rect 4212 23820 4712 23848
rect 4212 23808 4218 23820
rect 4706 23808 4712 23820
rect 4764 23848 4770 23860
rect 5353 23851 5411 23857
rect 5353 23848 5365 23851
rect 4764 23820 5365 23848
rect 4764 23808 4770 23820
rect 5353 23817 5365 23820
rect 5399 23817 5411 23851
rect 5353 23811 5411 23817
rect 6641 23851 6699 23857
rect 6641 23817 6653 23851
rect 6687 23848 6699 23851
rect 7926 23848 7932 23860
rect 6687 23820 7932 23848
rect 6687 23817 6699 23820
rect 6641 23811 6699 23817
rect 7926 23808 7932 23820
rect 7984 23848 7990 23860
rect 9125 23851 9183 23857
rect 9125 23848 9137 23851
rect 7984 23820 9137 23848
rect 7984 23808 7990 23820
rect 9125 23817 9137 23820
rect 9171 23817 9183 23851
rect 9125 23811 9183 23817
rect 9769 23851 9827 23857
rect 9769 23817 9781 23851
rect 9815 23848 9827 23851
rect 9858 23848 9864 23860
rect 9815 23820 9864 23848
rect 9815 23817 9827 23820
rect 9769 23811 9827 23817
rect 9858 23808 9864 23820
rect 9916 23848 9922 23860
rect 10134 23848 10140 23860
rect 9916 23820 10140 23848
rect 9916 23808 9922 23820
rect 10134 23808 10140 23820
rect 10192 23808 10198 23860
rect 10226 23808 10232 23860
rect 10284 23848 10290 23860
rect 10413 23851 10471 23857
rect 10413 23848 10425 23851
rect 10284 23820 10425 23848
rect 10284 23808 10290 23820
rect 10413 23817 10425 23820
rect 10459 23848 10471 23851
rect 11054 23848 11060 23860
rect 10459 23820 11060 23848
rect 10459 23817 10471 23820
rect 10413 23811 10471 23817
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 4341 23783 4399 23789
rect 4341 23749 4353 23783
rect 4387 23780 4399 23783
rect 4522 23780 4528 23792
rect 4387 23752 4528 23780
rect 4387 23749 4399 23752
rect 4341 23743 4399 23749
rect 4522 23740 4528 23752
rect 4580 23780 4586 23792
rect 5721 23783 5779 23789
rect 5721 23780 5733 23783
rect 4580 23752 5733 23780
rect 4580 23740 4586 23752
rect 5721 23749 5733 23752
rect 5767 23749 5779 23783
rect 5721 23743 5779 23749
rect 6730 23740 6736 23792
rect 6788 23780 6794 23792
rect 7285 23783 7343 23789
rect 7285 23780 7297 23783
rect 6788 23752 7297 23780
rect 6788 23740 6794 23752
rect 7285 23749 7297 23752
rect 7331 23780 7343 23783
rect 7558 23780 7564 23792
rect 7331 23752 7564 23780
rect 7331 23749 7343 23752
rect 7285 23743 7343 23749
rect 7558 23740 7564 23752
rect 7616 23740 7622 23792
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23712 2007 23715
rect 3234 23712 3240 23724
rect 1995 23684 3240 23712
rect 1995 23681 2007 23684
rect 1949 23675 2007 23681
rect 3234 23672 3240 23684
rect 3292 23712 3298 23724
rect 3421 23715 3479 23721
rect 3421 23712 3433 23715
rect 3292 23684 3433 23712
rect 3292 23672 3298 23684
rect 3421 23681 3433 23684
rect 3467 23712 3479 23715
rect 3881 23715 3939 23721
rect 3881 23712 3893 23715
rect 3467 23684 3893 23712
rect 3467 23681 3479 23684
rect 3421 23675 3479 23681
rect 3881 23681 3893 23684
rect 3927 23712 3939 23715
rect 4982 23712 4988 23724
rect 3927 23684 4988 23712
rect 3927 23681 3939 23684
rect 3881 23675 3939 23681
rect 4982 23672 4988 23684
rect 5040 23672 5046 23724
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 4709 23647 4767 23653
rect 4709 23644 4721 23647
rect 4295 23616 4721 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4709 23613 4721 23616
rect 4755 23644 4767 23647
rect 4890 23644 4896 23656
rect 4755 23616 4896 23644
rect 4755 23613 4767 23616
rect 4709 23607 4767 23613
rect 4890 23604 4896 23616
rect 4948 23644 4954 23656
rect 5074 23644 5080 23656
rect 4948 23616 5080 23644
rect 4948 23604 4954 23616
rect 5074 23604 5080 23616
rect 5132 23604 5138 23656
rect 8018 23653 8024 23656
rect 7745 23647 7803 23653
rect 7745 23644 7757 23647
rect 7576 23616 7757 23644
rect 2590 23536 2596 23588
rect 2648 23576 2654 23588
rect 2685 23579 2743 23585
rect 2685 23576 2697 23579
rect 2648 23548 2697 23576
rect 2648 23536 2654 23548
rect 2685 23545 2697 23548
rect 2731 23576 2743 23579
rect 4798 23576 4804 23588
rect 2731 23548 3188 23576
rect 4759 23548 4804 23576
rect 2731 23545 2743 23548
rect 2685 23539 2743 23545
rect 3160 23520 3188 23548
rect 4798 23536 4804 23548
rect 4856 23536 4862 23588
rect 2774 23468 2780 23520
rect 2832 23508 2838 23520
rect 3142 23508 3148 23520
rect 2832 23480 2877 23508
rect 3103 23480 3148 23508
rect 2832 23468 2838 23480
rect 3142 23468 3148 23480
rect 3200 23468 3206 23520
rect 3237 23511 3295 23517
rect 3237 23477 3249 23511
rect 3283 23508 3295 23511
rect 3510 23508 3516 23520
rect 3283 23480 3516 23508
rect 3283 23477 3295 23480
rect 3237 23471 3295 23477
rect 3510 23468 3516 23480
rect 3568 23468 3574 23520
rect 4246 23468 4252 23520
rect 4304 23508 4310 23520
rect 4522 23508 4528 23520
rect 4304 23480 4528 23508
rect 4304 23468 4310 23480
rect 4522 23468 4528 23480
rect 4580 23468 4586 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7576 23517 7604 23616
rect 7745 23613 7757 23616
rect 7791 23613 7803 23647
rect 8012 23644 8024 23653
rect 7979 23616 8024 23644
rect 7745 23607 7803 23613
rect 8012 23607 8024 23616
rect 8018 23604 8024 23607
rect 8076 23604 8082 23656
rect 7561 23511 7619 23517
rect 7561 23508 7573 23511
rect 6972 23480 7573 23508
rect 6972 23468 6978 23480
rect 7561 23477 7573 23480
rect 7607 23508 7619 23511
rect 8202 23508 8208 23520
rect 7607 23480 8208 23508
rect 7607 23477 7619 23480
rect 7561 23471 7619 23477
rect 8202 23468 8208 23480
rect 8260 23468 8266 23520
rect 10137 23511 10195 23517
rect 10137 23477 10149 23511
rect 10183 23508 10195 23511
rect 10318 23508 10324 23520
rect 10183 23480 10324 23508
rect 10183 23477 10195 23480
rect 10137 23471 10195 23477
rect 10318 23468 10324 23480
rect 10376 23468 10382 23520
rect 10962 23468 10968 23520
rect 11020 23508 11026 23520
rect 11241 23511 11299 23517
rect 11241 23508 11253 23511
rect 11020 23480 11253 23508
rect 11020 23468 11026 23480
rect 11241 23477 11253 23480
rect 11287 23477 11299 23511
rect 11241 23471 11299 23477
rect 11514 23468 11520 23520
rect 11572 23508 11578 23520
rect 11701 23511 11759 23517
rect 11701 23508 11713 23511
rect 11572 23480 11713 23508
rect 11572 23468 11578 23480
rect 11701 23477 11713 23480
rect 11747 23508 11759 23511
rect 12342 23508 12348 23520
rect 11747 23480 12348 23508
rect 11747 23477 11759 23480
rect 11701 23471 11759 23477
rect 12342 23468 12348 23480
rect 12400 23468 12406 23520
rect 1104 23418 14812 23440
rect 1104 23366 6315 23418
rect 6367 23366 6379 23418
rect 6431 23366 6443 23418
rect 6495 23366 6507 23418
rect 6559 23366 11648 23418
rect 11700 23366 11712 23418
rect 11764 23366 11776 23418
rect 11828 23366 11840 23418
rect 11892 23366 14812 23418
rect 1104 23344 14812 23366
rect 1578 23304 1584 23316
rect 1539 23276 1584 23304
rect 1578 23264 1584 23276
rect 1636 23264 1642 23316
rect 2317 23307 2375 23313
rect 2317 23273 2329 23307
rect 2363 23304 2375 23307
rect 2406 23304 2412 23316
rect 2363 23276 2412 23304
rect 2363 23273 2375 23276
rect 2317 23267 2375 23273
rect 2406 23264 2412 23276
rect 2464 23264 2470 23316
rect 3881 23307 3939 23313
rect 3881 23273 3893 23307
rect 3927 23304 3939 23307
rect 4062 23304 4068 23316
rect 3927 23276 4068 23304
rect 3927 23273 3939 23276
rect 3881 23267 3939 23273
rect 4062 23264 4068 23276
rect 4120 23264 4126 23316
rect 4433 23307 4491 23313
rect 4433 23273 4445 23307
rect 4479 23304 4491 23307
rect 4798 23304 4804 23316
rect 4479 23276 4804 23304
rect 4479 23273 4491 23276
rect 4433 23267 4491 23273
rect 4798 23264 4804 23276
rect 4856 23304 4862 23316
rect 5442 23304 5448 23316
rect 4856 23276 5448 23304
rect 4856 23264 4862 23276
rect 5442 23264 5448 23276
rect 5500 23264 5506 23316
rect 5905 23307 5963 23313
rect 5905 23304 5917 23307
rect 5543 23276 5917 23304
rect 1949 23239 2007 23245
rect 1949 23205 1961 23239
rect 1995 23236 2007 23239
rect 2682 23236 2688 23248
rect 1995 23208 2688 23236
rect 1995 23205 2007 23208
rect 1949 23199 2007 23205
rect 2682 23196 2688 23208
rect 2740 23196 2746 23248
rect 2777 23239 2835 23245
rect 2777 23205 2789 23239
rect 2823 23236 2835 23239
rect 2866 23236 2872 23248
rect 2823 23208 2872 23236
rect 2823 23205 2835 23208
rect 2777 23199 2835 23205
rect 2866 23196 2872 23208
rect 2924 23196 2930 23248
rect 4982 23196 4988 23248
rect 5040 23236 5046 23248
rect 5543 23236 5571 23276
rect 5905 23273 5917 23276
rect 5951 23273 5963 23307
rect 5905 23267 5963 23273
rect 7009 23307 7067 23313
rect 7009 23273 7021 23307
rect 7055 23273 7067 23307
rect 7009 23267 7067 23273
rect 5040 23208 5571 23236
rect 5040 23196 5046 23208
rect 5718 23196 5724 23248
rect 5776 23236 5782 23248
rect 7024 23236 7052 23267
rect 7190 23264 7196 23316
rect 7248 23304 7254 23316
rect 7377 23307 7435 23313
rect 7377 23304 7389 23307
rect 7248 23276 7389 23304
rect 7248 23264 7254 23276
rect 7377 23273 7389 23276
rect 7423 23304 7435 23307
rect 8389 23307 8447 23313
rect 8389 23304 8401 23307
rect 7423 23276 8401 23304
rect 7423 23273 7435 23276
rect 7377 23267 7435 23273
rect 8389 23273 8401 23276
rect 8435 23273 8447 23307
rect 11054 23304 11060 23316
rect 11015 23276 11060 23304
rect 8389 23267 8447 23273
rect 11054 23264 11060 23276
rect 11112 23264 11118 23316
rect 12618 23304 12624 23316
rect 12531 23276 12624 23304
rect 12618 23264 12624 23276
rect 12676 23304 12682 23316
rect 13078 23304 13084 23316
rect 12676 23276 13084 23304
rect 12676 23264 12682 23276
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 8018 23236 8024 23248
rect 5776 23208 7052 23236
rect 7979 23208 8024 23236
rect 5776 23196 5782 23208
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 10962 23236 10968 23248
rect 9692 23208 10968 23236
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 1670 23168 1676 23180
rect 1443 23140 1676 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 1670 23128 1676 23140
rect 1728 23128 1734 23180
rect 4798 23177 4804 23180
rect 4792 23131 4804 23177
rect 4856 23168 4862 23180
rect 4856 23140 4892 23168
rect 4798 23128 4804 23131
rect 4856 23128 4862 23140
rect 9582 23128 9588 23180
rect 9640 23168 9646 23180
rect 9692 23177 9720 23208
rect 10962 23196 10968 23208
rect 11020 23196 11026 23248
rect 12250 23196 12256 23248
rect 12308 23236 12314 23248
rect 12529 23239 12587 23245
rect 12529 23236 12541 23239
rect 12308 23208 12541 23236
rect 12308 23196 12314 23208
rect 12529 23205 12541 23208
rect 12575 23236 12587 23239
rect 12710 23236 12716 23248
rect 12575 23208 12716 23236
rect 12575 23205 12587 23208
rect 12529 23199 12587 23205
rect 12710 23196 12716 23208
rect 12768 23196 12774 23248
rect 9677 23171 9735 23177
rect 9677 23168 9689 23171
rect 9640 23140 9689 23168
rect 9640 23128 9646 23140
rect 9677 23137 9689 23140
rect 9723 23137 9735 23171
rect 9677 23131 9735 23137
rect 9944 23171 10002 23177
rect 9944 23137 9956 23171
rect 9990 23168 10002 23171
rect 10226 23168 10232 23180
rect 9990 23140 10232 23168
rect 9990 23137 10002 23140
rect 9944 23131 10002 23137
rect 10226 23128 10232 23140
rect 10284 23168 10290 23180
rect 10870 23168 10876 23180
rect 10284 23140 10876 23168
rect 10284 23128 10290 23140
rect 10870 23128 10876 23140
rect 10928 23128 10934 23180
rect 12342 23128 12348 23180
rect 12400 23168 12406 23180
rect 12400 23140 12848 23168
rect 12400 23128 12406 23140
rect 2774 23060 2780 23112
rect 2832 23100 2838 23112
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2832 23072 2881 23100
rect 2832 23060 2838 23072
rect 2869 23069 2881 23072
rect 2915 23100 2927 23103
rect 2958 23100 2964 23112
rect 2915 23072 2964 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 2958 23060 2964 23072
rect 3016 23060 3022 23112
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23100 3111 23103
rect 4062 23100 4068 23112
rect 3099 23072 4068 23100
rect 3099 23069 3111 23072
rect 3053 23063 3111 23069
rect 2222 22992 2228 23044
rect 2280 23032 2286 23044
rect 3068 23032 3096 23063
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 4525 23103 4583 23109
rect 4525 23069 4537 23103
rect 4571 23069 4583 23103
rect 4525 23063 4583 23069
rect 6549 23103 6607 23109
rect 6549 23069 6561 23103
rect 6595 23100 6607 23103
rect 7466 23100 7472 23112
rect 6595 23072 7472 23100
rect 6595 23069 6607 23072
rect 6549 23063 6607 23069
rect 2280 23004 3096 23032
rect 2280 22992 2286 23004
rect 4540 22964 4568 23063
rect 7466 23060 7472 23072
rect 7524 23060 7530 23112
rect 7561 23103 7619 23109
rect 7561 23069 7573 23103
rect 7607 23069 7619 23103
rect 7561 23063 7619 23069
rect 6914 23032 6920 23044
rect 6827 23004 6920 23032
rect 6914 22992 6920 23004
rect 6972 23032 6978 23044
rect 7576 23032 7604 23063
rect 11790 23060 11796 23112
rect 11848 23100 11854 23112
rect 12618 23100 12624 23112
rect 11848 23072 12624 23100
rect 11848 23060 11854 23072
rect 12618 23060 12624 23072
rect 12676 23060 12682 23112
rect 12820 23109 12848 23140
rect 12805 23103 12863 23109
rect 12805 23069 12817 23103
rect 12851 23100 12863 23103
rect 12851 23072 13308 23100
rect 12851 23069 12863 23072
rect 12805 23063 12863 23069
rect 6972 23004 7604 23032
rect 6972 22992 6978 23004
rect 13280 22976 13308 23072
rect 4706 22964 4712 22976
rect 4540 22936 4712 22964
rect 4706 22924 4712 22936
rect 4764 22964 4770 22976
rect 5166 22964 5172 22976
rect 4764 22936 5172 22964
rect 4764 22924 4770 22936
rect 5166 22924 5172 22936
rect 5224 22924 5230 22976
rect 12158 22964 12164 22976
rect 12119 22936 12164 22964
rect 12158 22924 12164 22936
rect 12216 22924 12222 22976
rect 13262 22964 13268 22976
rect 13223 22936 13268 22964
rect 13262 22924 13268 22936
rect 13320 22924 13326 22976
rect 1104 22874 14812 22896
rect 1104 22822 3648 22874
rect 3700 22822 3712 22874
rect 3764 22822 3776 22874
rect 3828 22822 3840 22874
rect 3892 22822 8982 22874
rect 9034 22822 9046 22874
rect 9098 22822 9110 22874
rect 9162 22822 9174 22874
rect 9226 22822 14315 22874
rect 14367 22822 14379 22874
rect 14431 22822 14443 22874
rect 14495 22822 14507 22874
rect 14559 22822 14812 22874
rect 1104 22800 14812 22822
rect 1857 22763 1915 22769
rect 1857 22729 1869 22763
rect 1903 22760 1915 22763
rect 2958 22760 2964 22772
rect 1903 22732 2964 22760
rect 1903 22729 1915 22732
rect 1857 22723 1915 22729
rect 2958 22720 2964 22732
rect 3016 22720 3022 22772
rect 4062 22760 4068 22772
rect 4023 22732 4068 22760
rect 4062 22720 4068 22732
rect 4120 22720 4126 22772
rect 8205 22763 8263 22769
rect 8205 22760 8217 22763
rect 5920 22732 8217 22760
rect 2222 22692 2228 22704
rect 2183 22664 2228 22692
rect 2222 22652 2228 22664
rect 2280 22652 2286 22704
rect 2498 22692 2504 22704
rect 2459 22664 2504 22692
rect 2498 22652 2504 22664
rect 2556 22652 2562 22704
rect 5077 22695 5135 22701
rect 5077 22661 5089 22695
rect 5123 22692 5135 22695
rect 5258 22692 5264 22704
rect 5123 22664 5264 22692
rect 5123 22661 5135 22664
rect 5077 22655 5135 22661
rect 5258 22652 5264 22664
rect 5316 22692 5322 22704
rect 5920 22692 5948 22732
rect 8205 22729 8217 22732
rect 8251 22729 8263 22763
rect 8205 22723 8263 22729
rect 8294 22720 8300 22772
rect 8352 22760 8358 22772
rect 8941 22763 8999 22769
rect 8941 22760 8953 22763
rect 8352 22732 8953 22760
rect 8352 22720 8358 22732
rect 8941 22729 8953 22732
rect 8987 22760 8999 22763
rect 9309 22763 9367 22769
rect 9309 22760 9321 22763
rect 8987 22732 9321 22760
rect 8987 22729 8999 22732
rect 8941 22723 8999 22729
rect 9309 22729 9321 22732
rect 9355 22729 9367 22763
rect 10870 22760 10876 22772
rect 10831 22732 10876 22760
rect 9309 22723 9367 22729
rect 5316 22664 5948 22692
rect 5316 22652 5322 22664
rect 2516 22624 2544 22652
rect 2685 22627 2743 22633
rect 2685 22624 2697 22627
rect 2516 22596 2697 22624
rect 2685 22593 2697 22596
rect 2731 22593 2743 22627
rect 2685 22587 2743 22593
rect 5350 22584 5356 22636
rect 5408 22624 5414 22636
rect 5629 22627 5687 22633
rect 5629 22624 5641 22627
rect 5408 22596 5641 22624
rect 5408 22584 5414 22596
rect 5629 22593 5641 22596
rect 5675 22624 5687 22627
rect 5718 22624 5724 22636
rect 5675 22596 5724 22624
rect 5675 22593 5687 22596
rect 5629 22587 5687 22593
rect 5718 22584 5724 22596
rect 5776 22584 5782 22636
rect 5813 22627 5871 22633
rect 5813 22593 5825 22627
rect 5859 22624 5871 22627
rect 5920 22624 5948 22664
rect 5859 22596 5948 22624
rect 9324 22624 9352 22723
rect 10870 22720 10876 22732
rect 10928 22760 10934 22772
rect 11425 22763 11483 22769
rect 11425 22760 11437 22763
rect 10928 22732 11437 22760
rect 10928 22720 10934 22732
rect 11425 22729 11437 22732
rect 11471 22729 11483 22763
rect 11425 22723 11483 22729
rect 11790 22692 11796 22704
rect 11751 22664 11796 22692
rect 11790 22652 11796 22664
rect 11848 22652 11854 22704
rect 9493 22627 9551 22633
rect 9493 22624 9505 22627
rect 9324 22596 9505 22624
rect 5859 22593 5871 22596
rect 5813 22587 5871 22593
rect 9493 22593 9505 22596
rect 9539 22593 9551 22627
rect 9493 22587 9551 22593
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 12584 22596 12940 22624
rect 12584 22584 12590 22596
rect 2952 22559 3010 22565
rect 2952 22525 2964 22559
rect 2998 22556 3010 22559
rect 3234 22556 3240 22568
rect 2998 22528 3240 22556
rect 2998 22525 3010 22528
rect 2952 22519 3010 22525
rect 3234 22516 3240 22528
rect 3292 22516 3298 22568
rect 5534 22556 5540 22568
rect 5495 22528 5540 22556
rect 5534 22516 5540 22528
rect 5592 22516 5598 22568
rect 6822 22556 6828 22568
rect 6564 22528 6828 22556
rect 4798 22448 4804 22500
rect 4856 22488 4862 22500
rect 6178 22488 6184 22500
rect 4856 22460 6184 22488
rect 4856 22448 4862 22460
rect 6178 22448 6184 22460
rect 6236 22448 6242 22500
rect 4706 22420 4712 22432
rect 4667 22392 4712 22420
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5166 22420 5172 22432
rect 5127 22392 5172 22420
rect 5166 22380 5172 22392
rect 5224 22380 5230 22432
rect 5718 22380 5724 22432
rect 5776 22420 5782 22432
rect 6564 22429 6592 22528
rect 6822 22516 6828 22528
rect 6880 22516 6886 22568
rect 6914 22516 6920 22568
rect 6972 22556 6978 22568
rect 7098 22565 7104 22568
rect 7081 22559 7104 22565
rect 7081 22556 7093 22559
rect 6972 22528 7093 22556
rect 6972 22516 6978 22528
rect 7081 22525 7093 22528
rect 7156 22556 7162 22568
rect 12253 22559 12311 22565
rect 7156 22528 7229 22556
rect 7081 22519 7104 22525
rect 7098 22516 7104 22519
rect 7156 22516 7162 22528
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 12710 22556 12716 22568
rect 12299 22528 12716 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 12710 22516 12716 22528
rect 12768 22516 12774 22568
rect 12912 22565 12940 22596
rect 12986 22584 12992 22636
rect 13044 22624 13050 22636
rect 13081 22627 13139 22633
rect 13081 22624 13093 22627
rect 13044 22596 13093 22624
rect 13044 22584 13050 22596
rect 13081 22593 13093 22596
rect 13127 22624 13139 22627
rect 13262 22624 13268 22636
rect 13127 22596 13268 22624
rect 13127 22593 13139 22596
rect 13081 22587 13139 22593
rect 13262 22584 13268 22596
rect 13320 22624 13326 22636
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13320 22596 13829 22624
rect 13320 22584 13326 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 12897 22559 12955 22565
rect 12897 22525 12909 22559
rect 12943 22556 12955 22559
rect 13630 22556 13636 22568
rect 12943 22528 13636 22556
rect 12943 22525 12955 22528
rect 12897 22519 12955 22525
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 9760 22491 9818 22497
rect 9760 22457 9772 22491
rect 9806 22488 9818 22491
rect 9858 22488 9864 22500
rect 9806 22460 9864 22488
rect 9806 22457 9818 22460
rect 9760 22451 9818 22457
rect 9858 22448 9864 22460
rect 9916 22448 9922 22500
rect 12802 22488 12808 22500
rect 12715 22460 12808 22488
rect 12802 22448 12808 22460
rect 12860 22488 12866 22500
rect 13449 22491 13507 22497
rect 13449 22488 13461 22491
rect 12860 22460 13461 22488
rect 12860 22448 12866 22460
rect 13449 22457 13461 22460
rect 13495 22457 13507 22491
rect 13449 22451 13507 22457
rect 6549 22423 6607 22429
rect 6549 22420 6561 22423
rect 5776 22392 6561 22420
rect 5776 22380 5782 22392
rect 6549 22389 6561 22392
rect 6595 22389 6607 22423
rect 12434 22420 12440 22432
rect 12395 22392 12440 22420
rect 6549 22383 6607 22389
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 1104 22330 14812 22352
rect 1104 22278 6315 22330
rect 6367 22278 6379 22330
rect 6431 22278 6443 22330
rect 6495 22278 6507 22330
rect 6559 22278 11648 22330
rect 11700 22278 11712 22330
rect 11764 22278 11776 22330
rect 11828 22278 11840 22330
rect 11892 22278 14812 22330
rect 1104 22256 14812 22278
rect 1670 22216 1676 22228
rect 1631 22188 1676 22216
rect 1670 22176 1676 22188
rect 1728 22176 1734 22228
rect 2777 22219 2835 22225
rect 2777 22185 2789 22219
rect 2823 22216 2835 22219
rect 3234 22216 3240 22228
rect 2823 22188 3240 22216
rect 2823 22185 2835 22188
rect 2777 22179 2835 22185
rect 3234 22176 3240 22188
rect 3292 22176 3298 22228
rect 4798 22216 4804 22228
rect 4759 22188 4804 22216
rect 4798 22176 4804 22188
rect 4856 22176 4862 22228
rect 6178 22176 6184 22228
rect 6236 22216 6242 22228
rect 6365 22219 6423 22225
rect 6365 22216 6377 22219
rect 6236 22188 6377 22216
rect 6236 22176 6242 22188
rect 6365 22185 6377 22188
rect 6411 22185 6423 22219
rect 6365 22179 6423 22185
rect 7466 22176 7472 22228
rect 7524 22216 7530 22228
rect 7561 22219 7619 22225
rect 7561 22216 7573 22219
rect 7524 22188 7573 22216
rect 7524 22176 7530 22188
rect 7561 22185 7573 22188
rect 7607 22185 7619 22219
rect 7561 22179 7619 22185
rect 10045 22219 10103 22225
rect 10045 22185 10057 22219
rect 10091 22216 10103 22219
rect 11241 22219 11299 22225
rect 11241 22216 11253 22219
rect 10091 22188 11253 22216
rect 10091 22185 10103 22188
rect 10045 22179 10103 22185
rect 11241 22185 11253 22188
rect 11287 22185 11299 22219
rect 12802 22216 12808 22228
rect 12763 22188 12808 22216
rect 11241 22179 11299 22185
rect 5258 22157 5264 22160
rect 5252 22148 5264 22157
rect 5219 22120 5264 22148
rect 5252 22111 5264 22120
rect 5258 22108 5264 22111
rect 5316 22108 5322 22160
rect 10060 22148 10088 22179
rect 12802 22176 12808 22188
rect 12860 22176 12866 22228
rect 9600 22120 10088 22148
rect 11701 22151 11759 22157
rect 2409 22083 2467 22089
rect 2409 22049 2421 22083
rect 2455 22080 2467 22083
rect 2866 22080 2872 22092
rect 2455 22052 2872 22080
rect 2455 22049 2467 22052
rect 2409 22043 2467 22049
rect 2866 22040 2872 22052
rect 2924 22040 2930 22092
rect 4706 22040 4712 22092
rect 4764 22080 4770 22092
rect 4985 22083 5043 22089
rect 4985 22080 4997 22083
rect 4764 22052 4997 22080
rect 4764 22040 4770 22052
rect 4985 22049 4997 22052
rect 5031 22080 5043 22083
rect 5718 22080 5724 22092
rect 5031 22052 5724 22080
rect 5031 22049 5043 22052
rect 4985 22043 5043 22049
rect 5718 22040 5724 22052
rect 5776 22040 5782 22092
rect 7926 22080 7932 22092
rect 7887 22052 7932 22080
rect 7926 22040 7932 22052
rect 7984 22040 7990 22092
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22080 9183 22083
rect 9600 22080 9628 22120
rect 11701 22117 11713 22151
rect 11747 22148 11759 22151
rect 12158 22148 12164 22160
rect 11747 22120 12164 22148
rect 11747 22117 11759 22120
rect 11701 22111 11759 22117
rect 12158 22108 12164 22120
rect 12216 22108 12222 22160
rect 9171 22052 9628 22080
rect 11149 22083 11207 22089
rect 9171 22049 9183 22052
rect 9125 22043 9183 22049
rect 11149 22049 11161 22083
rect 11195 22080 11207 22083
rect 11609 22083 11667 22089
rect 11609 22080 11621 22083
rect 11195 22052 11621 22080
rect 11195 22049 11207 22052
rect 11149 22043 11207 22049
rect 11609 22049 11621 22052
rect 11655 22080 11667 22083
rect 12434 22080 12440 22092
rect 11655 22052 12440 22080
rect 11655 22049 11667 22052
rect 11609 22043 11667 22049
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 7469 22015 7527 22021
rect 7469 21981 7481 22015
rect 7515 22012 7527 22015
rect 8018 22012 8024 22024
rect 7515 21984 8024 22012
rect 7515 21981 7527 21984
rect 7469 21975 7527 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 8113 22015 8171 22021
rect 8113 21981 8125 22015
rect 8159 21981 8171 22015
rect 8113 21975 8171 21981
rect 7834 21904 7840 21956
rect 7892 21944 7898 21956
rect 8128 21944 8156 21975
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10137 22015 10195 22021
rect 10137 22012 10149 22015
rect 10100 21984 10149 22012
rect 10100 21972 10106 21984
rect 10137 21981 10149 21984
rect 10183 21981 10195 22015
rect 10137 21975 10195 21981
rect 10226 21972 10232 22024
rect 10284 22012 10290 22024
rect 10284 21984 10329 22012
rect 10284 21972 10290 21984
rect 10594 21972 10600 22024
rect 10652 22012 10658 22024
rect 10778 22012 10784 22024
rect 10652 21984 10784 22012
rect 10652 21972 10658 21984
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 11330 21972 11336 22024
rect 11388 22012 11394 22024
rect 11885 22015 11943 22021
rect 11885 22012 11897 22015
rect 11388 21984 11897 22012
rect 11388 21972 11394 21984
rect 11885 21981 11897 21984
rect 11931 22012 11943 22015
rect 12342 22012 12348 22024
rect 11931 21984 12348 22012
rect 11931 21981 11943 21984
rect 11885 21975 11943 21981
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 7892 21916 8156 21944
rect 9493 21947 9551 21953
rect 7892 21904 7898 21916
rect 9493 21913 9505 21947
rect 9539 21944 9551 21947
rect 9858 21944 9864 21956
rect 9539 21916 9864 21944
rect 9539 21913 9551 21916
rect 9493 21907 9551 21913
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 4433 21879 4491 21885
rect 4433 21845 4445 21879
rect 4479 21876 4491 21879
rect 5350 21876 5356 21888
rect 4479 21848 5356 21876
rect 4479 21845 4491 21848
rect 4433 21839 4491 21845
rect 5350 21836 5356 21848
rect 5408 21836 5414 21888
rect 7098 21876 7104 21888
rect 7059 21848 7104 21876
rect 7098 21836 7104 21848
rect 7156 21836 7162 21888
rect 9674 21876 9680 21888
rect 9635 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 10778 21876 10784 21888
rect 10739 21848 10784 21876
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 12526 21876 12532 21888
rect 12487 21848 12532 21876
rect 12526 21836 12532 21848
rect 12584 21836 12590 21888
rect 1104 21786 14812 21808
rect 1104 21734 3648 21786
rect 3700 21734 3712 21786
rect 3764 21734 3776 21786
rect 3828 21734 3840 21786
rect 3892 21734 8982 21786
rect 9034 21734 9046 21786
rect 9098 21734 9110 21786
rect 9162 21734 9174 21786
rect 9226 21734 14315 21786
rect 14367 21734 14379 21786
rect 14431 21734 14443 21786
rect 14495 21734 14507 21786
rect 14559 21734 14812 21786
rect 1104 21712 14812 21734
rect 1578 21672 1584 21684
rect 1539 21644 1584 21672
rect 1578 21632 1584 21644
rect 1636 21632 1642 21684
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 3145 21675 3203 21681
rect 3145 21672 3157 21675
rect 2924 21644 3157 21672
rect 2924 21632 2930 21644
rect 3145 21641 3157 21644
rect 3191 21641 3203 21675
rect 3145 21635 3203 21641
rect 3510 21632 3516 21684
rect 3568 21672 3574 21684
rect 4709 21675 4767 21681
rect 4709 21672 4721 21675
rect 3568 21644 4721 21672
rect 3568 21632 3574 21644
rect 4709 21641 4721 21644
rect 4755 21641 4767 21675
rect 4709 21635 4767 21641
rect 7377 21675 7435 21681
rect 7377 21641 7389 21675
rect 7423 21672 7435 21675
rect 7834 21672 7840 21684
rect 7423 21644 7840 21672
rect 7423 21641 7435 21644
rect 7377 21635 7435 21641
rect 7834 21632 7840 21644
rect 7892 21632 7898 21684
rect 9769 21675 9827 21681
rect 9769 21641 9781 21675
rect 9815 21672 9827 21675
rect 10226 21672 10232 21684
rect 9815 21644 10232 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 10226 21632 10232 21644
rect 10284 21632 10290 21684
rect 11330 21672 11336 21684
rect 11291 21644 11336 21672
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 12434 21632 12440 21684
rect 12492 21672 12498 21684
rect 12492 21644 12537 21672
rect 12492 21632 12498 21644
rect 6641 21607 6699 21613
rect 6641 21573 6653 21607
rect 6687 21604 6699 21607
rect 7926 21604 7932 21616
rect 6687 21576 7932 21604
rect 6687 21573 6699 21576
rect 6641 21567 6699 21573
rect 7926 21564 7932 21576
rect 7984 21604 7990 21616
rect 8205 21607 8263 21613
rect 8205 21604 8217 21607
rect 7984 21576 8217 21604
rect 7984 21564 7990 21576
rect 8205 21573 8217 21576
rect 8251 21573 8263 21607
rect 8205 21567 8263 21573
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 3697 21539 3755 21545
rect 3697 21536 3709 21539
rect 3292 21508 3709 21536
rect 3292 21496 3298 21508
rect 3697 21505 3709 21508
rect 3743 21505 3755 21539
rect 3697 21499 3755 21505
rect 4798 21496 4804 21548
rect 4856 21536 4862 21548
rect 5261 21539 5319 21545
rect 5261 21536 5273 21539
rect 4856 21508 5273 21536
rect 4856 21496 4862 21508
rect 5261 21505 5273 21508
rect 5307 21505 5319 21539
rect 5261 21499 5319 21505
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21536 7803 21539
rect 8110 21536 8116 21548
rect 7791 21508 8116 21536
rect 7791 21505 7803 21508
rect 7745 21499 7803 21505
rect 8110 21496 8116 21508
rect 8168 21536 8174 21548
rect 8757 21539 8815 21545
rect 8757 21536 8769 21539
rect 8168 21508 8769 21536
rect 8168 21496 8174 21508
rect 8757 21505 8769 21508
rect 8803 21505 8815 21539
rect 8757 21499 8815 21505
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10689 21539 10747 21545
rect 10689 21536 10701 21539
rect 9916 21508 10701 21536
rect 9916 21496 9922 21508
rect 10689 21505 10701 21508
rect 10735 21536 10747 21539
rect 11348 21536 11376 21632
rect 10735 21508 11376 21536
rect 10735 21505 10747 21508
rect 10689 21499 10747 21505
rect 12618 21496 12624 21548
rect 12676 21536 12682 21548
rect 12986 21536 12992 21548
rect 12676 21508 12992 21536
rect 12676 21496 12682 21508
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 1397 21471 1455 21477
rect 1397 21437 1409 21471
rect 1443 21437 1455 21471
rect 1397 21431 1455 21437
rect 3053 21471 3111 21477
rect 3053 21437 3065 21471
rect 3099 21468 3111 21471
rect 3513 21471 3571 21477
rect 3513 21468 3525 21471
rect 3099 21440 3525 21468
rect 3099 21437 3111 21440
rect 3053 21431 3111 21437
rect 3513 21437 3525 21440
rect 3559 21468 3571 21471
rect 4062 21468 4068 21480
rect 3559 21440 4068 21468
rect 3559 21437 3571 21440
rect 3513 21431 3571 21437
rect 1412 21400 1440 21431
rect 4062 21428 4068 21440
rect 4120 21468 4126 21480
rect 4706 21468 4712 21480
rect 4120 21440 4712 21468
rect 4120 21428 4126 21440
rect 4706 21428 4712 21440
rect 4764 21428 4770 21480
rect 10413 21471 10471 21477
rect 10413 21437 10425 21471
rect 10459 21468 10471 21471
rect 10778 21468 10784 21480
rect 10459 21440 10784 21468
rect 10459 21437 10471 21440
rect 10413 21431 10471 21437
rect 10778 21428 10784 21440
rect 10836 21428 10842 21480
rect 11238 21428 11244 21480
rect 11296 21468 11302 21480
rect 12161 21471 12219 21477
rect 12161 21468 12173 21471
rect 11296 21440 12173 21468
rect 11296 21428 11302 21440
rect 12161 21437 12173 21440
rect 12207 21468 12219 21471
rect 12805 21471 12863 21477
rect 12805 21468 12817 21471
rect 12207 21440 12817 21468
rect 12207 21437 12219 21440
rect 12161 21431 12219 21437
rect 12805 21437 12817 21440
rect 12851 21468 12863 21471
rect 13078 21468 13084 21480
rect 12851 21440 13084 21468
rect 12851 21437 12863 21440
rect 12805 21431 12863 21437
rect 13078 21428 13084 21440
rect 13136 21428 13142 21480
rect 1946 21400 1952 21412
rect 1412 21372 1952 21400
rect 1946 21360 1952 21372
rect 2004 21360 2010 21412
rect 4617 21403 4675 21409
rect 4617 21369 4629 21403
rect 4663 21400 4675 21403
rect 8665 21403 8723 21409
rect 8665 21400 8677 21403
rect 4663 21372 5212 21400
rect 4663 21369 4675 21372
rect 4617 21363 4675 21369
rect 3418 21292 3424 21344
rect 3476 21332 3482 21344
rect 3605 21335 3663 21341
rect 3605 21332 3617 21335
rect 3476 21304 3617 21332
rect 3476 21292 3482 21304
rect 3605 21301 3617 21304
rect 3651 21301 3663 21335
rect 5074 21332 5080 21344
rect 5035 21304 5080 21332
rect 3605 21295 3663 21301
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 5184 21341 5212 21372
rect 8036 21372 8677 21400
rect 5169 21335 5227 21341
rect 5169 21301 5181 21335
rect 5215 21332 5227 21335
rect 5350 21332 5356 21344
rect 5215 21304 5356 21332
rect 5215 21301 5227 21304
rect 5169 21295 5227 21301
rect 5350 21292 5356 21304
rect 5408 21292 5414 21344
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 7650 21292 7656 21344
rect 7708 21332 7714 21344
rect 7926 21332 7932 21344
rect 7708 21304 7932 21332
rect 7708 21292 7714 21304
rect 7926 21292 7932 21304
rect 7984 21332 7990 21344
rect 8036 21341 8064 21372
rect 8665 21369 8677 21372
rect 8711 21369 8723 21403
rect 8665 21363 8723 21369
rect 9306 21360 9312 21412
rect 9364 21400 9370 21412
rect 9401 21403 9459 21409
rect 9401 21400 9413 21403
rect 9364 21372 9413 21400
rect 9364 21360 9370 21372
rect 9401 21369 9413 21372
rect 9447 21400 9459 21403
rect 10505 21403 10563 21409
rect 10505 21400 10517 21403
rect 9447 21372 10517 21400
rect 9447 21369 9459 21372
rect 9401 21363 9459 21369
rect 10505 21369 10517 21372
rect 10551 21369 10563 21403
rect 12897 21403 12955 21409
rect 12897 21400 12909 21403
rect 10505 21363 10563 21369
rect 11808 21372 12909 21400
rect 8021 21335 8079 21341
rect 8021 21332 8033 21335
rect 7984 21304 8033 21332
rect 7984 21292 7990 21304
rect 8021 21301 8033 21304
rect 8067 21301 8079 21335
rect 8021 21295 8079 21301
rect 8386 21292 8392 21344
rect 8444 21332 8450 21344
rect 8570 21332 8576 21344
rect 8444 21304 8576 21332
rect 8444 21292 8450 21304
rect 8570 21292 8576 21304
rect 8628 21292 8634 21344
rect 10042 21332 10048 21344
rect 10003 21304 10048 21332
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 11514 21292 11520 21344
rect 11572 21332 11578 21344
rect 11808 21341 11836 21372
rect 12897 21369 12909 21372
rect 12943 21369 12955 21403
rect 12897 21363 12955 21369
rect 11793 21335 11851 21341
rect 11793 21332 11805 21335
rect 11572 21304 11805 21332
rect 11572 21292 11578 21304
rect 11793 21301 11805 21304
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 1104 21242 14812 21264
rect 1104 21190 6315 21242
rect 6367 21190 6379 21242
rect 6431 21190 6443 21242
rect 6495 21190 6507 21242
rect 6559 21190 11648 21242
rect 11700 21190 11712 21242
rect 11764 21190 11776 21242
rect 11828 21190 11840 21242
rect 11892 21190 14812 21242
rect 1104 21168 14812 21190
rect 5169 21131 5227 21137
rect 5169 21097 5181 21131
rect 5215 21128 5227 21131
rect 5258 21128 5264 21140
rect 5215 21100 5264 21128
rect 5215 21097 5227 21100
rect 5169 21091 5227 21097
rect 5258 21088 5264 21100
rect 5316 21088 5322 21140
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 10042 21128 10048 21140
rect 9539 21100 10048 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 10042 21088 10048 21100
rect 10100 21088 10106 21140
rect 10502 21088 10508 21140
rect 10560 21128 10566 21140
rect 10597 21131 10655 21137
rect 10597 21128 10609 21131
rect 10560 21100 10609 21128
rect 10560 21088 10566 21100
rect 10597 21097 10609 21100
rect 10643 21128 10655 21131
rect 10778 21128 10784 21140
rect 10643 21100 10784 21128
rect 10643 21097 10655 21100
rect 10597 21091 10655 21097
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11057 21131 11115 21137
rect 11057 21097 11069 21131
rect 11103 21128 11115 21131
rect 11514 21128 11520 21140
rect 11103 21100 11520 21128
rect 11103 21097 11115 21100
rect 11057 21091 11115 21097
rect 11514 21088 11520 21100
rect 11572 21088 11578 21140
rect 12158 21128 12164 21140
rect 12119 21100 12164 21128
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21060 6975 21063
rect 7098 21060 7104 21072
rect 6963 21032 7104 21060
rect 6963 21029 6975 21032
rect 6917 21023 6975 21029
rect 7098 21020 7104 21032
rect 7156 21060 7162 21072
rect 7742 21060 7748 21072
rect 7156 21032 7748 21060
rect 7156 21020 7162 21032
rect 7742 21020 7748 21032
rect 7800 21020 7806 21072
rect 11422 21060 11428 21072
rect 11383 21032 11428 21060
rect 11422 21020 11428 21032
rect 11480 21020 11486 21072
rect 7006 20952 7012 21004
rect 7064 20992 7070 21004
rect 7190 20992 7196 21004
rect 7064 20964 7196 20992
rect 7064 20952 7070 20964
rect 7190 20952 7196 20964
rect 7248 20992 7254 21004
rect 7469 20995 7527 21001
rect 7469 20992 7481 20995
rect 7248 20964 7481 20992
rect 7248 20952 7254 20964
rect 7469 20961 7481 20964
rect 7515 20961 7527 20995
rect 7469 20955 7527 20961
rect 9858 20952 9864 21004
rect 9916 20992 9922 21004
rect 10045 20995 10103 21001
rect 10045 20992 10057 20995
rect 9916 20964 10057 20992
rect 9916 20952 9922 20964
rect 10045 20961 10057 20964
rect 10091 20961 10103 20995
rect 10045 20955 10103 20961
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 11572 20964 11617 20992
rect 11572 20952 11578 20964
rect 6822 20884 6828 20936
rect 6880 20924 6886 20936
rect 7558 20924 7564 20936
rect 6880 20896 7564 20924
rect 6880 20884 6886 20896
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 7745 20927 7803 20933
rect 7745 20893 7757 20927
rect 7791 20924 7803 20927
rect 7834 20924 7840 20936
rect 7791 20896 7840 20924
rect 7791 20893 7803 20896
rect 7745 20887 7803 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 11606 20924 11612 20936
rect 11567 20896 11612 20924
rect 11606 20884 11612 20896
rect 11664 20884 11670 20936
rect 6549 20859 6607 20865
rect 6549 20825 6561 20859
rect 6595 20856 6607 20859
rect 6914 20856 6920 20868
rect 6595 20828 6920 20856
rect 6595 20825 6607 20828
rect 6549 20819 6607 20825
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 3237 20791 3295 20797
rect 3237 20757 3249 20791
rect 3283 20788 3295 20791
rect 3418 20788 3424 20800
rect 3283 20760 3424 20788
rect 3283 20757 3295 20760
rect 3237 20751 3295 20757
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 3789 20791 3847 20797
rect 3789 20757 3801 20791
rect 3835 20788 3847 20791
rect 4062 20788 4068 20800
rect 3835 20760 4068 20788
rect 3835 20757 3847 20760
rect 3789 20751 3847 20757
rect 4062 20748 4068 20760
rect 4120 20748 4126 20800
rect 4801 20791 4859 20797
rect 4801 20757 4813 20791
rect 4847 20788 4859 20791
rect 5074 20788 5080 20800
rect 4847 20760 5080 20788
rect 4847 20757 4859 20760
rect 4801 20751 4859 20757
rect 5074 20748 5080 20760
rect 5132 20748 5138 20800
rect 7098 20788 7104 20800
rect 7059 20760 7104 20788
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 8297 20791 8355 20797
rect 8297 20757 8309 20791
rect 8343 20788 8355 20791
rect 8386 20788 8392 20800
rect 8343 20760 8392 20788
rect 8343 20757 8355 20760
rect 8297 20751 8355 20757
rect 8386 20748 8392 20760
rect 8444 20748 8450 20800
rect 9125 20791 9183 20797
rect 9125 20757 9137 20791
rect 9171 20788 9183 20791
rect 9398 20788 9404 20800
rect 9171 20760 9404 20788
rect 9171 20757 9183 20760
rect 9125 20751 9183 20757
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 12529 20791 12587 20797
rect 12529 20757 12541 20791
rect 12575 20788 12587 20791
rect 12618 20788 12624 20800
rect 12575 20760 12624 20788
rect 12575 20757 12587 20760
rect 12529 20751 12587 20757
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 1104 20698 14812 20720
rect 1104 20646 3648 20698
rect 3700 20646 3712 20698
rect 3764 20646 3776 20698
rect 3828 20646 3840 20698
rect 3892 20646 8982 20698
rect 9034 20646 9046 20698
rect 9098 20646 9110 20698
rect 9162 20646 9174 20698
rect 9226 20646 14315 20698
rect 14367 20646 14379 20698
rect 14431 20646 14443 20698
rect 14495 20646 14507 20698
rect 14559 20646 14812 20698
rect 1104 20624 14812 20646
rect 5534 20544 5540 20596
rect 5592 20584 5598 20596
rect 6825 20587 6883 20593
rect 6825 20584 6837 20587
rect 5592 20556 6837 20584
rect 5592 20544 5598 20556
rect 6825 20553 6837 20556
rect 6871 20553 6883 20587
rect 6825 20547 6883 20553
rect 9033 20587 9091 20593
rect 9033 20553 9045 20587
rect 9079 20584 9091 20587
rect 9306 20584 9312 20596
rect 9079 20556 9312 20584
rect 9079 20553 9091 20556
rect 9033 20547 9091 20553
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 6273 20519 6331 20525
rect 6273 20485 6285 20519
rect 6319 20516 6331 20519
rect 6638 20516 6644 20528
rect 6319 20488 6644 20516
rect 6319 20485 6331 20488
rect 6273 20479 6331 20485
rect 6638 20476 6644 20488
rect 6696 20516 6702 20528
rect 7834 20516 7840 20528
rect 6696 20488 7840 20516
rect 6696 20476 6702 20488
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 9398 20476 9404 20528
rect 9456 20516 9462 20528
rect 10597 20519 10655 20525
rect 10597 20516 10609 20519
rect 9456 20488 10609 20516
rect 9456 20476 9462 20488
rect 10597 20485 10609 20488
rect 10643 20485 10655 20519
rect 10597 20479 10655 20485
rect 4249 20451 4307 20457
rect 4249 20448 4261 20451
rect 3988 20420 4261 20448
rect 3988 20392 4016 20420
rect 4249 20417 4261 20420
rect 4295 20417 4307 20451
rect 4249 20411 4307 20417
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7285 20451 7343 20457
rect 7285 20448 7297 20451
rect 7156 20420 7297 20448
rect 7156 20408 7162 20420
rect 7285 20417 7297 20420
rect 7331 20417 7343 20451
rect 7285 20411 7343 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20448 7527 20451
rect 7742 20448 7748 20460
rect 7515 20420 7748 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 3605 20383 3663 20389
rect 3605 20349 3617 20383
rect 3651 20380 3663 20383
rect 3970 20380 3976 20392
rect 3651 20352 3976 20380
rect 3651 20349 3663 20352
rect 3605 20343 3663 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7193 20383 7251 20389
rect 7193 20380 7205 20383
rect 6972 20352 7205 20380
rect 6972 20340 6978 20352
rect 7193 20349 7205 20352
rect 7239 20349 7251 20383
rect 7300 20380 7328 20411
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 8941 20451 8999 20457
rect 8941 20417 8953 20451
rect 8987 20448 8999 20451
rect 9582 20448 9588 20460
rect 8987 20420 9588 20448
rect 8987 20417 8999 20420
rect 8941 20411 8999 20417
rect 9582 20408 9588 20420
rect 9640 20408 9646 20460
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 10520 20420 11161 20448
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 7300 20352 8217 20380
rect 7193 20343 7251 20349
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 9398 20380 9404 20392
rect 9359 20352 9404 20380
rect 8205 20343 8263 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 10520 20324 10548 20420
rect 11149 20417 11161 20420
rect 11195 20448 11207 20451
rect 11606 20448 11612 20460
rect 11195 20420 11612 20448
rect 11195 20417 11207 20420
rect 11149 20411 11207 20417
rect 11606 20408 11612 20420
rect 11664 20448 11670 20460
rect 11977 20451 12035 20457
rect 11977 20448 11989 20451
rect 11664 20420 11989 20448
rect 11664 20408 11670 20420
rect 11977 20417 11989 20420
rect 12023 20417 12035 20451
rect 11977 20411 12035 20417
rect 10778 20340 10784 20392
rect 10836 20380 10842 20392
rect 10965 20383 11023 20389
rect 10965 20380 10977 20383
rect 10836 20352 10977 20380
rect 10836 20340 10842 20352
rect 10965 20349 10977 20352
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 5721 20315 5779 20321
rect 5721 20281 5733 20315
rect 5767 20312 5779 20315
rect 7006 20312 7012 20324
rect 5767 20284 7012 20312
rect 5767 20281 5779 20284
rect 5721 20275 5779 20281
rect 7006 20272 7012 20284
rect 7064 20272 7070 20324
rect 10137 20315 10195 20321
rect 10137 20281 10149 20315
rect 10183 20312 10195 20315
rect 10502 20312 10508 20324
rect 10183 20284 10508 20312
rect 10183 20281 10195 20284
rect 10137 20275 10195 20281
rect 10502 20272 10508 20284
rect 10560 20272 10566 20324
rect 11057 20315 11115 20321
rect 11057 20312 11069 20315
rect 10888 20284 11069 20312
rect 3602 20204 3608 20256
rect 3660 20244 3666 20256
rect 3697 20247 3755 20253
rect 3697 20244 3709 20247
rect 3660 20216 3709 20244
rect 3660 20204 3666 20216
rect 3697 20213 3709 20216
rect 3743 20213 3755 20247
rect 4062 20244 4068 20256
rect 4023 20216 4068 20244
rect 3697 20207 3755 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4212 20216 4257 20244
rect 4212 20204 4218 20216
rect 6178 20204 6184 20256
rect 6236 20244 6242 20256
rect 6549 20247 6607 20253
rect 6549 20244 6561 20247
rect 6236 20216 6561 20244
rect 6236 20204 6242 20216
rect 6549 20213 6561 20216
rect 6595 20244 6607 20247
rect 6822 20244 6828 20256
rect 6595 20216 6828 20244
rect 6595 20213 6607 20216
rect 6549 20207 6607 20213
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7190 20204 7196 20256
rect 7248 20244 7254 20256
rect 7837 20247 7895 20253
rect 7837 20244 7849 20247
rect 7248 20216 7849 20244
rect 7248 20204 7254 20216
rect 7837 20213 7849 20216
rect 7883 20213 7895 20247
rect 7837 20207 7895 20213
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 9548 20216 9593 20244
rect 9548 20204 9554 20216
rect 10226 20204 10232 20256
rect 10284 20244 10290 20256
rect 10413 20247 10471 20253
rect 10413 20244 10425 20247
rect 10284 20216 10425 20244
rect 10284 20204 10290 20216
rect 10413 20213 10425 20216
rect 10459 20244 10471 20247
rect 10888 20244 10916 20284
rect 11057 20281 11069 20284
rect 11103 20281 11115 20315
rect 11057 20275 11115 20281
rect 10459 20216 10916 20244
rect 10459 20213 10471 20216
rect 10413 20207 10471 20213
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11572 20216 11621 20244
rect 11572 20204 11578 20216
rect 11609 20213 11621 20216
rect 11655 20213 11667 20247
rect 11609 20207 11667 20213
rect 1104 20154 14812 20176
rect 1104 20102 6315 20154
rect 6367 20102 6379 20154
rect 6431 20102 6443 20154
rect 6495 20102 6507 20154
rect 6559 20102 11648 20154
rect 11700 20102 11712 20154
rect 11764 20102 11776 20154
rect 11828 20102 11840 20154
rect 11892 20102 14812 20154
rect 1104 20080 14812 20102
rect 3789 20043 3847 20049
rect 3789 20009 3801 20043
rect 3835 20040 3847 20043
rect 4154 20040 4160 20052
rect 3835 20012 4160 20040
rect 3835 20009 3847 20012
rect 3789 20003 3847 20009
rect 4154 20000 4160 20012
rect 4212 20040 4218 20052
rect 4525 20043 4583 20049
rect 4525 20040 4537 20043
rect 4212 20012 4537 20040
rect 4212 20000 4218 20012
rect 4525 20009 4537 20012
rect 4571 20009 4583 20043
rect 4890 20040 4896 20052
rect 4851 20012 4896 20040
rect 4525 20003 4583 20009
rect 4890 20000 4896 20012
rect 4948 20000 4954 20052
rect 7742 20040 7748 20052
rect 7703 20012 7748 20040
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9490 20040 9496 20052
rect 9171 20012 9496 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9490 20000 9496 20012
rect 9548 20040 9554 20052
rect 9953 20043 10011 20049
rect 9953 20040 9965 20043
rect 9548 20012 9965 20040
rect 9548 20000 9554 20012
rect 9953 20009 9965 20012
rect 9999 20009 10011 20043
rect 9953 20003 10011 20009
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10686 20040 10692 20052
rect 10100 20012 10692 20040
rect 10100 20000 10106 20012
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 11146 20040 11152 20052
rect 11059 20012 11152 20040
rect 11146 20000 11152 20012
rect 11204 20040 11210 20052
rect 11422 20040 11428 20052
rect 11204 20012 11428 20040
rect 11204 20000 11210 20012
rect 11422 20000 11428 20012
rect 11480 20000 11486 20052
rect 12618 20000 12624 20052
rect 12676 20040 12682 20052
rect 12897 20043 12955 20049
rect 12897 20040 12909 20043
rect 12676 20012 12909 20040
rect 12676 20000 12682 20012
rect 12897 20009 12909 20012
rect 12943 20009 12955 20043
rect 12897 20003 12955 20009
rect 6638 19981 6644 19984
rect 6632 19972 6644 19981
rect 6599 19944 6644 19972
rect 6632 19935 6644 19944
rect 6638 19932 6644 19935
rect 6696 19932 6702 19984
rect 10410 19932 10416 19984
rect 10468 19932 10474 19984
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 6365 19907 6423 19913
rect 6365 19904 6377 19907
rect 5868 19876 6377 19904
rect 5868 19864 5874 19876
rect 6365 19873 6377 19876
rect 6411 19873 6423 19907
rect 6365 19867 6423 19873
rect 9950 19864 9956 19916
rect 10008 19904 10014 19916
rect 10321 19907 10379 19913
rect 10321 19904 10333 19907
rect 10008 19876 10333 19904
rect 10008 19864 10014 19876
rect 10321 19873 10333 19876
rect 10367 19904 10379 19907
rect 10428 19904 10456 19932
rect 11790 19913 11796 19916
rect 11784 19904 11796 19913
rect 10367 19876 10456 19904
rect 11751 19876 11796 19904
rect 10367 19873 10379 19876
rect 10321 19867 10379 19873
rect 11784 19867 11796 19876
rect 11790 19864 11796 19867
rect 11848 19864 11854 19916
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 4985 19839 5043 19845
rect 4985 19836 4997 19839
rect 4764 19808 4997 19836
rect 4764 19796 4770 19808
rect 4985 19805 4997 19808
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19805 5135 19839
rect 10410 19836 10416 19848
rect 10371 19808 10416 19836
rect 5077 19799 5135 19805
rect 4522 19728 4528 19780
rect 4580 19768 4586 19780
rect 5092 19768 5120 19799
rect 10410 19796 10416 19808
rect 10468 19796 10474 19848
rect 10502 19796 10508 19848
rect 10560 19836 10566 19848
rect 10560 19808 10605 19836
rect 10560 19796 10566 19808
rect 10962 19796 10968 19848
rect 11020 19836 11026 19848
rect 11422 19836 11428 19848
rect 11020 19808 11428 19836
rect 11020 19796 11026 19808
rect 11422 19796 11428 19808
rect 11480 19836 11486 19848
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 11480 19808 11529 19836
rect 11480 19796 11486 19808
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 4580 19740 5120 19768
rect 4580 19728 4586 19740
rect 1104 19610 14812 19632
rect 1104 19558 3648 19610
rect 3700 19558 3712 19610
rect 3764 19558 3776 19610
rect 3828 19558 3840 19610
rect 3892 19558 8982 19610
rect 9034 19558 9046 19610
rect 9098 19558 9110 19610
rect 9162 19558 9174 19610
rect 9226 19558 14315 19610
rect 14367 19558 14379 19610
rect 14431 19558 14443 19610
rect 14495 19558 14507 19610
rect 14559 19558 14812 19610
rect 1104 19536 14812 19558
rect 6089 19499 6147 19505
rect 6089 19465 6101 19499
rect 6135 19496 6147 19499
rect 6638 19496 6644 19508
rect 6135 19468 6644 19496
rect 6135 19465 6147 19468
rect 6089 19459 6147 19465
rect 6638 19456 6644 19468
rect 6696 19456 6702 19508
rect 6914 19456 6920 19508
rect 6972 19496 6978 19508
rect 7193 19499 7251 19505
rect 7193 19496 7205 19499
rect 6972 19468 7205 19496
rect 6972 19456 6978 19468
rect 7193 19465 7205 19468
rect 7239 19465 7251 19499
rect 10502 19496 10508 19508
rect 10463 19468 10508 19496
rect 7193 19459 7251 19465
rect 10502 19456 10508 19468
rect 10560 19496 10566 19508
rect 11057 19499 11115 19505
rect 11057 19496 11069 19499
rect 10560 19468 11069 19496
rect 10560 19456 10566 19468
rect 11057 19465 11069 19468
rect 11103 19496 11115 19499
rect 11790 19496 11796 19508
rect 11103 19468 11796 19496
rect 11103 19465 11115 19468
rect 11057 19459 11115 19465
rect 11790 19456 11796 19468
rect 11848 19496 11854 19508
rect 11885 19499 11943 19505
rect 11885 19496 11897 19499
rect 11848 19468 11897 19496
rect 11848 19456 11854 19468
rect 11885 19465 11897 19468
rect 11931 19465 11943 19499
rect 11885 19459 11943 19465
rect 4614 19320 4620 19372
rect 4672 19360 4678 19372
rect 4982 19360 4988 19372
rect 4672 19332 4988 19360
rect 4672 19320 4678 19332
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 5718 19360 5724 19372
rect 5684 19332 5724 19360
rect 5684 19320 5690 19332
rect 5718 19320 5724 19332
rect 5776 19320 5782 19372
rect 7834 19360 7840 19372
rect 7795 19332 7840 19360
rect 7834 19320 7840 19332
rect 7892 19320 7898 19372
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 11146 19360 11152 19372
rect 10836 19332 11152 19360
rect 10836 19320 10842 19332
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11422 19320 11428 19372
rect 11480 19360 11486 19372
rect 11517 19363 11575 19369
rect 11517 19360 11529 19363
rect 11480 19332 11529 19360
rect 11480 19320 11486 19332
rect 11517 19329 11529 19332
rect 11563 19329 11575 19363
rect 11517 19323 11575 19329
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 12066 19360 12072 19372
rect 12032 19332 12072 19360
rect 12032 19320 12038 19332
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 13354 19320 13360 19372
rect 13412 19360 13418 19372
rect 13446 19360 13452 19372
rect 13412 19332 13452 19360
rect 13412 19320 13418 19332
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19292 2835 19295
rect 2869 19295 2927 19301
rect 2869 19292 2881 19295
rect 2823 19264 2881 19292
rect 2823 19261 2835 19264
rect 2777 19255 2835 19261
rect 2869 19261 2881 19264
rect 2915 19292 2927 19295
rect 2915 19264 5764 19292
rect 2915 19261 2927 19264
rect 2869 19255 2927 19261
rect 5736 19236 5764 19264
rect 7006 19252 7012 19304
rect 7064 19292 7070 19304
rect 7561 19295 7619 19301
rect 7561 19292 7573 19295
rect 7064 19264 7573 19292
rect 7064 19252 7070 19264
rect 7561 19261 7573 19264
rect 7607 19261 7619 19295
rect 7561 19255 7619 19261
rect 8202 19252 8208 19304
rect 8260 19292 8266 19304
rect 8386 19292 8392 19304
rect 8260 19264 8392 19292
rect 8260 19252 8266 19264
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 9033 19295 9091 19301
rect 9033 19261 9045 19295
rect 9079 19292 9091 19295
rect 9122 19292 9128 19304
rect 9079 19264 9128 19292
rect 9079 19261 9091 19264
rect 9033 19255 9091 19261
rect 9122 19252 9128 19264
rect 9180 19252 9186 19304
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 3114 19227 3172 19233
rect 3114 19224 3126 19227
rect 3016 19196 3126 19224
rect 3016 19184 3022 19196
rect 3114 19193 3126 19196
rect 3160 19193 3172 19227
rect 3114 19187 3172 19193
rect 3970 19184 3976 19236
rect 4028 19224 4034 19236
rect 4614 19224 4620 19236
rect 4028 19196 4620 19224
rect 4028 19184 4034 19196
rect 4264 19165 4292 19196
rect 4614 19184 4620 19196
rect 4672 19184 4678 19236
rect 4706 19184 4712 19236
rect 4764 19224 4770 19236
rect 5169 19227 5227 19233
rect 5169 19224 5181 19227
rect 4764 19196 5181 19224
rect 4764 19184 4770 19196
rect 5169 19193 5181 19196
rect 5215 19193 5227 19227
rect 5169 19187 5227 19193
rect 5718 19184 5724 19236
rect 5776 19224 5782 19236
rect 6457 19227 6515 19233
rect 6457 19224 6469 19227
rect 5776 19196 6469 19224
rect 5776 19184 5782 19196
rect 6457 19193 6469 19196
rect 6503 19224 6515 19227
rect 8110 19224 8116 19236
rect 6503 19196 8116 19224
rect 6503 19193 6515 19196
rect 6457 19187 6515 19193
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 9306 19184 9312 19236
rect 9364 19233 9370 19236
rect 9364 19227 9428 19233
rect 9364 19193 9382 19227
rect 9416 19193 9428 19227
rect 9364 19187 9428 19193
rect 9364 19184 9370 19187
rect 4249 19159 4307 19165
rect 4249 19125 4261 19159
rect 4295 19125 4307 19159
rect 4890 19156 4896 19168
rect 4851 19128 4896 19156
rect 4249 19119 4307 19125
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5353 19159 5411 19165
rect 5353 19156 5365 19159
rect 5316 19128 5365 19156
rect 5316 19116 5322 19128
rect 5353 19125 5365 19128
rect 5399 19125 5411 19159
rect 7098 19156 7104 19168
rect 7059 19128 7104 19156
rect 5353 19119 5411 19125
rect 7098 19116 7104 19128
rect 7156 19156 7162 19168
rect 7650 19156 7656 19168
rect 7156 19128 7656 19156
rect 7156 19116 7162 19128
rect 7650 19116 7656 19128
rect 7708 19116 7714 19168
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8386 19156 8392 19168
rect 8343 19128 8392 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 8754 19116 8760 19168
rect 8812 19156 8818 19168
rect 9490 19156 9496 19168
rect 8812 19128 9496 19156
rect 8812 19116 8818 19128
rect 9490 19116 9496 19128
rect 9548 19116 9554 19168
rect 1104 19066 14812 19088
rect 1104 19014 6315 19066
rect 6367 19014 6379 19066
rect 6431 19014 6443 19066
rect 6495 19014 6507 19066
rect 6559 19014 11648 19066
rect 11700 19014 11712 19066
rect 11764 19014 11776 19066
rect 11828 19014 11840 19066
rect 11892 19014 14812 19066
rect 1104 18992 14812 19014
rect 3970 18912 3976 18964
rect 4028 18952 4034 18964
rect 4890 18952 4896 18964
rect 4028 18924 4896 18952
rect 4028 18912 4034 18924
rect 4890 18912 4896 18924
rect 4948 18912 4954 18964
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7193 18955 7251 18961
rect 7193 18952 7205 18955
rect 7064 18924 7205 18952
rect 7064 18912 7070 18924
rect 7193 18921 7205 18924
rect 7239 18921 7251 18955
rect 7193 18915 7251 18921
rect 7653 18955 7711 18961
rect 7653 18921 7665 18955
rect 7699 18952 7711 18955
rect 7834 18952 7840 18964
rect 7699 18924 7840 18952
rect 7699 18921 7711 18924
rect 7653 18915 7711 18921
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 5718 18884 5724 18896
rect 4908 18856 5724 18884
rect 4908 18828 4936 18856
rect 5718 18844 5724 18856
rect 5776 18844 5782 18896
rect 4890 18816 4896 18828
rect 4803 18788 4896 18816
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 5160 18819 5218 18825
rect 5160 18785 5172 18819
rect 5206 18816 5218 18819
rect 5534 18816 5540 18828
rect 5206 18788 5540 18816
rect 5206 18785 5218 18788
rect 5160 18779 5218 18785
rect 5534 18776 5540 18788
rect 5592 18776 5598 18828
rect 8386 18816 8392 18828
rect 8347 18788 8392 18816
rect 8386 18776 8392 18788
rect 8444 18776 8450 18828
rect 8478 18748 8484 18760
rect 8439 18720 8484 18748
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8628 18720 8673 18748
rect 8628 18708 8634 18720
rect 9950 18708 9956 18760
rect 10008 18748 10014 18760
rect 10321 18751 10379 18757
rect 10321 18748 10333 18751
rect 10008 18720 10333 18748
rect 10008 18708 10014 18720
rect 10321 18717 10333 18720
rect 10367 18717 10379 18751
rect 10321 18711 10379 18717
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18612 3022 18624
rect 4522 18612 4528 18624
rect 3016 18584 4528 18612
rect 3016 18572 3022 18584
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 6270 18612 6276 18624
rect 6231 18584 6276 18612
rect 6270 18572 6276 18584
rect 6328 18572 6334 18624
rect 8018 18612 8024 18624
rect 7979 18584 8024 18612
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 9217 18615 9275 18621
rect 9217 18581 9229 18615
rect 9263 18612 9275 18615
rect 9306 18612 9312 18624
rect 9263 18584 9312 18612
rect 9263 18581 9275 18584
rect 9217 18575 9275 18581
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 10045 18615 10103 18621
rect 10045 18581 10057 18615
rect 10091 18612 10103 18615
rect 10410 18612 10416 18624
rect 10091 18584 10416 18612
rect 10091 18581 10103 18584
rect 10045 18575 10103 18581
rect 10410 18572 10416 18584
rect 10468 18572 10474 18624
rect 1104 18522 14812 18544
rect 1104 18470 3648 18522
rect 3700 18470 3712 18522
rect 3764 18470 3776 18522
rect 3828 18470 3840 18522
rect 3892 18470 8982 18522
rect 9034 18470 9046 18522
rect 9098 18470 9110 18522
rect 9162 18470 9174 18522
rect 9226 18470 14315 18522
rect 14367 18470 14379 18522
rect 14431 18470 14443 18522
rect 14495 18470 14507 18522
rect 14559 18470 14812 18522
rect 1104 18448 14812 18470
rect 1578 18408 1584 18420
rect 1539 18380 1584 18408
rect 1578 18368 1584 18380
rect 1636 18368 1642 18420
rect 4154 18368 4160 18420
rect 4212 18408 4218 18420
rect 4801 18411 4859 18417
rect 4801 18408 4813 18411
rect 4212 18380 4813 18408
rect 4212 18368 4218 18380
rect 4801 18377 4813 18380
rect 4847 18377 4859 18411
rect 4801 18371 4859 18377
rect 4341 18343 4399 18349
rect 4341 18309 4353 18343
rect 4387 18340 4399 18343
rect 4890 18340 4896 18352
rect 4387 18312 4896 18340
rect 4387 18309 4399 18312
rect 4341 18303 4399 18309
rect 4890 18300 4896 18312
rect 4948 18300 4954 18352
rect 4522 18232 4528 18284
rect 4580 18272 4586 18284
rect 5353 18275 5411 18281
rect 5353 18272 5365 18275
rect 4580 18244 5365 18272
rect 4580 18232 4586 18244
rect 5353 18241 5365 18244
rect 5399 18272 5411 18275
rect 6181 18275 6239 18281
rect 6181 18272 6193 18275
rect 5399 18244 6193 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 6181 18241 6193 18244
rect 6227 18272 6239 18275
rect 6270 18272 6276 18284
rect 6227 18244 6276 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 6270 18232 6276 18244
rect 6328 18232 6334 18284
rect 1397 18207 1455 18213
rect 1397 18173 1409 18207
rect 1443 18204 1455 18207
rect 3973 18207 4031 18213
rect 1443 18176 1992 18204
rect 1443 18173 1455 18176
rect 1397 18167 1455 18173
rect 1964 18080 1992 18176
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 5169 18207 5227 18213
rect 5169 18204 5181 18207
rect 4019 18176 5181 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 5169 18173 5181 18176
rect 5215 18204 5227 18207
rect 5258 18204 5264 18216
rect 5215 18176 5264 18204
rect 5215 18173 5227 18176
rect 5169 18167 5227 18173
rect 5258 18164 5264 18176
rect 5316 18164 5322 18216
rect 7929 18207 7987 18213
rect 7929 18173 7941 18207
rect 7975 18204 7987 18207
rect 8021 18207 8079 18213
rect 8021 18204 8033 18207
rect 7975 18176 8033 18204
rect 7975 18173 7987 18176
rect 7929 18167 7987 18173
rect 8021 18173 8033 18176
rect 8067 18204 8079 18207
rect 8110 18204 8116 18216
rect 8067 18176 8116 18204
rect 8067 18173 8079 18176
rect 8021 18167 8079 18173
rect 8110 18164 8116 18176
rect 8168 18164 8174 18216
rect 8570 18164 8576 18216
rect 8628 18164 8634 18216
rect 7193 18139 7251 18145
rect 7193 18105 7205 18139
rect 7239 18136 7251 18139
rect 7561 18139 7619 18145
rect 7561 18136 7573 18139
rect 7239 18108 7573 18136
rect 7239 18105 7251 18108
rect 7193 18099 7251 18105
rect 7561 18105 7573 18108
rect 7607 18136 7619 18139
rect 8288 18139 8346 18145
rect 8288 18136 8300 18139
rect 7607 18108 8300 18136
rect 7607 18105 7619 18108
rect 7561 18099 7619 18105
rect 8288 18105 8300 18108
rect 8334 18136 8346 18139
rect 8588 18136 8616 18164
rect 9214 18136 9220 18148
rect 8334 18108 9220 18136
rect 8334 18105 8346 18108
rect 8288 18099 8346 18105
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 1946 18068 1952 18080
rect 1907 18040 1952 18068
rect 1946 18028 1952 18040
rect 2004 18028 2010 18080
rect 4430 18028 4436 18080
rect 4488 18068 4494 18080
rect 4709 18071 4767 18077
rect 4709 18068 4721 18071
rect 4488 18040 4721 18068
rect 4488 18028 4494 18040
rect 4709 18037 4721 18040
rect 4755 18068 4767 18071
rect 5258 18068 5264 18080
rect 4755 18040 5264 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 5534 18028 5540 18080
rect 5592 18068 5598 18080
rect 5813 18071 5871 18077
rect 5813 18068 5825 18071
rect 5592 18040 5825 18068
rect 5592 18028 5598 18040
rect 5813 18037 5825 18040
rect 5859 18037 5871 18071
rect 5813 18031 5871 18037
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 9306 18068 9312 18080
rect 8628 18040 9312 18068
rect 8628 18028 8634 18040
rect 9306 18028 9312 18040
rect 9364 18068 9370 18080
rect 9401 18071 9459 18077
rect 9401 18068 9413 18071
rect 9364 18040 9413 18068
rect 9364 18028 9370 18040
rect 9401 18037 9413 18040
rect 9447 18037 9459 18071
rect 9401 18031 9459 18037
rect 1104 17978 14812 18000
rect 1104 17926 6315 17978
rect 6367 17926 6379 17978
rect 6431 17926 6443 17978
rect 6495 17926 6507 17978
rect 6559 17926 11648 17978
rect 11700 17926 11712 17978
rect 11764 17926 11776 17978
rect 11828 17926 11840 17978
rect 11892 17926 14812 17978
rect 1104 17904 14812 17926
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 5166 17864 5172 17876
rect 4120 17836 5172 17864
rect 4120 17824 4126 17836
rect 5166 17824 5172 17836
rect 5224 17864 5230 17876
rect 5261 17867 5319 17873
rect 5261 17864 5273 17867
rect 5224 17836 5273 17864
rect 5224 17824 5230 17836
rect 5261 17833 5273 17836
rect 5307 17833 5319 17867
rect 7742 17864 7748 17876
rect 7703 17836 7748 17864
rect 5261 17827 5319 17833
rect 7742 17824 7748 17836
rect 7800 17824 7806 17876
rect 8018 17824 8024 17876
rect 8076 17864 8082 17876
rect 8205 17867 8263 17873
rect 8205 17864 8217 17867
rect 8076 17836 8217 17864
rect 8076 17824 8082 17836
rect 8205 17833 8217 17836
rect 8251 17833 8263 17867
rect 8205 17827 8263 17833
rect 8110 17728 8116 17740
rect 8071 17700 8116 17728
rect 8110 17688 8116 17700
rect 8168 17688 8174 17740
rect 9766 17688 9772 17740
rect 9824 17728 9830 17740
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9824 17700 10057 17728
rect 9824 17688 9830 17700
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 11422 17688 11428 17740
rect 11480 17728 11486 17740
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11480 17700 11621 17728
rect 11480 17688 11486 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 11876 17731 11934 17737
rect 11876 17697 11888 17731
rect 11922 17728 11934 17731
rect 12158 17728 12164 17740
rect 11922 17700 12164 17728
rect 11922 17697 11934 17700
rect 11876 17691 11934 17697
rect 12158 17688 12164 17700
rect 12216 17688 12222 17740
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 4304 17632 5365 17660
rect 4304 17620 4310 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5534 17660 5540 17672
rect 5495 17632 5540 17660
rect 5353 17623 5411 17629
rect 5534 17620 5540 17632
rect 5592 17620 5598 17672
rect 7926 17620 7932 17672
rect 7984 17660 7990 17672
rect 8297 17663 8355 17669
rect 8297 17660 8309 17663
rect 7984 17632 8309 17660
rect 7984 17620 7990 17632
rect 8297 17629 8309 17632
rect 8343 17660 8355 17663
rect 8570 17660 8576 17672
rect 8343 17632 8576 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 8570 17620 8576 17632
rect 8628 17620 8634 17672
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10229 17663 10287 17669
rect 10229 17629 10241 17663
rect 10275 17629 10287 17663
rect 10229 17623 10287 17629
rect 2774 17552 2780 17604
rect 2832 17592 2838 17604
rect 4893 17595 4951 17601
rect 4893 17592 4905 17595
rect 2832 17564 4905 17592
rect 2832 17552 2838 17564
rect 4893 17561 4905 17564
rect 4939 17561 4951 17595
rect 4893 17555 4951 17561
rect 7653 17595 7711 17601
rect 7653 17561 7665 17595
rect 7699 17592 7711 17595
rect 8478 17592 8484 17604
rect 7699 17564 8484 17592
rect 7699 17561 7711 17564
rect 7653 17555 7711 17561
rect 8478 17552 8484 17564
rect 8536 17592 8542 17604
rect 9677 17595 9735 17601
rect 9677 17592 9689 17595
rect 8536 17564 9689 17592
rect 8536 17552 8542 17564
rect 9677 17561 9689 17564
rect 9723 17561 9735 17595
rect 9677 17555 9735 17561
rect 3053 17527 3111 17533
rect 3053 17493 3065 17527
rect 3099 17524 3111 17527
rect 3418 17524 3424 17536
rect 3099 17496 3424 17524
rect 3099 17493 3111 17496
rect 3053 17487 3111 17493
rect 3418 17484 3424 17496
rect 3476 17484 3482 17536
rect 6914 17524 6920 17536
rect 6875 17496 6920 17524
rect 6914 17484 6920 17496
rect 6972 17484 6978 17536
rect 7285 17527 7343 17533
rect 7285 17493 7297 17527
rect 7331 17524 7343 17527
rect 7374 17524 7380 17536
rect 7331 17496 7380 17524
rect 7331 17493 7343 17496
rect 7285 17487 7343 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 8757 17527 8815 17533
rect 8757 17524 8769 17527
rect 8628 17496 8769 17524
rect 8628 17484 8634 17496
rect 8757 17493 8769 17496
rect 8803 17524 8815 17527
rect 10244 17524 10272 17623
rect 10686 17524 10692 17536
rect 8803 17496 10272 17524
rect 10647 17496 10692 17524
rect 8803 17493 8815 17496
rect 8757 17487 8815 17493
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 12986 17524 12992 17536
rect 12947 17496 12992 17524
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 1104 17434 14812 17456
rect 1104 17382 3648 17434
rect 3700 17382 3712 17434
rect 3764 17382 3776 17434
rect 3828 17382 3840 17434
rect 3892 17382 8982 17434
rect 9034 17382 9046 17434
rect 9098 17382 9110 17434
rect 9162 17382 9174 17434
rect 9226 17382 14315 17434
rect 14367 17382 14379 17434
rect 14431 17382 14443 17434
rect 14495 17382 14507 17434
rect 14559 17382 14812 17434
rect 1104 17360 14812 17382
rect 4062 17320 4068 17332
rect 4023 17292 4068 17320
rect 4062 17280 4068 17292
rect 4120 17280 4126 17332
rect 4246 17280 4252 17332
rect 4304 17320 4310 17332
rect 4341 17323 4399 17329
rect 4341 17320 4353 17323
rect 4304 17292 4353 17320
rect 4304 17280 4310 17292
rect 4341 17289 4353 17292
rect 4387 17289 4399 17323
rect 7926 17320 7932 17332
rect 7887 17292 7932 17320
rect 4341 17283 4399 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8573 17323 8631 17329
rect 8573 17320 8585 17323
rect 8444 17292 8585 17320
rect 8444 17280 8450 17292
rect 8573 17289 8585 17292
rect 8619 17289 8631 17323
rect 10134 17320 10140 17332
rect 10095 17292 10140 17320
rect 8573 17283 8631 17289
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 11422 17280 11428 17332
rect 11480 17320 11486 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 11480 17292 11621 17320
rect 11480 17280 11486 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 2682 17212 2688 17264
rect 2740 17252 2746 17264
rect 2961 17255 3019 17261
rect 2961 17252 2973 17255
rect 2740 17224 2973 17252
rect 2740 17212 2746 17224
rect 2961 17221 2973 17224
rect 3007 17221 3019 17255
rect 2961 17215 3019 17221
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 6086 17252 6092 17264
rect 5960 17224 6092 17252
rect 5960 17212 5966 17224
rect 6086 17212 6092 17224
rect 6144 17212 6150 17264
rect 10042 17252 10048 17264
rect 10003 17224 10048 17252
rect 10042 17212 10048 17224
rect 10100 17212 10106 17264
rect 3418 17184 3424 17196
rect 3379 17156 3424 17184
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 3513 17187 3571 17193
rect 3513 17153 3525 17187
rect 3559 17153 3571 17187
rect 5534 17184 5540 17196
rect 5447 17156 5540 17184
rect 3513 17147 3571 17153
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17116 2927 17119
rect 3528 17116 3556 17147
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 6914 17144 6920 17196
rect 6972 17184 6978 17196
rect 7285 17187 7343 17193
rect 7285 17184 7297 17187
rect 6972 17156 7297 17184
rect 6972 17144 6978 17156
rect 7285 17153 7297 17156
rect 7331 17153 7343 17187
rect 7285 17147 7343 17153
rect 7469 17187 7527 17193
rect 7469 17153 7481 17187
rect 7515 17184 7527 17187
rect 7650 17184 7656 17196
rect 7515 17156 7656 17184
rect 7515 17153 7527 17156
rect 7469 17147 7527 17153
rect 4062 17116 4068 17128
rect 2915 17088 4068 17116
rect 2915 17085 2927 17088
rect 2869 17079 2927 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 5350 17116 5356 17128
rect 4847 17088 5356 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 5442 17076 5448 17128
rect 5500 17116 5506 17128
rect 5552 17116 5580 17144
rect 5905 17119 5963 17125
rect 5905 17116 5917 17119
rect 5500 17088 5917 17116
rect 5500 17076 5506 17088
rect 5905 17085 5917 17088
rect 5951 17085 5963 17119
rect 5905 17079 5963 17085
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 7484 17116 7512 17147
rect 7650 17144 7656 17156
rect 7708 17144 7714 17196
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 9122 17184 9128 17196
rect 8628 17156 9128 17184
rect 8628 17144 8634 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 9674 17144 9680 17196
rect 9732 17184 9738 17196
rect 10686 17184 10692 17196
rect 9732 17156 10692 17184
rect 9732 17144 9738 17156
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 6687 17088 7512 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10100 17088 10609 17116
rect 10100 17076 10106 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 2501 17051 2559 17057
rect 2501 17017 2513 17051
rect 2547 17048 2559 17051
rect 3329 17051 3387 17057
rect 3329 17048 3341 17051
rect 2547 17020 3341 17048
rect 2547 17017 2559 17020
rect 2501 17011 2559 17017
rect 3329 17017 3341 17020
rect 3375 17048 3387 17051
rect 3510 17048 3516 17060
rect 3375 17020 3516 17048
rect 3375 17017 3387 17020
rect 3329 17011 3387 17017
rect 3510 17008 3516 17020
rect 3568 17008 3574 17060
rect 5074 17008 5080 17060
rect 5132 17048 5138 17060
rect 5261 17051 5319 17057
rect 5261 17048 5273 17051
rect 5132 17020 5273 17048
rect 5132 17008 5138 17020
rect 5261 17017 5273 17020
rect 5307 17048 5319 17051
rect 9950 17048 9956 17060
rect 5307 17020 9956 17048
rect 5307 17017 5319 17020
rect 5261 17011 5319 17017
rect 9950 17008 9956 17020
rect 10008 17008 10014 17060
rect 10318 17008 10324 17060
rect 10376 17048 10382 17060
rect 10505 17051 10563 17057
rect 10505 17048 10517 17051
rect 10376 17020 10517 17048
rect 10376 17008 10382 17020
rect 10505 17017 10517 17020
rect 10551 17048 10563 17051
rect 11149 17051 11207 17057
rect 11149 17048 11161 17051
rect 10551 17020 11161 17048
rect 10551 17017 10563 17020
rect 10505 17011 10563 17017
rect 11149 17017 11161 17020
rect 11195 17017 11207 17051
rect 11149 17011 11207 17017
rect 4890 16980 4896 16992
rect 4851 16952 4896 16980
rect 4890 16940 4896 16952
rect 4948 16940 4954 16992
rect 6638 16940 6644 16992
rect 6696 16980 6702 16992
rect 6825 16983 6883 16989
rect 6825 16980 6837 16983
rect 6696 16952 6837 16980
rect 6696 16940 6702 16952
rect 6825 16949 6837 16952
rect 6871 16949 6883 16983
rect 6825 16943 6883 16949
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7374 16980 7380 16992
rect 7239 16952 7380 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7374 16940 7380 16952
rect 7432 16940 7438 16992
rect 8481 16983 8539 16989
rect 8481 16949 8493 16983
rect 8527 16980 8539 16983
rect 8938 16980 8944 16992
rect 8527 16952 8944 16980
rect 8527 16949 8539 16952
rect 8481 16943 8539 16949
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9030 16940 9036 16992
rect 9088 16980 9094 16992
rect 9674 16980 9680 16992
rect 9088 16952 9133 16980
rect 9635 16952 9680 16980
rect 9088 16940 9094 16952
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 12069 16983 12127 16989
rect 12069 16949 12081 16983
rect 12115 16980 12127 16983
rect 12158 16980 12164 16992
rect 12115 16952 12164 16980
rect 12115 16949 12127 16952
rect 12069 16943 12127 16949
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 1104 16890 14812 16912
rect 1104 16838 6315 16890
rect 6367 16838 6379 16890
rect 6431 16838 6443 16890
rect 6495 16838 6507 16890
rect 6559 16838 11648 16890
rect 11700 16838 11712 16890
rect 11764 16838 11776 16890
rect 11828 16838 11840 16890
rect 11892 16838 14812 16890
rect 1104 16816 14812 16838
rect 2406 16776 2412 16788
rect 2367 16748 2412 16776
rect 2406 16736 2412 16748
rect 2464 16736 2470 16788
rect 2590 16736 2596 16788
rect 2648 16776 2654 16788
rect 2774 16776 2780 16788
rect 2648 16748 2780 16776
rect 2648 16736 2654 16748
rect 2774 16736 2780 16748
rect 2832 16776 2838 16788
rect 2832 16748 2877 16776
rect 2832 16736 2838 16748
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 4065 16779 4123 16785
rect 4065 16776 4077 16779
rect 3476 16748 4077 16776
rect 3476 16736 3482 16748
rect 4065 16745 4077 16748
rect 4111 16745 4123 16779
rect 4522 16776 4528 16788
rect 4483 16748 4528 16776
rect 4065 16739 4123 16745
rect 4522 16736 4528 16748
rect 4580 16736 4586 16788
rect 5074 16776 5080 16788
rect 5035 16748 5080 16776
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 7650 16776 7656 16788
rect 7611 16748 7656 16776
rect 7650 16736 7656 16748
rect 7708 16736 7714 16788
rect 8018 16736 8024 16788
rect 8076 16776 8082 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 8076 16748 8217 16776
rect 8076 16736 8082 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 9493 16779 9551 16785
rect 9493 16745 9505 16779
rect 9539 16776 9551 16779
rect 10134 16776 10140 16788
rect 9539 16748 10140 16776
rect 9539 16745 9551 16748
rect 9493 16739 9551 16745
rect 10134 16736 10140 16748
rect 10192 16736 10198 16788
rect 10686 16736 10692 16788
rect 10744 16776 10750 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 10744 16748 11621 16776
rect 10744 16736 10750 16748
rect 11609 16745 11621 16748
rect 11655 16745 11667 16779
rect 11609 16739 11667 16745
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 4890 16708 4896 16720
rect 2915 16680 4896 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2884 16572 2912 16671
rect 4890 16668 4896 16680
rect 4948 16668 4954 16720
rect 7282 16668 7288 16720
rect 7340 16708 7346 16720
rect 7926 16708 7932 16720
rect 7340 16680 7932 16708
rect 7340 16668 7346 16680
rect 7926 16668 7932 16680
rect 7984 16668 7990 16720
rect 8938 16668 8944 16720
rect 8996 16708 9002 16720
rect 9582 16708 9588 16720
rect 8996 16680 9588 16708
rect 8996 16668 9002 16680
rect 9582 16668 9588 16680
rect 9640 16668 9646 16720
rect 9674 16668 9680 16720
rect 9732 16708 9738 16720
rect 11422 16708 11428 16720
rect 9732 16680 11428 16708
rect 9732 16668 9738 16680
rect 4430 16640 4436 16652
rect 4391 16612 4436 16640
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6529 16643 6587 16649
rect 6529 16640 6541 16643
rect 6236 16612 6541 16640
rect 6236 16600 6242 16612
rect 6529 16609 6541 16612
rect 6575 16609 6587 16643
rect 8202 16640 8208 16652
rect 8115 16612 8208 16640
rect 6529 16603 6587 16609
rect 8202 16600 8208 16612
rect 8260 16640 8266 16652
rect 8573 16643 8631 16649
rect 8573 16640 8585 16643
rect 8260 16612 8585 16640
rect 8260 16600 8266 16612
rect 8573 16609 8585 16612
rect 8619 16640 8631 16643
rect 9030 16640 9036 16652
rect 8619 16612 9036 16640
rect 8619 16609 8631 16612
rect 8573 16603 8631 16609
rect 9030 16600 9036 16612
rect 9088 16600 9094 16652
rect 9122 16600 9128 16652
rect 9180 16640 9186 16652
rect 10244 16649 10272 16680
rect 11422 16668 11428 16680
rect 11480 16668 11486 16720
rect 10502 16649 10508 16652
rect 9861 16643 9919 16649
rect 9861 16640 9873 16643
rect 9180 16612 9873 16640
rect 9180 16600 9186 16612
rect 9861 16609 9873 16612
rect 9907 16609 9919 16643
rect 9861 16603 9919 16609
rect 10229 16643 10287 16649
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10496 16640 10508 16649
rect 10463 16612 10508 16640
rect 10229 16603 10287 16609
rect 10496 16603 10508 16612
rect 2096 16544 2912 16572
rect 2096 16532 2102 16544
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3053 16575 3111 16581
rect 3053 16572 3065 16575
rect 3016 16544 3065 16572
rect 3016 16532 3022 16544
rect 3053 16541 3065 16544
rect 3099 16572 3111 16575
rect 3510 16572 3516 16584
rect 3099 16544 3516 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3510 16532 3516 16544
rect 3568 16532 3574 16584
rect 4614 16572 4620 16584
rect 4575 16544 4620 16572
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 6270 16572 6276 16584
rect 6231 16544 6276 16572
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 8018 16532 8024 16584
rect 8076 16572 8082 16584
rect 8220 16572 8248 16600
rect 8076 16544 8248 16572
rect 8076 16532 8082 16544
rect 9876 16436 9904 16603
rect 10502 16600 10508 16603
rect 10560 16600 10566 16652
rect 10042 16436 10048 16448
rect 9876 16408 10048 16436
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 1104 16346 14812 16368
rect 1104 16294 3648 16346
rect 3700 16294 3712 16346
rect 3764 16294 3776 16346
rect 3828 16294 3840 16346
rect 3892 16294 8982 16346
rect 9034 16294 9046 16346
rect 9098 16294 9110 16346
rect 9162 16294 9174 16346
rect 9226 16294 14315 16346
rect 14367 16294 14379 16346
rect 14431 16294 14443 16346
rect 14495 16294 14507 16346
rect 14559 16294 14812 16346
rect 1104 16272 14812 16294
rect 1578 16232 1584 16244
rect 1539 16204 1584 16232
rect 1578 16192 1584 16204
rect 1636 16192 1642 16244
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 4154 16192 4160 16244
rect 4212 16232 4218 16244
rect 4249 16235 4307 16241
rect 4249 16232 4261 16235
rect 4212 16204 4261 16232
rect 4212 16192 4218 16204
rect 4249 16201 4261 16204
rect 4295 16201 4307 16235
rect 6822 16232 6828 16244
rect 6783 16204 6828 16232
rect 4249 16195 4307 16201
rect 6822 16192 6828 16204
rect 6880 16192 6886 16244
rect 9217 16235 9275 16241
rect 9217 16201 9229 16235
rect 9263 16232 9275 16235
rect 9674 16232 9680 16244
rect 9263 16204 9680 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 6641 16099 6699 16105
rect 6641 16065 6653 16099
rect 6687 16096 6699 16099
rect 7282 16096 7288 16108
rect 6687 16068 7288 16096
rect 6687 16065 6699 16068
rect 6641 16059 6699 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16096 7527 16099
rect 7558 16096 7564 16108
rect 7515 16068 7564 16096
rect 7515 16065 7527 16068
rect 7469 16059 7527 16065
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8478 16056 8484 16108
rect 8536 16096 8542 16108
rect 9324 16105 9352 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10042 16192 10048 16244
rect 10100 16232 10106 16244
rect 10689 16235 10747 16241
rect 10689 16232 10701 16235
rect 10100 16204 10701 16232
rect 10100 16192 10106 16204
rect 10689 16201 10701 16204
rect 10735 16201 10747 16235
rect 10689 16195 10747 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11422 16232 11428 16244
rect 11379 16204 11428 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 8536 16068 9321 16096
rect 8536 16056 8542 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 1394 16028 1400 16040
rect 1355 16000 1400 16028
rect 1394 15988 1400 16000
rect 1452 15988 1458 16040
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 2823 16000 2881 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 2869 15997 2881 16000
rect 2915 16028 2927 16031
rect 5905 16031 5963 16037
rect 2915 16000 5396 16028
rect 2915 15997 2927 16000
rect 2869 15991 2927 15997
rect 5368 15972 5396 16000
rect 5905 15997 5917 16031
rect 5951 16028 5963 16031
rect 6178 16028 6184 16040
rect 5951 16000 6184 16028
rect 5951 15997 5963 16000
rect 5905 15991 5963 15997
rect 6178 15988 6184 16000
rect 6236 15988 6242 16040
rect 6270 15988 6276 16040
rect 6328 16028 6334 16040
rect 6822 16028 6828 16040
rect 6328 16000 6828 16028
rect 6328 15988 6334 16000
rect 6822 15988 6828 16000
rect 6880 15988 6886 16040
rect 6914 15988 6920 16040
rect 6972 16028 6978 16040
rect 7193 16031 7251 16037
rect 7193 16028 7205 16031
rect 6972 16000 7205 16028
rect 6972 15988 6978 16000
rect 7193 15997 7205 16000
rect 7239 16028 7251 16031
rect 7742 16028 7748 16040
rect 7239 16000 7748 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 7742 15988 7748 16000
rect 7800 15988 7806 16040
rect 2409 15963 2467 15969
rect 2409 15929 2421 15963
rect 2455 15960 2467 15963
rect 2455 15932 2912 15960
rect 2455 15929 2467 15932
rect 2409 15923 2467 15929
rect 2884 15892 2912 15932
rect 2958 15920 2964 15972
rect 3016 15960 3022 15972
rect 3114 15963 3172 15969
rect 3114 15960 3126 15963
rect 3016 15932 3126 15960
rect 3016 15920 3022 15932
rect 3114 15929 3126 15932
rect 3160 15960 3172 15963
rect 4614 15960 4620 15972
rect 3160 15932 4620 15960
rect 3160 15929 3172 15932
rect 3114 15923 3172 15929
rect 4614 15920 4620 15932
rect 4672 15960 4678 15972
rect 4801 15963 4859 15969
rect 4801 15960 4813 15963
rect 4672 15932 4813 15960
rect 4672 15920 4678 15932
rect 4801 15929 4813 15932
rect 4847 15929 4859 15963
rect 4801 15923 4859 15929
rect 5350 15920 5356 15972
rect 5408 15960 5414 15972
rect 6288 15960 6316 15988
rect 5408 15932 6316 15960
rect 5408 15920 5414 15932
rect 9490 15920 9496 15972
rect 9548 15969 9554 15972
rect 9548 15963 9612 15969
rect 9548 15929 9566 15963
rect 9600 15929 9612 15963
rect 9548 15923 9612 15929
rect 9548 15920 9554 15923
rect 3510 15892 3516 15904
rect 2884 15864 3516 15892
rect 3510 15852 3516 15864
rect 3568 15852 3574 15904
rect 7929 15895 7987 15901
rect 7929 15861 7941 15895
rect 7975 15892 7987 15895
rect 8110 15892 8116 15904
rect 7975 15864 8116 15892
rect 7975 15861 7987 15864
rect 7929 15855 7987 15861
rect 8110 15852 8116 15864
rect 8168 15892 8174 15904
rect 8386 15892 8392 15904
rect 8168 15864 8392 15892
rect 8168 15852 8174 15864
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 1104 15802 14812 15824
rect 1104 15750 6315 15802
rect 6367 15750 6379 15802
rect 6431 15750 6443 15802
rect 6495 15750 6507 15802
rect 6559 15750 11648 15802
rect 11700 15750 11712 15802
rect 11764 15750 11776 15802
rect 11828 15750 11840 15802
rect 11892 15750 14812 15802
rect 1104 15728 14812 15750
rect 1394 15648 1400 15700
rect 1452 15688 1458 15700
rect 1581 15691 1639 15697
rect 1581 15688 1593 15691
rect 1452 15660 1593 15688
rect 1452 15648 1458 15660
rect 1581 15657 1593 15660
rect 1627 15657 1639 15691
rect 1581 15651 1639 15657
rect 2501 15691 2559 15697
rect 2501 15657 2513 15691
rect 2547 15688 2559 15691
rect 2590 15688 2596 15700
rect 2547 15660 2596 15688
rect 2547 15657 2559 15660
rect 2501 15651 2559 15657
rect 2590 15648 2596 15660
rect 2648 15648 2654 15700
rect 2958 15688 2964 15700
rect 2919 15660 2964 15688
rect 2958 15648 2964 15660
rect 3016 15648 3022 15700
rect 4062 15648 4068 15700
rect 4120 15688 4126 15700
rect 4430 15688 4436 15700
rect 4120 15660 4436 15688
rect 4120 15648 4126 15660
rect 4430 15648 4436 15660
rect 4488 15688 4494 15700
rect 4617 15691 4675 15697
rect 4617 15688 4629 15691
rect 4488 15660 4629 15688
rect 4488 15648 4494 15660
rect 4617 15657 4629 15660
rect 4663 15657 4675 15691
rect 6914 15688 6920 15700
rect 6875 15660 6920 15688
rect 4617 15651 4675 15657
rect 6914 15648 6920 15660
rect 6972 15648 6978 15700
rect 7374 15688 7380 15700
rect 7335 15660 7380 15688
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 9401 15691 9459 15697
rect 9401 15657 9413 15691
rect 9447 15688 9459 15691
rect 9490 15688 9496 15700
rect 9447 15660 9496 15688
rect 9447 15657 9459 15660
rect 9401 15651 9459 15657
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9858 15688 9864 15700
rect 9819 15660 9864 15688
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 10502 15648 10508 15700
rect 10560 15688 10566 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 10560 15660 10885 15688
rect 10560 15648 10566 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 10873 15651 10931 15657
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 13170 15688 13176 15700
rect 12575 15660 13176 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 4341 15623 4399 15629
rect 4341 15589 4353 15623
rect 4387 15620 4399 15623
rect 4522 15620 4528 15632
rect 4387 15592 4528 15620
rect 4387 15589 4399 15592
rect 4341 15583 4399 15589
rect 4522 15580 4528 15592
rect 4580 15580 4586 15632
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 11885 15623 11943 15629
rect 11112 15592 11836 15620
rect 11112 15580 11118 15592
rect 4154 15512 4160 15564
rect 4212 15552 4218 15564
rect 5149 15555 5207 15561
rect 5149 15552 5161 15555
rect 4212 15524 5161 15552
rect 4212 15512 4218 15524
rect 5149 15521 5161 15524
rect 5195 15552 5207 15555
rect 5534 15552 5540 15564
rect 5195 15524 5540 15552
rect 5195 15521 5207 15524
rect 5149 15515 5207 15521
rect 5534 15512 5540 15524
rect 5592 15512 5598 15564
rect 7098 15512 7104 15564
rect 7156 15552 7162 15564
rect 7745 15555 7803 15561
rect 7745 15552 7757 15555
rect 7156 15524 7757 15552
rect 7156 15512 7162 15524
rect 7745 15521 7757 15524
rect 7791 15552 7803 15555
rect 8018 15552 8024 15564
rect 7791 15524 8024 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 8018 15512 8024 15524
rect 8076 15512 8082 15564
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 11808 15561 11836 15592
rect 11885 15589 11897 15623
rect 11931 15620 11943 15623
rect 11974 15620 11980 15632
rect 11931 15592 11980 15620
rect 11931 15589 11943 15592
rect 11885 15583 11943 15589
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 9732 15524 10241 15552
rect 9732 15512 9738 15524
rect 10229 15521 10241 15524
rect 10275 15552 10287 15555
rect 11793 15555 11851 15561
rect 10275 15524 11468 15552
rect 10275 15521 10287 15524
rect 10229 15515 10287 15521
rect 4890 15484 4896 15496
rect 4851 15456 4896 15484
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 7834 15484 7840 15496
rect 7795 15456 7840 15484
rect 7834 15444 7840 15456
rect 7892 15444 7898 15496
rect 7929 15487 7987 15493
rect 7929 15453 7941 15487
rect 7975 15453 7987 15487
rect 10318 15484 10324 15496
rect 10279 15456 10324 15484
rect 7929 15447 7987 15453
rect 7193 15419 7251 15425
rect 7193 15416 7205 15419
rect 6288 15388 7205 15416
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 6288 15357 6316 15388
rect 7193 15385 7205 15388
rect 7239 15416 7251 15419
rect 7558 15416 7564 15428
rect 7239 15388 7564 15416
rect 7239 15385 7251 15388
rect 7193 15379 7251 15385
rect 7558 15376 7564 15388
rect 7616 15416 7622 15428
rect 7944 15416 7972 15447
rect 10318 15444 10324 15456
rect 10376 15444 10382 15496
rect 10502 15484 10508 15496
rect 10463 15456 10508 15484
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 11440 15425 11468 15524
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12342 15552 12348 15564
rect 11839 15524 12348 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 11977 15487 12035 15493
rect 11977 15484 11989 15487
rect 11756 15456 11989 15484
rect 11756 15444 11762 15456
rect 11977 15453 11989 15456
rect 12023 15484 12035 15487
rect 12158 15484 12164 15496
rect 12023 15456 12164 15484
rect 12023 15453 12035 15456
rect 11977 15447 12035 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 7616 15388 7972 15416
rect 11425 15419 11483 15425
rect 7616 15376 7622 15388
rect 11425 15385 11437 15419
rect 11471 15385 11483 15419
rect 11425 15379 11483 15385
rect 6273 15351 6331 15357
rect 6273 15348 6285 15351
rect 6236 15320 6285 15348
rect 6236 15308 6242 15320
rect 6273 15317 6285 15320
rect 6319 15317 6331 15351
rect 6273 15311 6331 15317
rect 1104 15258 14812 15280
rect 1104 15206 3648 15258
rect 3700 15206 3712 15258
rect 3764 15206 3776 15258
rect 3828 15206 3840 15258
rect 3892 15206 8982 15258
rect 9034 15206 9046 15258
rect 9098 15206 9110 15258
rect 9162 15206 9174 15258
rect 9226 15206 14315 15258
rect 14367 15206 14379 15258
rect 14431 15206 14443 15258
rect 14495 15206 14507 15258
rect 14559 15206 14812 15258
rect 1104 15184 14812 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 2682 15144 2688 15156
rect 1995 15116 2688 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 1397 14943 1455 14949
rect 1397 14909 1409 14943
rect 1443 14940 1455 14943
rect 1964 14940 1992 15107
rect 2682 15104 2688 15116
rect 2740 15104 2746 15156
rect 4062 15144 4068 15156
rect 4023 15116 4068 15144
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4614 15104 4620 15156
rect 4672 15144 4678 15156
rect 4890 15144 4896 15156
rect 4672 15116 4896 15144
rect 4672 15104 4678 15116
rect 4890 15104 4896 15116
rect 4948 15144 4954 15156
rect 5169 15147 5227 15153
rect 5169 15144 5181 15147
rect 4948 15116 5181 15144
rect 4948 15104 4954 15116
rect 5169 15113 5181 15116
rect 5215 15144 5227 15147
rect 5350 15144 5356 15156
rect 5215 15116 5356 15144
rect 5215 15113 5227 15116
rect 5169 15107 5227 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5534 15144 5540 15156
rect 5495 15116 5540 15144
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 10318 15144 10324 15156
rect 10279 15116 10324 15144
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 10962 15144 10968 15156
rect 10919 15116 10968 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 10962 15104 10968 15116
rect 11020 15104 11026 15156
rect 9953 15079 10011 15085
rect 9953 15045 9965 15079
rect 9999 15076 10011 15079
rect 10502 15076 10508 15088
rect 9999 15048 10508 15076
rect 9999 15045 10011 15048
rect 9953 15039 10011 15045
rect 10502 15036 10508 15048
rect 10560 15036 10566 15088
rect 3510 14968 3516 15020
rect 3568 15008 3574 15020
rect 3605 15011 3663 15017
rect 3605 15008 3617 15011
rect 3568 14980 3617 15008
rect 3568 14968 3574 14980
rect 3605 14977 3617 14980
rect 3651 15008 3663 15011
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 3651 14980 4629 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 4617 14971 4675 14977
rect 12158 14968 12164 15020
rect 12216 15008 12222 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12216 14980 13001 15008
rect 12216 14968 12222 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 1443 14912 1992 14940
rect 3973 14943 4031 14949
rect 1443 14909 1455 14912
rect 1397 14903 1455 14909
rect 3973 14909 3985 14943
rect 4019 14940 4031 14943
rect 4430 14940 4436 14952
rect 4019 14912 4436 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 6822 14900 6828 14952
rect 6880 14940 6886 14952
rect 7837 14943 7895 14949
rect 7837 14940 7849 14943
rect 6880 14912 7849 14940
rect 6880 14900 6886 14912
rect 7837 14909 7849 14912
rect 7883 14940 7895 14943
rect 8478 14940 8484 14952
rect 7883 14912 8484 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4580 14776 4625 14804
rect 4580 14764 4586 14776
rect 6178 14764 6184 14816
rect 6236 14804 6242 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 6236 14776 6561 14804
rect 6236 14764 6242 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 7098 14804 7104 14816
rect 7059 14776 7104 14804
rect 6549 14767 6607 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7742 14804 7748 14816
rect 7515 14776 7748 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 7944 14804 7972 14912
rect 8478 14900 8484 14912
rect 8536 14900 8542 14952
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 10778 14940 10784 14952
rect 10284 14912 10784 14940
rect 10284 14900 10290 14912
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 12894 14940 12900 14952
rect 12807 14912 12900 14940
rect 12894 14900 12900 14912
rect 12952 14940 12958 14952
rect 13170 14940 13176 14952
rect 12952 14912 13176 14940
rect 12952 14900 12958 14912
rect 13170 14900 13176 14912
rect 13228 14900 13234 14952
rect 8110 14881 8116 14884
rect 8104 14872 8116 14881
rect 8071 14844 8116 14872
rect 8104 14835 8116 14844
rect 8168 14872 8174 14884
rect 8570 14872 8576 14884
rect 8168 14844 8576 14872
rect 8110 14832 8116 14835
rect 8168 14832 8174 14844
rect 8570 14832 8576 14844
rect 8628 14832 8634 14884
rect 11698 14872 11704 14884
rect 11164 14844 11704 14872
rect 8018 14804 8024 14816
rect 7944 14776 8024 14804
rect 8018 14764 8024 14776
rect 8076 14764 8082 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9306 14804 9312 14816
rect 9263 14776 9312 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 11164 14813 11192 14844
rect 11698 14832 11704 14844
rect 11756 14832 11762 14884
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 12710 14872 12716 14884
rect 12299 14844 12716 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12710 14832 12716 14844
rect 12768 14872 12774 14884
rect 12805 14875 12863 14881
rect 12805 14872 12817 14875
rect 12768 14844 12817 14872
rect 12768 14832 12774 14844
rect 12805 14841 12817 14844
rect 12851 14872 12863 14875
rect 13998 14872 14004 14884
rect 12851 14844 14004 14872
rect 12851 14841 12863 14844
rect 12805 14835 12863 14841
rect 13998 14832 14004 14844
rect 14056 14832 14062 14884
rect 11149 14807 11207 14813
rect 11149 14804 11161 14807
rect 10836 14776 11161 14804
rect 10836 14764 10842 14776
rect 11149 14773 11161 14776
rect 11195 14773 11207 14807
rect 11330 14804 11336 14816
rect 11291 14776 11336 14804
rect 11149 14767 11207 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 11885 14807 11943 14813
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 12158 14804 12164 14816
rect 11931 14776 12164 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12492 14776 12537 14804
rect 12492 14764 12498 14776
rect 1104 14714 14812 14736
rect 1104 14662 6315 14714
rect 6367 14662 6379 14714
rect 6431 14662 6443 14714
rect 6495 14662 6507 14714
rect 6559 14662 11648 14714
rect 11700 14662 11712 14714
rect 11764 14662 11776 14714
rect 11828 14662 11840 14714
rect 11892 14662 14812 14714
rect 1104 14640 14812 14662
rect 4341 14603 4399 14609
rect 4341 14569 4353 14603
rect 4387 14600 4399 14603
rect 4522 14600 4528 14612
rect 4387 14572 4528 14600
rect 4387 14569 4399 14572
rect 4341 14563 4399 14569
rect 4522 14560 4528 14572
rect 4580 14600 4586 14612
rect 4709 14603 4767 14609
rect 4709 14600 4721 14603
rect 4580 14572 4721 14600
rect 4580 14560 4586 14572
rect 4709 14569 4721 14572
rect 4755 14569 4767 14603
rect 4709 14563 4767 14569
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 5132 14572 5181 14600
rect 5132 14560 5138 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 8018 14600 8024 14612
rect 7979 14572 8024 14600
rect 5169 14563 5227 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 9493 14603 9551 14609
rect 9493 14569 9505 14603
rect 9539 14600 9551 14603
rect 9582 14600 9588 14612
rect 9539 14572 9588 14600
rect 9539 14569 9551 14572
rect 9493 14563 9551 14569
rect 9582 14560 9588 14572
rect 9640 14560 9646 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 10318 14600 10324 14612
rect 10275 14572 10324 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 10318 14560 10324 14572
rect 10376 14560 10382 14612
rect 11517 14603 11575 14609
rect 11517 14569 11529 14603
rect 11563 14600 11575 14603
rect 11974 14600 11980 14612
rect 11563 14572 11980 14600
rect 11563 14569 11575 14572
rect 11517 14563 11575 14569
rect 11974 14560 11980 14572
rect 12032 14600 12038 14612
rect 12434 14600 12440 14612
rect 12032 14572 12440 14600
rect 12032 14560 12038 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 5350 14532 5356 14544
rect 5092 14504 5356 14532
rect 4890 14424 4896 14476
rect 4948 14464 4954 14476
rect 5092 14473 5120 14504
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 7282 14492 7288 14544
rect 7340 14532 7346 14544
rect 7469 14535 7527 14541
rect 7469 14532 7481 14535
rect 7340 14504 7481 14532
rect 7340 14492 7346 14504
rect 7469 14501 7481 14504
rect 7515 14532 7527 14535
rect 7834 14532 7840 14544
rect 7515 14504 7840 14532
rect 7515 14501 7527 14504
rect 7469 14495 7527 14501
rect 7834 14492 7840 14504
rect 7892 14492 7898 14544
rect 12158 14532 12164 14544
rect 12084 14504 12164 14532
rect 5077 14467 5135 14473
rect 5077 14464 5089 14467
rect 4948 14436 5089 14464
rect 4948 14424 4954 14436
rect 5077 14433 5089 14436
rect 5123 14433 5135 14467
rect 5077 14427 5135 14433
rect 6914 14424 6920 14476
rect 6972 14464 6978 14476
rect 7374 14464 7380 14476
rect 6972 14436 7380 14464
rect 6972 14424 6978 14436
rect 7374 14424 7380 14436
rect 7432 14424 7438 14476
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 9582 14464 9588 14476
rect 8812 14436 9588 14464
rect 8812 14424 8818 14436
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 10594 14464 10600 14476
rect 10555 14436 10600 14464
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11790 14464 11796 14476
rect 11480 14436 11796 14464
rect 11480 14424 11486 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 11882 14424 11888 14476
rect 11940 14464 11946 14476
rect 12084 14473 12112 14504
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 12049 14467 12112 14473
rect 12049 14464 12061 14467
rect 11940 14436 12061 14464
rect 11940 14424 11946 14436
rect 12049 14433 12061 14436
rect 12095 14436 12112 14467
rect 12095 14433 12107 14436
rect 12049 14427 12107 14433
rect 5353 14399 5411 14405
rect 5353 14365 5365 14399
rect 5399 14396 5411 14399
rect 5442 14396 5448 14408
rect 5399 14368 5448 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 7558 14396 7564 14408
rect 7519 14368 7564 14396
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10410 14396 10416 14408
rect 10183 14368 10416 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10410 14356 10416 14368
rect 10468 14396 10474 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10468 14368 10701 14396
rect 10468 14356 10474 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 10689 14359 10747 14365
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 10836 14368 10881 14396
rect 10836 14356 10842 14368
rect 6549 14331 6607 14337
rect 6549 14297 6561 14331
rect 6595 14328 6607 14331
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6595 14300 7021 14328
rect 6595 14297 6607 14300
rect 6549 14291 6607 14297
rect 7009 14297 7021 14300
rect 7055 14328 7067 14331
rect 7282 14328 7288 14340
rect 7055 14300 7288 14328
rect 7055 14297 7067 14300
rect 7009 14291 7067 14297
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 6917 14263 6975 14269
rect 6917 14229 6929 14263
rect 6963 14260 6975 14263
rect 7558 14260 7564 14272
rect 6963 14232 7564 14260
rect 6963 14229 6975 14232
rect 6917 14223 6975 14229
rect 7558 14220 7564 14232
rect 7616 14220 7622 14272
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8389 14263 8447 14269
rect 8389 14260 8401 14263
rect 8168 14232 8401 14260
rect 8168 14220 8174 14232
rect 8389 14229 8401 14232
rect 8435 14229 8447 14263
rect 8846 14260 8852 14272
rect 8807 14232 8852 14260
rect 8389 14223 8447 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 10778 14220 10784 14272
rect 10836 14260 10842 14272
rect 13173 14263 13231 14269
rect 13173 14260 13185 14263
rect 10836 14232 13185 14260
rect 10836 14220 10842 14232
rect 13173 14229 13185 14232
rect 13219 14229 13231 14263
rect 13173 14223 13231 14229
rect 1104 14170 14812 14192
rect 1104 14118 3648 14170
rect 3700 14118 3712 14170
rect 3764 14118 3776 14170
rect 3828 14118 3840 14170
rect 3892 14118 8982 14170
rect 9034 14118 9046 14170
rect 9098 14118 9110 14170
rect 9162 14118 9174 14170
rect 9226 14118 14315 14170
rect 14367 14118 14379 14170
rect 14431 14118 14443 14170
rect 14495 14118 14507 14170
rect 14559 14118 14812 14170
rect 1104 14096 14812 14118
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 5074 14056 5080 14068
rect 4847 14028 5080 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 5074 14016 5080 14028
rect 5132 14056 5138 14068
rect 5350 14056 5356 14068
rect 5132 14028 5356 14056
rect 5132 14016 5138 14028
rect 5350 14016 5356 14028
rect 5408 14016 5414 14068
rect 6178 14056 6184 14068
rect 6139 14028 6184 14056
rect 6178 14016 6184 14028
rect 6236 14016 6242 14068
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14056 6699 14059
rect 6730 14056 6736 14068
rect 6687 14028 6736 14056
rect 6687 14025 6699 14028
rect 6641 14019 6699 14025
rect 6730 14016 6736 14028
rect 6788 14016 6794 14068
rect 7834 14056 7840 14068
rect 7795 14028 7840 14056
rect 7834 14016 7840 14028
rect 7892 14016 7898 14068
rect 8386 14056 8392 14068
rect 8347 14028 8392 14056
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 10226 14056 10232 14068
rect 10187 14028 10232 14056
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10410 14056 10416 14068
rect 10371 14028 10416 14056
rect 10410 14016 10416 14028
rect 10468 14016 10474 14068
rect 11790 14056 11796 14068
rect 11751 14028 11796 14056
rect 11790 14016 11796 14028
rect 11848 14016 11854 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 12032 14028 12173 14056
rect 12032 14016 12038 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 8297 13991 8355 13997
rect 8297 13957 8309 13991
rect 8343 13988 8355 13991
rect 9306 13988 9312 14000
rect 8343 13960 9312 13988
rect 8343 13957 8355 13960
rect 8297 13951 8355 13957
rect 4890 13880 4896 13932
rect 4948 13920 4954 13932
rect 5077 13923 5135 13929
rect 5077 13920 5089 13923
rect 4948 13892 5089 13920
rect 4948 13880 4954 13892
rect 5077 13889 5089 13892
rect 5123 13889 5135 13923
rect 7282 13920 7288 13932
rect 7243 13892 7288 13920
rect 5077 13883 5135 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 8846 13920 8852 13932
rect 8807 13892 8852 13920
rect 8846 13880 8852 13892
rect 8904 13880 8910 13932
rect 8956 13929 8984 13960
rect 9306 13948 9312 13960
rect 9364 13948 9370 14000
rect 9585 13991 9643 13997
rect 9585 13957 9597 13991
rect 9631 13988 9643 13991
rect 10778 13988 10784 14000
rect 9631 13960 10784 13988
rect 9631 13957 9643 13960
rect 9585 13951 9643 13957
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 12176 13988 12204 14019
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 12437 14059 12495 14065
rect 12437 14056 12449 14059
rect 12400 14028 12449 14056
rect 12400 14016 12406 14028
rect 12437 14025 12449 14028
rect 12483 14025 12495 14059
rect 12437 14019 12495 14025
rect 12526 13988 12532 14000
rect 12176 13960 12532 13988
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 9953 13923 10011 13929
rect 9953 13889 9965 13923
rect 9999 13920 10011 13923
rect 10965 13923 11023 13929
rect 10965 13920 10977 13923
rect 9999 13892 10977 13920
rect 9999 13889 10011 13892
rect 9953 13883 10011 13889
rect 10965 13889 10977 13892
rect 11011 13920 11023 13923
rect 11425 13923 11483 13929
rect 11425 13920 11437 13923
rect 11011 13892 11437 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 11425 13889 11437 13892
rect 11471 13920 11483 13923
rect 11882 13920 11888 13932
rect 11471 13892 11888 13920
rect 11471 13889 11483 13892
rect 11425 13883 11483 13889
rect 11882 13880 11888 13892
rect 11940 13920 11946 13932
rect 12158 13920 12164 13932
rect 11940 13892 12164 13920
rect 11940 13880 11946 13892
rect 12158 13880 12164 13892
rect 12216 13920 12222 13932
rect 13081 13923 13139 13929
rect 13081 13920 13093 13923
rect 12216 13892 13093 13920
rect 12216 13880 12222 13892
rect 13081 13889 13093 13892
rect 13127 13920 13139 13923
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 13127 13892 13461 13920
rect 13127 13889 13139 13892
rect 13081 13883 13139 13889
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 5442 13852 5448 13864
rect 5403 13824 5448 13852
rect 5442 13812 5448 13824
rect 5500 13812 5506 13864
rect 6730 13812 6736 13864
rect 6788 13852 6794 13864
rect 8864 13852 8892 13880
rect 6788 13824 6868 13852
rect 6788 13812 6794 13824
rect 6840 13784 6868 13824
rect 8312 13824 8892 13852
rect 7193 13787 7251 13793
rect 7193 13784 7205 13787
rect 6840 13756 7205 13784
rect 7193 13753 7205 13756
rect 7239 13753 7251 13787
rect 7193 13747 7251 13753
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 7208 13716 7236 13747
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 8312 13784 8340 13824
rect 10226 13812 10232 13864
rect 10284 13852 10290 13864
rect 10781 13855 10839 13861
rect 10781 13852 10793 13855
rect 10284 13824 10793 13852
rect 10284 13812 10290 13824
rect 10781 13821 10793 13824
rect 10827 13821 10839 13855
rect 10781 13815 10839 13821
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12584 13824 12909 13852
rect 12584 13812 12590 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 8076 13756 8340 13784
rect 8076 13744 8082 13756
rect 8202 13716 8208 13728
rect 7208 13688 8208 13716
rect 8202 13676 8208 13688
rect 8260 13676 8266 13728
rect 8754 13716 8760 13728
rect 8715 13688 8760 13716
rect 8754 13676 8760 13688
rect 8812 13676 8818 13728
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 10928 13688 10973 13716
rect 10928 13676 10934 13688
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 12618 13716 12624 13728
rect 11388 13688 12624 13716
rect 11388 13676 11394 13688
rect 12618 13676 12624 13688
rect 12676 13716 12682 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12676 13688 12817 13716
rect 12676 13676 12682 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 12805 13679 12863 13685
rect 1104 13626 14812 13648
rect 1104 13574 6315 13626
rect 6367 13574 6379 13626
rect 6431 13574 6443 13626
rect 6495 13574 6507 13626
rect 6559 13574 11648 13626
rect 11700 13574 11712 13626
rect 11764 13574 11776 13626
rect 11828 13574 11840 13626
rect 11892 13574 14812 13626
rect 1104 13552 14812 13574
rect 1486 13472 1492 13524
rect 1544 13512 1550 13524
rect 1581 13515 1639 13521
rect 1581 13512 1593 13515
rect 1544 13484 1593 13512
rect 1544 13472 1550 13484
rect 1581 13481 1593 13484
rect 1627 13481 1639 13515
rect 1581 13475 1639 13481
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6144 13484 6285 13512
rect 6144 13472 6150 13484
rect 6273 13481 6285 13484
rect 6319 13512 6331 13515
rect 6822 13512 6828 13524
rect 6319 13484 6828 13512
rect 6319 13481 6331 13484
rect 6273 13475 6331 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 8662 13512 8668 13524
rect 8527 13484 8668 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 8662 13472 8668 13484
rect 8720 13472 8726 13524
rect 9953 13515 10011 13521
rect 9953 13481 9965 13515
rect 9999 13512 10011 13515
rect 10594 13512 10600 13524
rect 9999 13484 10600 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10594 13472 10600 13484
rect 10652 13512 10658 13524
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 10652 13484 11621 13512
rect 10652 13472 10658 13484
rect 11609 13481 11621 13484
rect 11655 13481 11667 13515
rect 11609 13475 11667 13481
rect 11977 13515 12035 13521
rect 11977 13481 11989 13515
rect 12023 13512 12035 13515
rect 12066 13512 12072 13524
rect 12023 13484 12072 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 12618 13512 12624 13524
rect 12579 13484 12624 13512
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 5810 13404 5816 13456
rect 5868 13444 5874 13456
rect 6365 13447 6423 13453
rect 6365 13444 6377 13447
rect 5868 13416 6377 13444
rect 5868 13404 5874 13416
rect 6365 13413 6377 13416
rect 6411 13444 6423 13447
rect 6638 13444 6644 13456
rect 6411 13416 6644 13444
rect 6411 13413 6423 13416
rect 6365 13407 6423 13413
rect 6638 13404 6644 13416
rect 6696 13404 6702 13456
rect 7374 13404 7380 13456
rect 7432 13444 7438 13456
rect 7929 13447 7987 13453
rect 7929 13444 7941 13447
rect 7432 13416 7941 13444
rect 7432 13404 7438 13416
rect 7929 13413 7941 13416
rect 7975 13444 7987 13447
rect 8754 13444 8760 13456
rect 7975 13416 8760 13444
rect 7975 13413 7987 13416
rect 7929 13407 7987 13413
rect 8754 13404 8760 13416
rect 8812 13404 8818 13456
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 8389 13379 8447 13385
rect 8389 13345 8401 13379
rect 8435 13376 8447 13379
rect 8846 13376 8852 13388
rect 8435 13348 8852 13376
rect 8435 13345 8447 13348
rect 8389 13339 8447 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 9950 13336 9956 13388
rect 10008 13376 10014 13388
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 10008 13348 10425 13376
rect 10008 13336 10014 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12069 13379 12127 13385
rect 12069 13376 12081 13379
rect 12032 13348 12081 13376
rect 12032 13336 12038 13348
rect 12069 13345 12081 13348
rect 12115 13345 12127 13379
rect 12069 13339 12127 13345
rect 6454 13308 6460 13320
rect 6415 13280 6460 13308
rect 6454 13268 6460 13280
rect 6512 13268 6518 13320
rect 8110 13268 8116 13320
rect 8168 13308 8174 13320
rect 8573 13311 8631 13317
rect 8573 13308 8585 13311
rect 8168 13280 8585 13308
rect 8168 13268 8174 13280
rect 8573 13277 8585 13280
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10505 13311 10563 13317
rect 10505 13308 10517 13311
rect 10376 13280 10517 13308
rect 10376 13268 10382 13280
rect 10505 13277 10517 13280
rect 10551 13277 10563 13311
rect 10686 13308 10692 13320
rect 10647 13280 10692 13308
rect 10505 13271 10563 13277
rect 10686 13268 10692 13280
rect 10744 13268 10750 13320
rect 12158 13308 12164 13320
rect 12119 13280 12164 13308
rect 12158 13268 12164 13280
rect 12216 13268 12222 13320
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 10870 13240 10876 13252
rect 10091 13212 10876 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 10870 13200 10876 13212
rect 10928 13240 10934 13252
rect 11057 13243 11115 13249
rect 11057 13240 11069 13243
rect 10928 13212 11069 13240
rect 10928 13200 10934 13212
rect 11057 13209 11069 13212
rect 11103 13209 11115 13243
rect 11057 13203 11115 13209
rect 2682 13172 2688 13184
rect 2643 13144 2688 13172
rect 2682 13132 2688 13144
rect 2740 13132 2746 13184
rect 5905 13175 5963 13181
rect 5905 13141 5917 13175
rect 5951 13172 5963 13175
rect 6638 13172 6644 13184
rect 5951 13144 6644 13172
rect 5951 13141 5963 13144
rect 5905 13135 5963 13141
rect 6638 13132 6644 13144
rect 6696 13132 6702 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7009 13175 7067 13181
rect 7009 13172 7021 13175
rect 6972 13144 7021 13172
rect 6972 13132 6978 13144
rect 7009 13141 7021 13144
rect 7055 13141 7067 13175
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7009 13135 7067 13141
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 9125 13175 9183 13181
rect 9125 13141 9137 13175
rect 9171 13172 9183 13175
rect 9306 13172 9312 13184
rect 9171 13144 9312 13172
rect 9171 13141 9183 13144
rect 9125 13135 9183 13141
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 1104 13082 14812 13104
rect 1104 13030 3648 13082
rect 3700 13030 3712 13082
rect 3764 13030 3776 13082
rect 3828 13030 3840 13082
rect 3892 13030 8982 13082
rect 9034 13030 9046 13082
rect 9098 13030 9110 13082
rect 9162 13030 9174 13082
rect 9226 13030 14315 13082
rect 14367 13030 14379 13082
rect 14431 13030 14443 13082
rect 14495 13030 14507 13082
rect 14559 13030 14812 13082
rect 1104 13008 14812 13030
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5997 12971 6055 12977
rect 5997 12968 6009 12971
rect 5776 12940 6009 12968
rect 5776 12928 5782 12940
rect 5997 12937 6009 12940
rect 6043 12968 6055 12971
rect 6454 12968 6460 12980
rect 6043 12940 6460 12968
rect 6043 12937 6055 12940
rect 5997 12931 6055 12937
rect 6454 12928 6460 12940
rect 6512 12968 6518 12980
rect 6822 12968 6828 12980
rect 6512 12940 6828 12968
rect 6512 12928 6518 12940
rect 6822 12928 6828 12940
rect 6880 12928 6886 12980
rect 7374 12968 7380 12980
rect 7335 12940 7380 12968
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 8757 12971 8815 12977
rect 8757 12968 8769 12971
rect 8720 12940 8769 12968
rect 8720 12928 8726 12940
rect 8757 12937 8769 12940
rect 8803 12968 8815 12971
rect 8846 12968 8852 12980
rect 8803 12940 8852 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 8846 12928 8852 12940
rect 8904 12928 8910 12980
rect 10321 12971 10379 12977
rect 10321 12937 10333 12971
rect 10367 12968 10379 12971
rect 10686 12968 10692 12980
rect 10367 12940 10692 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10686 12928 10692 12940
rect 10744 12968 10750 12980
rect 11241 12971 11299 12977
rect 11241 12968 11253 12971
rect 10744 12940 11253 12968
rect 10744 12928 10750 12940
rect 11241 12937 11253 12940
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 11701 12971 11759 12977
rect 11701 12937 11713 12971
rect 11747 12968 11759 12971
rect 12066 12968 12072 12980
rect 11747 12940 12072 12968
rect 11747 12937 11759 12940
rect 11701 12931 11759 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12158 12928 12164 12980
rect 12216 12968 12222 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12216 12940 12633 12968
rect 12216 12928 12222 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 12621 12931 12679 12937
rect 5629 12903 5687 12909
rect 5629 12869 5641 12903
rect 5675 12900 5687 12903
rect 5810 12900 5816 12912
rect 5675 12872 5816 12900
rect 5675 12869 5687 12872
rect 5629 12863 5687 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 11422 12900 11428 12912
rect 11204 12872 11428 12900
rect 11204 12860 11210 12872
rect 11422 12860 11428 12872
rect 11480 12900 11486 12912
rect 11974 12900 11980 12912
rect 11480 12872 11980 12900
rect 11480 12860 11486 12872
rect 11974 12860 11980 12872
rect 12032 12860 12038 12912
rect 12084 12900 12112 12928
rect 12526 12900 12532 12912
rect 12084 12872 12532 12900
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 6178 12832 6184 12844
rect 5828 12804 6184 12832
rect 5828 12776 5856 12804
rect 6178 12792 6184 12804
rect 6236 12792 6242 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7929 12835 7987 12841
rect 7929 12832 7941 12835
rect 6687 12804 7941 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7929 12801 7941 12804
rect 7975 12832 7987 12835
rect 8110 12832 8116 12844
rect 7975 12804 8116 12832
rect 7975 12801 7987 12804
rect 7929 12795 7987 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8478 12832 8484 12844
rect 8391 12804 8484 12832
rect 8478 12792 8484 12804
rect 8536 12832 8542 12844
rect 8754 12832 8760 12844
rect 8536 12804 8760 12832
rect 8536 12792 8542 12804
rect 8754 12792 8760 12804
rect 8812 12792 8818 12844
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2516 12736 2605 12764
rect 1670 12696 1676 12708
rect 1631 12668 1676 12696
rect 1670 12656 1676 12668
rect 1728 12656 1734 12708
rect 2516 12640 2544 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 2849 12767 2907 12773
rect 2849 12764 2861 12767
rect 2740 12736 2861 12764
rect 2740 12724 2746 12736
rect 2849 12733 2861 12736
rect 2895 12733 2907 12767
rect 2849 12727 2907 12733
rect 5810 12724 5816 12776
rect 5868 12724 5874 12776
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 7745 12767 7803 12773
rect 7745 12764 7757 12767
rect 7524 12736 7757 12764
rect 7524 12724 7530 12736
rect 7745 12733 7757 12736
rect 7791 12764 7803 12767
rect 8386 12764 8392 12776
rect 7791 12736 8392 12764
rect 7791 12733 7803 12736
rect 7745 12727 7803 12733
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 8938 12764 8944 12776
rect 8899 12736 8944 12764
rect 8938 12724 8944 12736
rect 8996 12724 9002 12776
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 7834 12696 7840 12708
rect 7331 12668 7840 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7834 12656 7840 12668
rect 7892 12656 7898 12708
rect 9208 12699 9266 12705
rect 9208 12665 9220 12699
rect 9254 12696 9266 12699
rect 9306 12696 9312 12708
rect 9254 12668 9312 12696
rect 9254 12665 9266 12668
rect 9208 12659 9266 12665
rect 9306 12656 9312 12668
rect 9364 12656 9370 12708
rect 2498 12628 2504 12640
rect 2459 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12588 2562 12640
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4062 12628 4068 12640
rect 4019 12600 4068 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 7466 12588 7472 12640
rect 7524 12628 7530 12640
rect 7650 12628 7656 12640
rect 7524 12600 7656 12628
rect 7524 12588 7530 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 10410 12588 10416 12640
rect 10468 12628 10474 12640
rect 10873 12631 10931 12637
rect 10873 12628 10885 12631
rect 10468 12600 10885 12628
rect 10468 12588 10474 12600
rect 10873 12597 10885 12600
rect 10919 12597 10931 12631
rect 10873 12591 10931 12597
rect 1104 12538 14812 12560
rect 1104 12486 6315 12538
rect 6367 12486 6379 12538
rect 6431 12486 6443 12538
rect 6495 12486 6507 12538
rect 6559 12486 11648 12538
rect 11700 12486 11712 12538
rect 11764 12486 11776 12538
rect 11828 12486 11840 12538
rect 11892 12486 14812 12538
rect 1104 12464 14812 12486
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 6086 12424 6092 12436
rect 6047 12396 6092 12424
rect 6086 12384 6092 12396
rect 6144 12384 6150 12436
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 6549 12427 6607 12433
rect 6549 12424 6561 12427
rect 6236 12396 6561 12424
rect 6236 12384 6242 12396
rect 6549 12393 6561 12396
rect 6595 12393 6607 12427
rect 6549 12387 6607 12393
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 7561 12427 7619 12433
rect 7561 12424 7573 12427
rect 6880 12396 7573 12424
rect 6880 12384 6886 12396
rect 7561 12393 7573 12396
rect 7607 12424 7619 12427
rect 7650 12424 7656 12436
rect 7607 12396 7656 12424
rect 7607 12393 7619 12396
rect 7561 12387 7619 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 8110 12424 8116 12436
rect 8071 12396 8116 12424
rect 8110 12384 8116 12396
rect 8168 12384 8174 12436
rect 8386 12384 8392 12436
rect 8444 12424 8450 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8444 12396 8585 12424
rect 8444 12384 8450 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 8573 12387 8631 12393
rect 9950 12384 9956 12436
rect 10008 12424 10014 12436
rect 10045 12427 10103 12433
rect 10045 12424 10057 12427
rect 10008 12396 10057 12424
rect 10008 12384 10014 12396
rect 10045 12393 10057 12396
rect 10091 12424 10103 12427
rect 10318 12424 10324 12436
rect 10091 12396 10324 12424
rect 10091 12393 10103 12396
rect 10045 12387 10103 12393
rect 10318 12384 10324 12396
rect 10376 12384 10382 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 12158 12424 12164 12436
rect 11747 12396 12164 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 4120 12328 4200 12356
rect 4120 12316 4126 12328
rect 4172 12288 4200 12328
rect 7006 12316 7012 12368
rect 7064 12356 7070 12368
rect 7190 12356 7196 12368
rect 7064 12328 7196 12356
rect 7064 12316 7070 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 11330 12356 11336 12368
rect 10428 12328 11336 12356
rect 4332 12291 4390 12297
rect 4332 12288 4344 12291
rect 4172 12260 4344 12288
rect 4332 12257 4344 12260
rect 4378 12288 4390 12291
rect 4614 12288 4620 12300
rect 4378 12260 4620 12288
rect 4378 12257 4390 12260
rect 4332 12251 4390 12257
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6380 12260 6929 12288
rect 2498 12180 2504 12232
rect 2556 12220 2562 12232
rect 4062 12220 4068 12232
rect 2556 12192 4068 12220
rect 2556 12180 2562 12192
rect 4062 12180 4068 12192
rect 4120 12180 4126 12232
rect 2590 12084 2596 12096
rect 2551 12056 2596 12084
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 6380 12093 6408 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 6638 12180 6644 12232
rect 6696 12220 6702 12232
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6696 12192 7021 12220
rect 6696 12180 6702 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7190 12220 7196 12232
rect 7103 12192 7196 12220
rect 7009 12183 7067 12189
rect 7190 12180 7196 12192
rect 7248 12220 7254 12232
rect 9306 12220 9312 12232
rect 7248 12192 9312 12220
rect 7248 12180 7254 12192
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10428 12220 10456 12328
rect 11330 12316 11336 12328
rect 11388 12316 11394 12368
rect 10594 12297 10600 12300
rect 10588 12288 10600 12297
rect 10555 12260 10600 12288
rect 10588 12251 10600 12260
rect 10594 12248 10600 12251
rect 10652 12248 10658 12300
rect 10367 12192 10456 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 8938 12112 8944 12164
rect 8996 12152 9002 12164
rect 9950 12152 9956 12164
rect 8996 12124 9956 12152
rect 8996 12112 9002 12124
rect 9950 12112 9956 12124
rect 10008 12152 10014 12164
rect 10336 12152 10364 12183
rect 10008 12124 10364 12152
rect 10008 12112 10014 12124
rect 6365 12087 6423 12093
rect 6365 12084 6377 12087
rect 5224 12056 6377 12084
rect 5224 12044 5230 12056
rect 6365 12053 6377 12056
rect 6411 12053 6423 12087
rect 6365 12047 6423 12053
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 8956 12084 8984 12112
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 7432 12056 9045 12084
rect 7432 12044 7438 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9033 12047 9091 12053
rect 1104 11994 14812 12016
rect 1104 11942 3648 11994
rect 3700 11942 3712 11994
rect 3764 11942 3776 11994
rect 3828 11942 3840 11994
rect 3892 11942 8982 11994
rect 9034 11942 9046 11994
rect 9098 11942 9110 11994
rect 9162 11942 9174 11994
rect 9226 11942 14315 11994
rect 14367 11942 14379 11994
rect 14431 11942 14443 11994
rect 14495 11942 14507 11994
rect 14559 11942 14812 11994
rect 1104 11920 14812 11942
rect 2409 11883 2467 11889
rect 2409 11849 2421 11883
rect 2455 11880 2467 11883
rect 2498 11880 2504 11892
rect 2455 11852 2504 11880
rect 2455 11849 2467 11852
rect 2409 11843 2467 11849
rect 2498 11840 2504 11852
rect 2556 11840 2562 11892
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 3881 11883 3939 11889
rect 3881 11880 3893 11883
rect 2740 11852 3893 11880
rect 2740 11840 2746 11852
rect 3881 11849 3893 11852
rect 3927 11849 3939 11883
rect 3881 11843 3939 11849
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4525 11883 4583 11889
rect 4525 11880 4537 11883
rect 4212 11852 4537 11880
rect 4212 11840 4218 11852
rect 4525 11849 4537 11852
rect 4571 11880 4583 11883
rect 4890 11880 4896 11892
rect 4571 11852 4896 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4890 11840 4896 11852
rect 4948 11840 4954 11892
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7190 11880 7196 11892
rect 6687 11852 7196 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 8757 11883 8815 11889
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 9306 11880 9312 11892
rect 8803 11852 9312 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9950 11840 9956 11892
rect 10008 11880 10014 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 10008 11852 10333 11880
rect 10008 11840 10014 11852
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 10321 11843 10379 11849
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10689 11883 10747 11889
rect 10689 11880 10701 11883
rect 10652 11852 10701 11880
rect 10652 11840 10658 11852
rect 10689 11849 10701 11852
rect 10735 11849 10747 11883
rect 10689 11843 10747 11849
rect 2516 11753 2544 11840
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 5629 11747 5687 11753
rect 5629 11744 5641 11747
rect 5500 11716 5641 11744
rect 5500 11704 5506 11716
rect 5629 11713 5641 11716
rect 5675 11744 5687 11747
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5675 11716 6009 11744
rect 5675 11713 5687 11716
rect 5629 11707 5687 11713
rect 5997 11713 6009 11716
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 2768 11679 2826 11685
rect 2768 11676 2780 11679
rect 2648 11648 2780 11676
rect 2648 11636 2654 11648
rect 2768 11645 2780 11648
rect 2814 11676 2826 11679
rect 5460 11676 5488 11704
rect 7374 11676 7380 11688
rect 2814 11648 5488 11676
rect 7208 11648 7380 11676
rect 2814 11645 2826 11648
rect 2768 11639 2826 11645
rect 3326 11568 3332 11620
rect 3384 11608 3390 11620
rect 4893 11611 4951 11617
rect 3384 11580 4016 11608
rect 3384 11568 3390 11580
rect 3988 11540 4016 11580
rect 4893 11577 4905 11611
rect 4939 11608 4951 11611
rect 5445 11611 5503 11617
rect 5445 11608 5457 11611
rect 4939 11580 5457 11608
rect 4939 11577 4951 11580
rect 4893 11571 4951 11577
rect 5445 11577 5457 11580
rect 5491 11608 5503 11611
rect 5626 11608 5632 11620
rect 5491 11580 5632 11608
rect 5491 11577 5503 11580
rect 5445 11571 5503 11577
rect 5626 11568 5632 11580
rect 5684 11608 5690 11620
rect 6178 11608 6184 11620
rect 5684 11580 6184 11608
rect 5684 11568 5690 11580
rect 6178 11568 6184 11580
rect 6236 11568 6242 11620
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 3988 11512 4997 11540
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5132 11512 5365 11540
rect 5132 11500 5138 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 7208 11549 7236 11648
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7650 11685 7656 11688
rect 7644 11676 7656 11685
rect 7611 11648 7656 11676
rect 7644 11639 7656 11648
rect 7650 11636 7656 11639
rect 7708 11636 7714 11688
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6788 11512 7205 11540
rect 6788 11500 6794 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 7193 11503 7251 11509
rect 1104 11450 14812 11472
rect 1104 11398 6315 11450
rect 6367 11398 6379 11450
rect 6431 11398 6443 11450
rect 6495 11398 6507 11450
rect 6559 11398 11648 11450
rect 11700 11398 11712 11450
rect 11764 11398 11776 11450
rect 11828 11398 11840 11450
rect 11892 11398 14812 11450
rect 1104 11376 14812 11398
rect 4157 11339 4215 11345
rect 4157 11305 4169 11339
rect 4203 11336 4215 11339
rect 5074 11336 5080 11348
rect 4203 11308 5080 11336
rect 4203 11305 4215 11308
rect 4157 11299 4215 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5166 11296 5172 11348
rect 5224 11336 5230 11348
rect 5224 11308 5269 11336
rect 5224 11296 5230 11308
rect 5350 11296 5356 11348
rect 5408 11296 5414 11348
rect 6638 11336 6644 11348
rect 6599 11308 6644 11336
rect 6638 11296 6644 11308
rect 6696 11296 6702 11348
rect 7650 11296 7656 11348
rect 7708 11336 7714 11348
rect 8113 11339 8171 11345
rect 8113 11336 8125 11339
rect 7708 11308 8125 11336
rect 7708 11296 7714 11308
rect 8113 11305 8125 11308
rect 8159 11305 8171 11339
rect 8113 11299 8171 11305
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11268 2835 11271
rect 2958 11268 2964 11280
rect 2823 11240 2964 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 4614 11268 4620 11280
rect 4575 11240 4620 11268
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 2556 11172 3096 11200
rect 2556 11160 2562 11172
rect 3068 11141 3096 11172
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 4632 11132 4660 11228
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 5368 11200 5396 11296
rect 7000 11271 7058 11277
rect 7000 11237 7012 11271
rect 7046 11268 7058 11271
rect 7558 11268 7564 11280
rect 7046 11240 7564 11268
rect 7046 11237 7058 11240
rect 7000 11231 7058 11237
rect 7558 11228 7564 11240
rect 7616 11228 7622 11280
rect 5534 11200 5540 11212
rect 5224 11172 5396 11200
rect 5495 11172 5540 11200
rect 5224 11160 5230 11172
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 5626 11132 5632 11144
rect 3099 11104 4660 11132
rect 5587 11104 5632 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 2774 11024 2780 11076
rect 2832 11064 2838 11076
rect 2884 11064 2912 11095
rect 5626 11092 5632 11104
rect 5684 11092 5690 11144
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 5776 11104 5821 11132
rect 5776 11092 5782 11104
rect 6086 11092 6092 11144
rect 6144 11132 6150 11144
rect 6730 11132 6736 11144
rect 6144 11104 6736 11132
rect 6144 11092 6150 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 2832 11036 2912 11064
rect 2832 11024 2838 11036
rect 5258 11024 5264 11076
rect 5316 11064 5322 11076
rect 5736 11064 5764 11092
rect 5316 11036 5764 11064
rect 5316 11024 5322 11036
rect 1394 10956 1400 11008
rect 1452 10996 1458 11008
rect 2409 10999 2467 11005
rect 2409 10996 2421 10999
rect 1452 10968 2421 10996
rect 1452 10956 1458 10968
rect 2409 10965 2421 10968
rect 2455 10965 2467 10999
rect 2409 10959 2467 10965
rect 1104 10906 14812 10928
rect 1104 10854 3648 10906
rect 3700 10854 3712 10906
rect 3764 10854 3776 10906
rect 3828 10854 3840 10906
rect 3892 10854 8982 10906
rect 9034 10854 9046 10906
rect 9098 10854 9110 10906
rect 9162 10854 9174 10906
rect 9226 10854 14315 10906
rect 14367 10854 14379 10906
rect 14431 10854 14443 10906
rect 14495 10854 14507 10906
rect 14559 10854 14812 10906
rect 1104 10832 14812 10854
rect 2498 10792 2504 10804
rect 2459 10764 2504 10792
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 2682 10752 2688 10804
rect 2740 10792 2746 10804
rect 2777 10795 2835 10801
rect 2777 10792 2789 10795
rect 2740 10764 2789 10792
rect 2740 10752 2746 10764
rect 2777 10761 2789 10764
rect 2823 10761 2835 10795
rect 2958 10792 2964 10804
rect 2919 10764 2964 10792
rect 2777 10755 2835 10761
rect 2958 10752 2964 10764
rect 3016 10752 3022 10804
rect 2133 10727 2191 10733
rect 2133 10693 2145 10727
rect 2179 10724 2191 10727
rect 4525 10727 4583 10733
rect 4525 10724 4537 10727
rect 2179 10696 4537 10724
rect 2179 10693 2191 10696
rect 2133 10687 2191 10693
rect 3326 10588 3332 10600
rect 3287 10560 3332 10588
rect 3326 10548 3332 10560
rect 3384 10548 3390 10600
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10588 3479 10591
rect 3528 10588 3556 10696
rect 4525 10693 4537 10696
rect 4571 10693 4583 10727
rect 4525 10687 4583 10693
rect 5626 10684 5632 10736
rect 5684 10724 5690 10736
rect 6825 10727 6883 10733
rect 6825 10724 6837 10727
rect 5684 10696 6837 10724
rect 5684 10684 5690 10696
rect 6825 10693 6837 10696
rect 6871 10693 6883 10727
rect 6825 10687 6883 10693
rect 3605 10659 3663 10665
rect 3605 10625 3617 10659
rect 3651 10656 3663 10659
rect 3694 10656 3700 10668
rect 3651 10628 3700 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5442 10656 5448 10668
rect 5215 10628 5448 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10656 5963 10659
rect 6086 10656 6092 10668
rect 5951 10628 6092 10656
rect 5951 10625 5963 10628
rect 5905 10619 5963 10625
rect 6086 10616 6092 10628
rect 6144 10616 6150 10668
rect 7469 10659 7527 10665
rect 7469 10625 7481 10659
rect 7515 10656 7527 10659
rect 7558 10656 7564 10668
rect 7515 10628 7564 10656
rect 7515 10625 7527 10628
rect 7469 10619 7527 10625
rect 7558 10616 7564 10628
rect 7616 10656 7622 10668
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7616 10628 7849 10656
rect 7616 10616 7622 10628
rect 7837 10625 7849 10628
rect 7883 10625 7895 10659
rect 7837 10619 7895 10625
rect 3467 10560 3556 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 4890 10548 4896 10600
rect 4948 10548 4954 10600
rect 4908 10520 4936 10548
rect 4985 10523 5043 10529
rect 4985 10520 4997 10523
rect 3988 10492 4997 10520
rect 1765 10455 1823 10461
rect 1765 10421 1777 10455
rect 1811 10452 1823 10455
rect 2406 10452 2412 10464
rect 1811 10424 2412 10452
rect 1811 10421 1823 10424
rect 1765 10415 1823 10421
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 3234 10412 3240 10464
rect 3292 10452 3298 10464
rect 3988 10461 4016 10492
rect 4985 10489 4997 10492
rect 5031 10489 5043 10523
rect 5902 10520 5908 10532
rect 4985 10483 5043 10489
rect 5736 10492 5908 10520
rect 3973 10455 4031 10461
rect 3973 10452 3985 10455
rect 3292 10424 3985 10452
rect 3292 10412 3298 10424
rect 3973 10421 3985 10424
rect 4019 10421 4031 10455
rect 3973 10415 4031 10421
rect 4433 10455 4491 10461
rect 4433 10421 4445 10455
rect 4479 10452 4491 10455
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 4479 10424 4905 10452
rect 4479 10421 4491 10424
rect 4433 10415 4491 10421
rect 4893 10421 4905 10424
rect 4939 10452 4951 10455
rect 5736 10452 5764 10492
rect 5902 10480 5908 10492
rect 5960 10520 5966 10532
rect 6641 10523 6699 10529
rect 6641 10520 6653 10523
rect 5960 10492 6653 10520
rect 5960 10480 5966 10492
rect 6641 10489 6653 10492
rect 6687 10520 6699 10523
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 6687 10492 7205 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7193 10489 7205 10492
rect 7239 10520 7251 10523
rect 7374 10520 7380 10532
rect 7239 10492 7380 10520
rect 7239 10489 7251 10492
rect 7193 10483 7251 10489
rect 7374 10480 7380 10492
rect 7432 10480 7438 10532
rect 4939 10424 5764 10452
rect 4939 10421 4951 10424
rect 4893 10415 4951 10421
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5868 10424 6285 10452
rect 5868 10412 5874 10424
rect 6273 10421 6285 10424
rect 6319 10452 6331 10455
rect 7282 10452 7288 10464
rect 6319 10424 7288 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 8386 10452 8392 10464
rect 8347 10424 8392 10452
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 12437 10455 12495 10461
rect 12437 10421 12449 10455
rect 12483 10452 12495 10455
rect 13354 10452 13360 10464
rect 12483 10424 13360 10452
rect 12483 10421 12495 10424
rect 12437 10415 12495 10421
rect 13354 10412 13360 10424
rect 13412 10412 13418 10464
rect 1104 10362 14812 10384
rect 1104 10310 6315 10362
rect 6367 10310 6379 10362
rect 6431 10310 6443 10362
rect 6495 10310 6507 10362
rect 6559 10310 11648 10362
rect 11700 10310 11712 10362
rect 11764 10310 11776 10362
rect 11828 10310 11840 10362
rect 11892 10310 14812 10362
rect 1104 10288 14812 10310
rect 1578 10248 1584 10260
rect 1539 10220 1584 10248
rect 1578 10208 1584 10220
rect 1636 10208 1642 10260
rect 2406 10248 2412 10260
rect 2367 10220 2412 10248
rect 2406 10208 2412 10220
rect 2464 10248 2470 10260
rect 2682 10248 2688 10260
rect 2464 10220 2688 10248
rect 2464 10208 2470 10220
rect 2682 10208 2688 10220
rect 2740 10208 2746 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 3421 10251 3479 10257
rect 3421 10248 3433 10251
rect 3384 10220 3433 10248
rect 3384 10208 3390 10220
rect 3421 10217 3433 10220
rect 3467 10217 3479 10251
rect 5258 10248 5264 10260
rect 5219 10220 5264 10248
rect 3421 10211 3479 10217
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5905 10251 5963 10257
rect 5905 10248 5917 10251
rect 5592 10220 5917 10248
rect 5592 10208 5598 10220
rect 5905 10217 5917 10220
rect 5951 10248 5963 10251
rect 6549 10251 6607 10257
rect 6549 10248 6561 10251
rect 5951 10220 6561 10248
rect 5951 10217 5963 10220
rect 5905 10211 5963 10217
rect 6549 10217 6561 10220
rect 6595 10217 6607 10251
rect 6549 10211 6607 10217
rect 6917 10251 6975 10257
rect 6917 10217 6929 10251
rect 6963 10248 6975 10251
rect 7098 10248 7104 10260
rect 6963 10220 7104 10248
rect 6963 10217 6975 10220
rect 6917 10211 6975 10217
rect 7098 10208 7104 10220
rect 7156 10248 7162 10260
rect 8386 10248 8392 10260
rect 7156 10220 8392 10248
rect 7156 10208 7162 10220
rect 8386 10208 8392 10220
rect 8444 10208 8450 10260
rect 9950 10208 9956 10260
rect 10008 10208 10014 10260
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10180 2375 10183
rect 2958 10180 2964 10192
rect 2363 10152 2964 10180
rect 2363 10149 2375 10152
rect 2317 10143 2375 10149
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 4893 10183 4951 10189
rect 4893 10149 4905 10183
rect 4939 10180 4951 10183
rect 5074 10180 5080 10192
rect 4939 10152 5080 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 5074 10140 5080 10152
rect 5132 10180 5138 10192
rect 5442 10180 5448 10192
rect 5132 10152 5448 10180
rect 5132 10140 5138 10152
rect 5442 10140 5448 10152
rect 5500 10140 5506 10192
rect 5626 10180 5632 10192
rect 5587 10152 5632 10180
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 7558 10180 7564 10192
rect 7519 10152 7564 10180
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 1394 10112 1400 10124
rect 1355 10084 1400 10112
rect 1394 10072 1400 10084
rect 1452 10072 1458 10124
rect 2774 10072 2780 10124
rect 2832 10112 2838 10124
rect 4062 10112 4068 10124
rect 2832 10084 4068 10112
rect 2832 10072 2838 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 6822 10072 6828 10124
rect 6880 10112 6886 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6880 10084 7021 10112
rect 6880 10072 6886 10084
rect 7009 10081 7021 10084
rect 7055 10112 7067 10115
rect 7374 10112 7380 10124
rect 7055 10084 7380 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7374 10072 7380 10084
rect 7432 10072 7438 10124
rect 2866 10044 2872 10056
rect 2827 10016 2872 10044
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3053 10047 3111 10053
rect 3053 10013 3065 10047
rect 3099 10044 3111 10047
rect 3694 10044 3700 10056
rect 3099 10016 3700 10044
rect 3099 10013 3111 10016
rect 3053 10007 3111 10013
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 2958 9976 2964 9988
rect 2648 9948 2964 9976
rect 2648 9936 2654 9948
rect 2958 9936 2964 9948
rect 3016 9976 3022 9988
rect 3068 9976 3096 10007
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 7193 10047 7251 10053
rect 7193 10013 7205 10047
rect 7239 10044 7251 10047
rect 7576 10044 7604 10140
rect 9968 10112 9996 10208
rect 10686 10140 10692 10192
rect 10744 10189 10750 10192
rect 10744 10183 10808 10189
rect 10744 10149 10762 10183
rect 10796 10149 10808 10183
rect 10744 10143 10808 10149
rect 10744 10140 10750 10143
rect 10505 10115 10563 10121
rect 10505 10112 10517 10115
rect 9968 10084 10517 10112
rect 10505 10081 10517 10084
rect 10551 10081 10563 10115
rect 13446 10112 13452 10124
rect 13407 10084 13452 10112
rect 10505 10075 10563 10081
rect 13446 10072 13452 10084
rect 13504 10072 13510 10124
rect 7239 10016 7604 10044
rect 7239 10013 7251 10016
rect 7193 10007 7251 10013
rect 12894 10004 12900 10056
rect 12952 10044 12958 10056
rect 13541 10047 13599 10053
rect 13541 10044 13553 10047
rect 12952 10016 13553 10044
rect 12952 10004 12958 10016
rect 13541 10013 13553 10016
rect 13587 10013 13599 10047
rect 13541 10007 13599 10013
rect 3016 9948 3096 9976
rect 3016 9936 3022 9948
rect 4522 9908 4528 9920
rect 4483 9880 4528 9908
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10870 9908 10876 9920
rect 10459 9880 10876 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 11885 9911 11943 9917
rect 11885 9877 11897 9911
rect 11931 9908 11943 9911
rect 11974 9908 11980 9920
rect 11931 9880 11980 9908
rect 11931 9877 11943 9880
rect 11885 9871 11943 9877
rect 11974 9868 11980 9880
rect 12032 9908 12038 9920
rect 12437 9911 12495 9917
rect 12437 9908 12449 9911
rect 12032 9880 12449 9908
rect 12032 9868 12038 9880
rect 12437 9877 12449 9880
rect 12483 9908 12495 9911
rect 12526 9908 12532 9920
rect 12483 9880 12532 9908
rect 12483 9877 12495 9880
rect 12437 9871 12495 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12802 9868 12808 9920
rect 12860 9908 12866 9920
rect 12897 9911 12955 9917
rect 12897 9908 12909 9911
rect 12860 9880 12909 9908
rect 12860 9868 12866 9880
rect 12897 9877 12909 9880
rect 12943 9908 12955 9911
rect 12989 9911 13047 9917
rect 12989 9908 13001 9911
rect 12943 9880 13001 9908
rect 12943 9877 12955 9880
rect 12897 9871 12955 9877
rect 12989 9877 13001 9880
rect 13035 9877 13047 9911
rect 12989 9871 13047 9877
rect 1104 9818 14812 9840
rect 1104 9766 3648 9818
rect 3700 9766 3712 9818
rect 3764 9766 3776 9818
rect 3828 9766 3840 9818
rect 3892 9766 8982 9818
rect 9034 9766 9046 9818
rect 9098 9766 9110 9818
rect 9162 9766 9174 9818
rect 9226 9766 14315 9818
rect 14367 9766 14379 9818
rect 14431 9766 14443 9818
rect 14495 9766 14507 9818
rect 14559 9766 14812 9818
rect 1104 9744 14812 9766
rect 2866 9704 2872 9716
rect 2827 9676 2872 9704
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 2958 9664 2964 9716
rect 3016 9664 3022 9716
rect 7098 9704 7104 9716
rect 7059 9676 7104 9704
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7469 9707 7527 9713
rect 7469 9673 7481 9707
rect 7515 9704 7527 9707
rect 7558 9704 7564 9716
rect 7515 9676 7564 9704
rect 7515 9673 7527 9676
rect 7469 9667 7527 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 9916 9676 10517 9704
rect 9916 9664 9922 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 12894 9704 12900 9716
rect 10505 9667 10563 9673
rect 12360 9676 12900 9704
rect 2976 9636 3004 9664
rect 2875 9608 3004 9636
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2875 9568 2903 9608
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4433 9639 4491 9645
rect 4433 9636 4445 9639
rect 4120 9608 4445 9636
rect 4120 9596 4126 9608
rect 4433 9605 4445 9608
rect 4479 9605 4491 9639
rect 4433 9599 4491 9605
rect 7006 9596 7012 9648
rect 7064 9596 7070 9648
rect 12253 9639 12311 9645
rect 12253 9605 12265 9639
rect 12299 9636 12311 9639
rect 12360 9636 12388 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13412 9676 13768 9704
rect 13412 9664 13418 9676
rect 12299 9608 12388 9636
rect 12437 9639 12495 9645
rect 12299 9605 12311 9608
rect 12253 9599 12311 9605
rect 12437 9605 12449 9639
rect 12483 9605 12495 9639
rect 13446 9636 13452 9648
rect 13407 9608 13452 9636
rect 12437 9599 12495 9605
rect 2455 9540 2903 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 2958 9528 2964 9580
rect 3016 9568 3022 9580
rect 3513 9571 3571 9577
rect 3513 9568 3525 9571
rect 3016 9540 3525 9568
rect 3016 9528 3022 9540
rect 3513 9537 3525 9540
rect 3559 9568 3571 9571
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3559 9540 3985 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3973 9537 3985 9540
rect 4019 9568 4031 9571
rect 5074 9568 5080 9580
rect 4019 9540 5080 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2682 9500 2688 9512
rect 1719 9472 2688 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 2823 9472 3249 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 3237 9469 3249 9472
rect 3283 9500 3295 9503
rect 3326 9500 3332 9512
rect 3283 9472 3332 9500
rect 3283 9469 3295 9472
rect 3237 9463 3295 9469
rect 3326 9460 3332 9472
rect 3384 9460 3390 9512
rect 3418 9460 3424 9512
rect 3476 9500 3482 9512
rect 6178 9500 6184 9512
rect 3476 9472 6184 9500
rect 3476 9460 3482 9472
rect 6178 9460 6184 9472
rect 6236 9500 6242 9512
rect 6549 9503 6607 9509
rect 6549 9500 6561 9503
rect 6236 9472 6561 9500
rect 6236 9460 6242 9472
rect 6549 9469 6561 9472
rect 6595 9500 6607 9503
rect 6822 9500 6828 9512
rect 6595 9472 6828 9500
rect 6595 9469 6607 9472
rect 6549 9463 6607 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 2041 9435 2099 9441
rect 2041 9401 2053 9435
rect 2087 9432 2099 9435
rect 2087 9404 3372 9432
rect 2087 9401 2099 9404
rect 2041 9395 2099 9401
rect 3344 9376 3372 9404
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4580 9404 4905 9432
rect 4580 9392 4586 9404
rect 4893 9401 4905 9404
rect 4939 9432 4951 9435
rect 7024 9432 7052 9596
rect 9306 9528 9312 9580
rect 9364 9568 9370 9580
rect 9674 9568 9680 9580
rect 9364 9540 9680 9568
rect 9364 9528 9370 9540
rect 9674 9528 9680 9540
rect 9732 9528 9738 9580
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 10686 9568 10692 9580
rect 9907 9540 10692 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 9125 9503 9183 9509
rect 9125 9469 9137 9503
rect 9171 9500 9183 9503
rect 9876 9500 9904 9531
rect 10686 9528 10692 9540
rect 10744 9528 10750 9580
rect 10962 9528 10968 9580
rect 11020 9568 11026 9580
rect 11333 9571 11391 9577
rect 11333 9568 11345 9571
rect 11020 9540 11345 9568
rect 11020 9528 11026 9540
rect 11333 9537 11345 9540
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 9171 9472 9904 9500
rect 9171 9469 9183 9472
rect 9125 9463 9183 9469
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 10928 9472 11161 9500
rect 10928 9460 10934 9472
rect 11149 9469 11161 9472
rect 11195 9500 11207 9503
rect 12452 9500 12480 9599
rect 13446 9596 13452 9608
rect 13504 9596 13510 9648
rect 13740 9636 13768 9676
rect 13817 9639 13875 9645
rect 13817 9636 13829 9639
rect 13740 9608 13829 9636
rect 13817 9605 13829 9608
rect 13863 9605 13875 9639
rect 13817 9599 13875 9605
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12584 9540 13001 9568
rect 12584 9528 12590 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 12802 9500 12808 9512
rect 11195 9472 12480 9500
rect 12763 9472 12808 9500
rect 11195 9469 11207 9472
rect 11149 9463 11207 9469
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 7558 9432 7564 9444
rect 4939 9404 7564 9432
rect 4939 9401 4951 9404
rect 4893 9395 4951 9401
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 9585 9435 9643 9441
rect 9585 9432 9597 9435
rect 8680 9404 9597 9432
rect 8680 9376 8708 9404
rect 9585 9401 9597 9404
rect 9631 9401 9643 9435
rect 9585 9395 9643 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11241 9435 11299 9441
rect 11241 9432 11253 9435
rect 11112 9404 11253 9432
rect 11112 9392 11118 9404
rect 11241 9401 11253 9404
rect 11287 9401 11299 9435
rect 11241 9395 11299 9401
rect 3326 9364 3332 9376
rect 3287 9336 3332 9364
rect 3326 9324 3332 9336
rect 3384 9324 3390 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4387 9336 4813 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4801 9333 4813 9336
rect 4847 9364 4859 9367
rect 5994 9364 6000 9376
rect 4847 9336 6000 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 5994 9324 6000 9336
rect 6052 9324 6058 9376
rect 8662 9364 8668 9376
rect 8623 9336 8668 9364
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9214 9364 9220 9376
rect 9175 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9324 9278 9376
rect 10778 9364 10784 9376
rect 10739 9336 10784 9364
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 12434 9364 12440 9376
rect 11931 9336 12440 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 12434 9324 12440 9336
rect 12492 9364 12498 9376
rect 12897 9367 12955 9373
rect 12897 9364 12909 9367
rect 12492 9336 12909 9364
rect 12492 9324 12498 9336
rect 12897 9333 12909 9336
rect 12943 9333 12955 9367
rect 12897 9327 12955 9333
rect 1104 9274 14812 9296
rect 1104 9222 6315 9274
rect 6367 9222 6379 9274
rect 6431 9222 6443 9274
rect 6495 9222 6507 9274
rect 6559 9222 11648 9274
rect 11700 9222 11712 9274
rect 11764 9222 11776 9274
rect 11828 9222 11840 9274
rect 11892 9222 14812 9274
rect 1104 9200 14812 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1452 9132 1593 9160
rect 1452 9120 1458 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2501 9163 2559 9169
rect 2501 9129 2513 9163
rect 2547 9160 2559 9163
rect 2866 9160 2872 9172
rect 2547 9132 2872 9160
rect 2547 9129 2559 9132
rect 2501 9123 2559 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 2958 9120 2964 9172
rect 3016 9160 3022 9172
rect 3016 9132 3061 9160
rect 3016 9120 3022 9132
rect 5074 9120 5080 9172
rect 5132 9160 5138 9172
rect 5445 9163 5503 9169
rect 5445 9160 5457 9163
rect 5132 9132 5457 9160
rect 5132 9120 5138 9132
rect 5445 9129 5457 9132
rect 5491 9129 5503 9163
rect 5445 9123 5503 9129
rect 8389 9163 8447 9169
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8846 9160 8852 9172
rect 8435 9132 8852 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 10134 9160 10140 9172
rect 10095 9132 10140 9160
rect 10134 9120 10140 9132
rect 10192 9120 10198 9172
rect 10226 9120 10232 9172
rect 10284 9160 10290 9172
rect 10778 9160 10784 9172
rect 10284 9132 10784 9160
rect 10284 9120 10290 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9092 3479 9095
rect 4246 9092 4252 9104
rect 3467 9064 4252 9092
rect 3467 9061 3479 9064
rect 3421 9055 3479 9061
rect 4246 9052 4252 9064
rect 4304 9101 4310 9104
rect 4304 9095 4368 9101
rect 4304 9061 4322 9095
rect 4356 9061 4368 9095
rect 4304 9055 4368 9061
rect 4304 9052 4310 9055
rect 9858 9052 9864 9104
rect 9916 9092 9922 9104
rect 11974 9101 11980 9104
rect 11968 9092 11980 9101
rect 9916 9064 11744 9092
rect 11935 9064 11980 9092
rect 9916 9052 9922 9064
rect 11716 9036 11744 9064
rect 11968 9055 11980 9064
rect 11974 9052 11980 9055
rect 12032 9052 12038 9104
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7742 9024 7748 9036
rect 7432 8996 7748 9024
rect 7432 8984 7438 8996
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 9950 8984 9956 9036
rect 10008 9024 10014 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 10008 8996 10057 9024
rect 10008 8984 10014 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 11698 9024 11704 9036
rect 11611 8996 11704 9024
rect 10045 8987 10103 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 4028 8928 4077 8956
rect 4028 8916 4034 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 8478 8956 8484 8968
rect 8439 8928 8484 8956
rect 4065 8919 4123 8925
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 8573 8959 8631 8965
rect 8573 8925 8585 8959
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 8588 8888 8616 8919
rect 9033 8891 9091 8897
rect 9033 8888 9045 8891
rect 7852 8860 9045 8888
rect 7852 8832 7880 8860
rect 9033 8857 9045 8860
rect 9079 8888 9091 8891
rect 10226 8888 10232 8900
rect 9079 8860 10232 8888
rect 9079 8857 9091 8860
rect 9033 8851 9091 8857
rect 10226 8848 10232 8860
rect 10284 8888 10290 8900
rect 10336 8888 10364 8919
rect 10284 8860 10364 8888
rect 10284 8848 10290 8860
rect 10686 8848 10692 8900
rect 10744 8888 10750 8900
rect 10744 8860 11008 8888
rect 10744 8848 10750 8860
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8820 7435 8823
rect 7558 8820 7564 8832
rect 7423 8792 7564 8820
rect 7423 8789 7435 8792
rect 7377 8783 7435 8789
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 7834 8820 7840 8832
rect 7795 8792 7840 8820
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 8018 8820 8024 8832
rect 7979 8792 8024 8820
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 10870 8820 10876 8832
rect 10831 8792 10876 8820
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 10980 8820 11008 8860
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 11517 8891 11575 8897
rect 11517 8888 11529 8891
rect 11112 8860 11529 8888
rect 11112 8848 11118 8860
rect 11517 8857 11529 8860
rect 11563 8857 11575 8891
rect 11517 8851 11575 8857
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 10980 8792 11253 8820
rect 11241 8789 11253 8792
rect 11287 8820 11299 8823
rect 12894 8820 12900 8832
rect 11287 8792 12900 8820
rect 11287 8789 11299 8792
rect 11241 8783 11299 8789
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13078 8820 13084 8832
rect 13039 8792 13084 8820
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 1104 8730 14812 8752
rect 1104 8678 3648 8730
rect 3700 8678 3712 8730
rect 3764 8678 3776 8730
rect 3828 8678 3840 8730
rect 3892 8678 8982 8730
rect 9034 8678 9046 8730
rect 9098 8678 9110 8730
rect 9162 8678 9174 8730
rect 9226 8678 14315 8730
rect 14367 8678 14379 8730
rect 14431 8678 14443 8730
rect 14495 8678 14507 8730
rect 14559 8678 14812 8730
rect 1104 8656 14812 8678
rect 3326 8616 3332 8628
rect 3287 8588 3332 8616
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 7285 8619 7343 8625
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 8662 8616 8668 8628
rect 7331 8588 8668 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 8662 8576 8668 8588
rect 8720 8576 8726 8628
rect 8757 8619 8815 8625
rect 8757 8585 8769 8619
rect 8803 8616 8815 8619
rect 8846 8616 8852 8628
rect 8803 8588 8852 8616
rect 8803 8585 8815 8588
rect 8757 8579 8815 8585
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8616 10287 8619
rect 10686 8616 10692 8628
rect 10275 8588 10692 8616
rect 10275 8585 10287 8588
rect 10229 8579 10287 8585
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 11425 8619 11483 8625
rect 11425 8616 11437 8619
rect 11388 8588 11437 8616
rect 11388 8576 11394 8588
rect 11425 8585 11437 8588
rect 11471 8616 11483 8619
rect 11974 8616 11980 8628
rect 11471 8588 11980 8616
rect 11471 8585 11483 8588
rect 11425 8579 11483 8585
rect 11974 8576 11980 8588
rect 12032 8576 12038 8628
rect 12434 8616 12440 8628
rect 12395 8588 12440 8616
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 9950 8508 9956 8560
rect 10008 8548 10014 8560
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10008 8520 10793 8548
rect 10008 8508 10014 8520
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 11698 8548 11704 8560
rect 11659 8520 11704 8548
rect 10781 8511 10839 8517
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8480 3295 8483
rect 3786 8480 3792 8492
rect 3283 8452 3792 8480
rect 3283 8449 3295 8452
rect 3237 8443 3295 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8480 4031 8483
rect 4246 8480 4252 8492
rect 4019 8452 4252 8480
rect 4019 8449 4031 8452
rect 3973 8443 4031 8449
rect 4246 8440 4252 8452
rect 4304 8480 4310 8492
rect 7834 8480 7840 8492
rect 4304 8452 4752 8480
rect 7747 8452 7840 8480
rect 4304 8440 4310 8452
rect 2682 8304 2688 8356
rect 2740 8344 2746 8356
rect 3970 8344 3976 8356
rect 2740 8316 3976 8344
rect 2740 8304 2746 8316
rect 3970 8304 3976 8316
rect 4028 8344 4034 8356
rect 4028 8316 4476 8344
rect 4028 8304 4034 8316
rect 3694 8276 3700 8288
rect 3655 8248 3700 8276
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4448 8285 4476 8316
rect 4724 8288 4752 8452
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 8389 8483 8447 8489
rect 8389 8449 8401 8483
rect 8435 8480 8447 8483
rect 8478 8480 8484 8492
rect 8435 8452 8484 8480
rect 8435 8449 8447 8452
rect 8389 8443 8447 8449
rect 8478 8440 8484 8452
rect 8536 8480 8542 8492
rect 8536 8452 8984 8480
rect 8536 8440 8542 8452
rect 6546 8412 6552 8424
rect 6507 8384 6552 8412
rect 6546 8372 6552 8384
rect 6604 8412 6610 8424
rect 7852 8412 7880 8440
rect 6604 8384 7880 8412
rect 6604 8372 6610 8384
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 6914 8344 6920 8356
rect 6319 8316 6920 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7193 8347 7251 8353
rect 7193 8313 7205 8347
rect 7239 8344 7251 8347
rect 7374 8344 7380 8356
rect 7239 8316 7380 8344
rect 7239 8313 7251 8316
rect 7193 8307 7251 8313
rect 7374 8304 7380 8316
rect 7432 8344 7438 8356
rect 7432 8316 7512 8344
rect 7432 8304 7438 8316
rect 4433 8279 4491 8285
rect 4433 8245 4445 8279
rect 4479 8276 4491 8279
rect 4522 8276 4528 8288
rect 4479 8248 4528 8276
rect 4479 8245 4491 8248
rect 4433 8239 4491 8245
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4706 8276 4712 8288
rect 4667 8248 4712 8276
rect 4706 8236 4712 8248
rect 4764 8236 4770 8288
rect 7484 8276 7512 8316
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7653 8347 7711 8353
rect 7653 8344 7665 8347
rect 7616 8316 7665 8344
rect 7616 8304 7622 8316
rect 7653 8313 7665 8316
rect 7699 8313 7711 8347
rect 7653 8307 7711 8313
rect 7745 8347 7803 8353
rect 7745 8313 7757 8347
rect 7791 8313 7803 8347
rect 7852 8344 7880 8384
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8720 8384 8861 8412
rect 8720 8372 8726 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8956 8412 8984 8452
rect 12894 8440 12900 8492
rect 12952 8480 12958 8492
rect 12989 8483 13047 8489
rect 12989 8480 13001 8483
rect 12952 8452 13001 8480
rect 12952 8440 12958 8452
rect 12989 8449 13001 8452
rect 13035 8449 13047 8483
rect 12989 8443 13047 8449
rect 9582 8412 9588 8424
rect 8956 8384 9588 8412
rect 8849 8375 8907 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 12253 8415 12311 8421
rect 12253 8412 12265 8415
rect 11296 8384 12265 8412
rect 11296 8372 11302 8384
rect 12253 8381 12265 8384
rect 12299 8412 12311 8415
rect 12299 8384 12848 8412
rect 12299 8381 12311 8384
rect 12253 8375 12311 8381
rect 12820 8353 12848 8384
rect 9094 8347 9152 8353
rect 9094 8344 9106 8347
rect 7852 8316 9106 8344
rect 7745 8307 7803 8313
rect 9094 8313 9106 8316
rect 9140 8313 9152 8347
rect 9094 8307 9152 8313
rect 12805 8347 12863 8353
rect 12805 8313 12817 8347
rect 12851 8344 12863 8347
rect 13170 8344 13176 8356
rect 12851 8316 13176 8344
rect 12851 8313 12863 8316
rect 12805 8307 12863 8313
rect 7760 8276 7788 8307
rect 13170 8304 13176 8316
rect 13228 8304 13234 8356
rect 8018 8276 8024 8288
rect 7484 8248 8024 8276
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 12894 8276 12900 8288
rect 12855 8248 12900 8276
rect 12894 8236 12900 8248
rect 12952 8236 12958 8288
rect 1104 8186 14812 8208
rect 1104 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 11648 8186
rect 11700 8134 11712 8186
rect 11764 8134 11776 8186
rect 11828 8134 11840 8186
rect 11892 8134 14812 8186
rect 1104 8112 14812 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 1857 8075 1915 8081
rect 1857 8072 1869 8075
rect 1820 8044 1869 8072
rect 1820 8032 1826 8044
rect 1857 8041 1869 8044
rect 1903 8072 1915 8075
rect 2682 8072 2688 8084
rect 1903 8044 2688 8072
rect 1903 8041 1915 8044
rect 1857 8035 1915 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 3418 8072 3424 8084
rect 3331 8044 3424 8072
rect 3418 8032 3424 8044
rect 3476 8072 3482 8084
rect 3694 8072 3700 8084
rect 3476 8044 3700 8072
rect 3476 8032 3482 8044
rect 3694 8032 3700 8044
rect 3752 8072 3758 8084
rect 8754 8072 8760 8084
rect 3752 8044 8760 8072
rect 3752 8032 3758 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 10134 8072 10140 8084
rect 9640 8044 10140 8072
rect 9640 8032 9646 8044
rect 10134 8032 10140 8044
rect 10192 8032 10198 8084
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 10284 8044 10517 8072
rect 10284 8032 10290 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 11054 8072 11060 8084
rect 10735 8044 11060 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 11054 8032 11060 8044
rect 11112 8032 11118 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 12529 8075 12587 8081
rect 11204 8044 11249 8072
rect 11204 8032 11210 8044
rect 12529 8041 12541 8075
rect 12575 8072 12587 8075
rect 12894 8072 12900 8084
rect 12575 8044 12900 8072
rect 12575 8041 12587 8044
rect 12529 8035 12587 8041
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 8662 8004 8668 8016
rect 7024 7976 8668 8004
rect 4798 7945 4804 7948
rect 4792 7936 4804 7945
rect 4759 7908 4804 7936
rect 4792 7899 4804 7908
rect 4798 7896 4804 7899
rect 4856 7896 4862 7948
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7024 7877 7052 7976
rect 8662 7964 8668 7976
rect 8720 8004 8726 8016
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 8720 7976 8953 8004
rect 8720 7964 8726 7976
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 12802 8004 12808 8016
rect 12763 7976 12808 8004
rect 8941 7967 8999 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 7282 7945 7288 7948
rect 7276 7936 7288 7945
rect 7243 7908 7288 7936
rect 7276 7899 7288 7908
rect 7282 7896 7288 7899
rect 7340 7896 7346 7948
rect 11054 7936 11060 7948
rect 11015 7908 11060 7936
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6880 7840 7021 7868
rect 6880 7828 6886 7840
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 8352 7840 9689 7868
rect 8352 7828 8358 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 11330 7868 11336 7880
rect 11291 7840 11336 7868
rect 9677 7831 9735 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 5534 7692 5540 7744
rect 5592 7732 5598 7744
rect 5905 7735 5963 7741
rect 5905 7732 5917 7735
rect 5592 7704 5917 7732
rect 5592 7692 5598 7704
rect 5905 7701 5917 7704
rect 5951 7701 5963 7735
rect 6546 7732 6552 7744
rect 6507 7704 6552 7732
rect 5905 7695 5963 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7006 7732 7012 7744
rect 6963 7704 7012 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7006 7692 7012 7704
rect 7064 7732 7070 7744
rect 7650 7732 7656 7744
rect 7064 7704 7656 7732
rect 7064 7692 7070 7704
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 8389 7735 8447 7741
rect 8389 7732 8401 7735
rect 7708 7704 8401 7732
rect 7708 7692 7714 7704
rect 8389 7701 8401 7704
rect 8435 7701 8447 7735
rect 8389 7695 8447 7701
rect 1104 7642 14812 7664
rect 1104 7590 3648 7642
rect 3700 7590 3712 7642
rect 3764 7590 3776 7642
rect 3828 7590 3840 7642
rect 3892 7590 8982 7642
rect 9034 7590 9046 7642
rect 9098 7590 9110 7642
rect 9162 7590 9174 7642
rect 9226 7590 14315 7642
rect 14367 7590 14379 7642
rect 14431 7590 14443 7642
rect 14495 7590 14507 7642
rect 14559 7590 14812 7642
rect 1104 7568 14812 7590
rect 3142 7528 3148 7540
rect 3103 7500 3148 7528
rect 3142 7488 3148 7500
rect 3200 7488 3206 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7800 7500 8033 7528
rect 7800 7488 7806 7500
rect 8021 7497 8033 7500
rect 8067 7528 8079 7531
rect 10321 7531 10379 7537
rect 8067 7500 8708 7528
rect 8067 7497 8079 7500
rect 8021 7491 8079 7497
rect 8573 7463 8631 7469
rect 8573 7460 8585 7463
rect 7484 7432 8585 7460
rect 1762 7392 1768 7404
rect 1723 7364 1768 7392
rect 1762 7352 1768 7364
rect 1820 7352 1826 7404
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4798 7392 4804 7404
rect 4295 7364 4804 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4798 7352 4804 7364
rect 4856 7392 4862 7404
rect 5442 7392 5448 7404
rect 4856 7364 5448 7392
rect 4856 7352 4862 7364
rect 5442 7352 5448 7364
rect 5500 7392 5506 7404
rect 5629 7395 5687 7401
rect 5629 7392 5641 7395
rect 5500 7364 5641 7392
rect 5500 7352 5506 7364
rect 5629 7361 5641 7364
rect 5675 7361 5687 7395
rect 5629 7355 5687 7361
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 7484 7401 7512 7432
rect 8573 7429 8585 7432
rect 8619 7429 8631 7463
rect 8573 7423 8631 7429
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 6604 7364 7481 7392
rect 6604 7352 6610 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7650 7392 7656 7404
rect 7611 7364 7656 7392
rect 7469 7355 7527 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6972 7296 7389 7324
rect 6972 7284 6978 7296
rect 7377 7293 7389 7296
rect 7423 7324 7435 7327
rect 7834 7324 7840 7336
rect 7423 7296 7840 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 8680 7324 8708 7500
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 11054 7528 11060 7540
rect 10367 7500 11060 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 11054 7488 11060 7500
rect 11112 7528 11118 7540
rect 11701 7531 11759 7537
rect 11701 7528 11713 7531
rect 11112 7500 11713 7528
rect 11112 7488 11118 7500
rect 11701 7497 11713 7500
rect 11747 7497 11759 7531
rect 11701 7491 11759 7497
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 15746 7528 15752 7540
rect 14056 7500 15752 7528
rect 14056 7488 14062 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 10686 7420 10692 7472
rect 10744 7460 10750 7472
rect 11330 7460 11336 7472
rect 10744 7432 10916 7460
rect 11291 7432 11336 7460
rect 10744 7420 10750 7432
rect 9122 7392 9128 7404
rect 9083 7364 9128 7392
rect 9122 7352 9128 7364
rect 9180 7392 9186 7404
rect 9585 7395 9643 7401
rect 9585 7392 9597 7395
rect 9180 7364 9597 7392
rect 9180 7352 9186 7364
rect 9585 7361 9597 7364
rect 9631 7361 9643 7395
rect 10778 7392 10784 7404
rect 10739 7364 10784 7392
rect 9585 7355 9643 7361
rect 10778 7352 10784 7364
rect 10836 7352 10842 7404
rect 10888 7401 10916 7432
rect 11330 7420 11336 7432
rect 11388 7420 11394 7472
rect 10873 7395 10931 7401
rect 10873 7361 10885 7395
rect 10919 7361 10931 7395
rect 10873 7355 10931 7361
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 8680 7296 9045 7324
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 2010 7259 2068 7265
rect 2010 7256 2022 7259
rect 1596 7228 2022 7256
rect 1486 7148 1492 7200
rect 1544 7188 1550 7200
rect 1596 7197 1624 7228
rect 2010 7225 2022 7228
rect 2056 7225 2068 7259
rect 2010 7219 2068 7225
rect 4893 7259 4951 7265
rect 4893 7225 4905 7259
rect 4939 7256 4951 7259
rect 5258 7256 5264 7268
rect 4939 7228 5264 7256
rect 4939 7225 4951 7228
rect 4893 7219 4951 7225
rect 5258 7216 5264 7228
rect 5316 7256 5322 7268
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5316 7228 5549 7256
rect 5316 7216 5322 7228
rect 5537 7225 5549 7228
rect 5583 7225 5595 7259
rect 5537 7219 5595 7225
rect 6273 7259 6331 7265
rect 6273 7225 6285 7259
rect 6319 7256 6331 7259
rect 7282 7256 7288 7268
rect 6319 7228 7288 7256
rect 6319 7225 6331 7228
rect 6273 7219 6331 7225
rect 7282 7216 7288 7228
rect 7340 7216 7346 7268
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 1544 7160 1593 7188
rect 1544 7148 1550 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 1581 7151 1639 7157
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 4982 7148 4988 7200
rect 5040 7188 5046 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 5040 7160 5089 7188
rect 5040 7148 5046 7160
rect 5077 7157 5089 7160
rect 5123 7157 5135 7191
rect 5077 7151 5135 7157
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 5626 7188 5632 7200
rect 5491 7160 5632 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6549 7191 6607 7197
rect 6549 7188 6561 7191
rect 6144 7160 6561 7188
rect 6144 7148 6150 7160
rect 6549 7157 6561 7160
rect 6595 7188 6607 7191
rect 6822 7188 6828 7200
rect 6595 7160 6828 7188
rect 6595 7157 6607 7160
rect 6549 7151 6607 7157
rect 6822 7148 6828 7160
rect 6880 7148 6886 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7009 7191 7067 7197
rect 7009 7188 7021 7191
rect 6972 7160 7021 7188
rect 6972 7148 6978 7160
rect 7009 7157 7021 7160
rect 7055 7157 7067 7191
rect 7009 7151 7067 7157
rect 8481 7191 8539 7197
rect 8481 7157 8493 7191
rect 8527 7188 8539 7191
rect 8938 7188 8944 7200
rect 8527 7160 8944 7188
rect 8527 7157 8539 7160
rect 8481 7151 8539 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 10226 7188 10232 7200
rect 10139 7160 10232 7188
rect 10226 7148 10232 7160
rect 10284 7188 10290 7200
rect 10689 7191 10747 7197
rect 10689 7188 10701 7191
rect 10284 7160 10701 7188
rect 10284 7148 10290 7160
rect 10689 7157 10701 7160
rect 10735 7188 10747 7191
rect 11974 7188 11980 7200
rect 10735 7160 11980 7188
rect 10735 7157 10747 7160
rect 10689 7151 10747 7157
rect 11974 7148 11980 7160
rect 12032 7148 12038 7200
rect 1104 7098 14812 7120
rect 1104 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 11648 7098
rect 11700 7046 11712 7098
rect 11764 7046 11776 7098
rect 11828 7046 11840 7098
rect 11892 7046 14812 7098
rect 1104 7024 14812 7046
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5258 6984 5264 6996
rect 5215 6956 5264 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5258 6944 5264 6956
rect 5316 6984 5322 6996
rect 5626 6984 5632 6996
rect 5316 6956 5632 6984
rect 5316 6944 5322 6956
rect 5626 6944 5632 6956
rect 5684 6944 5690 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7340 6956 7389 6984
rect 7340 6944 7346 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2314 6848 2320 6860
rect 1443 6820 2320 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2409 6851 2467 6857
rect 2409 6817 2421 6851
rect 2455 6848 2467 6851
rect 2498 6848 2504 6860
rect 2455 6820 2504 6848
rect 2455 6817 2467 6820
rect 2409 6811 2467 6817
rect 2498 6808 2504 6820
rect 2556 6848 2562 6860
rect 5718 6857 5724 6860
rect 2869 6851 2927 6857
rect 2869 6848 2881 6851
rect 2556 6820 2881 6848
rect 2556 6808 2562 6820
rect 2869 6817 2881 6820
rect 2915 6817 2927 6851
rect 2869 6811 2927 6817
rect 5712 6811 5724 6857
rect 5776 6848 5782 6860
rect 5776 6820 5812 6848
rect 5718 6808 5724 6811
rect 5776 6808 5782 6820
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 5132 6752 5457 6780
rect 5132 6740 5138 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 7392 6780 7420 6947
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7892 6956 7941 6984
rect 7892 6944 7898 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 8294 6984 8300 6996
rect 8255 6956 8300 6984
rect 7929 6947 7987 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8389 6987 8447 6993
rect 8389 6953 8401 6987
rect 8435 6984 8447 6987
rect 8478 6984 8484 6996
rect 8435 6956 8484 6984
rect 8435 6953 8447 6956
rect 8389 6947 8447 6953
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 10778 6984 10784 6996
rect 10739 6956 10784 6984
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11146 6984 11152 6996
rect 11107 6956 11152 6984
rect 11146 6944 11152 6956
rect 11204 6944 11210 6996
rect 8312 6916 8340 6944
rect 8220 6888 8340 6916
rect 10413 6919 10471 6925
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 8220 6848 8248 6888
rect 10413 6885 10425 6919
rect 10459 6916 10471 6919
rect 10686 6916 10692 6928
rect 10459 6888 10692 6916
rect 10459 6885 10471 6888
rect 10413 6879 10471 6885
rect 10686 6876 10692 6888
rect 10744 6876 10750 6928
rect 7883 6820 8248 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 9306 6848 9312 6860
rect 8904 6820 9312 6848
rect 8904 6808 8910 6820
rect 9306 6808 9312 6820
rect 9364 6848 9370 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9364 6820 9689 6848
rect 9364 6808 9370 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 12069 6851 12127 6857
rect 12069 6817 12081 6851
rect 12115 6848 12127 6851
rect 12158 6848 12164 6860
rect 12115 6820 12164 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 12336 6851 12394 6857
rect 12336 6817 12348 6851
rect 12382 6848 12394 6851
rect 12618 6848 12624 6860
rect 12382 6820 12624 6848
rect 12382 6817 12394 6820
rect 12336 6811 12394 6817
rect 12618 6808 12624 6820
rect 12676 6848 12682 6860
rect 13078 6848 13084 6860
rect 12676 6820 13084 6848
rect 12676 6808 12682 6820
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 8481 6783 8539 6789
rect 8481 6780 8493 6783
rect 7392 6752 8493 6780
rect 5445 6743 5503 6749
rect 8481 6749 8493 6752
rect 8527 6780 8539 6783
rect 9122 6780 9128 6792
rect 8527 6752 9128 6780
rect 8527 6749 8539 6752
rect 8481 6743 8539 6749
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9490 6780 9496 6792
rect 9180 6752 9496 6780
rect 9180 6740 9186 6752
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 2593 6715 2651 6721
rect 2593 6681 2605 6715
rect 2639 6712 2651 6715
rect 2682 6712 2688 6724
rect 2639 6684 2688 6712
rect 2639 6681 2651 6684
rect 2593 6675 2651 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 4617 6715 4675 6721
rect 4617 6681 4629 6715
rect 4663 6712 4675 6715
rect 4663 6684 5488 6712
rect 4663 6681 4675 6684
rect 4617 6675 4675 6681
rect 5460 6656 5488 6684
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 5500 6616 6837 6644
rect 5500 6604 5506 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 8904 6616 8953 6644
rect 8904 6604 8910 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9861 6647 9919 6653
rect 9861 6613 9873 6647
rect 9907 6644 9919 6647
rect 9950 6644 9956 6656
rect 9907 6616 9956 6644
rect 9907 6613 9919 6616
rect 9861 6607 9919 6613
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 13446 6644 13452 6656
rect 13407 6616 13452 6644
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 1104 6554 14812 6576
rect 1104 6502 3648 6554
rect 3700 6502 3712 6554
rect 3764 6502 3776 6554
rect 3828 6502 3840 6554
rect 3892 6502 8982 6554
rect 9034 6502 9046 6554
rect 9098 6502 9110 6554
rect 9162 6502 9174 6554
rect 9226 6502 14315 6554
rect 14367 6502 14379 6554
rect 14431 6502 14443 6554
rect 14495 6502 14507 6554
rect 14559 6502 14812 6554
rect 1104 6480 14812 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 3418 6440 3424 6452
rect 2087 6412 3424 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2056 6236 2084 6403
rect 3418 6400 3424 6412
rect 3476 6400 3482 6452
rect 5718 6400 5724 6452
rect 5776 6440 5782 6452
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 5776 6412 5917 6440
rect 5776 6400 5782 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 5905 6403 5963 6409
rect 7101 6443 7159 6449
rect 7101 6409 7113 6443
rect 7147 6440 7159 6443
rect 7466 6440 7472 6452
rect 7147 6412 7472 6440
rect 7147 6409 7159 6412
rect 7101 6403 7159 6409
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4522 6372 4528 6384
rect 4212 6344 4528 6372
rect 4212 6332 4218 6344
rect 4522 6332 4528 6344
rect 4580 6372 4586 6384
rect 5074 6372 5080 6384
rect 4580 6344 5080 6372
rect 4580 6332 4586 6344
rect 5074 6332 5080 6344
rect 5132 6372 5138 6384
rect 5537 6375 5595 6381
rect 5537 6372 5549 6375
rect 5132 6344 5549 6372
rect 5132 6332 5138 6344
rect 5537 6341 5549 6344
rect 5583 6372 5595 6375
rect 5626 6372 5632 6384
rect 5583 6344 5632 6372
rect 5583 6341 5595 6344
rect 5537 6335 5595 6341
rect 5626 6332 5632 6344
rect 5684 6372 5690 6384
rect 6086 6372 6092 6384
rect 5684 6344 6092 6372
rect 5684 6332 5690 6344
rect 6086 6332 6092 6344
rect 6144 6332 6150 6384
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4982 6304 4988 6316
rect 3743 6276 4988 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 4982 6264 4988 6276
rect 5040 6264 5046 6316
rect 5169 6307 5227 6313
rect 5169 6273 5181 6307
rect 5215 6304 5227 6307
rect 5442 6304 5448 6316
rect 5215 6276 5448 6304
rect 5215 6273 5227 6276
rect 5169 6267 5227 6273
rect 1443 6208 2084 6236
rect 2501 6239 2559 6245
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 4065 6239 4123 6245
rect 2547 6208 3096 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 3068 6112 3096 6208
rect 4065 6205 4077 6239
rect 4111 6236 4123 6239
rect 5184 6236 5212 6267
rect 5442 6264 5448 6276
rect 5500 6264 5506 6316
rect 7208 6245 7236 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 8478 6440 8484 6452
rect 7883 6412 8484 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 8478 6400 8484 6412
rect 8536 6400 8542 6452
rect 9306 6440 9312 6452
rect 9267 6412 9312 6440
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 12158 6440 12164 6452
rect 12119 6412 12164 6440
rect 12158 6400 12164 6412
rect 12216 6400 12222 6452
rect 12618 6440 12624 6452
rect 12579 6412 12624 6440
rect 12618 6400 12624 6412
rect 12676 6400 12682 6452
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8846 6304 8852 6316
rect 8536 6276 8852 6304
rect 8536 6264 8542 6276
rect 8846 6264 8852 6276
rect 8904 6304 8910 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 8904 6276 10425 6304
rect 8904 6264 8910 6276
rect 10413 6273 10425 6276
rect 10459 6304 10471 6307
rect 10873 6307 10931 6313
rect 10873 6304 10885 6307
rect 10459 6276 10885 6304
rect 10459 6273 10471 6276
rect 10413 6267 10471 6273
rect 10873 6273 10885 6276
rect 10919 6273 10931 6307
rect 10873 6267 10931 6273
rect 4111 6208 5212 6236
rect 7193 6239 7251 6245
rect 4111 6205 4123 6208
rect 4065 6199 4123 6205
rect 7193 6205 7205 6239
rect 7239 6205 7251 6239
rect 7193 6199 7251 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 9815 6208 10364 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 4893 6171 4951 6177
rect 4893 6168 4905 6171
rect 4479 6140 4905 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4893 6137 4905 6140
rect 4939 6168 4951 6171
rect 4982 6168 4988 6180
rect 4939 6140 4988 6168
rect 4939 6137 4951 6140
rect 4893 6131 4951 6137
rect 4982 6128 4988 6140
rect 5040 6128 5046 6180
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 7466 6168 7472 6180
rect 6052 6140 7472 6168
rect 6052 6128 6058 6140
rect 7466 6128 7472 6140
rect 7524 6128 7530 6180
rect 8018 6128 8024 6180
rect 8076 6168 8082 6180
rect 8205 6171 8263 6177
rect 8205 6168 8217 6171
rect 8076 6140 8217 6168
rect 8076 6128 8082 6140
rect 8205 6137 8217 6140
rect 8251 6168 8263 6171
rect 8251 6140 8800 6168
rect 8251 6137 8263 6140
rect 8205 6131 8263 6137
rect 1302 6060 1308 6112
rect 1360 6100 1366 6112
rect 1581 6103 1639 6109
rect 1581 6100 1593 6103
rect 1360 6072 1593 6100
rect 1360 6060 1366 6072
rect 1581 6069 1593 6072
rect 1627 6069 1639 6103
rect 2406 6100 2412 6112
rect 2367 6072 2412 6100
rect 1581 6063 1639 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3050 6100 3056 6112
rect 3011 6072 3056 6100
rect 3050 6060 3056 6072
rect 3108 6060 3114 6112
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 6641 6103 6699 6109
rect 6641 6069 6653 6103
rect 6687 6100 6699 6103
rect 6730 6100 6736 6112
rect 6687 6072 6736 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 7377 6103 7435 6109
rect 7377 6069 7389 6103
rect 7423 6100 7435 6103
rect 7650 6100 7656 6112
rect 7423 6072 7656 6100
rect 7423 6069 7435 6072
rect 7377 6063 7435 6069
rect 7650 6060 7656 6072
rect 7708 6060 7714 6112
rect 8294 6100 8300 6112
rect 8255 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 8662 6100 8668 6112
rect 8623 6072 8668 6100
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8772 6109 8800 6140
rect 9674 6128 9680 6180
rect 9732 6168 9738 6180
rect 10336 6177 10364 6208
rect 10229 6171 10287 6177
rect 10229 6168 10241 6171
rect 9732 6140 10241 6168
rect 9732 6128 9738 6140
rect 10229 6137 10241 6140
rect 10275 6137 10287 6171
rect 10229 6131 10287 6137
rect 10321 6171 10379 6177
rect 10321 6137 10333 6171
rect 10367 6168 10379 6171
rect 10502 6168 10508 6180
rect 10367 6140 10508 6168
rect 10367 6137 10379 6140
rect 10321 6131 10379 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 8757 6103 8815 6109
rect 8757 6069 8769 6103
rect 8803 6100 8815 6103
rect 8846 6100 8852 6112
rect 8803 6072 8852 6100
rect 8803 6069 8815 6072
rect 8757 6063 8815 6069
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 9858 6100 9864 6112
rect 9819 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10594 6100 10600 6112
rect 10192 6072 10600 6100
rect 10192 6060 10198 6072
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 1104 6010 14812 6032
rect 1104 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 11648 6010
rect 11700 5958 11712 6010
rect 11764 5958 11776 6010
rect 11828 5958 11840 6010
rect 11892 5958 14812 6010
rect 1104 5936 14812 5958
rect 4341 5899 4399 5905
rect 4341 5865 4353 5899
rect 4387 5896 4399 5899
rect 4522 5896 4528 5908
rect 4387 5868 4528 5896
rect 4387 5865 4399 5868
rect 4341 5859 4399 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 5718 5856 5724 5908
rect 5776 5896 5782 5908
rect 6638 5896 6644 5908
rect 5776 5868 6644 5896
rect 5776 5856 5782 5868
rect 6638 5856 6644 5868
rect 6696 5896 6702 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 6696 5868 7389 5896
rect 6696 5856 6702 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 7377 5859 7435 5865
rect 4801 5831 4859 5837
rect 4801 5797 4813 5831
rect 4847 5828 4859 5831
rect 4890 5828 4896 5840
rect 4847 5800 4896 5828
rect 4847 5797 4859 5800
rect 4801 5791 4859 5797
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6264 5831 6322 5837
rect 6264 5828 6276 5831
rect 6052 5800 6276 5828
rect 6052 5788 6058 5800
rect 6264 5797 6276 5800
rect 6310 5828 6322 5831
rect 7006 5828 7012 5840
rect 6310 5800 7012 5828
rect 6310 5797 6322 5800
rect 6264 5791 6322 5797
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 9674 5788 9680 5840
rect 9732 5828 9738 5840
rect 9861 5831 9919 5837
rect 9861 5828 9873 5831
rect 9732 5800 9873 5828
rect 9732 5788 9738 5800
rect 9861 5797 9873 5800
rect 9907 5797 9919 5831
rect 9861 5791 9919 5797
rect 12060 5831 12118 5837
rect 12060 5797 12072 5831
rect 12106 5828 12118 5831
rect 12342 5828 12348 5840
rect 12106 5800 12348 5828
rect 12106 5797 12118 5800
rect 12060 5791 12118 5797
rect 1394 5760 1400 5772
rect 1355 5732 1400 5760
rect 1394 5720 1400 5732
rect 1452 5720 1458 5772
rect 2866 5760 2872 5772
rect 2779 5732 2872 5760
rect 2866 5720 2872 5732
rect 2924 5760 2930 5772
rect 5258 5760 5264 5772
rect 2924 5732 5264 5760
rect 2924 5720 2930 5732
rect 5258 5720 5264 5732
rect 5316 5720 5322 5772
rect 7929 5763 7987 5769
rect 7929 5760 7941 5763
rect 6012 5732 7941 5760
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 4982 5692 4988 5704
rect 4939 5664 4988 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5692 5135 5695
rect 5442 5692 5448 5704
rect 5123 5664 5448 5692
rect 5123 5661 5135 5664
rect 5077 5655 5135 5661
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5626 5652 5632 5704
rect 5684 5692 5690 5704
rect 6012 5701 6040 5732
rect 7929 5729 7941 5732
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 5684 5664 6009 5692
rect 5684 5652 5690 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 7944 5692 7972 5723
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 8481 5763 8539 5769
rect 8481 5760 8493 5763
rect 8076 5732 8493 5760
rect 8076 5720 8082 5732
rect 8481 5729 8493 5732
rect 8527 5760 8539 5763
rect 8570 5760 8576 5772
rect 8527 5732 8576 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 9493 5763 9551 5769
rect 9493 5729 9505 5763
rect 9539 5760 9551 5763
rect 10594 5760 10600 5772
rect 9539 5732 10600 5760
rect 9539 5729 9551 5732
rect 9493 5723 9551 5729
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 11330 5760 11336 5772
rect 11243 5732 11336 5760
rect 11330 5720 11336 5732
rect 11388 5760 11394 5772
rect 12084 5760 12112 5791
rect 12342 5788 12348 5800
rect 12400 5828 12406 5840
rect 13446 5828 13452 5840
rect 12400 5800 13452 5828
rect 12400 5788 12406 5800
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 11388 5732 12112 5760
rect 11388 5720 11394 5732
rect 8110 5692 8116 5704
rect 7944 5664 8116 5692
rect 5997 5655 6055 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 10686 5692 10692 5704
rect 10647 5664 10692 5692
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 10778 5652 10784 5704
rect 10836 5692 10842 5704
rect 11793 5695 11851 5701
rect 10836 5664 10881 5692
rect 10836 5652 10842 5664
rect 11793 5661 11805 5695
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 7374 5584 7380 5636
rect 7432 5624 7438 5636
rect 8665 5627 8723 5633
rect 8665 5624 8677 5627
rect 7432 5596 8677 5624
rect 7432 5584 7438 5596
rect 8665 5593 8677 5596
rect 8711 5593 8723 5627
rect 8665 5587 8723 5593
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10229 5627 10287 5633
rect 10229 5624 10241 5627
rect 9732 5596 10241 5624
rect 9732 5584 9738 5596
rect 10229 5593 10241 5596
rect 10275 5593 10287 5627
rect 10229 5587 10287 5593
rect 11808 5568 11836 5655
rect 934 5516 940 5568
rect 992 5556 998 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 992 5528 1593 5556
rect 992 5516 998 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 2682 5556 2688 5568
rect 2547 5528 2688 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 3418 5556 3424 5568
rect 3379 5528 3424 5556
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 3881 5559 3939 5565
rect 3881 5525 3893 5559
rect 3927 5556 3939 5559
rect 3970 5556 3976 5568
rect 3927 5528 3976 5556
rect 3927 5525 3939 5528
rect 3881 5519 3939 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4430 5556 4436 5568
rect 4391 5528 4436 5556
rect 4430 5516 4436 5528
rect 4488 5516 4494 5568
rect 5534 5556 5540 5568
rect 5495 5528 5540 5556
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 7098 5556 7104 5568
rect 5951 5528 7104 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7650 5516 7656 5568
rect 7708 5556 7714 5568
rect 8297 5559 8355 5565
rect 8297 5556 8309 5559
rect 7708 5528 8309 5556
rect 7708 5516 7714 5528
rect 8297 5525 8309 5528
rect 8343 5556 8355 5559
rect 8570 5556 8576 5568
rect 8343 5528 8576 5556
rect 8343 5525 8355 5528
rect 8297 5519 8355 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 11790 5556 11796 5568
rect 11703 5528 11796 5556
rect 11790 5516 11796 5528
rect 11848 5556 11854 5568
rect 12158 5556 12164 5568
rect 11848 5528 12164 5556
rect 11848 5516 11854 5528
rect 12158 5516 12164 5528
rect 12216 5516 12222 5568
rect 13170 5556 13176 5568
rect 13131 5528 13176 5556
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 1104 5466 14812 5488
rect 1104 5414 3648 5466
rect 3700 5414 3712 5466
rect 3764 5414 3776 5466
rect 3828 5414 3840 5466
rect 3892 5414 8982 5466
rect 9034 5414 9046 5466
rect 9098 5414 9110 5466
rect 9162 5414 9174 5466
rect 9226 5414 14315 5466
rect 14367 5414 14379 5466
rect 14431 5414 14443 5466
rect 14495 5414 14507 5466
rect 14559 5414 14812 5466
rect 1104 5392 14812 5414
rect 1394 5312 1400 5364
rect 1452 5352 1458 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1452 5324 1593 5352
rect 1452 5312 1458 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 1581 5315 1639 5321
rect 1596 5284 1624 5315
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 4341 5355 4399 5361
rect 2976 5324 4292 5352
rect 2976 5284 3004 5324
rect 1596 5256 3004 5284
rect 4264 5284 4292 5324
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4706 5352 4712 5364
rect 4387 5324 4712 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6549 5355 6607 5361
rect 6549 5352 6561 5355
rect 5684 5324 6561 5352
rect 5684 5312 5690 5324
rect 6549 5321 6561 5324
rect 6595 5321 6607 5355
rect 6549 5315 6607 5321
rect 7190 5312 7196 5364
rect 7248 5352 7254 5364
rect 7377 5355 7435 5361
rect 7377 5352 7389 5355
rect 7248 5324 7389 5352
rect 7248 5312 7254 5324
rect 7377 5321 7389 5324
rect 7423 5321 7435 5355
rect 8018 5352 8024 5364
rect 7979 5324 8024 5352
rect 7377 5315 7435 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 9490 5352 9496 5364
rect 9451 5324 9496 5352
rect 9490 5312 9496 5324
rect 9548 5312 9554 5364
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10652 5324 10793 5352
rect 10652 5312 10658 5324
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 10781 5315 10839 5321
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11790 5352 11796 5364
rect 11204 5324 11796 5352
rect 11204 5312 11210 5324
rect 11790 5312 11796 5324
rect 11848 5312 11854 5364
rect 12253 5355 12311 5361
rect 12253 5321 12265 5355
rect 12299 5352 12311 5355
rect 12342 5352 12348 5364
rect 12299 5324 12348 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 7650 5284 7656 5296
rect 4264 5256 7656 5284
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 10689 5287 10747 5293
rect 10689 5253 10701 5287
rect 10735 5284 10747 5287
rect 10870 5284 10876 5296
rect 10735 5256 10876 5284
rect 10735 5253 10747 5256
rect 10689 5247 10747 5253
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 8110 5216 8116 5228
rect 8071 5188 8116 5216
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 11330 5216 11336 5228
rect 11291 5188 11336 5216
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 1765 5151 1823 5157
rect 1765 5117 1777 5151
rect 1811 5117 1823 5151
rect 1765 5111 1823 5117
rect 2961 5151 3019 5157
rect 2961 5117 2973 5151
rect 3007 5148 3019 5151
rect 3510 5148 3516 5160
rect 3007 5120 3516 5148
rect 3007 5117 3019 5120
rect 2961 5111 3019 5117
rect 1780 5080 1808 5111
rect 3510 5108 3516 5120
rect 3568 5148 3574 5160
rect 4154 5148 4160 5160
rect 3568 5120 4160 5148
rect 3568 5108 3574 5120
rect 4154 5108 4160 5120
rect 4212 5108 4218 5160
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5629 5151 5687 5157
rect 5629 5148 5641 5151
rect 5408 5120 5641 5148
rect 5408 5108 5414 5120
rect 5629 5117 5641 5120
rect 5675 5148 5687 5151
rect 6181 5151 6239 5157
rect 6181 5148 6193 5151
rect 5675 5120 6193 5148
rect 5675 5117 5687 5120
rect 5629 5111 5687 5117
rect 6181 5117 6193 5120
rect 6227 5117 6239 5151
rect 6181 5111 6239 5117
rect 6825 5151 6883 5157
rect 6825 5117 6837 5151
rect 6871 5148 6883 5151
rect 7190 5148 7196 5160
rect 6871 5120 7196 5148
rect 6871 5117 6883 5120
rect 6825 5111 6883 5117
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 10318 5148 10324 5160
rect 10231 5120 10324 5148
rect 10318 5108 10324 5120
rect 10376 5148 10382 5160
rect 11149 5151 11207 5157
rect 11149 5148 11161 5151
rect 10376 5120 11161 5148
rect 10376 5108 10382 5120
rect 11149 5117 11161 5120
rect 11195 5148 11207 5151
rect 11422 5148 11428 5160
rect 11195 5120 11428 5148
rect 11195 5117 11207 5120
rect 11149 5111 11207 5117
rect 11422 5108 11428 5120
rect 11480 5108 11486 5160
rect 2406 5080 2412 5092
rect 1780 5052 2412 5080
rect 2406 5040 2412 5052
rect 2464 5040 2470 5092
rect 3206 5083 3264 5089
rect 3206 5080 3218 5083
rect 2976 5052 3218 5080
rect 2976 5024 3004 5052
rect 3206 5049 3218 5052
rect 3252 5080 3264 5083
rect 3418 5080 3424 5092
rect 3252 5052 3424 5080
rect 3252 5049 3264 5052
rect 3206 5043 3264 5049
rect 3418 5040 3424 5052
rect 3476 5040 3482 5092
rect 8386 5089 8392 5092
rect 8380 5080 8392 5089
rect 8347 5052 8392 5080
rect 8380 5043 8392 5052
rect 8386 5040 8392 5043
rect 8444 5040 8450 5092
rect 9306 5040 9312 5092
rect 9364 5080 9370 5092
rect 10870 5080 10876 5092
rect 9364 5052 10876 5080
rect 9364 5040 9370 5052
rect 10870 5040 10876 5052
rect 10928 5080 10934 5092
rect 11241 5083 11299 5089
rect 11241 5080 11253 5083
rect 10928 5052 11253 5080
rect 10928 5040 10934 5052
rect 11241 5049 11253 5052
rect 11287 5049 11299 5083
rect 11241 5043 11299 5049
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1949 5015 2007 5021
rect 1949 5012 1961 5015
rect 1452 4984 1961 5012
rect 1452 4972 1458 4984
rect 1949 4981 1961 4984
rect 1995 4981 2007 5015
rect 1949 4975 2007 4981
rect 2958 4972 2964 5024
rect 3016 4972 3022 5024
rect 4890 5012 4896 5024
rect 4851 4984 4896 5012
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 4982 4972 4988 5024
rect 5040 5012 5046 5024
rect 5350 5012 5356 5024
rect 5040 4984 5356 5012
rect 5040 4972 5046 4984
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 6086 5012 6092 5024
rect 5859 4984 6092 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 7006 5012 7012 5024
rect 6967 4984 7012 5012
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 12986 5012 12992 5024
rect 12483 4984 12992 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 1104 4922 14812 4944
rect 1104 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 11648 4922
rect 11700 4870 11712 4922
rect 11764 4870 11776 4922
rect 11828 4870 11840 4922
rect 11892 4870 14812 4922
rect 1104 4848 14812 4870
rect 2409 4811 2467 4817
rect 2409 4777 2421 4811
rect 2455 4808 2467 4811
rect 2498 4808 2504 4820
rect 2455 4780 2504 4808
rect 2455 4777 2467 4780
rect 2409 4771 2467 4777
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2774 4808 2780 4820
rect 2740 4780 2780 4808
rect 2740 4768 2746 4780
rect 2774 4768 2780 4780
rect 2832 4768 2838 4820
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 4065 4811 4123 4817
rect 4065 4808 4077 4811
rect 2924 4780 4077 4808
rect 2924 4768 2930 4780
rect 4065 4777 4077 4780
rect 4111 4777 4123 4811
rect 4522 4808 4528 4820
rect 4483 4780 4528 4808
rect 4065 4771 4123 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4856 4780 5181 4808
rect 4856 4768 4862 4780
rect 5169 4777 5181 4780
rect 5215 4808 5227 4811
rect 5442 4808 5448 4820
rect 5215 4780 5448 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 5592 4780 6561 4808
rect 5592 4768 5598 4780
rect 6549 4777 6561 4780
rect 6595 4808 6607 4811
rect 6822 4808 6828 4820
rect 6595 4780 6828 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6822 4768 6828 4780
rect 6880 4768 6886 4820
rect 7193 4811 7251 4817
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 8202 4808 8208 4820
rect 7239 4780 8208 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 8202 4768 8208 4780
rect 8260 4768 8266 4820
rect 8389 4811 8447 4817
rect 8389 4777 8401 4811
rect 8435 4808 8447 4811
rect 8754 4808 8760 4820
rect 8435 4780 8760 4808
rect 8435 4777 8447 4780
rect 8389 4771 8447 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9493 4811 9551 4817
rect 9493 4777 9505 4811
rect 9539 4808 9551 4811
rect 10597 4811 10655 4817
rect 10597 4808 10609 4811
rect 9539 4780 10609 4808
rect 9539 4777 9551 4780
rect 9493 4771 9551 4777
rect 10597 4777 10609 4780
rect 10643 4808 10655 4811
rect 10686 4808 10692 4820
rect 10643 4780 10692 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 12526 4808 12532 4820
rect 12439 4780 12532 4808
rect 12526 4768 12532 4780
rect 12584 4808 12590 4820
rect 12710 4808 12716 4820
rect 12584 4780 12716 4808
rect 12584 4768 12590 4780
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 2317 4743 2375 4749
rect 2317 4709 2329 4743
rect 2363 4740 2375 4743
rect 4430 4740 4436 4752
rect 2363 4712 4436 4740
rect 2363 4709 2375 4712
rect 2317 4703 2375 4709
rect 4430 4700 4436 4712
rect 4488 4700 4494 4752
rect 5994 4740 6000 4752
rect 5955 4712 6000 4740
rect 5994 4700 6000 4712
rect 6052 4700 6058 4752
rect 6457 4743 6515 4749
rect 6457 4709 6469 4743
rect 6503 4740 6515 4743
rect 6914 4740 6920 4752
rect 6503 4712 6920 4740
rect 6503 4709 6515 4712
rect 6457 4703 6515 4709
rect 2774 4632 2780 4684
rect 2832 4672 2838 4684
rect 4062 4672 4068 4684
rect 2832 4644 4068 4672
rect 2832 4632 2838 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 6472 4672 6500 4703
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 9125 4743 9183 4749
rect 9125 4709 9137 4743
rect 9171 4740 9183 4743
rect 9582 4740 9588 4752
rect 9171 4712 9588 4740
rect 9171 4709 9183 4712
rect 9125 4703 9183 4709
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 10505 4743 10563 4749
rect 10505 4709 10517 4743
rect 10551 4740 10563 4743
rect 10778 4740 10784 4752
rect 10551 4712 10784 4740
rect 10551 4709 10563 4712
rect 10505 4703 10563 4709
rect 10778 4700 10784 4712
rect 10836 4740 10842 4752
rect 13170 4740 13176 4752
rect 10836 4712 13176 4740
rect 10836 4700 10842 4712
rect 4264 4644 6500 4672
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 1670 4604 1676 4616
rect 1443 4576 1676 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 1946 4604 1952 4616
rect 1907 4576 1952 4604
rect 1946 4564 1952 4576
rect 2004 4564 2010 4616
rect 2958 4604 2964 4616
rect 2919 4576 2964 4604
rect 2958 4564 2964 4576
rect 3016 4564 3022 4616
rect 3881 4607 3939 4613
rect 3881 4573 3893 4607
rect 3927 4604 3939 4607
rect 4264 4604 4292 4644
rect 8018 4632 8024 4684
rect 8076 4672 8082 4684
rect 8481 4675 8539 4681
rect 8481 4672 8493 4675
rect 8076 4644 8493 4672
rect 8076 4632 8082 4644
rect 8481 4641 8493 4644
rect 8527 4672 8539 4675
rect 9490 4672 9496 4684
rect 8527 4644 9496 4672
rect 8527 4641 8539 4644
rect 8481 4635 8539 4641
rect 9490 4632 9496 4644
rect 9548 4632 9554 4684
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10284 4644 10977 4672
rect 10284 4632 10290 4644
rect 10965 4641 10977 4644
rect 11011 4672 11023 4675
rect 11238 4672 11244 4684
rect 11011 4644 11244 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 3927 4576 4292 4604
rect 4709 4607 4767 4613
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 6638 4604 6644 4616
rect 4755 4576 5580 4604
rect 6599 4576 6644 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 2774 4428 2780 4480
rect 2832 4468 2838 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2832 4440 3433 4468
rect 2832 4428 2838 4440
rect 3421 4437 3433 4440
rect 3467 4468 3479 4471
rect 3510 4468 3516 4480
rect 3467 4440 3516 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 5552 4477 5580 4576
rect 6638 4564 6644 4576
rect 6696 4564 6702 4616
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9674 4604 9680 4616
rect 8711 4576 9680 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 5810 4496 5816 4548
rect 5868 4536 5874 4548
rect 6089 4539 6147 4545
rect 6089 4536 6101 4539
rect 5868 4508 6101 4536
rect 5868 4496 5874 4508
rect 6089 4505 6101 4508
rect 6135 4505 6147 4539
rect 6089 4499 6147 4505
rect 7561 4539 7619 4545
rect 7561 4505 7573 4539
rect 7607 4536 7619 4539
rect 7929 4539 7987 4545
rect 7929 4536 7941 4539
rect 7607 4508 7941 4536
rect 7607 4505 7619 4508
rect 7561 4499 7619 4505
rect 7929 4505 7941 4508
rect 7975 4536 7987 4539
rect 8386 4536 8392 4548
rect 7975 4508 8392 4536
rect 7975 4505 7987 4508
rect 7929 4499 7987 4505
rect 8386 4496 8392 4508
rect 8444 4536 8450 4548
rect 8680 4536 8708 4567
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 10410 4564 10416 4616
rect 10468 4604 10474 4616
rect 10870 4604 10876 4616
rect 10468 4576 10876 4604
rect 10468 4564 10474 4576
rect 10870 4564 10876 4576
rect 10928 4604 10934 4616
rect 11057 4607 11115 4613
rect 11057 4604 11069 4607
rect 10928 4576 11069 4604
rect 10928 4564 10934 4576
rect 11057 4573 11069 4576
rect 11103 4573 11115 4607
rect 11057 4567 11115 4573
rect 11149 4607 11207 4613
rect 11149 4573 11161 4607
rect 11195 4604 11207 4607
rect 11330 4604 11336 4616
rect 11195 4576 11336 4604
rect 11195 4573 11207 4576
rect 11149 4567 11207 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 12618 4604 12624 4616
rect 12579 4576 12624 4604
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12728 4613 12756 4712
rect 13170 4700 13176 4712
rect 13228 4700 13234 4752
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 8444 4508 8708 4536
rect 8444 4496 8450 4508
rect 5537 4471 5595 4477
rect 5537 4437 5549 4471
rect 5583 4468 5595 4471
rect 5626 4468 5632 4480
rect 5583 4440 5632 4468
rect 5583 4437 5595 4440
rect 5537 4431 5595 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8110 4468 8116 4480
rect 8067 4440 8116 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 10226 4468 10232 4480
rect 10183 4440 10232 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 12158 4468 12164 4480
rect 12119 4440 12164 4468
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 13170 4468 13176 4480
rect 13131 4440 13176 4468
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 1104 4378 14812 4400
rect 1104 4326 3648 4378
rect 3700 4326 3712 4378
rect 3764 4326 3776 4378
rect 3828 4326 3840 4378
rect 3892 4326 8982 4378
rect 9034 4326 9046 4378
rect 9098 4326 9110 4378
rect 9162 4326 9174 4378
rect 9226 4326 14315 4378
rect 14367 4326 14379 4378
rect 14431 4326 14443 4378
rect 14495 4326 14507 4378
rect 14559 4326 14812 4378
rect 1104 4304 14812 4326
rect 2130 4264 2136 4276
rect 2091 4236 2136 4264
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3973 4267 4031 4273
rect 3973 4264 3985 4267
rect 3016 4236 3985 4264
rect 3016 4224 3022 4236
rect 3973 4233 3985 4236
rect 4019 4233 4031 4267
rect 4798 4264 4804 4276
rect 4759 4236 4804 4264
rect 3973 4227 4031 4233
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 6181 4267 6239 4273
rect 6181 4233 6193 4267
rect 6227 4264 6239 4267
rect 6638 4264 6644 4276
rect 6227 4236 6644 4264
rect 6227 4233 6239 4236
rect 6181 4227 6239 4233
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 6822 4264 6828 4276
rect 6783 4236 6828 4264
rect 6822 4224 6828 4236
rect 6880 4224 6886 4276
rect 8018 4264 8024 4276
rect 7979 4236 8024 4264
rect 8018 4224 8024 4236
rect 8076 4264 8082 4276
rect 8386 4264 8392 4276
rect 8076 4236 8392 4264
rect 8076 4224 8082 4236
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 11057 4267 11115 4273
rect 11057 4264 11069 4267
rect 10928 4236 11069 4264
rect 10928 4224 10934 4236
rect 11057 4233 11069 4236
rect 11103 4233 11115 4267
rect 11057 4227 11115 4233
rect 12253 4267 12311 4273
rect 12253 4233 12265 4267
rect 12299 4264 12311 4267
rect 12526 4264 12532 4276
rect 12299 4236 12532 4264
rect 12299 4233 12311 4236
rect 12253 4227 12311 4233
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 13817 4267 13875 4273
rect 13817 4264 13829 4267
rect 12676 4236 13829 4264
rect 12676 4224 12682 4236
rect 13817 4233 13829 4236
rect 13863 4233 13875 4267
rect 13817 4227 13875 4233
rect 4080 4168 5672 4196
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 1302 4128 1308 4140
rect 256 4100 1308 4128
rect 256 4088 262 4100
rect 1302 4088 1308 4100
rect 1360 4088 1366 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 4080 4128 4108 4168
rect 5644 4140 5672 4168
rect 5994 4156 6000 4208
rect 6052 4196 6058 4208
rect 6546 4196 6552 4208
rect 6052 4168 6552 4196
rect 6052 4156 6058 4168
rect 6546 4156 6552 4168
rect 6604 4156 6610 4208
rect 7006 4196 7012 4208
rect 6840 4168 7012 4196
rect 5626 4128 5632 4140
rect 3936 4100 4108 4128
rect 5587 4100 5632 4128
rect 3936 4088 3942 4100
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 6840 4128 6868 4168
rect 7006 4156 7012 4168
rect 7064 4156 7070 4208
rect 5776 4100 6868 4128
rect 5776 4088 5782 4100
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6972 4100 7297 4128
rect 6972 4088 6978 4100
rect 7285 4097 7297 4100
rect 7331 4097 7343 4131
rect 7285 4091 7343 4097
rect 7377 4131 7435 4137
rect 7377 4097 7389 4131
rect 7423 4097 7435 4131
rect 9122 4128 9128 4140
rect 9083 4100 9128 4128
rect 7377 4091 7435 4097
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 2130 4060 2136 4072
rect 1535 4032 2136 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 2130 4020 2136 4032
rect 2188 4020 2194 4072
rect 2501 4063 2559 4069
rect 2501 4029 2513 4063
rect 2547 4060 2559 4063
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 2547 4032 2605 4060
rect 2547 4029 2559 4032
rect 2501 4023 2559 4029
rect 2593 4029 2605 4032
rect 2639 4060 2651 4063
rect 2682 4060 2688 4072
rect 2639 4032 2688 4060
rect 2639 4029 2651 4032
rect 2593 4023 2651 4029
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2860 4063 2918 4069
rect 2860 4029 2872 4063
rect 2906 4060 2918 4063
rect 3896 4060 3924 4088
rect 5442 4060 5448 4072
rect 2906 4032 3924 4060
rect 5403 4032 5448 4060
rect 2906 4029 2918 4032
rect 2860 4023 2918 4029
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7193 4063 7251 4069
rect 7193 4060 7205 4063
rect 7156 4032 7205 4060
rect 7156 4020 7162 4032
rect 7193 4029 7205 4032
rect 7239 4029 7251 4063
rect 7193 4023 7251 4029
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 4212 3964 5120 3992
rect 4212 3952 4218 3964
rect 1673 3927 1731 3933
rect 1673 3893 1685 3927
rect 1719 3924 1731 3927
rect 2590 3924 2596 3936
rect 1719 3896 2596 3924
rect 1719 3893 1731 3896
rect 1673 3887 1731 3893
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 5092 3933 5120 3964
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5537 3995 5595 4001
rect 5537 3992 5549 3995
rect 5408 3964 5549 3992
rect 5408 3952 5414 3964
rect 5537 3961 5549 3964
rect 5583 3961 5595 3995
rect 5537 3955 5595 3961
rect 6546 3952 6552 4004
rect 6604 3992 6610 4004
rect 7392 3992 7420 4091
rect 9122 4088 9128 4100
rect 9180 4088 9186 4140
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4128 9551 4131
rect 10594 4128 10600 4140
rect 9539 4100 10600 4128
rect 9539 4097 9551 4100
rect 9493 4091 9551 4097
rect 10594 4088 10600 4100
rect 10652 4128 10658 4140
rect 10689 4131 10747 4137
rect 10689 4128 10701 4131
rect 10652 4100 10701 4128
rect 10652 4088 10658 4100
rect 10689 4097 10701 4100
rect 10735 4128 10747 4131
rect 11330 4128 11336 4140
rect 10735 4100 11336 4128
rect 10735 4097 10747 4100
rect 10689 4091 10747 4097
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 13081 4131 13139 4137
rect 13081 4128 13093 4131
rect 12768 4100 13093 4128
rect 12768 4088 12774 4100
rect 13081 4097 13093 4100
rect 13127 4128 13139 4131
rect 13449 4131 13507 4137
rect 13449 4128 13461 4131
rect 13127 4100 13461 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13449 4097 13461 4100
rect 13495 4097 13507 4131
rect 13449 4091 13507 4097
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4060 8999 4063
rect 9582 4060 9588 4072
rect 8987 4032 9588 4060
rect 8987 4029 8999 4032
rect 8941 4023 8999 4029
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10134 4060 10140 4072
rect 9999 4032 10140 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10134 4020 10140 4032
rect 10192 4060 10198 4072
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 10192 4032 10517 4060
rect 10192 4020 10198 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11425 4063 11483 4069
rect 11425 4060 11437 4063
rect 11296 4032 11437 4060
rect 11296 4020 11302 4032
rect 11425 4029 11437 4032
rect 11471 4029 11483 4063
rect 11425 4023 11483 4029
rect 12618 4020 12624 4072
rect 12676 4060 12682 4072
rect 12805 4063 12863 4069
rect 12805 4060 12817 4063
rect 12676 4032 12817 4060
rect 12676 4020 12682 4032
rect 12805 4029 12817 4032
rect 12851 4060 12863 4063
rect 13170 4060 13176 4072
rect 12851 4032 13176 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 6604 3964 7420 3992
rect 6604 3952 6610 3964
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 10376 3964 12480 3992
rect 10376 3952 10382 3964
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8570 3924 8576 3936
rect 8527 3896 8576 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9398 3924 9404 3936
rect 8895 3896 9404 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9398 3884 9404 3896
rect 9456 3884 9462 3936
rect 10042 3924 10048 3936
rect 10003 3896 10048 3924
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10226 3884 10232 3936
rect 10284 3924 10290 3936
rect 10413 3927 10471 3933
rect 10413 3924 10425 3927
rect 10284 3896 10425 3924
rect 10284 3884 10290 3896
rect 10413 3893 10425 3896
rect 10459 3893 10471 3927
rect 10413 3887 10471 3893
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 12452 3933 12480 3964
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11296 3896 11805 3924
rect 11296 3884 11302 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3893 12495 3927
rect 12437 3887 12495 3893
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13078 3924 13084 3936
rect 12943 3896 13084 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13078 3884 13084 3896
rect 13136 3884 13142 3936
rect 1104 3834 14812 3856
rect 1104 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 11648 3834
rect 11700 3782 11712 3834
rect 11764 3782 11776 3834
rect 11828 3782 11840 3834
rect 11892 3782 14812 3834
rect 1104 3760 14812 3782
rect 1673 3723 1731 3729
rect 1673 3689 1685 3723
rect 1719 3720 1731 3723
rect 2866 3720 2872 3732
rect 1719 3692 2872 3720
rect 1719 3689 1731 3692
rect 1673 3683 1731 3689
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3513 3723 3571 3729
rect 3513 3689 3525 3723
rect 3559 3720 3571 3723
rect 3878 3720 3884 3732
rect 3559 3692 3884 3720
rect 3559 3689 3571 3692
rect 3513 3683 3571 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4709 3723 4767 3729
rect 4709 3720 4721 3723
rect 4212 3692 4721 3720
rect 4212 3680 4218 3692
rect 4709 3689 4721 3692
rect 4755 3720 4767 3723
rect 5350 3720 5356 3732
rect 4755 3692 5356 3720
rect 4755 3689 4767 3692
rect 4709 3683 4767 3689
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 6914 3680 6920 3732
rect 6972 3720 6978 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 6972 3692 7665 3720
rect 6972 3680 6978 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 8021 3723 8079 3729
rect 8021 3689 8033 3723
rect 8067 3720 8079 3723
rect 8202 3720 8208 3732
rect 8067 3692 8208 3720
rect 8067 3689 8079 3692
rect 8021 3683 8079 3689
rect 8202 3680 8208 3692
rect 8260 3680 8266 3732
rect 8754 3720 8760 3732
rect 8715 3692 8760 3720
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 9490 3720 9496 3732
rect 9451 3692 9496 3720
rect 9490 3680 9496 3692
rect 9548 3680 9554 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 10318 3720 10324 3732
rect 9640 3692 10324 3720
rect 9640 3680 9646 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10594 3720 10600 3732
rect 10555 3692 10600 3720
rect 10594 3680 10600 3692
rect 10652 3680 10658 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10836 3692 10977 3720
rect 10836 3680 10842 3692
rect 10965 3689 10977 3692
rect 11011 3720 11023 3723
rect 11238 3720 11244 3732
rect 11011 3692 11244 3720
rect 11011 3689 11023 3692
rect 10965 3683 11023 3689
rect 11238 3680 11244 3692
rect 11296 3680 11302 3732
rect 2501 3655 2559 3661
rect 2501 3621 2513 3655
rect 2547 3652 2559 3655
rect 2958 3652 2964 3664
rect 2547 3624 2964 3652
rect 2547 3621 2559 3624
rect 2501 3615 2559 3621
rect 2958 3612 2964 3624
rect 3016 3612 3022 3664
rect 4338 3612 4344 3664
rect 4396 3652 4402 3664
rect 4617 3655 4675 3661
rect 4617 3652 4629 3655
rect 4396 3624 4629 3652
rect 4396 3612 4402 3624
rect 4617 3621 4629 3624
rect 4663 3652 4675 3655
rect 5166 3652 5172 3664
rect 4663 3624 5172 3652
rect 4663 3621 4675 3624
rect 4617 3615 4675 3621
rect 5166 3612 5172 3624
rect 5224 3612 5230 3664
rect 6181 3655 6239 3661
rect 6181 3621 6193 3655
rect 6227 3652 6239 3655
rect 8110 3652 8116 3664
rect 6227 3624 8116 3652
rect 6227 3621 6239 3624
rect 6181 3615 6239 3621
rect 8110 3612 8116 3624
rect 8168 3612 8174 3664
rect 9122 3652 9128 3664
rect 9035 3624 9128 3652
rect 9122 3612 9128 3624
rect 9180 3652 9186 3664
rect 9398 3652 9404 3664
rect 9180 3624 9404 3652
rect 9180 3612 9186 3624
rect 9398 3612 9404 3624
rect 9456 3652 9462 3664
rect 12710 3652 12716 3664
rect 9456 3624 12716 3652
rect 9456 3612 9462 3624
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 1762 3584 1768 3596
rect 1723 3556 1768 3584
rect 1762 3544 1768 3556
rect 1820 3544 1826 3596
rect 2866 3584 2872 3596
rect 2827 3556 2872 3584
rect 2866 3544 2872 3556
rect 2924 3544 2930 3596
rect 5074 3584 5080 3596
rect 4264 3556 5080 3584
rect 4264 3528 4292 3556
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 6273 3587 6331 3593
rect 6273 3553 6285 3587
rect 6319 3584 6331 3587
rect 6638 3584 6644 3596
rect 6319 3556 6644 3584
rect 6319 3553 6331 3556
rect 6273 3547 6331 3553
rect 6638 3544 6644 3556
rect 6696 3544 6702 3596
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 7282 3584 7288 3596
rect 6963 3556 7288 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 7282 3544 7288 3556
rect 7340 3584 7346 3596
rect 8018 3584 8024 3596
rect 7340 3556 8024 3584
rect 7340 3544 7346 3556
rect 8018 3544 8024 3556
rect 8076 3584 8082 3596
rect 9677 3587 9735 3593
rect 8076 3556 8248 3584
rect 8076 3544 8082 3556
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 4798 3476 4804 3528
rect 4856 3516 4862 3528
rect 5261 3519 5319 3525
rect 5261 3516 5273 3519
rect 4856 3488 5273 3516
rect 4856 3476 4862 3488
rect 5261 3485 5273 3488
rect 5307 3485 5319 3519
rect 5261 3479 5319 3485
rect 5813 3519 5871 3525
rect 5813 3485 5825 3519
rect 5859 3516 5871 3519
rect 7650 3516 7656 3528
rect 5859 3488 7656 3516
rect 5859 3485 5871 3488
rect 5813 3479 5871 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8220 3525 8248 3556
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 10778 3584 10784 3596
rect 9723 3556 10784 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 10778 3544 10784 3556
rect 10836 3544 10842 3596
rect 11146 3584 11152 3596
rect 11107 3556 11152 3584
rect 11146 3544 11152 3556
rect 11204 3544 11210 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 11405 3587 11463 3593
rect 11405 3584 11417 3587
rect 11296 3556 11417 3584
rect 11296 3544 11302 3556
rect 11405 3553 11417 3556
rect 11451 3553 11463 3587
rect 11405 3547 11463 3553
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 10226 3516 10232 3528
rect 8812 3488 10232 3516
rect 8812 3476 8818 3488
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 3053 3451 3111 3457
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 3510 3448 3516 3460
rect 3099 3420 3516 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 3510 3408 3516 3420
rect 3568 3408 3574 3460
rect 4982 3408 4988 3460
rect 5040 3448 5046 3460
rect 6457 3451 6515 3457
rect 6457 3448 6469 3451
rect 5040 3420 6469 3448
rect 5040 3408 5046 3420
rect 6457 3417 6469 3420
rect 6503 3417 6515 3451
rect 6457 3411 6515 3417
rect 12529 3451 12587 3457
rect 12529 3417 12541 3451
rect 12575 3448 12587 3451
rect 12710 3448 12716 3460
rect 12575 3420 12716 3448
rect 12575 3417 12587 3420
rect 12529 3411 12587 3417
rect 12710 3408 12716 3420
rect 12768 3408 12774 3460
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2130 3380 2136 3392
rect 1995 3352 2136 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 9858 3380 9864 3392
rect 9819 3352 9864 3380
rect 9858 3340 9864 3352
rect 9916 3340 9922 3392
rect 13078 3380 13084 3392
rect 13039 3352 13084 3380
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 1104 3290 14812 3312
rect 1104 3238 3648 3290
rect 3700 3238 3712 3290
rect 3764 3238 3776 3290
rect 3828 3238 3840 3290
rect 3892 3238 8982 3290
rect 9034 3238 9046 3290
rect 9098 3238 9110 3290
rect 9162 3238 9174 3290
rect 9226 3238 14315 3290
rect 14367 3238 14379 3290
rect 14431 3238 14443 3290
rect 14495 3238 14507 3290
rect 14559 3238 14812 3290
rect 1104 3216 14812 3238
rect 1762 3176 1768 3188
rect 1723 3148 1768 3176
rect 1762 3136 1768 3148
rect 1820 3136 1826 3188
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2924 3148 2973 3176
rect 2924 3136 2930 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 5626 3176 5632 3188
rect 5587 3148 5632 3176
rect 2961 3139 3019 3145
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6638 3176 6644 3188
rect 6411 3148 6644 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 7156 3148 7205 3176
rect 7156 3136 7162 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 9674 3136 9680 3188
rect 9732 3176 9738 3188
rect 10137 3179 10195 3185
rect 10137 3176 10149 3179
rect 9732 3148 10149 3176
rect 9732 3136 9738 3148
rect 10137 3145 10149 3148
rect 10183 3145 10195 3179
rect 10778 3176 10784 3188
rect 10739 3148 10784 3176
rect 10137 3139 10195 3145
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11422 3176 11428 3188
rect 11383 3148 11428 3176
rect 11422 3136 11428 3148
rect 11480 3136 11486 3188
rect 12066 3176 12072 3188
rect 11979 3148 12072 3176
rect 12066 3136 12072 3148
rect 12124 3176 12130 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12124 3148 12173 3176
rect 12124 3136 12130 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12161 3139 12219 3145
rect 12437 3179 12495 3185
rect 12437 3145 12449 3179
rect 12483 3176 12495 3179
rect 13078 3176 13084 3188
rect 12483 3148 13084 3176
rect 12483 3145 12495 3148
rect 12437 3139 12495 3145
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 2222 3108 2228 3120
rect 2183 3080 2228 3108
rect 2222 3068 2228 3080
rect 2280 3068 2286 3120
rect 3326 3040 3332 3052
rect 2608 3012 3332 3040
rect 2608 2981 2636 3012
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4154 3000 4160 3052
rect 4212 3040 4218 3052
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4212 3012 4261 3040
rect 4212 3000 4218 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 7650 3040 7656 3052
rect 7611 3012 7656 3040
rect 4249 3003 4307 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8018 3040 8024 3052
rect 7883 3012 8024 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13262 3040 13268 3052
rect 13127 3012 13268 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13262 3000 13268 3012
rect 13320 3040 13326 3052
rect 13449 3043 13507 3049
rect 13449 3040 13461 3043
rect 13320 3012 13461 3040
rect 13320 3000 13326 3012
rect 13449 3009 13461 3012
rect 13495 3009 13507 3043
rect 13449 3003 13507 3009
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 2593 2975 2651 2981
rect 2593 2972 2605 2975
rect 2087 2944 2605 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 2593 2941 2605 2944
rect 2639 2941 2651 2975
rect 2593 2935 2651 2941
rect 3145 2975 3203 2981
rect 3145 2941 3157 2975
rect 3191 2972 3203 2975
rect 3234 2972 3240 2984
rect 3191 2944 3240 2972
rect 3191 2941 3203 2944
rect 3145 2935 3203 2941
rect 3234 2932 3240 2944
rect 3292 2972 3298 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3292 2944 3709 2972
rect 3292 2932 3298 2944
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 4516 2975 4574 2981
rect 4516 2941 4528 2975
rect 4562 2972 4574 2975
rect 4798 2972 4804 2984
rect 4562 2944 4804 2972
rect 4562 2941 4574 2944
rect 4516 2935 4574 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2972 7159 2975
rect 7561 2975 7619 2981
rect 7561 2972 7573 2975
rect 7147 2944 7573 2972
rect 7147 2941 7159 2944
rect 7101 2935 7159 2941
rect 7561 2941 7573 2944
rect 7607 2972 7619 2975
rect 7926 2972 7932 2984
rect 7607 2944 7932 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8757 2975 8815 2981
rect 8757 2941 8769 2975
rect 8803 2972 8815 2975
rect 11149 2975 11207 2981
rect 8803 2944 9251 2972
rect 8803 2941 8815 2944
rect 8757 2935 8815 2941
rect 4157 2907 4215 2913
rect 4157 2873 4169 2907
rect 4203 2904 4215 2907
rect 5074 2904 5080 2916
rect 4203 2876 5080 2904
rect 4203 2873 4215 2876
rect 4157 2867 4215 2873
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 9030 2913 9036 2916
rect 8297 2907 8355 2913
rect 8297 2873 8309 2907
rect 8343 2904 8355 2907
rect 9002 2907 9036 2913
rect 9002 2904 9014 2907
rect 8343 2876 9014 2904
rect 8343 2873 8355 2876
rect 8297 2867 8355 2873
rect 9002 2873 9014 2876
rect 9088 2904 9094 2916
rect 9088 2876 9150 2904
rect 9002 2867 9036 2873
rect 9030 2864 9036 2867
rect 9088 2864 9094 2876
rect 3326 2836 3332 2848
rect 3287 2808 3332 2836
rect 3326 2796 3332 2808
rect 3384 2796 3390 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9223 2836 9251 2944
rect 11149 2941 11161 2975
rect 11195 2972 11207 2975
rect 11241 2975 11299 2981
rect 11241 2972 11253 2975
rect 11195 2944 11253 2972
rect 11195 2941 11207 2944
rect 11149 2935 11207 2941
rect 11241 2941 11253 2944
rect 11287 2972 11299 2975
rect 11287 2944 11928 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11900 2913 11928 2944
rect 11885 2907 11943 2913
rect 11885 2873 11897 2907
rect 11931 2904 11943 2907
rect 12894 2904 12900 2916
rect 11931 2876 12900 2904
rect 11931 2873 11943 2876
rect 11885 2867 11943 2873
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 9490 2836 9496 2848
rect 8711 2808 9496 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9490 2796 9496 2808
rect 9548 2796 9554 2848
rect 12069 2839 12127 2845
rect 12069 2805 12081 2839
rect 12115 2836 12127 2839
rect 12805 2839 12863 2845
rect 12805 2836 12817 2839
rect 12115 2808 12817 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 12805 2805 12817 2808
rect 12851 2836 12863 2839
rect 14918 2836 14924 2848
rect 12851 2808 14924 2836
rect 12851 2805 12863 2808
rect 12805 2799 12863 2805
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 1104 2746 14812 2768
rect 1104 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 11648 2746
rect 11700 2694 11712 2746
rect 11764 2694 11776 2746
rect 11828 2694 11840 2746
rect 11892 2694 14812 2746
rect 1104 2672 14812 2694
rect 1946 2632 1952 2644
rect 1907 2604 1952 2632
rect 1946 2592 1952 2604
rect 2004 2592 2010 2644
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4709 2635 4767 2641
rect 4709 2601 4721 2635
rect 4755 2632 4767 2635
rect 5258 2632 5264 2644
rect 4755 2604 5264 2632
rect 4755 2601 4767 2604
rect 4709 2595 4767 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 7098 2632 7104 2644
rect 7059 2604 7104 2632
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7466 2632 7472 2644
rect 7427 2604 7472 2632
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 7650 2592 7656 2644
rect 7708 2632 7714 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7708 2604 8125 2632
rect 7708 2592 7714 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 8481 2635 8539 2641
rect 8481 2601 8493 2635
rect 8527 2632 8539 2635
rect 9582 2632 9588 2644
rect 8527 2604 9588 2632
rect 8527 2601 8539 2604
rect 8481 2595 8539 2601
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 11701 2635 11759 2641
rect 11701 2632 11713 2635
rect 11204 2604 11713 2632
rect 11204 2592 11210 2604
rect 11701 2601 11713 2604
rect 11747 2601 11759 2635
rect 11701 2595 11759 2601
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12618 2632 12624 2644
rect 12492 2604 12537 2632
rect 12579 2604 12624 2632
rect 12492 2592 12498 2604
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 3513 2567 3571 2573
rect 3513 2533 3525 2567
rect 3559 2564 3571 2567
rect 4338 2564 4344 2576
rect 3559 2536 4344 2564
rect 3559 2533 3571 2536
rect 3513 2527 3571 2533
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 2869 2499 2927 2505
rect 1811 2468 2452 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 2424 2369 2452 2468
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3528 2496 3556 2527
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 2915 2468 3556 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 4798 2456 4804 2508
rect 4856 2456 4862 2508
rect 5166 2496 5172 2508
rect 5127 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2496 5230 2508
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 5224 2468 5825 2496
rect 5224 2456 5230 2468
rect 5813 2465 5825 2468
rect 5859 2465 5871 2499
rect 5813 2459 5871 2465
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7484 2496 7512 2592
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 9398 2564 9404 2576
rect 9263 2536 9404 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 9398 2524 9404 2536
rect 9456 2564 9462 2576
rect 10014 2567 10072 2573
rect 10014 2564 10026 2567
rect 9456 2536 10026 2564
rect 9456 2524 9462 2536
rect 10014 2533 10026 2536
rect 10060 2533 10072 2567
rect 10014 2527 10072 2533
rect 6963 2468 7512 2496
rect 8021 2499 8079 2505
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8021 2465 8033 2499
rect 8067 2496 8079 2499
rect 8067 2468 8800 2496
rect 8067 2465 8079 2468
rect 8021 2459 8079 2465
rect 3881 2431 3939 2437
rect 3881 2397 3893 2431
rect 3927 2428 3939 2431
rect 4816 2428 4844 2456
rect 5353 2431 5411 2437
rect 5353 2428 5365 2431
rect 3927 2400 5365 2428
rect 3927 2397 3939 2400
rect 3881 2391 3939 2397
rect 5353 2397 5365 2400
rect 5399 2428 5411 2431
rect 6181 2431 6239 2437
rect 6181 2428 6193 2431
rect 5399 2400 6193 2428
rect 5399 2397 5411 2400
rect 5353 2391 5411 2397
rect 6181 2397 6193 2400
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 8570 2428 8576 2440
rect 6779 2400 8576 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 8772 2437 8800 2468
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9548 2468 9597 2496
rect 9548 2456 9554 2468
rect 9585 2465 9597 2468
rect 9631 2496 9643 2499
rect 9769 2499 9827 2505
rect 9769 2496 9781 2499
rect 9631 2468 9781 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 9769 2465 9781 2468
rect 9815 2496 9827 2499
rect 11164 2496 11192 2592
rect 12452 2564 12480 2592
rect 13081 2567 13139 2573
rect 13081 2564 13093 2567
rect 12452 2536 13093 2564
rect 13081 2533 13093 2536
rect 13127 2533 13139 2567
rect 13081 2527 13139 2533
rect 12986 2496 12992 2508
rect 9815 2468 11192 2496
rect 12899 2468 12992 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 12986 2456 12992 2468
rect 13044 2496 13050 2508
rect 13633 2499 13691 2505
rect 13633 2496 13645 2499
rect 13044 2468 13645 2496
rect 13044 2456 13050 2468
rect 13633 2465 13645 2468
rect 13679 2465 13691 2499
rect 13633 2459 13691 2465
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9030 2428 9036 2440
rect 8803 2400 9036 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 9030 2388 9036 2400
rect 9088 2428 9094 2440
rect 13262 2428 13268 2440
rect 9088 2400 9260 2428
rect 13223 2400 13268 2428
rect 9088 2388 9094 2400
rect 2409 2363 2467 2369
rect 2409 2329 2421 2363
rect 2455 2360 2467 2363
rect 4801 2363 4859 2369
rect 2455 2332 4016 2360
rect 2455 2329 2467 2332
rect 2409 2323 2467 2329
rect 2958 2252 2964 2304
rect 3016 2292 3022 2304
rect 3053 2295 3111 2301
rect 3053 2292 3065 2295
rect 3016 2264 3065 2292
rect 3016 2252 3022 2264
rect 3053 2261 3065 2264
rect 3099 2261 3111 2295
rect 3988 2292 4016 2332
rect 4801 2329 4813 2363
rect 4847 2360 4859 2363
rect 5442 2360 5448 2372
rect 4847 2332 5448 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 5442 2320 5448 2332
rect 5500 2320 5506 2372
rect 7834 2292 7840 2304
rect 3988 2264 7840 2292
rect 3053 2255 3111 2261
rect 7834 2252 7840 2264
rect 7892 2252 7898 2304
rect 9232 2292 9260 2400
rect 13262 2388 13268 2400
rect 13320 2428 13326 2440
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 13320 2400 14013 2428
rect 13320 2388 13326 2400
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 9232 2264 11161 2292
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 1104 2202 14812 2224
rect 1104 2150 3648 2202
rect 3700 2150 3712 2202
rect 3764 2150 3776 2202
rect 3828 2150 3840 2202
rect 3892 2150 8982 2202
rect 9034 2150 9046 2202
rect 9098 2150 9110 2202
rect 9162 2150 9174 2202
rect 9226 2150 14315 2202
rect 14367 2150 14379 2202
rect 14431 2150 14443 2202
rect 14495 2150 14507 2202
rect 14559 2150 14812 2202
rect 1104 2128 14812 2150
<< via1 >>
rect 6315 37510 6367 37562
rect 6379 37510 6431 37562
rect 6443 37510 6495 37562
rect 6507 37510 6559 37562
rect 11648 37510 11700 37562
rect 11712 37510 11764 37562
rect 11776 37510 11828 37562
rect 11840 37510 11892 37562
rect 3648 36966 3700 37018
rect 3712 36966 3764 37018
rect 3776 36966 3828 37018
rect 3840 36966 3892 37018
rect 8982 36966 9034 37018
rect 9046 36966 9098 37018
rect 9110 36966 9162 37018
rect 9174 36966 9226 37018
rect 14315 36966 14367 37018
rect 14379 36966 14431 37018
rect 14443 36966 14495 37018
rect 14507 36966 14559 37018
rect 6184 36864 6236 36916
rect 5264 36660 5316 36712
rect 6315 36422 6367 36474
rect 6379 36422 6431 36474
rect 6443 36422 6495 36474
rect 6507 36422 6559 36474
rect 11648 36422 11700 36474
rect 11712 36422 11764 36474
rect 11776 36422 11828 36474
rect 11840 36422 11892 36474
rect 5356 36320 5408 36372
rect 6644 36320 6696 36372
rect 4712 36227 4764 36236
rect 4712 36193 4721 36227
rect 4721 36193 4755 36227
rect 4755 36193 4764 36227
rect 4712 36184 4764 36193
rect 6000 36184 6052 36236
rect 3648 35878 3700 35930
rect 3712 35878 3764 35930
rect 3776 35878 3828 35930
rect 3840 35878 3892 35930
rect 8982 35878 9034 35930
rect 9046 35878 9098 35930
rect 9110 35878 9162 35930
rect 9174 35878 9226 35930
rect 14315 35878 14367 35930
rect 14379 35878 14431 35930
rect 14443 35878 14495 35930
rect 14507 35878 14559 35930
rect 3332 35776 3384 35828
rect 3424 35776 3476 35828
rect 4252 35776 4304 35828
rect 7380 35776 7432 35828
rect 9864 35751 9916 35760
rect 9864 35717 9873 35751
rect 9873 35717 9907 35751
rect 9907 35717 9916 35751
rect 9864 35708 9916 35717
rect 4712 35640 4764 35692
rect 5816 35640 5868 35692
rect 4068 35572 4120 35624
rect 3516 35436 3568 35488
rect 5632 35479 5684 35488
rect 5632 35445 5641 35479
rect 5641 35445 5675 35479
rect 5675 35445 5684 35479
rect 5632 35436 5684 35445
rect 6000 35479 6052 35488
rect 6000 35445 6009 35479
rect 6009 35445 6043 35479
rect 6043 35445 6052 35479
rect 6000 35436 6052 35445
rect 9588 35436 9640 35488
rect 10692 35436 10744 35488
rect 6315 35334 6367 35386
rect 6379 35334 6431 35386
rect 6443 35334 6495 35386
rect 6507 35334 6559 35386
rect 11648 35334 11700 35386
rect 11712 35334 11764 35386
rect 11776 35334 11828 35386
rect 11840 35334 11892 35386
rect 940 35232 992 35284
rect 2136 35232 2188 35284
rect 5080 35275 5132 35284
rect 5080 35241 5089 35275
rect 5089 35241 5123 35275
rect 5123 35241 5132 35275
rect 5080 35232 5132 35241
rect 5724 35232 5776 35284
rect 7564 35275 7616 35284
rect 7564 35241 7573 35275
rect 7573 35241 7607 35275
rect 7607 35241 7616 35275
rect 7564 35232 7616 35241
rect 1676 35096 1728 35148
rect 3424 35096 3476 35148
rect 4896 35139 4948 35148
rect 4896 35105 4905 35139
rect 4905 35105 4939 35139
rect 4939 35105 4948 35139
rect 4896 35096 4948 35105
rect 6276 35139 6328 35148
rect 6276 35105 6285 35139
rect 6285 35105 6319 35139
rect 6319 35105 6328 35139
rect 6276 35096 6328 35105
rect 7656 35096 7708 35148
rect 8760 35096 8812 35148
rect 9496 35096 9548 35148
rect 9680 35071 9732 35080
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 12348 35071 12400 35080
rect 9680 35028 9732 35037
rect 12348 35037 12357 35071
rect 12357 35037 12391 35071
rect 12391 35037 12400 35071
rect 12348 35028 12400 35037
rect 6920 34960 6972 35012
rect 7932 34935 7984 34944
rect 7932 34901 7941 34935
rect 7941 34901 7975 34935
rect 7975 34901 7984 34935
rect 7932 34892 7984 34901
rect 10784 34892 10836 34944
rect 12900 34935 12952 34944
rect 12900 34901 12909 34935
rect 12909 34901 12943 34935
rect 12943 34901 12952 34935
rect 12900 34892 12952 34901
rect 3648 34790 3700 34842
rect 3712 34790 3764 34842
rect 3776 34790 3828 34842
rect 3840 34790 3892 34842
rect 8982 34790 9034 34842
rect 9046 34790 9098 34842
rect 9110 34790 9162 34842
rect 9174 34790 9226 34842
rect 14315 34790 14367 34842
rect 14379 34790 14431 34842
rect 14443 34790 14495 34842
rect 14507 34790 14559 34842
rect 204 34688 256 34740
rect 2688 34731 2740 34740
rect 2688 34697 2697 34731
rect 2697 34697 2731 34731
rect 2731 34697 2740 34731
rect 2688 34688 2740 34697
rect 7656 34688 7708 34740
rect 9680 34731 9732 34740
rect 9680 34697 9689 34731
rect 9689 34697 9723 34731
rect 9723 34697 9732 34731
rect 9680 34688 9732 34697
rect 12348 34688 12400 34740
rect 9864 34595 9916 34604
rect 2228 34484 2280 34536
rect 2504 34527 2556 34536
rect 2504 34493 2513 34527
rect 2513 34493 2547 34527
rect 2547 34493 2556 34527
rect 2504 34484 2556 34493
rect 3424 34484 3476 34536
rect 9864 34561 9873 34595
rect 9873 34561 9907 34595
rect 9907 34561 9916 34595
rect 9864 34552 9916 34561
rect 12072 34552 12124 34604
rect 12900 34552 12952 34604
rect 3976 34416 4028 34468
rect 4896 34484 4948 34536
rect 5908 34484 5960 34536
rect 6276 34484 6328 34536
rect 6828 34484 6880 34536
rect 7380 34527 7432 34536
rect 7380 34493 7389 34527
rect 7389 34493 7423 34527
rect 7423 34493 7432 34527
rect 7380 34484 7432 34493
rect 7932 34484 7984 34536
rect 8760 34484 8812 34536
rect 12348 34484 12400 34536
rect 4712 34416 4764 34468
rect 10784 34416 10836 34468
rect 13176 34484 13228 34536
rect 4804 34348 4856 34400
rect 8852 34348 8904 34400
rect 9496 34348 9548 34400
rect 11244 34391 11296 34400
rect 11244 34357 11253 34391
rect 11253 34357 11287 34391
rect 11287 34357 11296 34391
rect 11244 34348 11296 34357
rect 12440 34391 12492 34400
rect 12440 34357 12449 34391
rect 12449 34357 12483 34391
rect 12483 34357 12492 34391
rect 12440 34348 12492 34357
rect 6315 34246 6367 34298
rect 6379 34246 6431 34298
rect 6443 34246 6495 34298
rect 6507 34246 6559 34298
rect 11648 34246 11700 34298
rect 11712 34246 11764 34298
rect 11776 34246 11828 34298
rect 11840 34246 11892 34298
rect 1400 34144 1452 34196
rect 9496 34187 9548 34196
rect 9496 34153 9505 34187
rect 9505 34153 9539 34187
rect 9539 34153 9548 34187
rect 9496 34144 9548 34153
rect 9864 34187 9916 34196
rect 9864 34153 9873 34187
rect 9873 34153 9907 34187
rect 9907 34153 9916 34187
rect 9864 34144 9916 34153
rect 1676 34119 1728 34128
rect 1676 34085 1685 34119
rect 1685 34085 1719 34119
rect 1719 34085 1728 34119
rect 1676 34076 1728 34085
rect 11244 34119 11296 34128
rect 11244 34085 11253 34119
rect 11253 34085 11287 34119
rect 11287 34085 11296 34119
rect 12072 34119 12124 34128
rect 11244 34076 11296 34085
rect 12072 34085 12106 34119
rect 12106 34085 12124 34119
rect 12072 34076 12124 34085
rect 2596 34008 2648 34060
rect 4804 34008 4856 34060
rect 6276 34008 6328 34060
rect 8484 34008 8536 34060
rect 8576 34008 8628 34060
rect 10232 34008 10284 34060
rect 11060 34008 11112 34060
rect 11796 34051 11848 34060
rect 11796 34017 11805 34051
rect 11805 34017 11839 34051
rect 11839 34017 11848 34051
rect 11796 34008 11848 34017
rect 4712 33983 4764 33992
rect 4712 33949 4721 33983
rect 4721 33949 4755 33983
rect 4755 33949 4764 33983
rect 4712 33940 4764 33949
rect 3976 33804 4028 33856
rect 6092 33847 6144 33856
rect 6092 33813 6101 33847
rect 6101 33813 6135 33847
rect 6135 33813 6144 33847
rect 6092 33804 6144 33813
rect 6920 33804 6972 33856
rect 8852 33940 8904 33992
rect 10324 33940 10376 33992
rect 10784 33983 10836 33992
rect 10784 33949 10793 33983
rect 10793 33949 10827 33983
rect 10827 33949 10836 33983
rect 10784 33940 10836 33949
rect 7380 33872 7432 33924
rect 7840 33872 7892 33924
rect 7564 33847 7616 33856
rect 7564 33813 7573 33847
rect 7573 33813 7607 33847
rect 7607 33813 7616 33847
rect 7564 33804 7616 33813
rect 10508 33804 10560 33856
rect 12900 33804 12952 33856
rect 3648 33702 3700 33754
rect 3712 33702 3764 33754
rect 3776 33702 3828 33754
rect 3840 33702 3892 33754
rect 8982 33702 9034 33754
rect 9046 33702 9098 33754
rect 9110 33702 9162 33754
rect 9174 33702 9226 33754
rect 14315 33702 14367 33754
rect 14379 33702 14431 33754
rect 14443 33702 14495 33754
rect 14507 33702 14559 33754
rect 1492 33600 1544 33652
rect 2964 33600 3016 33652
rect 4160 33643 4212 33652
rect 4160 33609 4169 33643
rect 4169 33609 4203 33643
rect 4203 33609 4212 33643
rect 4160 33600 4212 33609
rect 4988 33600 5040 33652
rect 6276 33643 6328 33652
rect 6276 33609 6285 33643
rect 6285 33609 6319 33643
rect 6319 33609 6328 33643
rect 6276 33600 6328 33609
rect 8852 33643 8904 33652
rect 8852 33609 8861 33643
rect 8861 33609 8895 33643
rect 8895 33609 8904 33643
rect 8852 33600 8904 33609
rect 10784 33600 10836 33652
rect 11796 33600 11848 33652
rect 9680 33575 9732 33584
rect 9680 33541 9689 33575
rect 9689 33541 9723 33575
rect 9723 33541 9732 33575
rect 9680 33532 9732 33541
rect 10324 33532 10376 33584
rect 4712 33464 4764 33516
rect 11244 33507 11296 33516
rect 1952 33371 2004 33380
rect 1952 33337 1961 33371
rect 1961 33337 1995 33371
rect 1995 33337 2004 33371
rect 1952 33328 2004 33337
rect 2596 33260 2648 33312
rect 6736 33396 6788 33448
rect 11244 33473 11253 33507
rect 11253 33473 11287 33507
rect 11287 33473 11296 33507
rect 11244 33464 11296 33473
rect 12900 33464 12952 33516
rect 7840 33396 7892 33448
rect 11152 33396 11204 33448
rect 12440 33396 12492 33448
rect 6092 33328 6144 33380
rect 7104 33371 7156 33380
rect 7104 33337 7116 33371
rect 7116 33337 7156 33371
rect 7104 33328 7156 33337
rect 10508 33328 10560 33380
rect 4068 33260 4120 33312
rect 4620 33303 4672 33312
rect 4620 33269 4629 33303
rect 4629 33269 4663 33303
rect 4663 33269 4672 33303
rect 4620 33260 4672 33269
rect 6828 33260 6880 33312
rect 7472 33260 7524 33312
rect 10600 33303 10652 33312
rect 10600 33269 10609 33303
rect 10609 33269 10643 33303
rect 10643 33269 10652 33303
rect 10600 33260 10652 33269
rect 10784 33260 10836 33312
rect 12348 33260 12400 33312
rect 12900 33303 12952 33312
rect 12900 33269 12909 33303
rect 12909 33269 12943 33303
rect 12943 33269 12952 33303
rect 12900 33260 12952 33269
rect 6315 33158 6367 33210
rect 6379 33158 6431 33210
rect 6443 33158 6495 33210
rect 6507 33158 6559 33210
rect 11648 33158 11700 33210
rect 11712 33158 11764 33210
rect 11776 33158 11828 33210
rect 11840 33158 11892 33210
rect 1584 33099 1636 33108
rect 1584 33065 1593 33099
rect 1593 33065 1627 33099
rect 1627 33065 1636 33099
rect 1584 33056 1636 33065
rect 5448 33056 5500 33108
rect 7380 33056 7432 33108
rect 8024 33056 8076 33108
rect 9956 33056 10008 33108
rect 10232 33099 10284 33108
rect 10232 33065 10241 33099
rect 10241 33065 10275 33099
rect 10275 33065 10284 33099
rect 10232 33056 10284 33065
rect 10508 33099 10560 33108
rect 10508 33065 10517 33099
rect 10517 33065 10551 33099
rect 10551 33065 10560 33099
rect 10508 33056 10560 33065
rect 10600 33056 10652 33108
rect 12716 33099 12768 33108
rect 12716 33065 12725 33099
rect 12725 33065 12759 33099
rect 12759 33065 12768 33099
rect 12716 33056 12768 33065
rect 7104 32988 7156 33040
rect 1400 32963 1452 32972
rect 1400 32929 1409 32963
rect 1409 32929 1443 32963
rect 1443 32929 1452 32963
rect 1400 32920 1452 32929
rect 11520 32988 11572 33040
rect 12348 32988 12400 33040
rect 12624 32963 12676 32972
rect 6184 32895 6236 32904
rect 6184 32861 6193 32895
rect 6193 32861 6227 32895
rect 6227 32861 6236 32895
rect 6184 32852 6236 32861
rect 6368 32895 6420 32904
rect 6368 32861 6377 32895
rect 6377 32861 6411 32895
rect 6411 32861 6420 32895
rect 6368 32852 6420 32861
rect 6828 32852 6880 32904
rect 7288 32852 7340 32904
rect 7748 32895 7800 32904
rect 7748 32861 7757 32895
rect 7757 32861 7791 32895
rect 7791 32861 7800 32895
rect 7748 32852 7800 32861
rect 12624 32929 12633 32963
rect 12633 32929 12667 32963
rect 12667 32929 12676 32963
rect 12624 32920 12676 32929
rect 10048 32852 10100 32904
rect 10324 32852 10376 32904
rect 12348 32852 12400 32904
rect 12808 32895 12860 32904
rect 12808 32861 12817 32895
rect 12817 32861 12851 32895
rect 12851 32861 12860 32895
rect 12808 32852 12860 32861
rect 9864 32784 9916 32836
rect 11152 32784 11204 32836
rect 12072 32784 12124 32836
rect 3332 32759 3384 32768
rect 3332 32725 3341 32759
rect 3341 32725 3375 32759
rect 3375 32725 3384 32759
rect 3332 32716 3384 32725
rect 4160 32716 4212 32768
rect 4804 32716 4856 32768
rect 5724 32759 5776 32768
rect 5724 32725 5733 32759
rect 5733 32725 5767 32759
rect 5767 32725 5776 32759
rect 5724 32716 5776 32725
rect 8300 32759 8352 32768
rect 8300 32725 8309 32759
rect 8309 32725 8343 32759
rect 8343 32725 8352 32759
rect 8300 32716 8352 32725
rect 11244 32716 11296 32768
rect 11796 32759 11848 32768
rect 11796 32725 11805 32759
rect 11805 32725 11839 32759
rect 11839 32725 11848 32759
rect 11796 32716 11848 32725
rect 12440 32716 12492 32768
rect 12900 32716 12952 32768
rect 3648 32614 3700 32666
rect 3712 32614 3764 32666
rect 3776 32614 3828 32666
rect 3840 32614 3892 32666
rect 8982 32614 9034 32666
rect 9046 32614 9098 32666
rect 9110 32614 9162 32666
rect 9174 32614 9226 32666
rect 14315 32614 14367 32666
rect 14379 32614 14431 32666
rect 14443 32614 14495 32666
rect 14507 32614 14559 32666
rect 1400 32512 1452 32564
rect 5448 32555 5500 32564
rect 5448 32521 5457 32555
rect 5457 32521 5491 32555
rect 5491 32521 5500 32555
rect 5448 32512 5500 32521
rect 6184 32555 6236 32564
rect 6184 32521 6193 32555
rect 6193 32521 6227 32555
rect 6227 32521 6236 32555
rect 6184 32512 6236 32521
rect 7380 32512 7432 32564
rect 7932 32512 7984 32564
rect 8392 32512 8444 32564
rect 10600 32512 10652 32564
rect 10784 32555 10836 32564
rect 10784 32521 10793 32555
rect 10793 32521 10827 32555
rect 10827 32521 10836 32555
rect 10784 32512 10836 32521
rect 11796 32555 11848 32564
rect 11796 32521 11805 32555
rect 11805 32521 11839 32555
rect 11839 32521 11848 32555
rect 11796 32512 11848 32521
rect 12072 32512 12124 32564
rect 12256 32512 12308 32564
rect 12440 32555 12492 32564
rect 12440 32521 12449 32555
rect 12449 32521 12483 32555
rect 12483 32521 12492 32555
rect 12440 32512 12492 32521
rect 12624 32512 12676 32564
rect 6368 32444 6420 32496
rect 10324 32487 10376 32496
rect 10324 32453 10333 32487
rect 10333 32453 10367 32487
rect 10367 32453 10376 32487
rect 10324 32444 10376 32453
rect 3332 32376 3384 32428
rect 3792 32419 3844 32428
rect 3792 32385 3801 32419
rect 3801 32385 3835 32419
rect 3835 32385 3844 32419
rect 3792 32376 3844 32385
rect 10784 32376 10836 32428
rect 12716 32444 12768 32496
rect 3700 32351 3752 32360
rect 3700 32317 3709 32351
rect 3709 32317 3743 32351
rect 3743 32317 3752 32351
rect 3700 32308 3752 32317
rect 7288 32351 7340 32360
rect 7288 32317 7297 32351
rect 7297 32317 7331 32351
rect 7331 32317 7340 32351
rect 7288 32308 7340 32317
rect 7840 32308 7892 32360
rect 8024 32351 8076 32360
rect 8024 32317 8058 32351
rect 8058 32317 8076 32351
rect 8024 32308 8076 32317
rect 8300 32308 8352 32360
rect 12532 32308 12584 32360
rect 13176 32308 13228 32360
rect 3240 32215 3292 32224
rect 3240 32181 3249 32215
rect 3249 32181 3283 32215
rect 3283 32181 3292 32215
rect 3240 32172 3292 32181
rect 3608 32215 3660 32224
rect 3608 32181 3617 32215
rect 3617 32181 3651 32215
rect 3651 32181 3660 32215
rect 3608 32172 3660 32181
rect 4988 32172 5040 32224
rect 10692 32215 10744 32224
rect 10692 32181 10701 32215
rect 10701 32181 10735 32215
rect 10735 32181 10744 32215
rect 11152 32215 11204 32224
rect 10692 32172 10744 32181
rect 11152 32181 11161 32215
rect 11161 32181 11195 32215
rect 11195 32181 11204 32215
rect 11152 32172 11204 32181
rect 12256 32172 12308 32224
rect 6315 32070 6367 32122
rect 6379 32070 6431 32122
rect 6443 32070 6495 32122
rect 6507 32070 6559 32122
rect 11648 32070 11700 32122
rect 11712 32070 11764 32122
rect 11776 32070 11828 32122
rect 11840 32070 11892 32122
rect 3700 31968 3752 32020
rect 6184 31968 6236 32020
rect 6644 31968 6696 32020
rect 8852 31968 8904 32020
rect 10048 32011 10100 32020
rect 10048 31977 10057 32011
rect 10057 31977 10091 32011
rect 10091 31977 10100 32011
rect 10048 31968 10100 31977
rect 3792 31900 3844 31952
rect 4804 31900 4856 31952
rect 6828 31900 6880 31952
rect 7196 31900 7248 31952
rect 9680 31832 9732 31884
rect 10232 31968 10284 32020
rect 10324 31968 10376 32020
rect 10784 32011 10836 32020
rect 10784 31977 10793 32011
rect 10793 31977 10827 32011
rect 10827 31977 10836 32011
rect 10784 31968 10836 31977
rect 11244 32011 11296 32020
rect 11244 31977 11253 32011
rect 11253 31977 11287 32011
rect 11287 31977 11296 32011
rect 11244 31968 11296 31977
rect 11520 32011 11572 32020
rect 11520 31977 11529 32011
rect 11529 31977 11563 32011
rect 11563 31977 11572 32011
rect 11520 31968 11572 31977
rect 12532 32011 12584 32020
rect 12532 31977 12541 32011
rect 12541 31977 12575 32011
rect 12575 31977 12584 32011
rect 12532 31968 12584 31977
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 7932 31764 7984 31816
rect 9588 31764 9640 31816
rect 12808 31807 12860 31816
rect 7380 31696 7432 31748
rect 9772 31696 9824 31748
rect 9956 31696 10008 31748
rect 10600 31696 10652 31748
rect 4252 31628 4304 31680
rect 4712 31628 4764 31680
rect 5080 31628 5132 31680
rect 7840 31671 7892 31680
rect 7840 31637 7849 31671
rect 7849 31637 7883 31671
rect 7883 31637 7892 31671
rect 7840 31628 7892 31637
rect 9588 31628 9640 31680
rect 10692 31628 10744 31680
rect 12072 31628 12124 31680
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 12808 31764 12860 31773
rect 3648 31526 3700 31578
rect 3712 31526 3764 31578
rect 3776 31526 3828 31578
rect 3840 31526 3892 31578
rect 8982 31526 9034 31578
rect 9046 31526 9098 31578
rect 9110 31526 9162 31578
rect 9174 31526 9226 31578
rect 14315 31526 14367 31578
rect 14379 31526 14431 31578
rect 14443 31526 14495 31578
rect 14507 31526 14559 31578
rect 4252 31424 4304 31476
rect 6920 31467 6972 31476
rect 6920 31433 6929 31467
rect 6929 31433 6963 31467
rect 6963 31433 6972 31467
rect 6920 31424 6972 31433
rect 7932 31467 7984 31476
rect 7932 31433 7941 31467
rect 7941 31433 7975 31467
rect 7975 31433 7984 31467
rect 7932 31424 7984 31433
rect 8300 31424 8352 31476
rect 9680 31424 9732 31476
rect 13544 31467 13596 31476
rect 3516 31356 3568 31408
rect 6828 31356 6880 31408
rect 4068 31288 4120 31340
rect 5080 31331 5132 31340
rect 5080 31297 5089 31331
rect 5089 31297 5123 31331
rect 5123 31297 5132 31331
rect 5080 31288 5132 31297
rect 7564 31331 7616 31340
rect 7564 31297 7573 31331
rect 7573 31297 7607 31331
rect 7607 31297 7616 31331
rect 7564 31288 7616 31297
rect 8208 31288 8260 31340
rect 4804 31152 4856 31204
rect 8576 31288 8628 31340
rect 8852 31263 8904 31272
rect 8852 31229 8861 31263
rect 8861 31229 8895 31263
rect 8895 31229 8904 31263
rect 8852 31220 8904 31229
rect 13544 31433 13553 31467
rect 13553 31433 13587 31467
rect 13587 31433 13596 31467
rect 13544 31424 13596 31433
rect 10600 31331 10652 31340
rect 10600 31297 10609 31331
rect 10609 31297 10643 31331
rect 10643 31297 10652 31331
rect 10600 31288 10652 31297
rect 13452 31220 13504 31272
rect 2872 31084 2924 31136
rect 3332 31127 3384 31136
rect 3332 31093 3341 31127
rect 3341 31093 3375 31127
rect 3375 31093 3384 31127
rect 3332 31084 3384 31093
rect 3516 31084 3568 31136
rect 4896 31127 4948 31136
rect 4896 31093 4905 31127
rect 4905 31093 4939 31127
rect 4939 31093 4948 31127
rect 4896 31084 4948 31093
rect 4988 31127 5040 31136
rect 4988 31093 4997 31127
rect 4997 31093 5031 31127
rect 5031 31093 5040 31127
rect 6644 31127 6696 31136
rect 4988 31084 5040 31093
rect 6644 31093 6653 31127
rect 6653 31093 6687 31127
rect 6687 31093 6696 31127
rect 6644 31084 6696 31093
rect 7288 31127 7340 31136
rect 7288 31093 7297 31127
rect 7297 31093 7331 31127
rect 7331 31093 7340 31127
rect 7288 31084 7340 31093
rect 7380 31127 7432 31136
rect 7380 31093 7389 31127
rect 7389 31093 7423 31127
rect 7423 31093 7432 31127
rect 7380 31084 7432 31093
rect 7748 31084 7800 31136
rect 8484 31084 8536 31136
rect 9772 31084 9824 31136
rect 10508 31127 10560 31136
rect 10508 31093 10517 31127
rect 10517 31093 10551 31127
rect 10551 31093 10560 31127
rect 10508 31084 10560 31093
rect 6315 30982 6367 31034
rect 6379 30982 6431 31034
rect 6443 30982 6495 31034
rect 6507 30982 6559 31034
rect 11648 30982 11700 31034
rect 11712 30982 11764 31034
rect 11776 30982 11828 31034
rect 11840 30982 11892 31034
rect 3332 30880 3384 30932
rect 6828 30923 6880 30932
rect 6828 30889 6837 30923
rect 6837 30889 6871 30923
rect 6871 30889 6880 30923
rect 6828 30880 6880 30889
rect 7564 30923 7616 30932
rect 7564 30889 7573 30923
rect 7573 30889 7607 30923
rect 7607 30889 7616 30923
rect 7564 30880 7616 30889
rect 8576 30923 8628 30932
rect 8576 30889 8585 30923
rect 8585 30889 8619 30923
rect 8619 30889 8628 30923
rect 8576 30880 8628 30889
rect 10048 30880 10100 30932
rect 10600 30880 10652 30932
rect 12440 30880 12492 30932
rect 3240 30812 3292 30864
rect 4896 30812 4948 30864
rect 12072 30812 12124 30864
rect 4436 30787 4488 30796
rect 4436 30753 4445 30787
rect 4445 30753 4479 30787
rect 4479 30753 4488 30787
rect 4436 30744 4488 30753
rect 6184 30744 6236 30796
rect 7104 30744 7156 30796
rect 11060 30744 11112 30796
rect 11612 30787 11664 30796
rect 11612 30753 11621 30787
rect 11621 30753 11655 30787
rect 11655 30753 11664 30787
rect 11612 30744 11664 30753
rect 4160 30676 4212 30728
rect 4528 30719 4580 30728
rect 4528 30685 4537 30719
rect 4537 30685 4571 30719
rect 4571 30685 4580 30719
rect 4528 30676 4580 30685
rect 4712 30719 4764 30728
rect 4712 30685 4721 30719
rect 4721 30685 4755 30719
rect 4755 30685 4764 30719
rect 5080 30719 5132 30728
rect 4712 30676 4764 30685
rect 5080 30685 5089 30719
rect 5089 30685 5123 30719
rect 5123 30685 5132 30719
rect 5080 30676 5132 30685
rect 6828 30676 6880 30728
rect 7288 30608 7340 30660
rect 6920 30540 6972 30592
rect 9772 30540 9824 30592
rect 10508 30540 10560 30592
rect 3648 30438 3700 30490
rect 3712 30438 3764 30490
rect 3776 30438 3828 30490
rect 3840 30438 3892 30490
rect 8982 30438 9034 30490
rect 9046 30438 9098 30490
rect 9110 30438 9162 30490
rect 9174 30438 9226 30490
rect 14315 30438 14367 30490
rect 14379 30438 14431 30490
rect 14443 30438 14495 30490
rect 14507 30438 14559 30490
rect 3976 30336 4028 30388
rect 4712 30336 4764 30388
rect 6828 30336 6880 30388
rect 11612 30379 11664 30388
rect 11612 30345 11621 30379
rect 11621 30345 11655 30379
rect 11655 30345 11664 30379
rect 11612 30336 11664 30345
rect 12072 30379 12124 30388
rect 12072 30345 12081 30379
rect 12081 30345 12115 30379
rect 12115 30345 12124 30379
rect 12072 30336 12124 30345
rect 4436 30268 4488 30320
rect 4068 30200 4120 30252
rect 4804 30200 4856 30252
rect 6920 30200 6972 30252
rect 7472 30243 7524 30252
rect 5816 30132 5868 30184
rect 7472 30209 7481 30243
rect 7481 30209 7515 30243
rect 7515 30209 7524 30243
rect 7472 30200 7524 30209
rect 10232 30243 10284 30252
rect 10232 30209 10241 30243
rect 10241 30209 10275 30243
rect 10275 30209 10284 30243
rect 10232 30200 10284 30209
rect 4160 30064 4212 30116
rect 6184 30107 6236 30116
rect 6184 30073 6193 30107
rect 6193 30073 6227 30107
rect 6227 30073 6236 30107
rect 6184 30064 6236 30073
rect 8116 30132 8168 30184
rect 9956 30132 10008 30184
rect 8852 30064 8904 30116
rect 5080 30039 5132 30048
rect 5080 30005 5089 30039
rect 5089 30005 5123 30039
rect 5123 30005 5132 30039
rect 5080 29996 5132 30005
rect 6828 30039 6880 30048
rect 6828 30005 6837 30039
rect 6837 30005 6871 30039
rect 6871 30005 6880 30039
rect 6828 29996 6880 30005
rect 7196 30039 7248 30048
rect 7196 30005 7205 30039
rect 7205 30005 7239 30039
rect 7239 30005 7248 30039
rect 7196 29996 7248 30005
rect 9680 30039 9732 30048
rect 9680 30005 9689 30039
rect 9689 30005 9723 30039
rect 9723 30005 9732 30039
rect 9680 29996 9732 30005
rect 6315 29894 6367 29946
rect 6379 29894 6431 29946
rect 6443 29894 6495 29946
rect 6507 29894 6559 29946
rect 11648 29894 11700 29946
rect 11712 29894 11764 29946
rect 11776 29894 11828 29946
rect 11840 29894 11892 29946
rect 1584 29835 1636 29844
rect 1584 29801 1593 29835
rect 1593 29801 1627 29835
rect 1627 29801 1636 29835
rect 1584 29792 1636 29801
rect 4528 29792 4580 29844
rect 5724 29835 5776 29844
rect 5724 29801 5733 29835
rect 5733 29801 5767 29835
rect 5767 29801 5776 29835
rect 5724 29792 5776 29801
rect 6736 29792 6788 29844
rect 7288 29792 7340 29844
rect 8024 29792 8076 29844
rect 10232 29792 10284 29844
rect 4160 29724 4212 29776
rect 7472 29724 7524 29776
rect 2320 29656 2372 29708
rect 6828 29656 6880 29708
rect 8024 29699 8076 29708
rect 8024 29665 8033 29699
rect 8033 29665 8067 29699
rect 8067 29665 8076 29699
rect 8024 29656 8076 29665
rect 5816 29631 5868 29640
rect 5816 29597 5825 29631
rect 5825 29597 5859 29631
rect 5859 29597 5868 29631
rect 5816 29588 5868 29597
rect 5264 29495 5316 29504
rect 5264 29461 5273 29495
rect 5273 29461 5307 29495
rect 5307 29461 5316 29495
rect 5264 29452 5316 29461
rect 8208 29631 8260 29640
rect 8208 29597 8217 29631
rect 8217 29597 8251 29631
rect 8251 29597 8260 29631
rect 10968 29724 11020 29776
rect 11060 29656 11112 29708
rect 8208 29588 8260 29597
rect 9588 29452 9640 29504
rect 10232 29452 10284 29504
rect 3648 29350 3700 29402
rect 3712 29350 3764 29402
rect 3776 29350 3828 29402
rect 3840 29350 3892 29402
rect 8982 29350 9034 29402
rect 9046 29350 9098 29402
rect 9110 29350 9162 29402
rect 9174 29350 9226 29402
rect 14315 29350 14367 29402
rect 14379 29350 14431 29402
rect 14443 29350 14495 29402
rect 14507 29350 14559 29402
rect 1584 29291 1636 29300
rect 1584 29257 1593 29291
rect 1593 29257 1627 29291
rect 1627 29257 1636 29291
rect 1584 29248 1636 29257
rect 2688 29248 2740 29300
rect 4068 29291 4120 29300
rect 4068 29257 4077 29291
rect 4077 29257 4111 29291
rect 4111 29257 4120 29291
rect 4068 29248 4120 29257
rect 4528 29248 4580 29300
rect 5724 29248 5776 29300
rect 6828 29248 6880 29300
rect 10968 29248 11020 29300
rect 8116 29180 8168 29232
rect 5080 29112 5132 29164
rect 5816 29112 5868 29164
rect 9036 29112 9088 29164
rect 9680 29112 9732 29164
rect 10048 29155 10100 29164
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 10232 29155 10284 29164
rect 10232 29121 10241 29155
rect 10241 29121 10275 29155
rect 10275 29121 10284 29155
rect 10232 29112 10284 29121
rect 7288 29087 7340 29096
rect 7288 29053 7297 29087
rect 7297 29053 7331 29087
rect 7331 29053 7340 29087
rect 7288 29044 7340 29053
rect 7840 29044 7892 29096
rect 11152 29044 11204 29096
rect 2320 29019 2372 29028
rect 2320 28985 2329 29019
rect 2329 28985 2363 29019
rect 2363 28985 2372 29019
rect 2320 28976 2372 28985
rect 6000 28976 6052 29028
rect 7012 28976 7064 29028
rect 8024 28976 8076 29028
rect 8576 28976 8628 29028
rect 11980 28976 12032 29028
rect 4252 28908 4304 28960
rect 5172 28908 5224 28960
rect 5356 28908 5408 28960
rect 9036 28951 9088 28960
rect 9036 28917 9045 28951
rect 9045 28917 9079 28951
rect 9079 28917 9088 28951
rect 9036 28908 9088 28917
rect 9588 28951 9640 28960
rect 9588 28917 9597 28951
rect 9597 28917 9631 28951
rect 9631 28917 9640 28951
rect 9588 28908 9640 28917
rect 11060 28951 11112 28960
rect 11060 28917 11069 28951
rect 11069 28917 11103 28951
rect 11103 28917 11112 28951
rect 11060 28908 11112 28917
rect 12532 28908 12584 28960
rect 6315 28806 6367 28858
rect 6379 28806 6431 28858
rect 6443 28806 6495 28858
rect 6507 28806 6559 28858
rect 11648 28806 11700 28858
rect 11712 28806 11764 28858
rect 11776 28806 11828 28858
rect 11840 28806 11892 28858
rect 2412 28747 2464 28756
rect 2412 28713 2421 28747
rect 2421 28713 2455 28747
rect 2455 28713 2464 28747
rect 2412 28704 2464 28713
rect 4896 28747 4948 28756
rect 4896 28713 4905 28747
rect 4905 28713 4939 28747
rect 4939 28713 4948 28747
rect 4896 28704 4948 28713
rect 10048 28704 10100 28756
rect 1676 28636 1728 28688
rect 2596 28636 2648 28688
rect 6092 28636 6144 28688
rect 12348 28636 12400 28688
rect 7288 28568 7340 28620
rect 10232 28568 10284 28620
rect 2872 28543 2924 28552
rect 2872 28509 2881 28543
rect 2881 28509 2915 28543
rect 2915 28509 2924 28543
rect 2872 28500 2924 28509
rect 2964 28500 3016 28552
rect 5080 28500 5132 28552
rect 5356 28543 5408 28552
rect 5356 28509 5365 28543
rect 5365 28509 5399 28543
rect 5399 28509 5408 28543
rect 5356 28500 5408 28509
rect 5540 28543 5592 28552
rect 5540 28509 5549 28543
rect 5549 28509 5583 28543
rect 5583 28509 5592 28543
rect 5540 28500 5592 28509
rect 6552 28543 6604 28552
rect 6552 28509 6561 28543
rect 6561 28509 6595 28543
rect 6595 28509 6604 28543
rect 6552 28500 6604 28509
rect 10968 28500 11020 28552
rect 8392 28432 8444 28484
rect 9036 28432 9088 28484
rect 12532 28475 12584 28484
rect 12532 28441 12541 28475
rect 12541 28441 12575 28475
rect 12575 28441 12584 28475
rect 12532 28432 12584 28441
rect 4252 28364 4304 28416
rect 8576 28407 8628 28416
rect 8576 28373 8585 28407
rect 8585 28373 8619 28407
rect 8619 28373 8628 28407
rect 8576 28364 8628 28373
rect 10692 28407 10744 28416
rect 10692 28373 10701 28407
rect 10701 28373 10735 28407
rect 10735 28373 10744 28407
rect 10692 28364 10744 28373
rect 3648 28262 3700 28314
rect 3712 28262 3764 28314
rect 3776 28262 3828 28314
rect 3840 28262 3892 28314
rect 8982 28262 9034 28314
rect 9046 28262 9098 28314
rect 9110 28262 9162 28314
rect 9174 28262 9226 28314
rect 14315 28262 14367 28314
rect 14379 28262 14431 28314
rect 14443 28262 14495 28314
rect 14507 28262 14559 28314
rect 2596 28160 2648 28212
rect 2872 28160 2924 28212
rect 5080 28203 5132 28212
rect 5080 28169 5089 28203
rect 5089 28169 5123 28203
rect 5123 28169 5132 28203
rect 5080 28160 5132 28169
rect 5540 28160 5592 28212
rect 7288 28203 7340 28212
rect 7288 28169 7297 28203
rect 7297 28169 7331 28203
rect 7331 28169 7340 28203
rect 7288 28160 7340 28169
rect 9680 28160 9732 28212
rect 12348 28160 12400 28212
rect 2964 28024 3016 28076
rect 10692 28024 10744 28076
rect 8392 27999 8444 28008
rect 8392 27965 8426 27999
rect 8426 27965 8444 27999
rect 2688 27820 2740 27872
rect 3792 27888 3844 27940
rect 5172 27888 5224 27940
rect 6552 27931 6604 27940
rect 6552 27897 6561 27931
rect 6561 27897 6595 27931
rect 6595 27897 6604 27931
rect 7932 27931 7984 27940
rect 6552 27888 6604 27897
rect 7932 27897 7941 27931
rect 7941 27897 7975 27931
rect 7975 27897 7984 27931
rect 8392 27956 8444 27965
rect 10968 27956 11020 28008
rect 7932 27888 7984 27897
rect 10048 27888 10100 27940
rect 4068 27820 4120 27872
rect 6092 27863 6144 27872
rect 6092 27829 6101 27863
rect 6101 27829 6135 27863
rect 6135 27829 6144 27863
rect 6092 27820 6144 27829
rect 6828 27863 6880 27872
rect 6828 27829 6837 27863
rect 6837 27829 6871 27863
rect 6871 27829 6880 27863
rect 6828 27820 6880 27829
rect 8300 27820 8352 27872
rect 10508 27820 10560 27872
rect 11336 27820 11388 27872
rect 6315 27718 6367 27770
rect 6379 27718 6431 27770
rect 6443 27718 6495 27770
rect 6507 27718 6559 27770
rect 11648 27718 11700 27770
rect 11712 27718 11764 27770
rect 11776 27718 11828 27770
rect 11840 27718 11892 27770
rect 3792 27659 3844 27668
rect 3792 27625 3801 27659
rect 3801 27625 3835 27659
rect 3835 27625 3844 27659
rect 3792 27616 3844 27625
rect 5356 27616 5408 27668
rect 7288 27616 7340 27668
rect 8392 27616 8444 27668
rect 10232 27616 10284 27668
rect 10508 27616 10560 27668
rect 11152 27616 11204 27668
rect 12164 27616 12216 27668
rect 2228 27548 2280 27600
rect 5816 27548 5868 27600
rect 2136 27480 2188 27532
rect 2780 27523 2832 27532
rect 2780 27489 2789 27523
rect 2789 27489 2823 27523
rect 2823 27489 2832 27523
rect 2780 27480 2832 27489
rect 8300 27480 8352 27532
rect 8760 27548 8812 27600
rect 9036 27591 9088 27600
rect 9036 27557 9045 27591
rect 9045 27557 9079 27591
rect 9079 27557 9088 27591
rect 9036 27548 9088 27557
rect 11336 27548 11388 27600
rect 3792 27412 3844 27464
rect 4160 27412 4212 27464
rect 5172 27412 5224 27464
rect 7932 27412 7984 27464
rect 2872 27344 2924 27396
rect 8852 27344 8904 27396
rect 8024 27319 8076 27328
rect 8024 27285 8033 27319
rect 8033 27285 8067 27319
rect 8067 27285 8076 27319
rect 8024 27276 8076 27285
rect 8300 27276 8352 27328
rect 8484 27276 8536 27328
rect 9956 27480 10008 27532
rect 10968 27455 11020 27464
rect 10968 27421 10977 27455
rect 10977 27421 11011 27455
rect 11011 27421 11020 27455
rect 10968 27412 11020 27421
rect 9772 27276 9824 27328
rect 10048 27276 10100 27328
rect 12164 27276 12216 27328
rect 12808 27276 12860 27328
rect 3648 27174 3700 27226
rect 3712 27174 3764 27226
rect 3776 27174 3828 27226
rect 3840 27174 3892 27226
rect 8982 27174 9034 27226
rect 9046 27174 9098 27226
rect 9110 27174 9162 27226
rect 9174 27174 9226 27226
rect 14315 27174 14367 27226
rect 14379 27174 14431 27226
rect 14443 27174 14495 27226
rect 14507 27174 14559 27226
rect 3976 27115 4028 27124
rect 3976 27081 3985 27115
rect 3985 27081 4019 27115
rect 4019 27081 4028 27115
rect 3976 27072 4028 27081
rect 5816 27072 5868 27124
rect 6092 27072 6144 27124
rect 9496 27115 9548 27124
rect 2136 27047 2188 27056
rect 2136 27013 2145 27047
rect 2145 27013 2179 27047
rect 2179 27013 2188 27047
rect 2136 27004 2188 27013
rect 2228 27004 2280 27056
rect 6184 27004 6236 27056
rect 9496 27081 9505 27115
rect 9505 27081 9539 27115
rect 9539 27081 9548 27115
rect 9496 27072 9548 27081
rect 8944 26979 8996 26988
rect 8944 26945 8953 26979
rect 8953 26945 8987 26979
rect 8987 26945 8996 26979
rect 8944 26936 8996 26945
rect 2412 26868 2464 26920
rect 2688 26868 2740 26920
rect 6828 26868 6880 26920
rect 7932 26868 7984 26920
rect 8760 26911 8812 26920
rect 8760 26877 8769 26911
rect 8769 26877 8803 26911
rect 8803 26877 8812 26911
rect 8760 26868 8812 26877
rect 2964 26800 3016 26852
rect 6000 26800 6052 26852
rect 6368 26800 6420 26852
rect 7196 26843 7248 26852
rect 7196 26809 7205 26843
rect 7205 26809 7239 26843
rect 7239 26809 7248 26843
rect 9956 27072 10008 27124
rect 10140 27072 10192 27124
rect 10784 27072 10836 27124
rect 11336 27115 11388 27124
rect 11336 27081 11345 27115
rect 11345 27081 11379 27115
rect 11379 27081 11388 27115
rect 11336 27072 11388 27081
rect 9772 27004 9824 27056
rect 10416 27004 10468 27056
rect 10876 26936 10928 26988
rect 12164 26936 12216 26988
rect 9864 26868 9916 26920
rect 10416 26868 10468 26920
rect 7196 26800 7248 26809
rect 5172 26732 5224 26784
rect 12808 26843 12860 26852
rect 12808 26809 12817 26843
rect 12817 26809 12851 26843
rect 12851 26809 12860 26843
rect 12808 26800 12860 26809
rect 9956 26775 10008 26784
rect 9956 26741 9965 26775
rect 9965 26741 9999 26775
rect 9999 26741 10008 26775
rect 9956 26732 10008 26741
rect 10508 26732 10560 26784
rect 10968 26775 11020 26784
rect 10968 26741 10977 26775
rect 10977 26741 11011 26775
rect 11011 26741 11020 26775
rect 10968 26732 11020 26741
rect 11520 26732 11572 26784
rect 12164 26775 12216 26784
rect 12164 26741 12173 26775
rect 12173 26741 12207 26775
rect 12207 26741 12216 26775
rect 12164 26732 12216 26741
rect 12440 26775 12492 26784
rect 12440 26741 12449 26775
rect 12449 26741 12483 26775
rect 12483 26741 12492 26775
rect 12900 26775 12952 26784
rect 12440 26732 12492 26741
rect 12900 26741 12909 26775
rect 12909 26741 12943 26775
rect 12943 26741 12952 26775
rect 12900 26732 12952 26741
rect 6315 26630 6367 26682
rect 6379 26630 6431 26682
rect 6443 26630 6495 26682
rect 6507 26630 6559 26682
rect 11648 26630 11700 26682
rect 11712 26630 11764 26682
rect 11776 26630 11828 26682
rect 11840 26630 11892 26682
rect 2964 26571 3016 26580
rect 2964 26537 2973 26571
rect 2973 26537 3007 26571
rect 3007 26537 3016 26571
rect 2964 26528 3016 26537
rect 6184 26528 6236 26580
rect 7196 26571 7248 26580
rect 7196 26537 7205 26571
rect 7205 26537 7239 26571
rect 7239 26537 7248 26571
rect 7196 26528 7248 26537
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 8024 26528 8076 26580
rect 8300 26528 8352 26580
rect 8944 26528 8996 26580
rect 10324 26571 10376 26580
rect 10324 26537 10333 26571
rect 10333 26537 10367 26571
rect 10367 26537 10376 26571
rect 10324 26528 10376 26537
rect 10692 26528 10744 26580
rect 11520 26528 11572 26580
rect 12900 26528 12952 26580
rect 8116 26503 8168 26512
rect 8116 26469 8125 26503
rect 8125 26469 8159 26503
rect 8159 26469 8168 26503
rect 8116 26460 8168 26469
rect 5448 26435 5500 26444
rect 5448 26401 5482 26435
rect 5482 26401 5500 26435
rect 5448 26392 5500 26401
rect 10692 26435 10744 26444
rect 10692 26401 10701 26435
rect 10701 26401 10735 26435
rect 10735 26401 10744 26435
rect 10692 26392 10744 26401
rect 12164 26435 12216 26444
rect 12164 26401 12198 26435
rect 12198 26401 12216 26435
rect 12164 26392 12216 26401
rect 5172 26367 5224 26376
rect 5172 26333 5181 26367
rect 5181 26333 5215 26367
rect 5215 26333 5224 26367
rect 5172 26324 5224 26333
rect 7932 26324 7984 26376
rect 8208 26324 8260 26376
rect 9864 26324 9916 26376
rect 10508 26324 10560 26376
rect 10876 26367 10928 26376
rect 10876 26333 10885 26367
rect 10885 26333 10919 26367
rect 10919 26333 10928 26367
rect 10876 26324 10928 26333
rect 11888 26367 11940 26376
rect 11888 26333 11897 26367
rect 11897 26333 11931 26367
rect 11931 26333 11940 26367
rect 11888 26324 11940 26333
rect 2412 26256 2464 26308
rect 8484 26256 8536 26308
rect 9496 26256 9548 26308
rect 13268 26299 13320 26308
rect 13268 26265 13277 26299
rect 13277 26265 13311 26299
rect 13311 26265 13320 26299
rect 13268 26256 13320 26265
rect 3648 26086 3700 26138
rect 3712 26086 3764 26138
rect 3776 26086 3828 26138
rect 3840 26086 3892 26138
rect 8982 26086 9034 26138
rect 9046 26086 9098 26138
rect 9110 26086 9162 26138
rect 9174 26086 9226 26138
rect 14315 26086 14367 26138
rect 14379 26086 14431 26138
rect 14443 26086 14495 26138
rect 14507 26086 14559 26138
rect 6828 26027 6880 26036
rect 6828 25993 6837 26027
rect 6837 25993 6871 26027
rect 6871 25993 6880 26027
rect 6828 25984 6880 25993
rect 7932 26027 7984 26036
rect 7932 25993 7941 26027
rect 7941 25993 7975 26027
rect 7975 25993 7984 26027
rect 7932 25984 7984 25993
rect 8300 26027 8352 26036
rect 8300 25993 8309 26027
rect 8309 25993 8343 26027
rect 8343 25993 8352 26027
rect 8300 25984 8352 25993
rect 10600 26027 10652 26036
rect 10600 25993 10609 26027
rect 10609 25993 10643 26027
rect 10643 25993 10652 26027
rect 10600 25984 10652 25993
rect 10692 25984 10744 26036
rect 5540 25848 5592 25900
rect 7472 25891 7524 25900
rect 7472 25857 7481 25891
rect 7481 25857 7515 25891
rect 7515 25857 7524 25891
rect 7472 25848 7524 25857
rect 8300 25848 8352 25900
rect 12164 25916 12216 25968
rect 8668 25780 8720 25832
rect 9956 25780 10008 25832
rect 11888 25823 11940 25832
rect 10968 25712 11020 25764
rect 11888 25789 11897 25823
rect 11897 25789 11931 25823
rect 11931 25789 11940 25823
rect 11888 25780 11940 25789
rect 5172 25687 5224 25696
rect 5172 25653 5181 25687
rect 5181 25653 5215 25687
rect 5215 25653 5224 25687
rect 5172 25644 5224 25653
rect 7288 25687 7340 25696
rect 7288 25653 7297 25687
rect 7297 25653 7331 25687
rect 7331 25653 7340 25687
rect 9496 25687 9548 25696
rect 7288 25644 7340 25653
rect 9496 25653 9505 25687
rect 9505 25653 9539 25687
rect 9539 25653 9548 25687
rect 9496 25644 9548 25653
rect 9588 25644 9640 25696
rect 6315 25542 6367 25594
rect 6379 25542 6431 25594
rect 6443 25542 6495 25594
rect 6507 25542 6559 25594
rect 11648 25542 11700 25594
rect 11712 25542 11764 25594
rect 11776 25542 11828 25594
rect 11840 25542 11892 25594
rect 1584 25483 1636 25492
rect 1584 25449 1593 25483
rect 1593 25449 1627 25483
rect 1627 25449 1636 25483
rect 1584 25440 1636 25449
rect 7288 25440 7340 25492
rect 9956 25440 10008 25492
rect 10876 25440 10928 25492
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 11060 25304 11112 25356
rect 4528 25279 4580 25288
rect 4528 25245 4537 25279
rect 4537 25245 4571 25279
rect 4571 25245 4580 25279
rect 4528 25236 4580 25245
rect 9496 25236 9548 25288
rect 10324 25279 10376 25288
rect 10324 25245 10333 25279
rect 10333 25245 10367 25279
rect 10367 25245 10376 25279
rect 10324 25236 10376 25245
rect 10600 25236 10652 25288
rect 10784 25236 10836 25288
rect 9680 25211 9732 25220
rect 9680 25177 9689 25211
rect 9689 25177 9723 25211
rect 9723 25177 9732 25211
rect 9680 25168 9732 25177
rect 8208 25100 8260 25152
rect 10232 25100 10284 25152
rect 10508 25100 10560 25152
rect 3648 24998 3700 25050
rect 3712 24998 3764 25050
rect 3776 24998 3828 25050
rect 3840 24998 3892 25050
rect 8982 24998 9034 25050
rect 9046 24998 9098 25050
rect 9110 24998 9162 25050
rect 9174 24998 9226 25050
rect 14315 24998 14367 25050
rect 14379 24998 14431 25050
rect 14443 24998 14495 25050
rect 14507 24998 14559 25050
rect 9496 24896 9548 24948
rect 10324 24896 10376 24948
rect 4896 24803 4948 24812
rect 4896 24769 4905 24803
rect 4905 24769 4939 24803
rect 4939 24769 4948 24803
rect 4896 24760 4948 24769
rect 4988 24760 5040 24812
rect 8024 24760 8076 24812
rect 9312 24803 9364 24812
rect 9312 24769 9321 24803
rect 9321 24769 9355 24803
rect 9355 24769 9364 24803
rect 9312 24760 9364 24769
rect 11520 24828 11572 24880
rect 10232 24760 10284 24812
rect 10876 24760 10928 24812
rect 11060 24760 11112 24812
rect 12348 24760 12400 24812
rect 4528 24692 4580 24744
rect 7656 24692 7708 24744
rect 8760 24692 8812 24744
rect 8852 24692 8904 24744
rect 2228 24667 2280 24676
rect 2228 24633 2262 24667
rect 2262 24633 2280 24667
rect 2228 24624 2280 24633
rect 2412 24556 2464 24608
rect 2964 24556 3016 24608
rect 4436 24599 4488 24608
rect 4436 24565 4445 24599
rect 4445 24565 4479 24599
rect 4479 24565 4488 24599
rect 4436 24556 4488 24565
rect 7932 24599 7984 24608
rect 7932 24565 7941 24599
rect 7941 24565 7975 24599
rect 7975 24565 7984 24599
rect 7932 24556 7984 24565
rect 8208 24556 8260 24608
rect 8484 24556 8536 24608
rect 10140 24556 10192 24608
rect 6315 24454 6367 24506
rect 6379 24454 6431 24506
rect 6443 24454 6495 24506
rect 6507 24454 6559 24506
rect 11648 24454 11700 24506
rect 11712 24454 11764 24506
rect 11776 24454 11828 24506
rect 11840 24454 11892 24506
rect 1400 24352 1452 24404
rect 2688 24395 2740 24404
rect 2688 24361 2697 24395
rect 2697 24361 2731 24395
rect 2731 24361 2740 24395
rect 2688 24352 2740 24361
rect 7932 24352 7984 24404
rect 9864 24352 9916 24404
rect 10876 24352 10928 24404
rect 7564 24327 7616 24336
rect 7564 24293 7573 24327
rect 7573 24293 7607 24327
rect 7607 24293 7616 24327
rect 7564 24284 7616 24293
rect 4068 24216 4120 24268
rect 4436 24259 4488 24268
rect 4436 24225 4445 24259
rect 4445 24225 4479 24259
rect 4479 24225 4488 24259
rect 4436 24216 4488 24225
rect 9680 24216 9732 24268
rect 10324 24216 10376 24268
rect 11520 24259 11572 24268
rect 11520 24225 11554 24259
rect 11554 24225 11572 24259
rect 11520 24216 11572 24225
rect 2412 24148 2464 24200
rect 2964 24191 3016 24200
rect 2964 24157 2973 24191
rect 2973 24157 3007 24191
rect 3007 24157 3016 24191
rect 2964 24148 3016 24157
rect 4528 24191 4580 24200
rect 4528 24157 4537 24191
rect 4537 24157 4571 24191
rect 4571 24157 4580 24191
rect 4528 24148 4580 24157
rect 4712 24191 4764 24200
rect 4712 24157 4721 24191
rect 4721 24157 4755 24191
rect 4755 24157 4764 24191
rect 4712 24148 4764 24157
rect 7932 24148 7984 24200
rect 10232 24191 10284 24200
rect 10232 24157 10241 24191
rect 10241 24157 10275 24191
rect 10275 24157 10284 24191
rect 10232 24148 10284 24157
rect 10968 24148 11020 24200
rect 2228 24012 2280 24064
rect 3516 24012 3568 24064
rect 4436 24012 4488 24064
rect 4896 24012 4948 24064
rect 5540 24012 5592 24064
rect 7196 24055 7248 24064
rect 7196 24021 7205 24055
rect 7205 24021 7239 24055
rect 7239 24021 7248 24055
rect 7196 24012 7248 24021
rect 9680 24055 9732 24064
rect 9680 24021 9689 24055
rect 9689 24021 9723 24055
rect 9723 24021 9732 24055
rect 9680 24012 9732 24021
rect 12440 24012 12492 24064
rect 3648 23910 3700 23962
rect 3712 23910 3764 23962
rect 3776 23910 3828 23962
rect 3840 23910 3892 23962
rect 8982 23910 9034 23962
rect 9046 23910 9098 23962
rect 9110 23910 9162 23962
rect 9174 23910 9226 23962
rect 14315 23910 14367 23962
rect 14379 23910 14431 23962
rect 14443 23910 14495 23962
rect 14507 23910 14559 23962
rect 2964 23808 3016 23860
rect 4160 23808 4212 23860
rect 4712 23808 4764 23860
rect 7932 23808 7984 23860
rect 9864 23808 9916 23860
rect 10140 23808 10192 23860
rect 10232 23808 10284 23860
rect 11060 23808 11112 23860
rect 4528 23740 4580 23792
rect 6736 23740 6788 23792
rect 7564 23740 7616 23792
rect 3240 23672 3292 23724
rect 4988 23715 5040 23724
rect 4988 23681 4997 23715
rect 4997 23681 5031 23715
rect 5031 23681 5040 23715
rect 4988 23672 5040 23681
rect 4896 23604 4948 23656
rect 5080 23604 5132 23656
rect 2596 23536 2648 23588
rect 4804 23579 4856 23588
rect 4804 23545 4813 23579
rect 4813 23545 4847 23579
rect 4847 23545 4856 23579
rect 4804 23536 4856 23545
rect 2780 23511 2832 23520
rect 2780 23477 2789 23511
rect 2789 23477 2823 23511
rect 2823 23477 2832 23511
rect 3148 23511 3200 23520
rect 2780 23468 2832 23477
rect 3148 23477 3157 23511
rect 3157 23477 3191 23511
rect 3191 23477 3200 23511
rect 3148 23468 3200 23477
rect 3516 23468 3568 23520
rect 4252 23468 4304 23520
rect 4528 23468 4580 23520
rect 6920 23468 6972 23520
rect 8024 23647 8076 23656
rect 8024 23613 8058 23647
rect 8058 23613 8076 23647
rect 8024 23604 8076 23613
rect 8208 23468 8260 23520
rect 10324 23468 10376 23520
rect 10968 23468 11020 23520
rect 11520 23468 11572 23520
rect 12348 23468 12400 23520
rect 6315 23366 6367 23418
rect 6379 23366 6431 23418
rect 6443 23366 6495 23418
rect 6507 23366 6559 23418
rect 11648 23366 11700 23418
rect 11712 23366 11764 23418
rect 11776 23366 11828 23418
rect 11840 23366 11892 23418
rect 1584 23307 1636 23316
rect 1584 23273 1593 23307
rect 1593 23273 1627 23307
rect 1627 23273 1636 23307
rect 1584 23264 1636 23273
rect 2412 23307 2464 23316
rect 2412 23273 2421 23307
rect 2421 23273 2455 23307
rect 2455 23273 2464 23307
rect 2412 23264 2464 23273
rect 4068 23264 4120 23316
rect 4804 23264 4856 23316
rect 5448 23264 5500 23316
rect 2688 23196 2740 23248
rect 2872 23196 2924 23248
rect 4988 23196 5040 23248
rect 5724 23196 5776 23248
rect 7196 23264 7248 23316
rect 11060 23307 11112 23316
rect 11060 23273 11069 23307
rect 11069 23273 11103 23307
rect 11103 23273 11112 23307
rect 11060 23264 11112 23273
rect 12624 23307 12676 23316
rect 12624 23273 12633 23307
rect 12633 23273 12667 23307
rect 12667 23273 12676 23307
rect 12624 23264 12676 23273
rect 13084 23264 13136 23316
rect 8024 23239 8076 23248
rect 8024 23205 8033 23239
rect 8033 23205 8067 23239
rect 8067 23205 8076 23239
rect 8024 23196 8076 23205
rect 1676 23128 1728 23180
rect 4804 23171 4856 23180
rect 4804 23137 4838 23171
rect 4838 23137 4856 23171
rect 4804 23128 4856 23137
rect 9588 23128 9640 23180
rect 10968 23196 11020 23248
rect 12256 23196 12308 23248
rect 12716 23196 12768 23248
rect 10232 23128 10284 23180
rect 10876 23128 10928 23180
rect 12348 23128 12400 23180
rect 2780 23060 2832 23112
rect 2964 23060 3016 23112
rect 2228 22992 2280 23044
rect 4068 23060 4120 23112
rect 7472 23103 7524 23112
rect 7472 23069 7481 23103
rect 7481 23069 7515 23103
rect 7515 23069 7524 23103
rect 7472 23060 7524 23069
rect 6920 23035 6972 23044
rect 6920 23001 6929 23035
rect 6929 23001 6963 23035
rect 6963 23001 6972 23035
rect 11796 23060 11848 23112
rect 12624 23060 12676 23112
rect 6920 22992 6972 23001
rect 4712 22924 4764 22976
rect 5172 22924 5224 22976
rect 12164 22967 12216 22976
rect 12164 22933 12173 22967
rect 12173 22933 12207 22967
rect 12207 22933 12216 22967
rect 12164 22924 12216 22933
rect 13268 22967 13320 22976
rect 13268 22933 13277 22967
rect 13277 22933 13311 22967
rect 13311 22933 13320 22967
rect 13268 22924 13320 22933
rect 3648 22822 3700 22874
rect 3712 22822 3764 22874
rect 3776 22822 3828 22874
rect 3840 22822 3892 22874
rect 8982 22822 9034 22874
rect 9046 22822 9098 22874
rect 9110 22822 9162 22874
rect 9174 22822 9226 22874
rect 14315 22822 14367 22874
rect 14379 22822 14431 22874
rect 14443 22822 14495 22874
rect 14507 22822 14559 22874
rect 2964 22720 3016 22772
rect 4068 22763 4120 22772
rect 4068 22729 4077 22763
rect 4077 22729 4111 22763
rect 4111 22729 4120 22763
rect 4068 22720 4120 22729
rect 2228 22695 2280 22704
rect 2228 22661 2237 22695
rect 2237 22661 2271 22695
rect 2271 22661 2280 22695
rect 2228 22652 2280 22661
rect 2504 22695 2556 22704
rect 2504 22661 2513 22695
rect 2513 22661 2547 22695
rect 2547 22661 2556 22695
rect 2504 22652 2556 22661
rect 5264 22652 5316 22704
rect 8300 22720 8352 22772
rect 10876 22763 10928 22772
rect 5356 22584 5408 22636
rect 5724 22584 5776 22636
rect 10876 22729 10885 22763
rect 10885 22729 10919 22763
rect 10919 22729 10928 22763
rect 10876 22720 10928 22729
rect 11796 22695 11848 22704
rect 11796 22661 11805 22695
rect 11805 22661 11839 22695
rect 11839 22661 11848 22695
rect 11796 22652 11848 22661
rect 12532 22584 12584 22636
rect 3240 22516 3292 22568
rect 5540 22559 5592 22568
rect 5540 22525 5549 22559
rect 5549 22525 5583 22559
rect 5583 22525 5592 22559
rect 5540 22516 5592 22525
rect 6828 22559 6880 22568
rect 4804 22448 4856 22500
rect 6184 22491 6236 22500
rect 6184 22457 6193 22491
rect 6193 22457 6227 22491
rect 6227 22457 6236 22491
rect 6184 22448 6236 22457
rect 4712 22423 4764 22432
rect 4712 22389 4721 22423
rect 4721 22389 4755 22423
rect 4755 22389 4764 22423
rect 4712 22380 4764 22389
rect 5172 22423 5224 22432
rect 5172 22389 5181 22423
rect 5181 22389 5215 22423
rect 5215 22389 5224 22423
rect 5172 22380 5224 22389
rect 5724 22380 5776 22432
rect 6828 22525 6837 22559
rect 6837 22525 6871 22559
rect 6871 22525 6880 22559
rect 6828 22516 6880 22525
rect 6920 22516 6972 22568
rect 7104 22559 7156 22568
rect 7104 22525 7127 22559
rect 7127 22525 7156 22559
rect 7104 22516 7156 22525
rect 12716 22516 12768 22568
rect 12992 22584 13044 22636
rect 13268 22584 13320 22636
rect 13636 22516 13688 22568
rect 9864 22448 9916 22500
rect 12808 22491 12860 22500
rect 12808 22457 12817 22491
rect 12817 22457 12851 22491
rect 12851 22457 12860 22491
rect 12808 22448 12860 22457
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 12440 22380 12492 22389
rect 6315 22278 6367 22330
rect 6379 22278 6431 22330
rect 6443 22278 6495 22330
rect 6507 22278 6559 22330
rect 11648 22278 11700 22330
rect 11712 22278 11764 22330
rect 11776 22278 11828 22330
rect 11840 22278 11892 22330
rect 1676 22219 1728 22228
rect 1676 22185 1685 22219
rect 1685 22185 1719 22219
rect 1719 22185 1728 22219
rect 1676 22176 1728 22185
rect 3240 22219 3292 22228
rect 3240 22185 3249 22219
rect 3249 22185 3283 22219
rect 3283 22185 3292 22219
rect 3240 22176 3292 22185
rect 4804 22219 4856 22228
rect 4804 22185 4813 22219
rect 4813 22185 4847 22219
rect 4847 22185 4856 22219
rect 4804 22176 4856 22185
rect 6184 22176 6236 22228
rect 7472 22176 7524 22228
rect 12808 22219 12860 22228
rect 5264 22151 5316 22160
rect 5264 22117 5298 22151
rect 5298 22117 5316 22151
rect 5264 22108 5316 22117
rect 12808 22185 12817 22219
rect 12817 22185 12851 22219
rect 12851 22185 12860 22219
rect 12808 22176 12860 22185
rect 2872 22040 2924 22092
rect 4712 22040 4764 22092
rect 5724 22040 5776 22092
rect 7932 22083 7984 22092
rect 7932 22049 7941 22083
rect 7941 22049 7975 22083
rect 7975 22049 7984 22083
rect 7932 22040 7984 22049
rect 12164 22108 12216 22160
rect 12440 22040 12492 22092
rect 8024 22015 8076 22024
rect 8024 21981 8033 22015
rect 8033 21981 8067 22015
rect 8067 21981 8076 22015
rect 8024 21972 8076 21981
rect 7840 21904 7892 21956
rect 10048 21972 10100 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10600 21972 10652 22024
rect 10784 21972 10836 22024
rect 11336 21972 11388 22024
rect 12348 21972 12400 22024
rect 9864 21904 9916 21956
rect 5356 21836 5408 21888
rect 7104 21879 7156 21888
rect 7104 21845 7113 21879
rect 7113 21845 7147 21879
rect 7147 21845 7156 21879
rect 7104 21836 7156 21845
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 10784 21879 10836 21888
rect 10784 21845 10793 21879
rect 10793 21845 10827 21879
rect 10827 21845 10836 21879
rect 10784 21836 10836 21845
rect 12532 21879 12584 21888
rect 12532 21845 12541 21879
rect 12541 21845 12575 21879
rect 12575 21845 12584 21879
rect 12532 21836 12584 21845
rect 3648 21734 3700 21786
rect 3712 21734 3764 21786
rect 3776 21734 3828 21786
rect 3840 21734 3892 21786
rect 8982 21734 9034 21786
rect 9046 21734 9098 21786
rect 9110 21734 9162 21786
rect 9174 21734 9226 21786
rect 14315 21734 14367 21786
rect 14379 21734 14431 21786
rect 14443 21734 14495 21786
rect 14507 21734 14559 21786
rect 1584 21675 1636 21684
rect 1584 21641 1593 21675
rect 1593 21641 1627 21675
rect 1627 21641 1636 21675
rect 1584 21632 1636 21641
rect 2872 21632 2924 21684
rect 3516 21632 3568 21684
rect 7840 21632 7892 21684
rect 10232 21632 10284 21684
rect 11336 21675 11388 21684
rect 11336 21641 11345 21675
rect 11345 21641 11379 21675
rect 11379 21641 11388 21675
rect 11336 21632 11388 21641
rect 12440 21675 12492 21684
rect 12440 21641 12449 21675
rect 12449 21641 12483 21675
rect 12483 21641 12492 21675
rect 12440 21632 12492 21641
rect 7932 21564 7984 21616
rect 3240 21496 3292 21548
rect 4804 21496 4856 21548
rect 8116 21496 8168 21548
rect 9864 21496 9916 21548
rect 12624 21496 12676 21548
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 4068 21428 4120 21480
rect 4712 21428 4764 21480
rect 10784 21428 10836 21480
rect 11244 21428 11296 21480
rect 13084 21428 13136 21480
rect 1952 21403 2004 21412
rect 1952 21369 1961 21403
rect 1961 21369 1995 21403
rect 1995 21369 2004 21403
rect 1952 21360 2004 21369
rect 3424 21292 3476 21344
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 5356 21292 5408 21344
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 7656 21292 7708 21344
rect 7932 21292 7984 21344
rect 9312 21360 9364 21412
rect 8392 21292 8444 21344
rect 8576 21335 8628 21344
rect 8576 21301 8585 21335
rect 8585 21301 8619 21335
rect 8619 21301 8628 21335
rect 8576 21292 8628 21301
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 11520 21292 11572 21344
rect 6315 21190 6367 21242
rect 6379 21190 6431 21242
rect 6443 21190 6495 21242
rect 6507 21190 6559 21242
rect 11648 21190 11700 21242
rect 11712 21190 11764 21242
rect 11776 21190 11828 21242
rect 11840 21190 11892 21242
rect 5264 21088 5316 21140
rect 10048 21088 10100 21140
rect 10508 21088 10560 21140
rect 10784 21088 10836 21140
rect 11520 21088 11572 21140
rect 12164 21131 12216 21140
rect 12164 21097 12173 21131
rect 12173 21097 12207 21131
rect 12207 21097 12216 21131
rect 12164 21088 12216 21097
rect 7104 21020 7156 21072
rect 7748 21020 7800 21072
rect 11428 21063 11480 21072
rect 11428 21029 11437 21063
rect 11437 21029 11471 21063
rect 11471 21029 11480 21063
rect 11428 21020 11480 21029
rect 7012 20952 7064 21004
rect 7196 20952 7248 21004
rect 9864 20952 9916 21004
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 6828 20884 6880 20936
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 7840 20884 7892 20936
rect 11612 20927 11664 20936
rect 11612 20893 11621 20927
rect 11621 20893 11655 20927
rect 11655 20893 11664 20927
rect 11612 20884 11664 20893
rect 6920 20816 6972 20868
rect 3424 20748 3476 20800
rect 4068 20748 4120 20800
rect 5080 20748 5132 20800
rect 7104 20791 7156 20800
rect 7104 20757 7113 20791
rect 7113 20757 7147 20791
rect 7147 20757 7156 20791
rect 7104 20748 7156 20757
rect 8392 20748 8444 20800
rect 9404 20748 9456 20800
rect 12624 20748 12676 20800
rect 3648 20646 3700 20698
rect 3712 20646 3764 20698
rect 3776 20646 3828 20698
rect 3840 20646 3892 20698
rect 8982 20646 9034 20698
rect 9046 20646 9098 20698
rect 9110 20646 9162 20698
rect 9174 20646 9226 20698
rect 14315 20646 14367 20698
rect 14379 20646 14431 20698
rect 14443 20646 14495 20698
rect 14507 20646 14559 20698
rect 5540 20544 5592 20596
rect 9312 20544 9364 20596
rect 6644 20476 6696 20528
rect 7840 20476 7892 20528
rect 9404 20476 9456 20528
rect 7104 20408 7156 20460
rect 3976 20340 4028 20392
rect 6920 20340 6972 20392
rect 7748 20408 7800 20460
rect 9588 20451 9640 20460
rect 9588 20417 9597 20451
rect 9597 20417 9631 20451
rect 9631 20417 9640 20451
rect 9588 20408 9640 20417
rect 9404 20383 9456 20392
rect 9404 20349 9413 20383
rect 9413 20349 9447 20383
rect 9447 20349 9456 20383
rect 9404 20340 9456 20349
rect 11612 20408 11664 20460
rect 10784 20340 10836 20392
rect 7012 20272 7064 20324
rect 10508 20272 10560 20324
rect 3608 20204 3660 20256
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4160 20247 4212 20256
rect 4160 20213 4169 20247
rect 4169 20213 4203 20247
rect 4203 20213 4212 20247
rect 4160 20204 4212 20213
rect 6184 20204 6236 20256
rect 6828 20204 6880 20256
rect 7196 20204 7248 20256
rect 9496 20247 9548 20256
rect 9496 20213 9505 20247
rect 9505 20213 9539 20247
rect 9539 20213 9548 20247
rect 9496 20204 9548 20213
rect 10232 20204 10284 20256
rect 11520 20204 11572 20256
rect 6315 20102 6367 20154
rect 6379 20102 6431 20154
rect 6443 20102 6495 20154
rect 6507 20102 6559 20154
rect 11648 20102 11700 20154
rect 11712 20102 11764 20154
rect 11776 20102 11828 20154
rect 11840 20102 11892 20154
rect 4160 20000 4212 20052
rect 4896 20043 4948 20052
rect 4896 20009 4905 20043
rect 4905 20009 4939 20043
rect 4939 20009 4948 20043
rect 4896 20000 4948 20009
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 9496 20000 9548 20052
rect 10048 20000 10100 20052
rect 10692 20000 10744 20052
rect 11152 20043 11204 20052
rect 11152 20009 11161 20043
rect 11161 20009 11195 20043
rect 11195 20009 11204 20043
rect 11152 20000 11204 20009
rect 11428 20000 11480 20052
rect 12624 20000 12676 20052
rect 6644 19975 6696 19984
rect 6644 19941 6678 19975
rect 6678 19941 6696 19975
rect 6644 19932 6696 19941
rect 10416 19932 10468 19984
rect 5816 19864 5868 19916
rect 9956 19864 10008 19916
rect 11796 19907 11848 19916
rect 11796 19873 11830 19907
rect 11830 19873 11848 19907
rect 11796 19864 11848 19873
rect 4712 19796 4764 19848
rect 10416 19839 10468 19848
rect 4528 19728 4580 19780
rect 10416 19805 10425 19839
rect 10425 19805 10459 19839
rect 10459 19805 10468 19839
rect 10416 19796 10468 19805
rect 10508 19839 10560 19848
rect 10508 19805 10517 19839
rect 10517 19805 10551 19839
rect 10551 19805 10560 19839
rect 10508 19796 10560 19805
rect 10968 19796 11020 19848
rect 11428 19796 11480 19848
rect 3648 19558 3700 19610
rect 3712 19558 3764 19610
rect 3776 19558 3828 19610
rect 3840 19558 3892 19610
rect 8982 19558 9034 19610
rect 9046 19558 9098 19610
rect 9110 19558 9162 19610
rect 9174 19558 9226 19610
rect 14315 19558 14367 19610
rect 14379 19558 14431 19610
rect 14443 19558 14495 19610
rect 14507 19558 14559 19610
rect 6644 19456 6696 19508
rect 6920 19456 6972 19508
rect 10508 19499 10560 19508
rect 10508 19465 10517 19499
rect 10517 19465 10551 19499
rect 10551 19465 10560 19499
rect 10508 19456 10560 19465
rect 11796 19456 11848 19508
rect 4620 19320 4672 19372
rect 4988 19320 5040 19372
rect 5632 19320 5684 19372
rect 5724 19320 5776 19372
rect 7840 19363 7892 19372
rect 7840 19329 7849 19363
rect 7849 19329 7883 19363
rect 7883 19329 7892 19363
rect 7840 19320 7892 19329
rect 10784 19320 10836 19372
rect 11152 19320 11204 19372
rect 11428 19320 11480 19372
rect 11980 19320 12032 19372
rect 12072 19320 12124 19372
rect 13360 19320 13412 19372
rect 13452 19320 13504 19372
rect 7012 19252 7064 19304
rect 8208 19252 8260 19304
rect 8392 19252 8444 19304
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 2964 19184 3016 19236
rect 3976 19184 4028 19236
rect 4620 19184 4672 19236
rect 4712 19184 4764 19236
rect 5724 19184 5776 19236
rect 8116 19184 8168 19236
rect 9312 19184 9364 19236
rect 4896 19159 4948 19168
rect 4896 19125 4905 19159
rect 4905 19125 4939 19159
rect 4939 19125 4948 19159
rect 4896 19116 4948 19125
rect 5264 19116 5316 19168
rect 7104 19159 7156 19168
rect 7104 19125 7113 19159
rect 7113 19125 7147 19159
rect 7147 19125 7156 19159
rect 7656 19159 7708 19168
rect 7104 19116 7156 19125
rect 7656 19125 7665 19159
rect 7665 19125 7699 19159
rect 7699 19125 7708 19159
rect 7656 19116 7708 19125
rect 8392 19116 8444 19168
rect 8760 19116 8812 19168
rect 9496 19116 9548 19168
rect 6315 19014 6367 19066
rect 6379 19014 6431 19066
rect 6443 19014 6495 19066
rect 6507 19014 6559 19066
rect 11648 19014 11700 19066
rect 11712 19014 11764 19066
rect 11776 19014 11828 19066
rect 11840 19014 11892 19066
rect 3976 18912 4028 18964
rect 4896 18912 4948 18964
rect 7012 18912 7064 18964
rect 7840 18912 7892 18964
rect 5724 18844 5776 18896
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 5540 18776 5592 18828
rect 8392 18819 8444 18828
rect 8392 18785 8401 18819
rect 8401 18785 8435 18819
rect 8435 18785 8444 18819
rect 8392 18776 8444 18785
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 8576 18751 8628 18760
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 9956 18708 10008 18760
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 4528 18615 4580 18624
rect 2964 18572 3016 18581
rect 4528 18581 4537 18615
rect 4537 18581 4571 18615
rect 4571 18581 4580 18615
rect 4528 18572 4580 18581
rect 6276 18615 6328 18624
rect 6276 18581 6285 18615
rect 6285 18581 6319 18615
rect 6319 18581 6328 18615
rect 6276 18572 6328 18581
rect 8024 18615 8076 18624
rect 8024 18581 8033 18615
rect 8033 18581 8067 18615
rect 8067 18581 8076 18615
rect 8024 18572 8076 18581
rect 9312 18572 9364 18624
rect 10416 18572 10468 18624
rect 3648 18470 3700 18522
rect 3712 18470 3764 18522
rect 3776 18470 3828 18522
rect 3840 18470 3892 18522
rect 8982 18470 9034 18522
rect 9046 18470 9098 18522
rect 9110 18470 9162 18522
rect 9174 18470 9226 18522
rect 14315 18470 14367 18522
rect 14379 18470 14431 18522
rect 14443 18470 14495 18522
rect 14507 18470 14559 18522
rect 1584 18411 1636 18420
rect 1584 18377 1593 18411
rect 1593 18377 1627 18411
rect 1627 18377 1636 18411
rect 1584 18368 1636 18377
rect 4160 18368 4212 18420
rect 4896 18300 4948 18352
rect 4528 18232 4580 18284
rect 6276 18232 6328 18284
rect 5264 18164 5316 18216
rect 8116 18164 8168 18216
rect 8576 18164 8628 18216
rect 9220 18096 9272 18148
rect 1952 18071 2004 18080
rect 1952 18037 1961 18071
rect 1961 18037 1995 18071
rect 1995 18037 2004 18071
rect 1952 18028 2004 18037
rect 4436 18028 4488 18080
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 5540 18028 5592 18080
rect 8576 18028 8628 18080
rect 9312 18028 9364 18080
rect 6315 17926 6367 17978
rect 6379 17926 6431 17978
rect 6443 17926 6495 17978
rect 6507 17926 6559 17978
rect 11648 17926 11700 17978
rect 11712 17926 11764 17978
rect 11776 17926 11828 17978
rect 11840 17926 11892 17978
rect 4068 17824 4120 17876
rect 5172 17824 5224 17876
rect 7748 17867 7800 17876
rect 7748 17833 7757 17867
rect 7757 17833 7791 17867
rect 7791 17833 7800 17867
rect 7748 17824 7800 17833
rect 8024 17824 8076 17876
rect 8116 17731 8168 17740
rect 8116 17697 8125 17731
rect 8125 17697 8159 17731
rect 8159 17697 8168 17731
rect 8116 17688 8168 17697
rect 9772 17688 9824 17740
rect 11428 17688 11480 17740
rect 12164 17688 12216 17740
rect 4252 17620 4304 17672
rect 5540 17663 5592 17672
rect 5540 17629 5549 17663
rect 5549 17629 5583 17663
rect 5583 17629 5592 17663
rect 5540 17620 5592 17629
rect 7932 17620 7984 17672
rect 8576 17620 8628 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 2780 17552 2832 17604
rect 8484 17552 8536 17604
rect 3424 17484 3476 17536
rect 6920 17527 6972 17536
rect 6920 17493 6929 17527
rect 6929 17493 6963 17527
rect 6963 17493 6972 17527
rect 6920 17484 6972 17493
rect 7380 17484 7432 17536
rect 8576 17484 8628 17536
rect 10692 17527 10744 17536
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 12992 17527 13044 17536
rect 12992 17493 13001 17527
rect 13001 17493 13035 17527
rect 13035 17493 13044 17527
rect 12992 17484 13044 17493
rect 3648 17382 3700 17434
rect 3712 17382 3764 17434
rect 3776 17382 3828 17434
rect 3840 17382 3892 17434
rect 8982 17382 9034 17434
rect 9046 17382 9098 17434
rect 9110 17382 9162 17434
rect 9174 17382 9226 17434
rect 14315 17382 14367 17434
rect 14379 17382 14431 17434
rect 14443 17382 14495 17434
rect 14507 17382 14559 17434
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 4252 17280 4304 17332
rect 7932 17323 7984 17332
rect 7932 17289 7941 17323
rect 7941 17289 7975 17323
rect 7975 17289 7984 17323
rect 7932 17280 7984 17289
rect 8392 17280 8444 17332
rect 10140 17323 10192 17332
rect 10140 17289 10149 17323
rect 10149 17289 10183 17323
rect 10183 17289 10192 17323
rect 10140 17280 10192 17289
rect 11428 17280 11480 17332
rect 2688 17212 2740 17264
rect 5908 17212 5960 17264
rect 6092 17212 6144 17264
rect 10048 17255 10100 17264
rect 10048 17221 10057 17255
rect 10057 17221 10091 17255
rect 10091 17221 10100 17255
rect 10048 17212 10100 17221
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 5540 17187 5592 17196
rect 5540 17153 5549 17187
rect 5549 17153 5583 17187
rect 5583 17153 5592 17187
rect 5540 17144 5592 17153
rect 6920 17144 6972 17196
rect 4068 17076 4120 17128
rect 5356 17119 5408 17128
rect 5356 17085 5365 17119
rect 5365 17085 5399 17119
rect 5399 17085 5408 17119
rect 5356 17076 5408 17085
rect 5448 17076 5500 17128
rect 7656 17144 7708 17196
rect 8576 17144 8628 17196
rect 9128 17187 9180 17196
rect 9128 17153 9137 17187
rect 9137 17153 9171 17187
rect 9171 17153 9180 17187
rect 9128 17144 9180 17153
rect 9680 17144 9732 17196
rect 10692 17187 10744 17196
rect 10692 17153 10701 17187
rect 10701 17153 10735 17187
rect 10735 17153 10744 17187
rect 10692 17144 10744 17153
rect 10048 17076 10100 17128
rect 3516 17008 3568 17060
rect 5080 17008 5132 17060
rect 9956 17008 10008 17060
rect 10324 17008 10376 17060
rect 4896 16983 4948 16992
rect 4896 16949 4905 16983
rect 4905 16949 4939 16983
rect 4939 16949 4948 16983
rect 4896 16940 4948 16949
rect 6644 16940 6696 16992
rect 7380 16940 7432 16992
rect 8944 16983 8996 16992
rect 8944 16949 8953 16983
rect 8953 16949 8987 16983
rect 8987 16949 8996 16983
rect 8944 16940 8996 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9680 16983 9732 16992
rect 9036 16940 9088 16949
rect 9680 16949 9689 16983
rect 9689 16949 9723 16983
rect 9723 16949 9732 16983
rect 9680 16940 9732 16949
rect 12164 16940 12216 16992
rect 6315 16838 6367 16890
rect 6379 16838 6431 16890
rect 6443 16838 6495 16890
rect 6507 16838 6559 16890
rect 11648 16838 11700 16890
rect 11712 16838 11764 16890
rect 11776 16838 11828 16890
rect 11840 16838 11892 16890
rect 2412 16779 2464 16788
rect 2412 16745 2421 16779
rect 2421 16745 2455 16779
rect 2455 16745 2464 16779
rect 2412 16736 2464 16745
rect 2596 16736 2648 16788
rect 2780 16779 2832 16788
rect 2780 16745 2789 16779
rect 2789 16745 2823 16779
rect 2823 16745 2832 16779
rect 2780 16736 2832 16745
rect 3424 16736 3476 16788
rect 4528 16779 4580 16788
rect 4528 16745 4537 16779
rect 4537 16745 4571 16779
rect 4571 16745 4580 16779
rect 4528 16736 4580 16745
rect 5080 16779 5132 16788
rect 5080 16745 5089 16779
rect 5089 16745 5123 16779
rect 5123 16745 5132 16779
rect 5080 16736 5132 16745
rect 7656 16779 7708 16788
rect 7656 16745 7665 16779
rect 7665 16745 7699 16779
rect 7699 16745 7708 16779
rect 7656 16736 7708 16745
rect 8024 16736 8076 16788
rect 10140 16736 10192 16788
rect 10692 16736 10744 16788
rect 2044 16532 2096 16584
rect 4896 16668 4948 16720
rect 7288 16668 7340 16720
rect 7932 16668 7984 16720
rect 8944 16668 8996 16720
rect 9588 16668 9640 16720
rect 9680 16668 9732 16720
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 6184 16600 6236 16652
rect 8208 16600 8260 16652
rect 9036 16600 9088 16652
rect 9128 16600 9180 16652
rect 11428 16668 11480 16720
rect 10508 16643 10560 16652
rect 10508 16609 10542 16643
rect 10542 16609 10560 16643
rect 2964 16532 3016 16584
rect 3516 16532 3568 16584
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 6276 16575 6328 16584
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 8024 16532 8076 16584
rect 10508 16600 10560 16609
rect 10048 16396 10100 16448
rect 3648 16294 3700 16346
rect 3712 16294 3764 16346
rect 3776 16294 3828 16346
rect 3840 16294 3892 16346
rect 8982 16294 9034 16346
rect 9046 16294 9098 16346
rect 9110 16294 9162 16346
rect 9174 16294 9226 16346
rect 14315 16294 14367 16346
rect 14379 16294 14431 16346
rect 14443 16294 14495 16346
rect 14507 16294 14559 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 4160 16192 4212 16244
rect 6828 16235 6880 16244
rect 6828 16201 6837 16235
rect 6837 16201 6871 16235
rect 6871 16201 6880 16235
rect 6828 16192 6880 16201
rect 7288 16099 7340 16108
rect 7288 16065 7297 16099
rect 7297 16065 7331 16099
rect 7331 16065 7340 16099
rect 7288 16056 7340 16065
rect 7564 16056 7616 16108
rect 8484 16056 8536 16108
rect 9680 16192 9732 16244
rect 10048 16192 10100 16244
rect 11428 16192 11480 16244
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 6184 15988 6236 16040
rect 6276 16031 6328 16040
rect 6276 15997 6285 16031
rect 6285 15997 6319 16031
rect 6319 15997 6328 16031
rect 6276 15988 6328 15997
rect 6828 15988 6880 16040
rect 6920 15988 6972 16040
rect 7748 15988 7800 16040
rect 2964 15920 3016 15972
rect 4620 15920 4672 15972
rect 5356 15920 5408 15972
rect 9496 15920 9548 15972
rect 3516 15852 3568 15904
rect 8116 15852 8168 15904
rect 8392 15852 8444 15904
rect 6315 15750 6367 15802
rect 6379 15750 6431 15802
rect 6443 15750 6495 15802
rect 6507 15750 6559 15802
rect 11648 15750 11700 15802
rect 11712 15750 11764 15802
rect 11776 15750 11828 15802
rect 11840 15750 11892 15802
rect 1400 15648 1452 15700
rect 2596 15648 2648 15700
rect 2964 15691 3016 15700
rect 2964 15657 2973 15691
rect 2973 15657 3007 15691
rect 3007 15657 3016 15691
rect 2964 15648 3016 15657
rect 4068 15648 4120 15700
rect 4436 15648 4488 15700
rect 6920 15691 6972 15700
rect 6920 15657 6929 15691
rect 6929 15657 6963 15691
rect 6963 15657 6972 15691
rect 6920 15648 6972 15657
rect 7380 15691 7432 15700
rect 7380 15657 7389 15691
rect 7389 15657 7423 15691
rect 7423 15657 7432 15691
rect 7380 15648 7432 15657
rect 9496 15648 9548 15700
rect 9864 15691 9916 15700
rect 9864 15657 9873 15691
rect 9873 15657 9907 15691
rect 9907 15657 9916 15691
rect 9864 15648 9916 15657
rect 10508 15648 10560 15700
rect 13176 15648 13228 15700
rect 4528 15580 4580 15632
rect 11060 15580 11112 15632
rect 4160 15512 4212 15564
rect 5540 15512 5592 15564
rect 7104 15512 7156 15564
rect 8024 15512 8076 15564
rect 9680 15512 9732 15564
rect 11980 15580 12032 15632
rect 4896 15487 4948 15496
rect 4896 15453 4905 15487
rect 4905 15453 4939 15487
rect 4939 15453 4948 15487
rect 4896 15444 4948 15453
rect 7840 15487 7892 15496
rect 7840 15453 7849 15487
rect 7849 15453 7883 15487
rect 7883 15453 7892 15487
rect 7840 15444 7892 15453
rect 10324 15487 10376 15496
rect 6184 15308 6236 15360
rect 7564 15376 7616 15428
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 10508 15487 10560 15496
rect 10508 15453 10517 15487
rect 10517 15453 10551 15487
rect 10551 15453 10560 15487
rect 10508 15444 10560 15453
rect 12348 15512 12400 15564
rect 11704 15444 11756 15496
rect 12164 15444 12216 15496
rect 3648 15206 3700 15258
rect 3712 15206 3764 15258
rect 3776 15206 3828 15258
rect 3840 15206 3892 15258
rect 8982 15206 9034 15258
rect 9046 15206 9098 15258
rect 9110 15206 9162 15258
rect 9174 15206 9226 15258
rect 14315 15206 14367 15258
rect 14379 15206 14431 15258
rect 14443 15206 14495 15258
rect 14507 15206 14559 15258
rect 2688 15104 2740 15156
rect 4068 15147 4120 15156
rect 4068 15113 4077 15147
rect 4077 15113 4111 15147
rect 4111 15113 4120 15147
rect 4068 15104 4120 15113
rect 4620 15104 4672 15156
rect 4896 15104 4948 15156
rect 5356 15104 5408 15156
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 10968 15104 11020 15156
rect 10508 15036 10560 15088
rect 3516 14968 3568 15020
rect 12164 14968 12216 15020
rect 4436 14943 4488 14952
rect 4436 14909 4445 14943
rect 4445 14909 4479 14943
rect 4479 14909 4488 14943
rect 4436 14900 4488 14909
rect 6828 14900 6880 14952
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 6184 14764 6236 14816
rect 7104 14807 7156 14816
rect 7104 14773 7113 14807
rect 7113 14773 7147 14807
rect 7147 14773 7156 14807
rect 7104 14764 7156 14773
rect 7748 14764 7800 14816
rect 8484 14900 8536 14952
rect 10232 14900 10284 14952
rect 10784 14900 10836 14952
rect 12900 14943 12952 14952
rect 12900 14909 12909 14943
rect 12909 14909 12943 14943
rect 12943 14909 12952 14943
rect 12900 14900 12952 14909
rect 13176 14900 13228 14952
rect 8116 14875 8168 14884
rect 8116 14841 8150 14875
rect 8150 14841 8168 14875
rect 8116 14832 8168 14841
rect 8576 14832 8628 14884
rect 8024 14764 8076 14816
rect 9312 14764 9364 14816
rect 10784 14764 10836 14816
rect 11704 14832 11756 14884
rect 12716 14832 12768 14884
rect 14004 14832 14056 14884
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 12164 14764 12216 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 6315 14662 6367 14714
rect 6379 14662 6431 14714
rect 6443 14662 6495 14714
rect 6507 14662 6559 14714
rect 11648 14662 11700 14714
rect 11712 14662 11764 14714
rect 11776 14662 11828 14714
rect 11840 14662 11892 14714
rect 4528 14560 4580 14612
rect 5080 14560 5132 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 9588 14560 9640 14612
rect 10324 14560 10376 14612
rect 11980 14560 12032 14612
rect 12440 14560 12492 14612
rect 4896 14424 4948 14476
rect 5356 14492 5408 14544
rect 7288 14492 7340 14544
rect 7840 14492 7892 14544
rect 6920 14424 6972 14476
rect 7380 14467 7432 14476
rect 7380 14433 7389 14467
rect 7389 14433 7423 14467
rect 7423 14433 7432 14467
rect 7380 14424 7432 14433
rect 8760 14424 8812 14476
rect 9588 14424 9640 14476
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 11428 14424 11480 14476
rect 11796 14467 11848 14476
rect 11796 14433 11805 14467
rect 11805 14433 11839 14467
rect 11839 14433 11848 14467
rect 11796 14424 11848 14433
rect 11888 14424 11940 14476
rect 12164 14492 12216 14544
rect 5448 14356 5500 14408
rect 7564 14399 7616 14408
rect 7564 14365 7573 14399
rect 7573 14365 7607 14399
rect 7607 14365 7616 14399
rect 7564 14356 7616 14365
rect 10416 14356 10468 14408
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 7288 14288 7340 14340
rect 7564 14220 7616 14272
rect 8116 14220 8168 14272
rect 8852 14263 8904 14272
rect 8852 14229 8861 14263
rect 8861 14229 8895 14263
rect 8895 14229 8904 14263
rect 8852 14220 8904 14229
rect 10784 14220 10836 14272
rect 3648 14118 3700 14170
rect 3712 14118 3764 14170
rect 3776 14118 3828 14170
rect 3840 14118 3892 14170
rect 8982 14118 9034 14170
rect 9046 14118 9098 14170
rect 9110 14118 9162 14170
rect 9174 14118 9226 14170
rect 14315 14118 14367 14170
rect 14379 14118 14431 14170
rect 14443 14118 14495 14170
rect 14507 14118 14559 14170
rect 5080 14016 5132 14068
rect 5356 14016 5408 14068
rect 6184 14059 6236 14068
rect 6184 14025 6193 14059
rect 6193 14025 6227 14059
rect 6227 14025 6236 14059
rect 6184 14016 6236 14025
rect 6736 14016 6788 14068
rect 7840 14059 7892 14068
rect 7840 14025 7849 14059
rect 7849 14025 7883 14059
rect 7883 14025 7892 14059
rect 7840 14016 7892 14025
rect 8392 14059 8444 14068
rect 8392 14025 8401 14059
rect 8401 14025 8435 14059
rect 8435 14025 8444 14059
rect 8392 14016 8444 14025
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 10416 14059 10468 14068
rect 10416 14025 10425 14059
rect 10425 14025 10459 14059
rect 10459 14025 10468 14059
rect 10416 14016 10468 14025
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 11980 14016 12032 14068
rect 4896 13880 4948 13932
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 7564 13880 7616 13932
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9312 13948 9364 14000
rect 10784 13948 10836 14000
rect 12348 14016 12400 14068
rect 12532 13948 12584 14000
rect 11888 13880 11940 13932
rect 12164 13880 12216 13932
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 6736 13812 6788 13864
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8024 13744 8076 13796
rect 10232 13812 10284 13864
rect 12532 13812 12584 13864
rect 8208 13676 8260 13728
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 10876 13719 10928 13728
rect 10876 13685 10885 13719
rect 10885 13685 10919 13719
rect 10919 13685 10928 13719
rect 10876 13676 10928 13685
rect 11336 13676 11388 13728
rect 12624 13676 12676 13728
rect 6315 13574 6367 13626
rect 6379 13574 6431 13626
rect 6443 13574 6495 13626
rect 6507 13574 6559 13626
rect 11648 13574 11700 13626
rect 11712 13574 11764 13626
rect 11776 13574 11828 13626
rect 11840 13574 11892 13626
rect 1492 13472 1544 13524
rect 6092 13472 6144 13524
rect 6828 13472 6880 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8668 13472 8720 13524
rect 10600 13472 10652 13524
rect 12072 13472 12124 13524
rect 12624 13515 12676 13524
rect 12624 13481 12633 13515
rect 12633 13481 12667 13515
rect 12667 13481 12676 13515
rect 12624 13472 12676 13481
rect 5816 13404 5868 13456
rect 6644 13404 6696 13456
rect 7380 13404 7432 13456
rect 8760 13404 8812 13456
rect 1676 13336 1728 13388
rect 8852 13336 8904 13388
rect 9956 13336 10008 13388
rect 11980 13336 12032 13388
rect 6460 13311 6512 13320
rect 6460 13277 6469 13311
rect 6469 13277 6503 13311
rect 6503 13277 6512 13311
rect 6460 13268 6512 13277
rect 8116 13268 8168 13320
rect 10324 13268 10376 13320
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 12164 13268 12216 13277
rect 10876 13200 10928 13252
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 6644 13132 6696 13184
rect 6920 13132 6972 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 9312 13132 9364 13184
rect 3648 13030 3700 13082
rect 3712 13030 3764 13082
rect 3776 13030 3828 13082
rect 3840 13030 3892 13082
rect 8982 13030 9034 13082
rect 9046 13030 9098 13082
rect 9110 13030 9162 13082
rect 9174 13030 9226 13082
rect 14315 13030 14367 13082
rect 14379 13030 14431 13082
rect 14443 13030 14495 13082
rect 14507 13030 14559 13082
rect 5724 12928 5776 12980
rect 6460 12928 6512 12980
rect 6828 12928 6880 12980
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8668 12928 8720 12980
rect 8852 12928 8904 12980
rect 10692 12928 10744 12980
rect 12072 12928 12124 12980
rect 12164 12928 12216 12980
rect 5816 12860 5868 12912
rect 11152 12860 11204 12912
rect 11428 12860 11480 12912
rect 11980 12903 12032 12912
rect 11980 12869 11989 12903
rect 11989 12869 12023 12903
rect 12023 12869 12032 12903
rect 11980 12860 12032 12869
rect 12532 12860 12584 12912
rect 6184 12792 6236 12844
rect 8116 12792 8168 12844
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 8760 12792 8812 12844
rect 1676 12699 1728 12708
rect 1676 12665 1685 12699
rect 1685 12665 1719 12699
rect 1719 12665 1728 12699
rect 1676 12656 1728 12665
rect 2688 12724 2740 12776
rect 5816 12724 5868 12776
rect 7472 12724 7524 12776
rect 8392 12724 8444 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 7840 12699 7892 12708
rect 7840 12665 7849 12699
rect 7849 12665 7883 12699
rect 7883 12665 7892 12699
rect 7840 12656 7892 12665
rect 9312 12656 9364 12708
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 4068 12588 4120 12640
rect 7472 12588 7524 12640
rect 7656 12588 7708 12640
rect 10416 12588 10468 12640
rect 6315 12486 6367 12538
rect 6379 12486 6431 12538
rect 6443 12486 6495 12538
rect 6507 12486 6559 12538
rect 11648 12486 11700 12538
rect 11712 12486 11764 12538
rect 11776 12486 11828 12538
rect 11840 12486 11892 12538
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 6092 12427 6144 12436
rect 6092 12393 6101 12427
rect 6101 12393 6135 12427
rect 6135 12393 6144 12427
rect 6092 12384 6144 12393
rect 6184 12384 6236 12436
rect 6828 12384 6880 12436
rect 7656 12384 7708 12436
rect 8116 12427 8168 12436
rect 8116 12393 8125 12427
rect 8125 12393 8159 12427
rect 8159 12393 8168 12427
rect 8116 12384 8168 12393
rect 8392 12384 8444 12436
rect 9956 12384 10008 12436
rect 10324 12384 10376 12436
rect 12164 12384 12216 12436
rect 4068 12316 4120 12368
rect 7012 12316 7064 12368
rect 7196 12316 7248 12368
rect 4620 12248 4672 12300
rect 2504 12180 2556 12232
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 5172 12044 5224 12096
rect 6644 12180 6696 12232
rect 7196 12223 7248 12232
rect 7196 12189 7205 12223
rect 7205 12189 7239 12223
rect 7239 12189 7248 12223
rect 7196 12180 7248 12189
rect 9312 12180 9364 12232
rect 11336 12316 11388 12368
rect 10600 12291 10652 12300
rect 10600 12257 10634 12291
rect 10634 12257 10652 12291
rect 10600 12248 10652 12257
rect 8944 12112 8996 12164
rect 9956 12112 10008 12164
rect 7380 12044 7432 12096
rect 3648 11942 3700 11994
rect 3712 11942 3764 11994
rect 3776 11942 3828 11994
rect 3840 11942 3892 11994
rect 8982 11942 9034 11994
rect 9046 11942 9098 11994
rect 9110 11942 9162 11994
rect 9174 11942 9226 11994
rect 14315 11942 14367 11994
rect 14379 11942 14431 11994
rect 14443 11942 14495 11994
rect 14507 11942 14559 11994
rect 2504 11840 2556 11892
rect 2688 11840 2740 11892
rect 4160 11840 4212 11892
rect 4896 11840 4948 11892
rect 7196 11840 7248 11892
rect 9312 11840 9364 11892
rect 9956 11840 10008 11892
rect 10600 11840 10652 11892
rect 5448 11704 5500 11756
rect 2596 11636 2648 11688
rect 7380 11679 7432 11688
rect 3332 11568 3384 11620
rect 5632 11568 5684 11620
rect 6184 11568 6236 11620
rect 5080 11500 5132 11552
rect 6736 11500 6788 11552
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 7656 11679 7708 11688
rect 7656 11645 7690 11679
rect 7690 11645 7708 11679
rect 7656 11636 7708 11645
rect 6315 11398 6367 11450
rect 6379 11398 6431 11450
rect 6443 11398 6495 11450
rect 6507 11398 6559 11450
rect 11648 11398 11700 11450
rect 11712 11398 11764 11450
rect 11776 11398 11828 11450
rect 11840 11398 11892 11450
rect 5080 11339 5132 11348
rect 5080 11305 5089 11339
rect 5089 11305 5123 11339
rect 5123 11305 5132 11339
rect 5080 11296 5132 11305
rect 5172 11339 5224 11348
rect 5172 11305 5181 11339
rect 5181 11305 5215 11339
rect 5215 11305 5224 11339
rect 5172 11296 5224 11305
rect 5356 11296 5408 11348
rect 6644 11339 6696 11348
rect 6644 11305 6653 11339
rect 6653 11305 6687 11339
rect 6687 11305 6696 11339
rect 6644 11296 6696 11305
rect 7656 11296 7708 11348
rect 2964 11228 3016 11280
rect 4620 11271 4672 11280
rect 4620 11237 4629 11271
rect 4629 11237 4663 11271
rect 4663 11237 4672 11271
rect 4620 11228 4672 11237
rect 2504 11160 2556 11212
rect 5172 11160 5224 11212
rect 7564 11228 7616 11280
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 5632 11135 5684 11144
rect 2780 11024 2832 11076
rect 5632 11101 5641 11135
rect 5641 11101 5675 11135
rect 5675 11101 5684 11135
rect 5632 11092 5684 11101
rect 5724 11135 5776 11144
rect 5724 11101 5733 11135
rect 5733 11101 5767 11135
rect 5767 11101 5776 11135
rect 5724 11092 5776 11101
rect 6092 11092 6144 11144
rect 6736 11135 6788 11144
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 5264 11024 5316 11076
rect 1400 10956 1452 11008
rect 3648 10854 3700 10906
rect 3712 10854 3764 10906
rect 3776 10854 3828 10906
rect 3840 10854 3892 10906
rect 8982 10854 9034 10906
rect 9046 10854 9098 10906
rect 9110 10854 9162 10906
rect 9174 10854 9226 10906
rect 14315 10854 14367 10906
rect 14379 10854 14431 10906
rect 14443 10854 14495 10906
rect 14507 10854 14559 10906
rect 2504 10795 2556 10804
rect 2504 10761 2513 10795
rect 2513 10761 2547 10795
rect 2547 10761 2556 10795
rect 2504 10752 2556 10761
rect 2688 10752 2740 10804
rect 2964 10795 3016 10804
rect 2964 10761 2973 10795
rect 2973 10761 3007 10795
rect 3007 10761 3016 10795
rect 2964 10752 3016 10761
rect 3332 10591 3384 10600
rect 3332 10557 3341 10591
rect 3341 10557 3375 10591
rect 3375 10557 3384 10591
rect 3332 10548 3384 10557
rect 5632 10684 5684 10736
rect 3700 10616 3752 10668
rect 5448 10616 5500 10668
rect 6092 10616 6144 10668
rect 7564 10616 7616 10668
rect 4896 10548 4948 10600
rect 2412 10412 2464 10464
rect 3240 10412 3292 10464
rect 5908 10480 5960 10532
rect 7380 10480 7432 10532
rect 5816 10412 5868 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 13360 10412 13412 10464
rect 6315 10310 6367 10362
rect 6379 10310 6431 10362
rect 6443 10310 6495 10362
rect 6507 10310 6559 10362
rect 11648 10310 11700 10362
rect 11712 10310 11764 10362
rect 11776 10310 11828 10362
rect 11840 10310 11892 10362
rect 1584 10251 1636 10260
rect 1584 10217 1593 10251
rect 1593 10217 1627 10251
rect 1627 10217 1636 10251
rect 1584 10208 1636 10217
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 2688 10208 2740 10260
rect 3332 10208 3384 10260
rect 5264 10251 5316 10260
rect 5264 10217 5273 10251
rect 5273 10217 5307 10251
rect 5307 10217 5316 10251
rect 5264 10208 5316 10217
rect 5540 10208 5592 10260
rect 7104 10208 7156 10260
rect 8392 10208 8444 10260
rect 9956 10208 10008 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 2964 10140 3016 10192
rect 5080 10140 5132 10192
rect 5448 10140 5500 10192
rect 5632 10183 5684 10192
rect 5632 10149 5641 10183
rect 5641 10149 5675 10183
rect 5675 10149 5684 10183
rect 5632 10140 5684 10149
rect 7564 10183 7616 10192
rect 7564 10149 7573 10183
rect 7573 10149 7607 10183
rect 7607 10149 7616 10183
rect 7564 10140 7616 10149
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2780 10115 2832 10124
rect 2780 10081 2789 10115
rect 2789 10081 2823 10115
rect 2823 10081 2832 10115
rect 2780 10072 2832 10081
rect 4068 10072 4120 10124
rect 6828 10072 6880 10124
rect 7380 10072 7432 10124
rect 2872 10047 2924 10056
rect 2872 10013 2881 10047
rect 2881 10013 2915 10047
rect 2915 10013 2924 10047
rect 2872 10004 2924 10013
rect 2596 9936 2648 9988
rect 2964 9936 3016 9988
rect 3700 10004 3752 10056
rect 10692 10140 10744 10192
rect 13452 10115 13504 10124
rect 13452 10081 13461 10115
rect 13461 10081 13495 10115
rect 13495 10081 13504 10115
rect 13452 10072 13504 10081
rect 12900 10004 12952 10056
rect 4528 9911 4580 9920
rect 4528 9877 4537 9911
rect 4537 9877 4571 9911
rect 4571 9877 4580 9911
rect 4528 9868 4580 9877
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 10876 9868 10928 9920
rect 11980 9868 12032 9920
rect 12532 9868 12584 9920
rect 12808 9868 12860 9920
rect 3648 9766 3700 9818
rect 3712 9766 3764 9818
rect 3776 9766 3828 9818
rect 3840 9766 3892 9818
rect 8982 9766 9034 9818
rect 9046 9766 9098 9818
rect 9110 9766 9162 9818
rect 9174 9766 9226 9818
rect 14315 9766 14367 9818
rect 14379 9766 14431 9818
rect 14443 9766 14495 9818
rect 14507 9766 14559 9818
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 2964 9664 3016 9716
rect 7104 9707 7156 9716
rect 7104 9673 7113 9707
rect 7113 9673 7147 9707
rect 7147 9673 7156 9707
rect 7104 9664 7156 9673
rect 7564 9664 7616 9716
rect 9864 9664 9916 9716
rect 4068 9596 4120 9648
rect 7012 9596 7064 9648
rect 12900 9664 12952 9716
rect 13360 9664 13412 9716
rect 13452 9639 13504 9648
rect 2964 9528 3016 9580
rect 5080 9571 5132 9580
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 2688 9460 2740 9512
rect 3332 9460 3384 9512
rect 3424 9460 3476 9512
rect 6184 9460 6236 9512
rect 6828 9460 6880 9512
rect 4528 9392 4580 9444
rect 9312 9528 9364 9580
rect 9680 9571 9732 9580
rect 9680 9537 9689 9571
rect 9689 9537 9723 9571
rect 9723 9537 9732 9571
rect 9680 9528 9732 9537
rect 10692 9528 10744 9580
rect 10968 9528 11020 9580
rect 10876 9460 10928 9512
rect 13452 9605 13461 9639
rect 13461 9605 13495 9639
rect 13495 9605 13504 9639
rect 13452 9596 13504 9605
rect 12532 9528 12584 9580
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 7564 9392 7616 9444
rect 11060 9392 11112 9444
rect 3332 9367 3384 9376
rect 3332 9333 3341 9367
rect 3341 9333 3375 9367
rect 3375 9333 3384 9367
rect 3332 9324 3384 9333
rect 6000 9324 6052 9376
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 9220 9367 9272 9376
rect 9220 9333 9229 9367
rect 9229 9333 9263 9367
rect 9263 9333 9272 9367
rect 9220 9324 9272 9333
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 12440 9324 12492 9376
rect 6315 9222 6367 9274
rect 6379 9222 6431 9274
rect 6443 9222 6495 9274
rect 6507 9222 6559 9274
rect 11648 9222 11700 9274
rect 11712 9222 11764 9274
rect 11776 9222 11828 9274
rect 11840 9222 11892 9274
rect 1400 9120 1452 9172
rect 2872 9120 2924 9172
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 5080 9120 5132 9172
rect 8852 9120 8904 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 10140 9163 10192 9172
rect 10140 9129 10149 9163
rect 10149 9129 10183 9163
rect 10183 9129 10192 9163
rect 10140 9120 10192 9129
rect 10232 9120 10284 9172
rect 10784 9120 10836 9172
rect 4252 9052 4304 9104
rect 9864 9052 9916 9104
rect 11980 9095 12032 9104
rect 11980 9061 12014 9095
rect 12014 9061 12032 9095
rect 11980 9052 12032 9061
rect 7380 8984 7432 9036
rect 7748 8984 7800 9036
rect 9956 8984 10008 9036
rect 11704 9027 11756 9036
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 3976 8916 4028 8968
rect 8484 8959 8536 8968
rect 8484 8925 8493 8959
rect 8493 8925 8527 8959
rect 8527 8925 8536 8959
rect 8484 8916 8536 8925
rect 10232 8848 10284 8900
rect 10692 8848 10744 8900
rect 7564 8780 7616 8832
rect 7840 8823 7892 8832
rect 7840 8789 7849 8823
rect 7849 8789 7883 8823
rect 7883 8789 7892 8823
rect 7840 8780 7892 8789
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 10876 8823 10928 8832
rect 10876 8789 10885 8823
rect 10885 8789 10919 8823
rect 10919 8789 10928 8823
rect 10876 8780 10928 8789
rect 11060 8848 11112 8900
rect 12900 8780 12952 8832
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 3648 8678 3700 8730
rect 3712 8678 3764 8730
rect 3776 8678 3828 8730
rect 3840 8678 3892 8730
rect 8982 8678 9034 8730
rect 9046 8678 9098 8730
rect 9110 8678 9162 8730
rect 9174 8678 9226 8730
rect 14315 8678 14367 8730
rect 14379 8678 14431 8730
rect 14443 8678 14495 8730
rect 14507 8678 14559 8730
rect 3332 8619 3384 8628
rect 3332 8585 3341 8619
rect 3341 8585 3375 8619
rect 3375 8585 3384 8619
rect 3332 8576 3384 8585
rect 8668 8576 8720 8628
rect 8852 8576 8904 8628
rect 10692 8576 10744 8628
rect 11336 8576 11388 8628
rect 11980 8576 12032 8628
rect 12440 8619 12492 8628
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 9956 8508 10008 8560
rect 11704 8551 11756 8560
rect 11704 8517 11713 8551
rect 11713 8517 11747 8551
rect 11747 8517 11756 8551
rect 11704 8508 11756 8517
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4252 8440 4304 8492
rect 7840 8483 7892 8492
rect 2688 8304 2740 8356
rect 3976 8304 4028 8356
rect 3700 8279 3752 8288
rect 3700 8245 3709 8279
rect 3709 8245 3743 8279
rect 3743 8245 3752 8279
rect 3700 8236 3752 8245
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 8484 8440 8536 8492
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 6920 8304 6972 8356
rect 7380 8304 7432 8356
rect 4528 8236 4580 8288
rect 4712 8279 4764 8288
rect 4712 8245 4721 8279
rect 4721 8245 4755 8279
rect 4755 8245 4764 8279
rect 4712 8236 4764 8245
rect 7564 8304 7616 8356
rect 8668 8372 8720 8424
rect 12900 8440 12952 8492
rect 9588 8372 9640 8424
rect 11244 8372 11296 8424
rect 13176 8304 13228 8356
rect 8024 8236 8076 8288
rect 12900 8279 12952 8288
rect 12900 8245 12909 8279
rect 12909 8245 12943 8279
rect 12943 8245 12952 8279
rect 12900 8236 12952 8245
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 11648 8134 11700 8186
rect 11712 8134 11764 8186
rect 11776 8134 11828 8186
rect 11840 8134 11892 8186
rect 1768 8032 1820 8084
rect 2688 8032 2740 8084
rect 3424 8075 3476 8084
rect 3424 8041 3433 8075
rect 3433 8041 3467 8075
rect 3467 8041 3476 8075
rect 3424 8032 3476 8041
rect 3700 8032 3752 8084
rect 8760 8032 8812 8084
rect 9588 8032 9640 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 10232 8032 10284 8084
rect 11060 8032 11112 8084
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 12900 8032 12952 8084
rect 4804 7939 4856 7948
rect 4804 7905 4838 7939
rect 4838 7905 4856 7939
rect 4804 7896 4856 7905
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 6828 7828 6880 7880
rect 8668 7964 8720 8016
rect 12808 8007 12860 8016
rect 12808 7973 12817 8007
rect 12817 7973 12851 8007
rect 12851 7973 12860 8007
rect 12808 7964 12860 7973
rect 7288 7939 7340 7948
rect 7288 7905 7322 7939
rect 7322 7905 7340 7939
rect 7288 7896 7340 7905
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 8300 7828 8352 7880
rect 11336 7871 11388 7880
rect 11336 7837 11345 7871
rect 11345 7837 11379 7871
rect 11379 7837 11388 7871
rect 11336 7828 11388 7837
rect 5540 7692 5592 7744
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 7012 7692 7064 7744
rect 7656 7692 7708 7744
rect 3648 7590 3700 7642
rect 3712 7590 3764 7642
rect 3776 7590 3828 7642
rect 3840 7590 3892 7642
rect 8982 7590 9034 7642
rect 9046 7590 9098 7642
rect 9110 7590 9162 7642
rect 9174 7590 9226 7642
rect 14315 7590 14367 7642
rect 14379 7590 14431 7642
rect 14443 7590 14495 7642
rect 14507 7590 14559 7642
rect 3148 7531 3200 7540
rect 3148 7497 3157 7531
rect 3157 7497 3191 7531
rect 3191 7497 3200 7531
rect 3148 7488 3200 7497
rect 7748 7488 7800 7540
rect 1768 7395 1820 7404
rect 1768 7361 1777 7395
rect 1777 7361 1811 7395
rect 1811 7361 1820 7395
rect 1768 7352 1820 7361
rect 4804 7352 4856 7404
rect 5448 7352 5500 7404
rect 6552 7352 6604 7404
rect 7656 7395 7708 7404
rect 7656 7361 7665 7395
rect 7665 7361 7699 7395
rect 7699 7361 7708 7395
rect 7656 7352 7708 7361
rect 6920 7284 6972 7336
rect 7840 7284 7892 7336
rect 11060 7488 11112 7540
rect 14004 7488 14056 7540
rect 15752 7488 15804 7540
rect 10692 7420 10744 7472
rect 11336 7463 11388 7472
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 10784 7395 10836 7404
rect 10784 7361 10793 7395
rect 10793 7361 10827 7395
rect 10827 7361 10836 7395
rect 10784 7352 10836 7361
rect 11336 7429 11345 7463
rect 11345 7429 11379 7463
rect 11379 7429 11388 7463
rect 11336 7420 11388 7429
rect 1492 7148 1544 7200
rect 5264 7216 5316 7268
rect 7288 7216 7340 7268
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 4988 7148 5040 7200
rect 5632 7148 5684 7200
rect 6092 7148 6144 7200
rect 6828 7148 6880 7200
rect 6920 7148 6972 7200
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 10232 7191 10284 7200
rect 10232 7157 10241 7191
rect 10241 7157 10275 7191
rect 10275 7157 10284 7191
rect 10232 7148 10284 7157
rect 11980 7148 12032 7200
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 11648 7046 11700 7098
rect 11712 7046 11764 7098
rect 11776 7046 11828 7098
rect 11840 7046 11892 7098
rect 5264 6944 5316 6996
rect 5632 6944 5684 6996
rect 7288 6944 7340 6996
rect 2320 6808 2372 6860
rect 2504 6808 2556 6860
rect 5724 6851 5776 6860
rect 5724 6817 5758 6851
rect 5758 6817 5776 6851
rect 5724 6808 5776 6817
rect 5080 6740 5132 6792
rect 7840 6944 7892 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8484 6944 8536 6996
rect 10784 6987 10836 6996
rect 10784 6953 10793 6987
rect 10793 6953 10827 6987
rect 10827 6953 10836 6987
rect 10784 6944 10836 6953
rect 11152 6987 11204 6996
rect 11152 6953 11161 6987
rect 11161 6953 11195 6987
rect 11195 6953 11204 6987
rect 11152 6944 11204 6953
rect 10692 6876 10744 6928
rect 8852 6808 8904 6860
rect 9312 6808 9364 6860
rect 12164 6808 12216 6860
rect 12624 6808 12676 6860
rect 13084 6808 13136 6860
rect 9128 6740 9180 6792
rect 9496 6740 9548 6792
rect 2688 6672 2740 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 5448 6604 5500 6656
rect 8852 6604 8904 6656
rect 9956 6604 10008 6656
rect 13452 6647 13504 6656
rect 13452 6613 13461 6647
rect 13461 6613 13495 6647
rect 13495 6613 13504 6647
rect 13452 6604 13504 6613
rect 3648 6502 3700 6554
rect 3712 6502 3764 6554
rect 3776 6502 3828 6554
rect 3840 6502 3892 6554
rect 8982 6502 9034 6554
rect 9046 6502 9098 6554
rect 9110 6502 9162 6554
rect 9174 6502 9226 6554
rect 14315 6502 14367 6554
rect 14379 6502 14431 6554
rect 14443 6502 14495 6554
rect 14507 6502 14559 6554
rect 3424 6400 3476 6452
rect 5724 6400 5776 6452
rect 4160 6332 4212 6384
rect 4528 6332 4580 6384
rect 5080 6332 5132 6384
rect 5632 6332 5684 6384
rect 6092 6332 6144 6384
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5448 6264 5500 6316
rect 7472 6400 7524 6452
rect 8484 6400 8536 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 12164 6443 12216 6452
rect 12164 6409 12173 6443
rect 12173 6409 12207 6443
rect 12207 6409 12216 6443
rect 12164 6400 12216 6409
rect 12624 6443 12676 6452
rect 12624 6409 12633 6443
rect 12633 6409 12667 6443
rect 12667 6409 12676 6443
rect 12624 6400 12676 6409
rect 8484 6264 8536 6316
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 4988 6128 5040 6180
rect 6000 6128 6052 6180
rect 7472 6128 7524 6180
rect 8024 6128 8076 6180
rect 1308 6060 1360 6112
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 6736 6060 6788 6112
rect 7656 6060 7708 6112
rect 8300 6103 8352 6112
rect 8300 6069 8309 6103
rect 8309 6069 8343 6103
rect 8343 6069 8352 6103
rect 8300 6060 8352 6069
rect 8668 6103 8720 6112
rect 8668 6069 8677 6103
rect 8677 6069 8711 6103
rect 8711 6069 8720 6103
rect 8668 6060 8720 6069
rect 9680 6128 9732 6180
rect 10508 6128 10560 6180
rect 8852 6060 8904 6112
rect 9864 6103 9916 6112
rect 9864 6069 9873 6103
rect 9873 6069 9907 6103
rect 9907 6069 9916 6103
rect 9864 6060 9916 6069
rect 10140 6060 10192 6112
rect 10600 6060 10652 6112
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 11648 5958 11700 6010
rect 11712 5958 11764 6010
rect 11776 5958 11828 6010
rect 11840 5958 11892 6010
rect 4528 5856 4580 5908
rect 5724 5856 5776 5908
rect 6644 5856 6696 5908
rect 4896 5788 4948 5840
rect 6000 5788 6052 5840
rect 7012 5788 7064 5840
rect 9680 5788 9732 5840
rect 1400 5763 1452 5772
rect 1400 5729 1409 5763
rect 1409 5729 1443 5763
rect 1443 5729 1452 5763
rect 1400 5720 1452 5729
rect 2872 5763 2924 5772
rect 2872 5729 2881 5763
rect 2881 5729 2915 5763
rect 2915 5729 2924 5763
rect 2872 5720 2924 5729
rect 5264 5720 5316 5772
rect 4988 5652 5040 5704
rect 5448 5652 5500 5704
rect 5632 5652 5684 5704
rect 8024 5720 8076 5772
rect 8576 5720 8628 5772
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 11336 5763 11388 5772
rect 11336 5729 11345 5763
rect 11345 5729 11379 5763
rect 11379 5729 11388 5763
rect 12348 5788 12400 5840
rect 13452 5788 13504 5840
rect 11336 5720 11388 5729
rect 8116 5652 8168 5704
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 7380 5584 7432 5636
rect 9680 5584 9732 5636
rect 940 5516 992 5568
rect 2688 5516 2740 5568
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 3976 5516 4028 5568
rect 4436 5559 4488 5568
rect 4436 5525 4445 5559
rect 4445 5525 4479 5559
rect 4479 5525 4488 5559
rect 4436 5516 4488 5525
rect 5540 5559 5592 5568
rect 5540 5525 5549 5559
rect 5549 5525 5583 5559
rect 5583 5525 5592 5559
rect 5540 5516 5592 5525
rect 7104 5516 7156 5568
rect 7656 5516 7708 5568
rect 8576 5516 8628 5568
rect 11796 5516 11848 5568
rect 12164 5516 12216 5568
rect 13176 5559 13228 5568
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 3648 5414 3700 5466
rect 3712 5414 3764 5466
rect 3776 5414 3828 5466
rect 3840 5414 3892 5466
rect 8982 5414 9034 5466
rect 9046 5414 9098 5466
rect 9110 5414 9162 5466
rect 9174 5414 9226 5466
rect 14315 5414 14367 5466
rect 14379 5414 14431 5466
rect 14443 5414 14495 5466
rect 14507 5414 14559 5466
rect 1400 5312 1452 5364
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 4712 5312 4764 5364
rect 5632 5312 5684 5364
rect 7196 5312 7248 5364
rect 8024 5355 8076 5364
rect 8024 5321 8033 5355
rect 8033 5321 8067 5355
rect 8067 5321 8076 5355
rect 8024 5312 8076 5321
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 10600 5312 10652 5364
rect 11152 5312 11204 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12348 5312 12400 5364
rect 7656 5244 7708 5296
rect 10876 5244 10928 5296
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 3516 5108 3568 5160
rect 4160 5108 4212 5160
rect 5356 5108 5408 5160
rect 7196 5108 7248 5160
rect 10324 5151 10376 5160
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 11428 5108 11480 5160
rect 2412 5083 2464 5092
rect 2412 5049 2421 5083
rect 2421 5049 2455 5083
rect 2455 5049 2464 5083
rect 2412 5040 2464 5049
rect 3424 5040 3476 5092
rect 8392 5083 8444 5092
rect 8392 5049 8426 5083
rect 8426 5049 8444 5083
rect 8392 5040 8444 5049
rect 9312 5040 9364 5092
rect 10876 5040 10928 5092
rect 1400 4972 1452 5024
rect 2964 4972 3016 5024
rect 4896 5015 4948 5024
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 4988 4972 5040 5024
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 6092 4972 6144 5024
rect 7012 5015 7064 5024
rect 7012 4981 7021 5015
rect 7021 4981 7055 5015
rect 7055 4981 7064 5015
rect 7012 4972 7064 4981
rect 12992 4972 13044 5024
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 11648 4870 11700 4922
rect 11712 4870 11764 4922
rect 11776 4870 11828 4922
rect 11840 4870 11892 4922
rect 2504 4768 2556 4820
rect 2688 4768 2740 4820
rect 2780 4768 2832 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 4804 4768 4856 4820
rect 5448 4768 5500 4820
rect 5540 4768 5592 4820
rect 6828 4768 6880 4820
rect 8208 4768 8260 4820
rect 8760 4768 8812 4820
rect 10692 4768 10744 4820
rect 12532 4811 12584 4820
rect 12532 4777 12541 4811
rect 12541 4777 12575 4811
rect 12575 4777 12584 4811
rect 12532 4768 12584 4777
rect 12716 4768 12768 4820
rect 4436 4743 4488 4752
rect 4436 4709 4445 4743
rect 4445 4709 4479 4743
rect 4479 4709 4488 4743
rect 4436 4700 4488 4709
rect 6000 4743 6052 4752
rect 6000 4709 6009 4743
rect 6009 4709 6043 4743
rect 6043 4709 6052 4743
rect 6000 4700 6052 4709
rect 2780 4675 2832 4684
rect 2780 4641 2789 4675
rect 2789 4641 2823 4675
rect 2823 4641 2832 4675
rect 2780 4632 2832 4641
rect 4068 4632 4120 4684
rect 6920 4700 6972 4752
rect 9588 4700 9640 4752
rect 10784 4700 10836 4752
rect 1676 4564 1728 4616
rect 1952 4607 2004 4616
rect 1952 4573 1961 4607
rect 1961 4573 1995 4607
rect 1995 4573 2004 4607
rect 1952 4564 2004 4573
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 8024 4632 8076 4684
rect 9496 4632 9548 4684
rect 10232 4632 10284 4684
rect 11244 4632 11296 4684
rect 6644 4607 6696 4616
rect 2780 4428 2832 4480
rect 3516 4428 3568 4480
rect 6644 4573 6653 4607
rect 6653 4573 6687 4607
rect 6687 4573 6696 4607
rect 6644 4564 6696 4573
rect 5816 4496 5868 4548
rect 8392 4496 8444 4548
rect 9680 4564 9732 4616
rect 10416 4564 10468 4616
rect 10876 4564 10928 4616
rect 11336 4564 11388 4616
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 13176 4700 13228 4752
rect 5632 4428 5684 4480
rect 8116 4428 8168 4480
rect 10232 4428 10284 4480
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 13176 4428 13228 4437
rect 3648 4326 3700 4378
rect 3712 4326 3764 4378
rect 3776 4326 3828 4378
rect 3840 4326 3892 4378
rect 8982 4326 9034 4378
rect 9046 4326 9098 4378
rect 9110 4326 9162 4378
rect 9174 4326 9226 4378
rect 14315 4326 14367 4378
rect 14379 4326 14431 4378
rect 14443 4326 14495 4378
rect 14507 4326 14559 4378
rect 2136 4267 2188 4276
rect 2136 4233 2145 4267
rect 2145 4233 2179 4267
rect 2179 4233 2188 4267
rect 2136 4224 2188 4233
rect 2964 4224 3016 4276
rect 4804 4267 4856 4276
rect 4804 4233 4813 4267
rect 4813 4233 4847 4267
rect 4847 4233 4856 4267
rect 4804 4224 4856 4233
rect 6644 4224 6696 4276
rect 6828 4267 6880 4276
rect 6828 4233 6837 4267
rect 6837 4233 6871 4267
rect 6871 4233 6880 4267
rect 6828 4224 6880 4233
rect 8024 4267 8076 4276
rect 8024 4233 8033 4267
rect 8033 4233 8067 4267
rect 8067 4233 8076 4267
rect 8024 4224 8076 4233
rect 8392 4224 8444 4276
rect 10876 4224 10928 4276
rect 12532 4224 12584 4276
rect 12624 4224 12676 4276
rect 204 4088 256 4140
rect 1308 4088 1360 4140
rect 3884 4088 3936 4140
rect 6000 4156 6052 4208
rect 6552 4199 6604 4208
rect 6552 4165 6561 4199
rect 6561 4165 6595 4199
rect 6595 4165 6604 4199
rect 6552 4156 6604 4165
rect 5632 4131 5684 4140
rect 5632 4097 5641 4131
rect 5641 4097 5675 4131
rect 5675 4097 5684 4131
rect 5632 4088 5684 4097
rect 5724 4088 5776 4140
rect 7012 4156 7064 4208
rect 6920 4088 6972 4140
rect 9128 4131 9180 4140
rect 2136 4020 2188 4072
rect 2688 4020 2740 4072
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 7104 4020 7156 4072
rect 4160 3952 4212 4004
rect 2596 3884 2648 3936
rect 5356 3952 5408 4004
rect 6552 3952 6604 4004
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 10600 4088 10652 4140
rect 11336 4088 11388 4140
rect 12716 4088 12768 4140
rect 9588 4020 9640 4072
rect 10140 4020 10192 4072
rect 11244 4020 11296 4072
rect 12624 4020 12676 4072
rect 13176 4020 13228 4072
rect 10324 3952 10376 4004
rect 8576 3884 8628 3936
rect 9404 3884 9456 3936
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10232 3884 10284 3936
rect 11244 3884 11296 3936
rect 13084 3884 13136 3936
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 11648 3782 11700 3834
rect 11712 3782 11764 3834
rect 11776 3782 11828 3834
rect 11840 3782 11892 3834
rect 2872 3680 2924 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 4160 3680 4212 3732
rect 5356 3680 5408 3732
rect 6920 3680 6972 3732
rect 8208 3680 8260 3732
rect 8760 3723 8812 3732
rect 8760 3689 8769 3723
rect 8769 3689 8803 3723
rect 8803 3689 8812 3723
rect 8760 3680 8812 3689
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 9588 3680 9640 3732
rect 10324 3723 10376 3732
rect 10324 3689 10333 3723
rect 10333 3689 10367 3723
rect 10367 3689 10376 3723
rect 10324 3680 10376 3689
rect 10600 3723 10652 3732
rect 10600 3689 10609 3723
rect 10609 3689 10643 3723
rect 10643 3689 10652 3723
rect 10600 3680 10652 3689
rect 10784 3680 10836 3732
rect 11244 3680 11296 3732
rect 2964 3612 3016 3664
rect 4344 3612 4396 3664
rect 5172 3655 5224 3664
rect 5172 3621 5181 3655
rect 5181 3621 5215 3655
rect 5215 3621 5224 3655
rect 5172 3612 5224 3621
rect 8116 3655 8168 3664
rect 8116 3621 8125 3655
rect 8125 3621 8159 3655
rect 8159 3621 8168 3655
rect 8116 3612 8168 3621
rect 9128 3655 9180 3664
rect 9128 3621 9137 3655
rect 9137 3621 9171 3655
rect 9171 3621 9180 3655
rect 9128 3612 9180 3621
rect 9404 3612 9456 3664
rect 12716 3612 12768 3664
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 6644 3544 6696 3596
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 8024 3544 8076 3596
rect 4252 3476 4304 3528
rect 4804 3476 4856 3528
rect 7656 3476 7708 3528
rect 10784 3544 10836 3596
rect 11152 3587 11204 3596
rect 11152 3553 11161 3587
rect 11161 3553 11195 3587
rect 11195 3553 11204 3587
rect 11152 3544 11204 3553
rect 11244 3544 11296 3596
rect 8760 3476 8812 3528
rect 10232 3476 10284 3528
rect 3516 3408 3568 3460
rect 4988 3408 5040 3460
rect 12716 3408 12768 3460
rect 2136 3340 2188 3392
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 13084 3383 13136 3392
rect 13084 3349 13093 3383
rect 13093 3349 13127 3383
rect 13127 3349 13136 3383
rect 13084 3340 13136 3349
rect 3648 3238 3700 3290
rect 3712 3238 3764 3290
rect 3776 3238 3828 3290
rect 3840 3238 3892 3290
rect 8982 3238 9034 3290
rect 9046 3238 9098 3290
rect 9110 3238 9162 3290
rect 9174 3238 9226 3290
rect 14315 3238 14367 3290
rect 14379 3238 14431 3290
rect 14443 3238 14495 3290
rect 14507 3238 14559 3290
rect 1768 3179 1820 3188
rect 1768 3145 1777 3179
rect 1777 3145 1811 3179
rect 1811 3145 1820 3179
rect 1768 3136 1820 3145
rect 2872 3136 2924 3188
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 6644 3136 6696 3188
rect 7104 3136 7156 3188
rect 9680 3136 9732 3188
rect 10784 3179 10836 3188
rect 10784 3145 10793 3179
rect 10793 3145 10827 3179
rect 10827 3145 10836 3179
rect 10784 3136 10836 3145
rect 11428 3179 11480 3188
rect 11428 3145 11437 3179
rect 11437 3145 11471 3179
rect 11471 3145 11480 3179
rect 11428 3136 11480 3145
rect 12072 3179 12124 3188
rect 12072 3145 12081 3179
rect 12081 3145 12115 3179
rect 12115 3145 12124 3179
rect 12072 3136 12124 3145
rect 13084 3136 13136 3188
rect 2228 3111 2280 3120
rect 2228 3077 2237 3111
rect 2237 3077 2271 3111
rect 2271 3077 2280 3111
rect 2228 3068 2280 3077
rect 3332 3000 3384 3052
rect 4160 3000 4212 3052
rect 7656 3043 7708 3052
rect 7656 3009 7665 3043
rect 7665 3009 7699 3043
rect 7699 3009 7708 3043
rect 7656 3000 7708 3009
rect 8024 3000 8076 3052
rect 13268 3000 13320 3052
rect 3240 2932 3292 2984
rect 4804 2932 4856 2984
rect 7932 2932 7984 2984
rect 5080 2864 5132 2916
rect 9036 2907 9088 2916
rect 9036 2873 9048 2907
rect 9048 2873 9088 2907
rect 9036 2864 9088 2873
rect 3332 2839 3384 2848
rect 3332 2805 3341 2839
rect 3341 2805 3375 2839
rect 3375 2805 3384 2839
rect 3332 2796 3384 2805
rect 12900 2907 12952 2916
rect 12900 2873 12909 2907
rect 12909 2873 12943 2907
rect 12943 2873 12952 2907
rect 12900 2864 12952 2873
rect 9496 2796 9548 2848
rect 14924 2796 14976 2848
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 11648 2694 11700 2746
rect 11712 2694 11764 2746
rect 11776 2694 11828 2746
rect 11840 2694 11892 2746
rect 1952 2635 2004 2644
rect 1952 2601 1961 2635
rect 1961 2601 1995 2635
rect 1995 2601 2004 2635
rect 1952 2592 2004 2601
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 5264 2635 5316 2644
rect 5264 2601 5273 2635
rect 5273 2601 5307 2635
rect 5307 2601 5316 2635
rect 5264 2592 5316 2601
rect 7104 2635 7156 2644
rect 7104 2601 7113 2635
rect 7113 2601 7147 2635
rect 7147 2601 7156 2635
rect 7104 2592 7156 2601
rect 7472 2635 7524 2644
rect 7472 2601 7481 2635
rect 7481 2601 7515 2635
rect 7515 2601 7524 2635
rect 7472 2592 7524 2601
rect 7656 2592 7708 2644
rect 9588 2592 9640 2644
rect 11152 2592 11204 2644
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 12624 2635 12676 2644
rect 12440 2592 12492 2601
rect 12624 2601 12633 2635
rect 12633 2601 12667 2635
rect 12667 2601 12676 2635
rect 12624 2592 12676 2601
rect 4344 2524 4396 2576
rect 4804 2456 4856 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 9404 2524 9456 2576
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9496 2456 9548 2508
rect 12992 2499 13044 2508
rect 12992 2465 13001 2499
rect 13001 2465 13035 2499
rect 13035 2465 13044 2499
rect 12992 2456 13044 2465
rect 9036 2388 9088 2440
rect 13268 2431 13320 2440
rect 2964 2252 3016 2304
rect 5448 2320 5500 2372
rect 7840 2252 7892 2304
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 3648 2150 3700 2202
rect 3712 2150 3764 2202
rect 3776 2150 3828 2202
rect 3840 2150 3892 2202
rect 8982 2150 9034 2202
rect 9046 2150 9098 2202
rect 9110 2150 9162 2202
rect 9174 2150 9226 2202
rect 14315 2150 14367 2202
rect 14379 2150 14431 2202
rect 14443 2150 14495 2202
rect 14507 2150 14559 2202
<< metal2 >>
rect 202 39520 258 40000
rect 570 39520 626 40000
rect 938 39520 994 40000
rect 1398 39520 1454 40000
rect 1766 39520 1822 40000
rect 2134 39520 2190 40000
rect 2594 39520 2650 40000
rect 2962 39520 3018 40000
rect 3330 39520 3386 40000
rect 3790 39520 3846 40000
rect 4158 39520 4214 40000
rect 4526 39520 4582 40000
rect 4986 39520 5042 40000
rect 5354 39520 5410 40000
rect 5722 39520 5778 40000
rect 6182 39520 6238 40000
rect 6550 39520 6606 40000
rect 6918 39520 6974 40000
rect 7378 39520 7434 40000
rect 7746 39520 7802 40000
rect 8206 39520 8262 40000
rect 8574 39520 8630 40000
rect 8942 39520 8998 40000
rect 9402 39520 9458 40000
rect 9770 39520 9826 40000
rect 10138 39520 10194 40000
rect 10598 39520 10654 40000
rect 10966 39520 11022 40000
rect 11334 39520 11390 40000
rect 11794 39520 11850 40000
rect 12162 39520 12218 40000
rect 12530 39520 12586 40000
rect 12990 39520 13046 40000
rect 13358 39520 13414 40000
rect 13726 39520 13782 40000
rect 14186 39522 14242 40000
rect 14108 39520 14242 39522
rect 14554 39520 14610 40000
rect 14922 39522 14978 40000
rect 14922 39520 15056 39522
rect 15382 39520 15438 40000
rect 15750 39520 15806 40000
rect 216 34746 244 39520
rect 584 35873 612 39520
rect 570 35864 626 35873
rect 570 35799 626 35808
rect 952 35290 980 39520
rect 940 35284 992 35290
rect 940 35226 992 35232
rect 204 34740 256 34746
rect 204 34682 256 34688
rect 1412 34202 1440 39520
rect 1490 36408 1546 36417
rect 1490 36343 1546 36352
rect 1400 34196 1452 34202
rect 1400 34138 1452 34144
rect 1504 33658 1532 36343
rect 1780 35193 1808 39520
rect 2148 35290 2176 39520
rect 2608 35329 2636 39520
rect 2686 38720 2742 38729
rect 2686 38655 2742 38664
rect 2594 35320 2650 35329
rect 2136 35284 2188 35290
rect 2594 35255 2650 35264
rect 2136 35226 2188 35232
rect 1766 35184 1822 35193
rect 1676 35148 1728 35154
rect 1766 35119 1822 35128
rect 1676 35090 1728 35096
rect 1688 34134 1716 35090
rect 2700 34746 2728 38655
rect 2688 34740 2740 34746
rect 2688 34682 2740 34688
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2504 34536 2556 34542
rect 2504 34478 2556 34484
rect 1676 34128 1728 34134
rect 1582 34096 1638 34105
rect 1676 34070 1728 34076
rect 1582 34031 1638 34040
rect 1492 33652 1544 33658
rect 1492 33594 1544 33600
rect 1398 33552 1454 33561
rect 1398 33487 1454 33496
rect 1412 32978 1440 33487
rect 1596 33114 1624 34031
rect 1584 33108 1636 33114
rect 1584 33050 1636 33056
rect 1400 32972 1452 32978
rect 1400 32914 1452 32920
rect 1412 32570 1440 32914
rect 1400 32564 1452 32570
rect 1400 32506 1452 32512
rect 1582 31648 1638 31657
rect 1582 31583 1638 31592
rect 1596 29850 1624 31583
rect 1584 29844 1636 29850
rect 1584 29786 1636 29792
rect 1582 29336 1638 29345
rect 1582 29271 1584 29280
rect 1636 29271 1638 29280
rect 1584 29242 1636 29248
rect 1688 28694 1716 34070
rect 1950 33416 2006 33425
rect 1950 33351 1952 33360
rect 2004 33351 2006 33360
rect 1952 33322 2004 33328
rect 1676 28688 1728 28694
rect 1676 28630 1728 28636
rect 2240 27606 2268 34478
rect 2410 30288 2466 30297
rect 2410 30223 2466 30232
rect 2320 29708 2372 29714
rect 2320 29650 2372 29656
rect 2332 29073 2360 29650
rect 2318 29064 2374 29073
rect 2318 28999 2320 29008
rect 2372 28999 2374 29008
rect 2320 28970 2372 28976
rect 2424 28762 2452 30223
rect 2412 28756 2464 28762
rect 2412 28698 2464 28704
rect 2228 27600 2280 27606
rect 2228 27542 2280 27548
rect 2136 27532 2188 27538
rect 2136 27474 2188 27480
rect 2148 27062 2176 27474
rect 2240 27062 2268 27542
rect 2136 27056 2188 27062
rect 1582 27024 1638 27033
rect 2136 26998 2188 27004
rect 2228 27056 2280 27062
rect 2228 26998 2280 27004
rect 1582 26959 1638 26968
rect 1596 25498 1624 26959
rect 2240 26897 2268 26998
rect 2412 26920 2464 26926
rect 2226 26888 2282 26897
rect 2412 26862 2464 26868
rect 2226 26823 2282 26832
rect 2424 26314 2452 26862
rect 2412 26308 2464 26314
rect 2412 26250 2464 26256
rect 1584 25492 1636 25498
rect 1584 25434 1636 25440
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1412 24410 1440 25298
rect 2228 24676 2280 24682
rect 2228 24618 2280 24624
rect 1582 24576 1638 24585
rect 1582 24511 1638 24520
rect 1400 24404 1452 24410
rect 1400 24346 1452 24352
rect 1596 23322 1624 24511
rect 2240 24070 2268 24618
rect 2424 24614 2452 26250
rect 2516 25265 2544 34478
rect 2596 34060 2648 34066
rect 2596 34002 2648 34008
rect 2608 33318 2636 34002
rect 2976 33658 3004 39520
rect 3344 35834 3372 39520
rect 3804 37210 3832 39520
rect 3804 37182 4108 37210
rect 3622 37020 3918 37040
rect 3678 37018 3702 37020
rect 3758 37018 3782 37020
rect 3838 37018 3862 37020
rect 3700 36966 3702 37018
rect 3764 36966 3776 37018
rect 3838 36966 3840 37018
rect 3678 36964 3702 36966
rect 3758 36964 3782 36966
rect 3838 36964 3862 36966
rect 3622 36944 3918 36964
rect 3622 35932 3918 35952
rect 3678 35930 3702 35932
rect 3758 35930 3782 35932
rect 3838 35930 3862 35932
rect 3700 35878 3702 35930
rect 3764 35878 3776 35930
rect 3838 35878 3840 35930
rect 3678 35876 3702 35878
rect 3758 35876 3782 35878
rect 3838 35876 3862 35878
rect 3422 35864 3478 35873
rect 3332 35828 3384 35834
rect 3622 35856 3918 35876
rect 4080 35850 4108 37182
rect 4172 35986 4200 39520
rect 4172 35958 4292 35986
rect 4080 35822 4200 35850
rect 4264 35834 4292 35958
rect 3422 35799 3424 35808
rect 3332 35770 3384 35776
rect 3476 35799 3478 35808
rect 3424 35770 3476 35776
rect 4068 35624 4120 35630
rect 4068 35566 4120 35572
rect 3516 35488 3568 35494
rect 3516 35430 3568 35436
rect 3424 35148 3476 35154
rect 3424 35090 3476 35096
rect 3436 34542 3464 35090
rect 3424 34536 3476 34542
rect 3424 34478 3476 34484
rect 2964 33652 3016 33658
rect 2964 33594 3016 33600
rect 2596 33312 2648 33318
rect 2596 33254 2648 33260
rect 2608 32337 2636 33254
rect 3332 32768 3384 32774
rect 3332 32710 3384 32716
rect 3344 32434 3372 32710
rect 3332 32428 3384 32434
rect 3332 32370 3384 32376
rect 2594 32328 2650 32337
rect 2594 32263 2650 32272
rect 2608 29186 2636 32263
rect 3240 32224 3292 32230
rect 3240 32166 3292 32172
rect 2872 31136 2924 31142
rect 2872 31078 2924 31084
rect 2884 29322 2912 31078
rect 3252 30870 3280 32166
rect 3332 31136 3384 31142
rect 3332 31078 3384 31084
rect 3344 30938 3372 31078
rect 3332 30932 3384 30938
rect 3332 30874 3384 30880
rect 3240 30864 3292 30870
rect 3240 30806 3292 30812
rect 2700 29306 2912 29322
rect 2688 29300 2912 29306
rect 2740 29294 2912 29300
rect 2688 29242 2740 29248
rect 2608 29158 2728 29186
rect 2594 28928 2650 28937
rect 2594 28863 2650 28872
rect 2608 28694 2636 28863
rect 2596 28688 2648 28694
rect 2596 28630 2648 28636
rect 2608 28218 2636 28630
rect 2596 28212 2648 28218
rect 2596 28154 2648 28160
rect 2700 28098 2728 29158
rect 2872 28552 2924 28558
rect 2872 28494 2924 28500
rect 2964 28552 3016 28558
rect 2964 28494 3016 28500
rect 2884 28218 2912 28494
rect 2872 28212 2924 28218
rect 2872 28154 2924 28160
rect 2608 28070 2728 28098
rect 2502 25256 2558 25265
rect 2502 25191 2558 25200
rect 2412 24608 2464 24614
rect 2412 24550 2464 24556
rect 2424 24290 2452 24550
rect 2424 24262 2544 24290
rect 2412 24200 2464 24206
rect 2412 24142 2464 24148
rect 2228 24064 2280 24070
rect 2228 24006 2280 24012
rect 1584 23316 1636 23322
rect 1584 23258 1636 23264
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1688 22273 1716 23122
rect 2240 23050 2268 24006
rect 2424 23322 2452 24142
rect 2412 23316 2464 23322
rect 2412 23258 2464 23264
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22710 2268 22986
rect 2516 22710 2544 24262
rect 2608 23594 2636 28070
rect 2688 27872 2740 27878
rect 2688 27814 2740 27820
rect 2700 26926 2728 27814
rect 2778 27568 2834 27577
rect 2778 27503 2780 27512
rect 2832 27503 2834 27512
rect 2780 27474 2832 27480
rect 2884 27402 2912 28154
rect 2976 28082 3004 28494
rect 2964 28076 3016 28082
rect 2964 28018 3016 28024
rect 2872 27396 2924 27402
rect 2872 27338 2924 27344
rect 2688 26920 2740 26926
rect 2688 26862 2740 26868
rect 2964 26852 3016 26858
rect 2964 26794 3016 26800
rect 2976 26586 3004 26794
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 2976 24614 3004 26522
rect 2964 24608 3016 24614
rect 2964 24550 3016 24556
rect 2688 24404 2740 24410
rect 2688 24346 2740 24352
rect 2596 23588 2648 23594
rect 2596 23530 2648 23536
rect 2700 23254 2728 24346
rect 2976 24206 3004 24550
rect 2964 24200 3016 24206
rect 2964 24142 3016 24148
rect 2976 23866 3004 24142
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 3240 23724 3292 23730
rect 3240 23666 3292 23672
rect 2780 23520 2832 23526
rect 2780 23462 2832 23468
rect 3148 23520 3200 23526
rect 3148 23462 3200 23468
rect 2688 23248 2740 23254
rect 2688 23190 2740 23196
rect 2792 23118 2820 23462
rect 2872 23248 2924 23254
rect 2872 23190 2924 23196
rect 2780 23112 2832 23118
rect 2780 23054 2832 23060
rect 2228 22704 2280 22710
rect 2228 22646 2280 22652
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 1674 22264 1730 22273
rect 1674 22199 1676 22208
rect 1728 22199 1730 22208
rect 1676 22170 1728 22176
rect 2884 22098 2912 23190
rect 2964 23112 3016 23118
rect 2964 23054 3016 23060
rect 2976 22778 3004 23054
rect 2964 22772 3016 22778
rect 2964 22714 3016 22720
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 1582 21992 1638 22001
rect 1582 21927 1638 21936
rect 1596 21690 1624 21927
rect 2884 21690 2912 22034
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 1950 21448 2006 21457
rect 1950 21383 1952 21392
rect 2004 21383 2006 21392
rect 1952 21354 2004 21360
rect 1582 19952 1638 19961
rect 1582 19887 1638 19896
rect 1596 18426 1624 19887
rect 2964 19236 3016 19242
rect 2964 19178 3016 19184
rect 2976 18630 3004 19178
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 1584 18420 1636 18426
rect 1584 18362 1636 18368
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1964 17785 1992 18022
rect 1950 17776 2006 17785
rect 1950 17711 2006 17720
rect 1582 17640 1638 17649
rect 1582 17575 1638 17584
rect 2780 17604 2832 17610
rect 1596 16250 1624 17575
rect 2780 17546 2832 17552
rect 2688 17264 2740 17270
rect 2688 17206 2740 17212
rect 2410 16824 2466 16833
rect 2410 16759 2412 16768
rect 2464 16759 2466 16768
rect 2596 16788 2648 16794
rect 2412 16730 2464 16736
rect 2596 16730 2648 16736
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16250 2084 16526
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1398 16144 1454 16153
rect 1398 16079 1454 16088
rect 1412 16046 1440 16079
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1412 15706 1440 15982
rect 2608 15706 2636 16730
rect 1400 15700 1452 15706
rect 1400 15642 1452 15648
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 1490 15192 1546 15201
rect 2700 15162 2728 17206
rect 2792 16794 2820 17546
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2976 16590 3004 18566
rect 3160 17649 3188 23462
rect 3252 22574 3280 23666
rect 3240 22568 3292 22574
rect 3240 22510 3292 22516
rect 3252 22234 3280 22510
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3252 21554 3280 22170
rect 3436 22114 3464 34478
rect 3528 32552 3556 35430
rect 3622 34844 3918 34864
rect 3678 34842 3702 34844
rect 3758 34842 3782 34844
rect 3838 34842 3862 34844
rect 3700 34790 3702 34842
rect 3764 34790 3776 34842
rect 3838 34790 3840 34842
rect 3678 34788 3702 34790
rect 3758 34788 3782 34790
rect 3838 34788 3862 34790
rect 3622 34768 3918 34788
rect 3976 34468 4028 34474
rect 3976 34410 4028 34416
rect 3988 33862 4016 34410
rect 3976 33856 4028 33862
rect 3976 33798 4028 33804
rect 3622 33756 3918 33776
rect 3678 33754 3702 33756
rect 3758 33754 3782 33756
rect 3838 33754 3862 33756
rect 3700 33702 3702 33754
rect 3764 33702 3776 33754
rect 3838 33702 3840 33754
rect 3678 33700 3702 33702
rect 3758 33700 3782 33702
rect 3838 33700 3862 33702
rect 3622 33680 3918 33700
rect 3622 32668 3918 32688
rect 3678 32666 3702 32668
rect 3758 32666 3782 32668
rect 3838 32666 3862 32668
rect 3700 32614 3702 32666
rect 3764 32614 3776 32666
rect 3838 32614 3840 32666
rect 3678 32612 3702 32614
rect 3758 32612 3782 32614
rect 3838 32612 3862 32614
rect 3622 32592 3918 32612
rect 3528 32524 3648 32552
rect 3620 32230 3648 32524
rect 3698 32464 3754 32473
rect 3698 32399 3754 32408
rect 3792 32428 3844 32434
rect 3712 32366 3740 32399
rect 3792 32370 3844 32376
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3608 32224 3660 32230
rect 3606 32192 3608 32201
rect 3660 32192 3662 32201
rect 3606 32127 3662 32136
rect 3712 32026 3740 32302
rect 3700 32020 3752 32026
rect 3700 31962 3752 31968
rect 3804 31958 3832 32370
rect 3792 31952 3844 31958
rect 3792 31894 3844 31900
rect 3622 31580 3918 31600
rect 3678 31578 3702 31580
rect 3758 31578 3782 31580
rect 3838 31578 3862 31580
rect 3700 31526 3702 31578
rect 3764 31526 3776 31578
rect 3838 31526 3840 31578
rect 3678 31524 3702 31526
rect 3758 31524 3782 31526
rect 3838 31524 3862 31526
rect 3622 31504 3918 31524
rect 3516 31408 3568 31414
rect 3516 31350 3568 31356
rect 3528 31142 3556 31350
rect 3516 31136 3568 31142
rect 3516 31078 3568 31084
rect 3622 30492 3918 30512
rect 3678 30490 3702 30492
rect 3758 30490 3782 30492
rect 3838 30490 3862 30492
rect 3700 30438 3702 30490
rect 3764 30438 3776 30490
rect 3838 30438 3840 30490
rect 3678 30436 3702 30438
rect 3758 30436 3782 30438
rect 3838 30436 3862 30438
rect 3622 30416 3918 30436
rect 3988 30394 4016 33798
rect 4080 33697 4108 35566
rect 4066 33688 4122 33697
rect 4172 33658 4200 35822
rect 4252 35828 4304 35834
rect 4252 35770 4304 35776
rect 4540 35737 4568 39520
rect 4712 36236 4764 36242
rect 4712 36178 4764 36184
rect 4526 35728 4582 35737
rect 4724 35698 4752 36178
rect 4526 35663 4582 35672
rect 4712 35692 4764 35698
rect 4712 35634 4764 35640
rect 4896 35148 4948 35154
rect 4896 35090 4948 35096
rect 4908 34542 4936 35090
rect 4896 34536 4948 34542
rect 4896 34478 4948 34484
rect 4712 34468 4764 34474
rect 4712 34410 4764 34416
rect 4724 33998 4752 34410
rect 4804 34400 4856 34406
rect 4804 34342 4856 34348
rect 4816 34066 4844 34342
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 4066 33623 4122 33632
rect 4160 33652 4212 33658
rect 4160 33594 4212 33600
rect 4724 33522 4752 33934
rect 4712 33516 4764 33522
rect 4712 33458 4764 33464
rect 4068 33312 4120 33318
rect 4620 33312 4672 33318
rect 4120 33260 4384 33266
rect 4068 33254 4384 33260
rect 4620 33254 4672 33260
rect 4080 33238 4384 33254
rect 4160 32768 4212 32774
rect 4080 32728 4160 32756
rect 4080 31346 4108 32728
rect 4160 32710 4212 32716
rect 4252 31680 4304 31686
rect 4252 31622 4304 31628
rect 4264 31482 4292 31622
rect 4252 31476 4304 31482
rect 4252 31418 4304 31424
rect 4068 31340 4120 31346
rect 4068 31282 4120 31288
rect 4160 30728 4212 30734
rect 4160 30670 4212 30676
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 3622 29404 3918 29424
rect 3678 29402 3702 29404
rect 3758 29402 3782 29404
rect 3838 29402 3862 29404
rect 3700 29350 3702 29402
rect 3764 29350 3776 29402
rect 3838 29350 3840 29402
rect 3678 29348 3702 29350
rect 3758 29348 3782 29350
rect 3838 29348 3862 29350
rect 3622 29328 3918 29348
rect 4080 29306 4108 30194
rect 4172 30122 4200 30670
rect 4356 30161 4384 33238
rect 4436 30796 4488 30802
rect 4436 30738 4488 30744
rect 4448 30326 4476 30738
rect 4528 30728 4580 30734
rect 4528 30670 4580 30676
rect 4436 30320 4488 30326
rect 4436 30262 4488 30268
rect 4342 30152 4398 30161
rect 4160 30116 4212 30122
rect 4342 30087 4398 30096
rect 4160 30058 4212 30064
rect 4172 29782 4200 30058
rect 4160 29776 4212 29782
rect 4160 29718 4212 29724
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4252 28960 4304 28966
rect 4252 28902 4304 28908
rect 4264 28422 4292 28902
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 3622 28316 3918 28336
rect 3678 28314 3702 28316
rect 3758 28314 3782 28316
rect 3838 28314 3862 28316
rect 3700 28262 3702 28314
rect 3764 28262 3776 28314
rect 3838 28262 3840 28314
rect 3678 28260 3702 28262
rect 3758 28260 3782 28262
rect 3838 28260 3862 28262
rect 3622 28240 3918 28260
rect 4264 28121 4292 28358
rect 4250 28112 4306 28121
rect 4250 28047 4306 28056
rect 3792 27940 3844 27946
rect 3792 27882 3844 27888
rect 3804 27674 3832 27882
rect 4068 27872 4120 27878
rect 4120 27832 4200 27860
rect 4068 27814 4120 27820
rect 3792 27668 3844 27674
rect 3792 27610 3844 27616
rect 3804 27470 3832 27610
rect 4172 27470 4200 27832
rect 3792 27464 3844 27470
rect 4160 27464 4212 27470
rect 3844 27412 4016 27418
rect 3792 27406 4016 27412
rect 4160 27406 4212 27412
rect 3804 27390 4016 27406
rect 3804 27341 3832 27390
rect 3622 27228 3918 27248
rect 3678 27226 3702 27228
rect 3758 27226 3782 27228
rect 3838 27226 3862 27228
rect 3700 27174 3702 27226
rect 3764 27174 3776 27226
rect 3838 27174 3840 27226
rect 3678 27172 3702 27174
rect 3758 27172 3782 27174
rect 3838 27172 3862 27174
rect 3622 27152 3918 27172
rect 3988 27130 4016 27390
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 3622 26140 3918 26160
rect 3678 26138 3702 26140
rect 3758 26138 3782 26140
rect 3838 26138 3862 26140
rect 3700 26086 3702 26138
rect 3764 26086 3776 26138
rect 3838 26086 3840 26138
rect 3678 26084 3702 26086
rect 3758 26084 3782 26086
rect 3838 26084 3862 26086
rect 3622 26064 3918 26084
rect 3622 25052 3918 25072
rect 3678 25050 3702 25052
rect 3758 25050 3782 25052
rect 3838 25050 3862 25052
rect 3700 24998 3702 25050
rect 3764 24998 3776 25050
rect 3838 24998 3840 25050
rect 3678 24996 3702 24998
rect 3758 24996 3782 24998
rect 3838 24996 3862 24998
rect 3622 24976 3918 24996
rect 4068 24268 4120 24274
rect 4068 24210 4120 24216
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3528 23526 3556 24006
rect 3622 23964 3918 23984
rect 3678 23962 3702 23964
rect 3758 23962 3782 23964
rect 3838 23962 3862 23964
rect 3700 23910 3702 23962
rect 3764 23910 3776 23962
rect 3838 23910 3840 23962
rect 3678 23908 3702 23910
rect 3758 23908 3782 23910
rect 3838 23908 3862 23910
rect 3622 23888 3918 23908
rect 3516 23520 3568 23526
rect 3516 23462 3568 23468
rect 3344 22086 3464 22114
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3146 17640 3202 17649
rect 3146 17575 3202 17584
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2964 15972 3016 15978
rect 2964 15914 3016 15920
rect 2976 15706 3004 15914
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 1490 15127 1546 15136
rect 2688 15156 2740 15162
rect 1504 13530 1532 15127
rect 2688 15098 2740 15104
rect 1584 14816 1636 14822
rect 1584 14758 1636 14764
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 1596 12889 1624 14758
rect 3344 14657 3372 22086
rect 3528 21690 3556 23462
rect 4080 23322 4108 24210
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4172 23202 4200 23802
rect 4264 23526 4292 28047
rect 4252 23520 4304 23526
rect 4252 23462 4304 23468
rect 4080 23174 4200 23202
rect 4080 23118 4108 23174
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 3622 22876 3918 22896
rect 3678 22874 3702 22876
rect 3758 22874 3782 22876
rect 3838 22874 3862 22876
rect 3700 22822 3702 22874
rect 3764 22822 3776 22874
rect 3838 22822 3840 22874
rect 3678 22820 3702 22822
rect 3758 22820 3782 22822
rect 3838 22820 3862 22822
rect 3622 22800 3918 22820
rect 4080 22778 4108 23054
rect 4068 22772 4120 22778
rect 4068 22714 4120 22720
rect 4356 22114 4384 30087
rect 4540 29850 4568 30670
rect 4528 29844 4580 29850
rect 4528 29786 4580 29792
rect 4540 29306 4568 29786
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4528 25288 4580 25294
rect 4528 25230 4580 25236
rect 4540 24750 4568 25230
rect 4528 24744 4580 24750
rect 4528 24686 4580 24692
rect 4436 24608 4488 24614
rect 4436 24550 4488 24556
rect 4448 24274 4476 24550
rect 4436 24268 4488 24274
rect 4436 24210 4488 24216
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4436 24064 4488 24070
rect 4436 24006 4488 24012
rect 4080 22086 4384 22114
rect 3622 21788 3918 21808
rect 3678 21786 3702 21788
rect 3758 21786 3782 21788
rect 3838 21786 3862 21788
rect 3700 21734 3702 21786
rect 3764 21734 3776 21786
rect 3838 21734 3840 21786
rect 3678 21732 3702 21734
rect 3758 21732 3782 21734
rect 3838 21732 3862 21734
rect 3622 21712 3918 21732
rect 3516 21684 3568 21690
rect 3516 21626 3568 21632
rect 4080 21486 4108 22086
rect 4068 21480 4120 21486
rect 4068 21422 4120 21428
rect 3424 21344 3476 21350
rect 3424 21286 3476 21292
rect 3436 20806 3464 21286
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3436 19417 3464 20742
rect 3622 20700 3918 20720
rect 3678 20698 3702 20700
rect 3758 20698 3782 20700
rect 3838 20698 3862 20700
rect 3700 20646 3702 20698
rect 3764 20646 3776 20698
rect 3838 20646 3840 20698
rect 3678 20644 3702 20646
rect 3758 20644 3782 20646
rect 3838 20644 3862 20646
rect 3622 20624 3918 20644
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3620 19802 3648 20198
rect 3528 19774 3648 19802
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17202 3464 17478
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3436 16794 3464 17138
rect 3528 17066 3556 19774
rect 3622 19612 3918 19632
rect 3678 19610 3702 19612
rect 3758 19610 3782 19612
rect 3838 19610 3862 19612
rect 3700 19558 3702 19610
rect 3764 19558 3776 19610
rect 3838 19558 3840 19610
rect 3678 19556 3702 19558
rect 3758 19556 3782 19558
rect 3838 19556 3862 19558
rect 3622 19536 3918 19556
rect 3988 19242 4016 20334
rect 4080 20262 4108 20742
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4080 19666 4108 20198
rect 4172 20058 4200 20198
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4080 19638 4200 19666
rect 3976 19236 4028 19242
rect 3976 19178 4028 19184
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3622 18524 3918 18544
rect 3678 18522 3702 18524
rect 3758 18522 3782 18524
rect 3838 18522 3862 18524
rect 3700 18470 3702 18522
rect 3764 18470 3776 18522
rect 3838 18470 3840 18522
rect 3678 18468 3702 18470
rect 3758 18468 3782 18470
rect 3838 18468 3862 18470
rect 3622 18448 3918 18468
rect 3622 17436 3918 17456
rect 3678 17434 3702 17436
rect 3758 17434 3782 17436
rect 3838 17434 3862 17436
rect 3700 17382 3702 17434
rect 3764 17382 3776 17434
rect 3838 17382 3840 17434
rect 3678 17380 3702 17382
rect 3758 17380 3782 17382
rect 3838 17380 3862 17382
rect 3622 17360 3918 17380
rect 3516 17060 3568 17066
rect 3516 17002 3568 17008
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15910 3556 16526
rect 3622 16348 3918 16368
rect 3678 16346 3702 16348
rect 3758 16346 3782 16348
rect 3838 16346 3862 16348
rect 3700 16294 3702 16346
rect 3764 16294 3776 16346
rect 3838 16294 3840 16346
rect 3678 16292 3702 16294
rect 3758 16292 3782 16294
rect 3838 16292 3862 16294
rect 3622 16272 3918 16292
rect 3516 15904 3568 15910
rect 3516 15846 3568 15852
rect 3528 15026 3556 15846
rect 3622 15260 3918 15280
rect 3678 15258 3702 15260
rect 3758 15258 3782 15260
rect 3838 15258 3862 15260
rect 3700 15206 3702 15258
rect 3764 15206 3776 15258
rect 3838 15206 3840 15258
rect 3678 15204 3702 15206
rect 3758 15204 3782 15206
rect 3838 15204 3862 15206
rect 3622 15184 3918 15204
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3330 14648 3386 14657
rect 3330 14583 3386 14592
rect 3622 14172 3918 14192
rect 3678 14170 3702 14172
rect 3758 14170 3782 14172
rect 3838 14170 3862 14172
rect 3700 14118 3702 14170
rect 3764 14118 3776 14170
rect 3838 14118 3840 14170
rect 3678 14116 3702 14118
rect 3758 14116 3782 14118
rect 3838 14116 3862 14118
rect 3622 14096 3918 14116
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1582 12880 1638 12889
rect 1582 12815 1638 12824
rect 1688 12753 1716 13330
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12782 2728 13126
rect 3622 13084 3918 13104
rect 3678 13082 3702 13084
rect 3758 13082 3782 13084
rect 3838 13082 3862 13084
rect 3700 13030 3702 13082
rect 3764 13030 3776 13082
rect 3838 13030 3840 13082
rect 3678 13028 3702 13030
rect 3758 13028 3782 13030
rect 3838 13028 3862 13030
rect 3622 13008 3918 13028
rect 2688 12776 2740 12782
rect 1674 12744 1730 12753
rect 2688 12718 2740 12724
rect 1674 12679 1676 12688
rect 1728 12679 1730 12688
rect 1676 12650 1728 12656
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2516 12238 2544 12582
rect 2504 12232 2556 12238
rect 2504 12174 2556 12180
rect 2516 11898 2544 12174
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2608 11694 2636 12038
rect 2700 11898 2728 12718
rect 3622 11996 3918 12016
rect 3678 11994 3702 11996
rect 3758 11994 3782 11996
rect 3838 11994 3862 11996
rect 3700 11942 3702 11994
rect 3764 11942 3776 11994
rect 3838 11942 3840 11994
rect 3678 11940 3702 11942
rect 3758 11940 3782 11942
rect 3838 11940 3862 11942
rect 3622 11920 3918 11940
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 1412 10130 1440 10950
rect 2516 10810 2544 11154
rect 2700 10810 2728 11834
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2780 11076 2832 11082
rect 2780 11018 2832 11024
rect 2504 10804 2556 10810
rect 2688 10804 2740 10810
rect 2504 10746 2556 10752
rect 2608 10764 2688 10792
rect 1582 10568 1638 10577
rect 1582 10503 1638 10512
rect 1596 10266 1624 10503
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10266 2452 10406
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 9178 1440 10066
rect 2608 9994 2636 10764
rect 2688 10746 2740 10752
rect 2688 10260 2740 10266
rect 2792 10248 2820 11018
rect 2976 10810 3004 11222
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2740 10220 2820 10248
rect 2688 10202 2740 10208
rect 2976 10198 3004 10746
rect 3344 10606 3372 11562
rect 3622 10908 3918 10928
rect 3678 10906 3702 10908
rect 3758 10906 3782 10908
rect 3838 10906 3862 10908
rect 3700 10854 3702 10906
rect 3764 10854 3776 10906
rect 3838 10854 3840 10906
rect 3678 10852 3702 10854
rect 3758 10852 3782 10854
rect 3838 10852 3862 10854
rect 3622 10832 3918 10852
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3332 10600 3384 10606
rect 3332 10542 3384 10548
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 2964 10192 3016 10198
rect 2964 10134 3016 10140
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2792 9602 2820 10066
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9722 2912 9998
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2976 9722 3004 9930
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2700 9574 2820 9602
rect 2700 9518 2728 9574
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2884 9178 2912 9658
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9178 3004 9522
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3146 8392 3202 8401
rect 2688 8356 2740 8362
rect 3146 8327 3202 8336
rect 2688 8298 2740 8304
rect 2700 8090 2728 8298
rect 2778 8120 2834 8129
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 2688 8084 2740 8090
rect 2778 8055 2834 8064
rect 2688 8026 2740 8032
rect 1780 7410 1808 8026
rect 1768 7404 1820 7410
rect 1768 7346 1820 7352
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 940 5568 992 5574
rect 940 5510 992 5516
rect 570 4176 626 4185
rect 204 4140 256 4146
rect 570 4111 626 4120
rect 204 4082 256 4088
rect 216 480 244 4082
rect 584 480 612 4111
rect 952 480 980 5510
rect 1320 4146 1348 6054
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1412 5370 1440 5714
rect 1400 5364 1452 5370
rect 1400 5306 1452 5312
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1308 4140 1360 4146
rect 1308 4082 1360 4088
rect 1412 480 1440 4966
rect 1504 1193 1532 7142
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1596 3505 1624 6598
rect 2332 6100 2360 6802
rect 2412 6112 2464 6118
rect 2332 6072 2412 6100
rect 2412 6054 2464 6060
rect 2134 5672 2190 5681
rect 2134 5607 2190 5616
rect 1676 4616 1728 4622
rect 1952 4616 2004 4622
rect 1676 4558 1728 4564
rect 1950 4584 1952 4593
rect 2004 4584 2006 4593
rect 1582 3496 1638 3505
rect 1582 3431 1638 3440
rect 1688 2553 1716 4558
rect 1950 4519 2006 4528
rect 2148 4282 2176 5607
rect 2424 5273 2452 6054
rect 2410 5264 2466 5273
rect 2410 5199 2466 5208
rect 2410 5128 2466 5137
rect 2410 5063 2412 5072
rect 2464 5063 2466 5072
rect 2412 5034 2464 5040
rect 2516 4826 2544 6802
rect 2792 6746 2820 8055
rect 3160 7546 3188 8327
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2700 6730 2820 6746
rect 2688 6724 2820 6730
rect 2740 6718 2820 6724
rect 2688 6666 2740 6672
rect 2688 6112 2740 6118
rect 3056 6112 3108 6118
rect 2688 6054 2740 6060
rect 3054 6080 3056 6089
rect 3108 6080 3110 6089
rect 2700 5817 2728 6054
rect 3054 6015 3110 6024
rect 2686 5808 2742 5817
rect 2686 5743 2742 5752
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 4826 2728 5510
rect 2884 5370 2912 5714
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2792 4690 2820 4762
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2148 4078 2176 4218
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 2688 4072 2740 4078
rect 2792 4060 2820 4422
rect 2740 4032 2820 4060
rect 2688 4014 2740 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 1858 3768 1914 3777
rect 1858 3703 1914 3712
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 1780 3505 1808 3538
rect 1766 3496 1822 3505
rect 1766 3431 1822 3440
rect 1780 3194 1808 3431
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1674 2544 1730 2553
rect 1674 2479 1730 2488
rect 1872 1714 1900 3703
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 1950 2816 2006 2825
rect 1950 2751 2006 2760
rect 1964 2650 1992 2751
rect 1952 2644 2004 2650
rect 1952 2586 2004 2592
rect 1780 1686 1900 1714
rect 1490 1184 1546 1193
rect 1490 1119 1546 1128
rect 1780 480 1808 1686
rect 2148 480 2176 3334
rect 2228 3120 2280 3126
rect 2226 3088 2228 3097
rect 2280 3088 2282 3097
rect 2226 3023 2282 3032
rect 2608 480 2636 3878
rect 2884 3738 2912 4762
rect 2976 4622 3004 4966
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2976 4282 3004 4558
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2976 3670 3004 4218
rect 3068 4185 3096 5510
rect 3054 4176 3110 4185
rect 3054 4111 3110 4120
rect 2964 3664 3016 3670
rect 2870 3632 2926 3641
rect 2964 3606 3016 3612
rect 2870 3567 2872 3576
rect 2924 3567 2926 3576
rect 2872 3538 2924 3544
rect 2884 3194 2912 3538
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3252 2990 3280 10406
rect 3344 10266 3372 10542
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3712 10062 3740 10610
rect 3988 10452 4016 18906
rect 4172 18426 4200 19638
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4448 18086 4476 24006
rect 4540 23798 4568 24142
rect 4528 23792 4580 23798
rect 4528 23734 4580 23740
rect 4528 23520 4580 23526
rect 4528 23462 4580 23468
rect 4540 20788 4568 23462
rect 4632 20913 4660 33254
rect 4724 31686 4752 33458
rect 4816 32774 4844 34002
rect 5000 33658 5028 39520
rect 5264 36712 5316 36718
rect 5264 36654 5316 36660
rect 5078 35320 5134 35329
rect 5078 35255 5080 35264
rect 5132 35255 5134 35264
rect 5080 35226 5132 35232
rect 4988 33652 5040 33658
rect 4988 33594 5040 33600
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 4804 31952 4856 31958
rect 4804 31894 4856 31900
rect 4712 31680 4764 31686
rect 4712 31622 4764 31628
rect 4816 31210 4844 31894
rect 4804 31204 4856 31210
rect 4804 31146 4856 31152
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4724 30394 4752 30670
rect 4712 30388 4764 30394
rect 4712 30330 4764 30336
rect 4816 30258 4844 31146
rect 5000 31142 5028 32166
rect 5080 31680 5132 31686
rect 5276 31668 5304 36654
rect 5368 36378 5396 39520
rect 5356 36372 5408 36378
rect 5356 36314 5408 36320
rect 5632 35488 5684 35494
rect 5632 35430 5684 35436
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 5460 32570 5488 33050
rect 5448 32564 5500 32570
rect 5448 32506 5500 32512
rect 5276 31640 5396 31668
rect 5080 31622 5132 31628
rect 5092 31346 5120 31622
rect 5080 31340 5132 31346
rect 5080 31282 5132 31288
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4988 31136 5040 31142
rect 4988 31078 5040 31084
rect 4908 30870 4936 31078
rect 4896 30864 4948 30870
rect 4896 30806 4948 30812
rect 5000 30297 5028 31078
rect 5092 30734 5120 31282
rect 5080 30728 5132 30734
rect 5080 30670 5132 30676
rect 4986 30288 5042 30297
rect 4804 30252 4856 30258
rect 4986 30223 5042 30232
rect 4804 30194 4856 30200
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 5092 29753 5120 29990
rect 5078 29744 5134 29753
rect 5078 29679 5134 29688
rect 5264 29504 5316 29510
rect 5264 29446 5316 29452
rect 5080 29164 5132 29170
rect 5080 29106 5132 29112
rect 4894 29064 4950 29073
rect 4894 28999 4950 29008
rect 4908 28762 4936 28999
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 5092 28558 5120 29106
rect 5172 28960 5224 28966
rect 5172 28902 5224 28908
rect 5080 28552 5132 28558
rect 5080 28494 5132 28500
rect 5092 28218 5120 28494
rect 5080 28212 5132 28218
rect 5080 28154 5132 28160
rect 5184 28064 5212 28902
rect 5276 28540 5304 29446
rect 5368 28966 5396 31640
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 5356 28552 5408 28558
rect 5276 28512 5356 28540
rect 5356 28494 5408 28500
rect 5540 28552 5592 28558
rect 5540 28494 5592 28500
rect 5092 28036 5212 28064
rect 4894 24848 4950 24857
rect 4894 24783 4896 24792
rect 4948 24783 4950 24792
rect 4988 24812 5040 24818
rect 4896 24754 4948 24760
rect 4988 24754 5040 24760
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4724 23866 4752 24142
rect 4908 24070 4936 24754
rect 4896 24064 4948 24070
rect 4896 24006 4948 24012
rect 4802 23896 4858 23905
rect 4712 23860 4764 23866
rect 4802 23831 4858 23840
rect 4712 23802 4764 23808
rect 4816 23594 4844 23831
rect 5000 23730 5028 24754
rect 4988 23724 5040 23730
rect 4988 23666 5040 23672
rect 4896 23656 4948 23662
rect 4896 23598 4948 23604
rect 4804 23588 4856 23594
rect 4804 23530 4856 23536
rect 4816 23322 4844 23530
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4804 23180 4856 23186
rect 4804 23122 4856 23128
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4724 22438 4752 22918
rect 4816 22506 4844 23122
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 22098 4752 22374
rect 4816 22234 4844 22442
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4816 21554 4844 22170
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4712 21480 4764 21486
rect 4764 21428 4844 21434
rect 4712 21422 4844 21428
rect 4724 21406 4844 21422
rect 4618 20904 4674 20913
rect 4618 20839 4674 20848
rect 4540 20760 4660 20788
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 18630 4568 19722
rect 4632 19378 4660 20760
rect 4712 19848 4764 19854
rect 4710 19816 4712 19825
rect 4764 19816 4766 19825
rect 4710 19751 4766 19760
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4724 19242 4752 19751
rect 4620 19236 4672 19242
rect 4620 19178 4672 19184
rect 4712 19236 4764 19242
rect 4712 19178 4764 19184
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4540 18290 4568 18566
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4080 17338 4108 17818
rect 4264 17678 4292 17709
rect 4252 17672 4304 17678
rect 4250 17640 4252 17649
rect 4304 17640 4306 17649
rect 4250 17575 4306 17584
rect 4264 17338 4292 17575
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16266 4108 17070
rect 4526 16824 4582 16833
rect 4526 16759 4528 16768
rect 4580 16759 4582 16768
rect 4528 16730 4580 16736
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4080 16250 4200 16266
rect 4080 16244 4212 16250
rect 4080 16238 4160 16244
rect 4160 16186 4212 16192
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 4080 15162 4108 15642
rect 4172 15570 4200 16186
rect 4448 15706 4476 16594
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4540 15638 4568 16730
rect 4632 16590 4660 19178
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4632 15978 4660 16526
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4620 15156 4672 15162
rect 4620 15098 4672 15104
rect 4434 15056 4490 15065
rect 4434 14991 4490 15000
rect 4448 14958 4476 14991
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4540 14618 4568 14758
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4632 13841 4660 15098
rect 4618 13832 4674 13841
rect 4618 13767 4674 13776
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12374 4108 12582
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4068 12232 4120 12238
rect 4120 12192 4200 12220
rect 4068 12174 4120 12180
rect 4172 11898 4200 12192
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4632 11286 4660 12242
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 3988 10424 4200 10452
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3622 9820 3918 9840
rect 3678 9818 3702 9820
rect 3758 9818 3782 9820
rect 3838 9818 3862 9820
rect 3700 9766 3702 9818
rect 3764 9766 3776 9818
rect 3838 9766 3840 9818
rect 3678 9764 3702 9766
rect 3758 9764 3782 9766
rect 3838 9764 3862 9766
rect 3622 9744 3918 9764
rect 4080 9654 4108 10066
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 3332 9512 3384 9518
rect 3330 9480 3332 9489
rect 3424 9512 3476 9518
rect 3384 9480 3386 9489
rect 3424 9454 3476 9460
rect 3330 9415 3386 9424
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 3344 8634 3372 9318
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3436 8514 3464 9454
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3622 8732 3918 8752
rect 3678 8730 3702 8732
rect 3758 8730 3782 8732
rect 3838 8730 3862 8732
rect 3700 8678 3702 8730
rect 3764 8678 3776 8730
rect 3838 8678 3840 8730
rect 3678 8676 3702 8678
rect 3758 8676 3782 8678
rect 3838 8676 3862 8678
rect 3622 8656 3918 8676
rect 3344 8486 3464 8514
rect 3790 8528 3846 8537
rect 3344 3058 3372 8486
rect 3790 8463 3792 8472
rect 3844 8463 3846 8472
rect 3792 8434 3844 8440
rect 3988 8362 4016 8910
rect 4172 8378 4200 10424
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4540 9450 4568 9862
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4252 9104 4304 9110
rect 4252 9046 4304 9052
rect 4264 8498 4292 9046
rect 4724 8514 4752 19178
rect 4252 8492 4304 8498
rect 4252 8434 4304 8440
rect 4632 8486 4752 8514
rect 3976 8356 4028 8362
rect 4172 8350 4292 8378
rect 3976 8298 4028 8304
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3712 8090 3740 8230
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3436 6458 3464 8026
rect 3622 7644 3918 7664
rect 3678 7642 3702 7644
rect 3758 7642 3782 7644
rect 3838 7642 3862 7644
rect 3700 7590 3702 7642
rect 3764 7590 3776 7642
rect 3838 7590 3840 7642
rect 3678 7588 3702 7590
rect 3758 7588 3782 7590
rect 3838 7588 3862 7590
rect 3622 7568 3918 7588
rect 3622 6556 3918 6576
rect 3678 6554 3702 6556
rect 3758 6554 3782 6556
rect 3838 6554 3862 6556
rect 3700 6502 3702 6554
rect 3764 6502 3776 6554
rect 3838 6502 3840 6554
rect 3678 6500 3702 6502
rect 3758 6500 3782 6502
rect 3838 6500 3862 6502
rect 3622 6480 3918 6500
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3436 5098 3464 5510
rect 3622 5468 3918 5488
rect 3678 5466 3702 5468
rect 3758 5466 3782 5468
rect 3838 5466 3862 5468
rect 3700 5414 3702 5466
rect 3764 5414 3776 5466
rect 3838 5414 3840 5466
rect 3678 5412 3702 5414
rect 3758 5412 3782 5414
rect 3838 5412 3862 5414
rect 3622 5392 3918 5412
rect 3516 5160 3568 5166
rect 3516 5102 3568 5108
rect 3424 5092 3476 5098
rect 3424 5034 3476 5040
rect 3528 4486 3556 5102
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3528 4128 3556 4422
rect 3622 4380 3918 4400
rect 3678 4378 3702 4380
rect 3758 4378 3782 4380
rect 3838 4378 3862 4380
rect 3700 4326 3702 4378
rect 3764 4326 3776 4378
rect 3838 4326 3840 4378
rect 3678 4324 3702 4326
rect 3758 4324 3782 4326
rect 3838 4324 3862 4326
rect 3622 4304 3918 4324
rect 3884 4140 3936 4146
rect 3528 4100 3832 4128
rect 3804 3482 3832 4100
rect 3884 4082 3936 4088
rect 3896 3738 3924 4082
rect 3988 3890 4016 5510
rect 4172 5166 4200 6326
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 4080 4570 4108 4626
rect 4080 4542 4200 4570
rect 4172 4010 4200 4542
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 3988 3862 4200 3890
rect 4172 3738 4200 3862
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3534 4292 8350
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4540 7886 4568 8230
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7206 4568 7822
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 6390 4568 7142
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4540 5914 4568 6054
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4448 4758 4476 5510
rect 4540 4826 4568 5850
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4344 3664 4396 3670
rect 4632 3641 4660 8486
rect 4712 8288 4764 8294
rect 4712 8230 4764 8236
rect 4724 5370 4752 8230
rect 4816 8072 4844 21406
rect 4908 20058 4936 23598
rect 5000 23254 5028 23666
rect 5092 23662 5120 28036
rect 5172 27940 5224 27946
rect 5172 27882 5224 27888
rect 5184 27470 5212 27882
rect 5368 27674 5396 28494
rect 5552 28218 5580 28494
rect 5540 28212 5592 28218
rect 5540 28154 5592 28160
rect 5356 27668 5408 27674
rect 5356 27610 5408 27616
rect 5172 27464 5224 27470
rect 5172 27406 5224 27412
rect 5184 26790 5212 27406
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 5184 26382 5212 26726
rect 5448 26444 5500 26450
rect 5448 26386 5500 26392
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5460 26330 5488 26386
rect 5184 25702 5212 26318
rect 5460 26302 5580 26330
rect 5552 25906 5580 26302
rect 5540 25900 5592 25906
rect 5540 25842 5592 25848
rect 5172 25696 5224 25702
rect 5172 25638 5224 25644
rect 5080 23656 5132 23662
rect 5080 23598 5132 23604
rect 4988 23248 5040 23254
rect 5184 23225 5212 25638
rect 5644 24721 5672 35430
rect 5736 35290 5764 39520
rect 6196 36922 6224 39520
rect 6564 37754 6592 39520
rect 6564 37726 6684 37754
rect 6289 37564 6585 37584
rect 6345 37562 6369 37564
rect 6425 37562 6449 37564
rect 6505 37562 6529 37564
rect 6367 37510 6369 37562
rect 6431 37510 6443 37562
rect 6505 37510 6507 37562
rect 6345 37508 6369 37510
rect 6425 37508 6449 37510
rect 6505 37508 6529 37510
rect 6289 37488 6585 37508
rect 6184 36916 6236 36922
rect 6184 36858 6236 36864
rect 6289 36476 6585 36496
rect 6345 36474 6369 36476
rect 6425 36474 6449 36476
rect 6505 36474 6529 36476
rect 6367 36422 6369 36474
rect 6431 36422 6443 36474
rect 6505 36422 6507 36474
rect 6345 36420 6369 36422
rect 6425 36420 6449 36422
rect 6505 36420 6529 36422
rect 6289 36400 6585 36420
rect 6656 36378 6684 37726
rect 6644 36372 6696 36378
rect 6644 36314 6696 36320
rect 6000 36236 6052 36242
rect 6000 36178 6052 36184
rect 5816 35692 5868 35698
rect 5816 35634 5868 35640
rect 5724 35284 5776 35290
rect 5724 35226 5776 35232
rect 5724 32768 5776 32774
rect 5724 32710 5776 32716
rect 5736 29850 5764 32710
rect 5828 30190 5856 35634
rect 6012 35494 6040 36178
rect 6000 35488 6052 35494
rect 6000 35430 6052 35436
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5816 30184 5868 30190
rect 5816 30126 5868 30132
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 5736 29306 5764 29786
rect 5816 29640 5868 29646
rect 5816 29582 5868 29588
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5722 29200 5778 29209
rect 5828 29170 5856 29582
rect 5722 29135 5778 29144
rect 5816 29164 5868 29170
rect 5736 24993 5764 29135
rect 5816 29106 5868 29112
rect 5828 27606 5856 29106
rect 5816 27600 5868 27606
rect 5816 27542 5868 27548
rect 5828 27130 5856 27542
rect 5816 27124 5868 27130
rect 5816 27066 5868 27072
rect 5722 24984 5778 24993
rect 5722 24919 5778 24928
rect 5630 24712 5686 24721
rect 5630 24647 5686 24656
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 4988 23190 5040 23196
rect 5170 23216 5226 23225
rect 5170 23151 5226 23160
rect 5184 22982 5212 23151
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 5184 22273 5212 22374
rect 5170 22264 5226 22273
rect 5170 22199 5226 22208
rect 5276 22166 5304 22646
rect 5356 22636 5408 22642
rect 5356 22578 5408 22584
rect 5264 22160 5316 22166
rect 5264 22102 5316 22108
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5092 20806 5120 21286
rect 5276 21146 5304 22102
rect 5368 21894 5396 22578
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5354 21584 5410 21593
rect 5354 21519 5410 21528
rect 5368 21350 5396 21519
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5264 21140 5316 21146
rect 5264 21082 5316 21088
rect 5080 20800 5132 20806
rect 5080 20742 5132 20748
rect 4896 20052 4948 20058
rect 4896 19994 4948 20000
rect 4908 19174 4936 19994
rect 4988 19372 5040 19378
rect 4988 19314 5040 19320
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18970 4936 19110
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4908 18358 4936 18770
rect 4896 18352 4948 18358
rect 4896 18294 4948 18300
rect 4896 16992 4948 16998
rect 4896 16934 4948 16940
rect 4908 16726 4936 16934
rect 4896 16720 4948 16726
rect 4896 16662 4948 16668
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4908 15162 4936 15438
rect 4896 15156 4948 15162
rect 4896 15098 4948 15104
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4908 13938 4936 14418
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4894 13832 4950 13841
rect 4894 13767 4950 13776
rect 4908 11898 4936 13767
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5000 11778 5028 19314
rect 5092 17066 5120 20742
rect 5170 19408 5226 19417
rect 5170 19343 5226 19352
rect 5184 17882 5212 19343
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5276 18222 5304 19110
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5080 17060 5132 17066
rect 5080 17002 5132 17008
rect 5092 16794 5120 17002
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5078 14648 5134 14657
rect 5078 14583 5080 14592
rect 5132 14583 5134 14592
rect 5080 14554 5132 14560
rect 5092 14074 5120 14554
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4908 11750 5028 11778
rect 4908 10606 4936 11750
rect 4986 11656 5042 11665
rect 4986 11591 5042 11600
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4816 8044 4936 8072
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7410 4844 7890
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4908 5846 4936 8044
rect 5000 7290 5028 11591
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5092 11354 5120 11494
rect 5184 11354 5212 12038
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5172 11212 5224 11218
rect 5276 11200 5304 18022
rect 5368 17134 5396 21286
rect 5460 17241 5488 23258
rect 5552 22574 5580 24006
rect 5724 23248 5776 23254
rect 5724 23190 5776 23196
rect 5736 22642 5764 23190
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5540 22568 5592 22574
rect 5540 22510 5592 22516
rect 5552 20602 5580 22510
rect 5724 22432 5776 22438
rect 5724 22374 5776 22380
rect 5736 22098 5764 22374
rect 5724 22092 5776 22098
rect 5724 22034 5776 22040
rect 5736 21434 5764 22034
rect 5736 21406 5856 21434
rect 5828 21350 5856 21406
rect 5816 21344 5868 21350
rect 5722 21312 5778 21321
rect 5816 21286 5868 21292
rect 5722 21247 5778 21256
rect 5540 20596 5592 20602
rect 5540 20538 5592 20544
rect 5736 19378 5764 21247
rect 5828 19922 5856 21286
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5552 18086 5580 18770
rect 5540 18080 5592 18086
rect 5540 18022 5592 18028
rect 5552 17678 5580 18022
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5446 17232 5502 17241
rect 5552 17202 5580 17614
rect 5446 17167 5502 17176
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5356 17128 5408 17134
rect 5354 17096 5356 17105
rect 5448 17128 5500 17134
rect 5408 17096 5410 17105
rect 5448 17070 5500 17076
rect 5354 17031 5410 17040
rect 5460 16658 5488 17070
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5368 15162 5396 15914
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5356 14544 5408 14550
rect 5354 14512 5356 14521
rect 5408 14512 5410 14521
rect 5354 14447 5410 14456
rect 5460 14414 5488 16594
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5552 15162 5580 15506
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5368 11354 5396 14010
rect 5460 13870 5488 14350
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5460 12442 5488 13806
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5276 11172 5396 11200
rect 5172 11154 5224 11160
rect 5080 10192 5132 10198
rect 5080 10134 5132 10140
rect 5092 9586 5120 10134
rect 5184 10033 5212 11154
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 5276 10266 5304 11018
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5170 10024 5226 10033
rect 5170 9959 5226 9968
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 5092 9178 5120 9522
rect 5080 9172 5132 9178
rect 5080 9114 5132 9120
rect 5262 7304 5318 7313
rect 5000 7262 5212 7290
rect 4988 7200 5040 7206
rect 4988 7142 5040 7148
rect 5000 6322 5028 7142
rect 5080 6792 5132 6798
rect 5080 6734 5132 6740
rect 5092 6390 5120 6734
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 4986 6216 5042 6225
rect 4986 6151 4988 6160
rect 5040 6151 5042 6160
rect 4988 6122 5040 6128
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4908 5030 4936 5782
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5000 5030 5028 5646
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 4816 4282 4844 4762
rect 4908 4729 4936 4966
rect 4894 4720 4950 4729
rect 4894 4655 4950 4664
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4344 3606 4396 3612
rect 4618 3632 4674 3641
rect 4252 3528 4304 3534
rect 3516 3460 3568 3466
rect 3804 3454 4200 3482
rect 4252 3470 4304 3476
rect 3516 3402 3568 3408
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 2976 480 3004 2246
rect 3344 480 3372 2790
rect 3528 1442 3556 3402
rect 3622 3292 3918 3312
rect 3678 3290 3702 3292
rect 3758 3290 3782 3292
rect 3838 3290 3862 3292
rect 3700 3238 3702 3290
rect 3764 3238 3776 3290
rect 3838 3238 3840 3290
rect 3678 3236 3702 3238
rect 3758 3236 3782 3238
rect 3838 3236 3862 3238
rect 3622 3216 3918 3236
rect 4172 3074 4200 3454
rect 4172 3058 4292 3074
rect 4160 3052 4292 3058
rect 4212 3046 4292 3052
rect 4160 2994 4212 3000
rect 4158 2952 4214 2961
rect 4158 2887 4214 2896
rect 3622 2204 3918 2224
rect 3678 2202 3702 2204
rect 3758 2202 3782 2204
rect 3838 2202 3862 2204
rect 3700 2150 3702 2202
rect 3764 2150 3776 2202
rect 3838 2150 3840 2202
rect 3678 2148 3702 2150
rect 3758 2148 3782 2150
rect 3838 2148 3862 2150
rect 3622 2128 3918 2148
rect 3528 1414 3832 1442
rect 3804 480 3832 1414
rect 4172 480 4200 2887
rect 4264 2650 4292 3046
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4356 2582 4384 3606
rect 4618 3567 4674 3576
rect 4816 3534 4844 4218
rect 5184 3670 5212 7262
rect 5262 7239 5264 7248
rect 5316 7239 5318 7248
rect 5264 7210 5316 7216
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5276 6769 5304 6938
rect 5262 6760 5318 6769
rect 5262 6695 5318 6704
rect 5276 5778 5304 6695
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5368 5166 5396 11172
rect 5460 10674 5488 11698
rect 5644 11626 5672 19314
rect 5724 19236 5776 19242
rect 5724 19178 5776 19184
rect 5736 18902 5764 19178
rect 5724 18896 5776 18902
rect 5724 18838 5776 18844
rect 5920 17354 5948 34478
rect 6012 29034 6040 35430
rect 6289 35388 6585 35408
rect 6345 35386 6369 35388
rect 6425 35386 6449 35388
rect 6505 35386 6529 35388
rect 6367 35334 6369 35386
rect 6431 35334 6443 35386
rect 6505 35334 6507 35386
rect 6345 35332 6369 35334
rect 6425 35332 6449 35334
rect 6505 35332 6529 35334
rect 6289 35312 6585 35332
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6288 34542 6316 35090
rect 6932 35018 6960 39520
rect 7392 35834 7420 39520
rect 7380 35828 7432 35834
rect 7380 35770 7432 35776
rect 7564 35284 7616 35290
rect 7564 35226 7616 35232
rect 7576 35193 7604 35226
rect 7562 35184 7618 35193
rect 7562 35119 7618 35128
rect 7656 35148 7708 35154
rect 7656 35090 7708 35096
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 7668 34746 7696 35090
rect 7656 34740 7708 34746
rect 7656 34682 7708 34688
rect 6276 34536 6328 34542
rect 6276 34478 6328 34484
rect 6828 34536 6880 34542
rect 7380 34536 7432 34542
rect 6880 34496 7052 34524
rect 6828 34478 6880 34484
rect 6289 34300 6585 34320
rect 6345 34298 6369 34300
rect 6425 34298 6449 34300
rect 6505 34298 6529 34300
rect 6367 34246 6369 34298
rect 6431 34246 6443 34298
rect 6505 34246 6507 34298
rect 6345 34244 6369 34246
rect 6425 34244 6449 34246
rect 6505 34244 6529 34246
rect 6289 34224 6585 34244
rect 6276 34060 6328 34066
rect 6276 34002 6328 34008
rect 6092 33856 6144 33862
rect 6092 33798 6144 33804
rect 6104 33386 6132 33798
rect 6288 33658 6316 34002
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6642 33688 6698 33697
rect 6276 33652 6328 33658
rect 6642 33623 6698 33632
rect 6276 33594 6328 33600
rect 6092 33380 6144 33386
rect 6092 33322 6144 33328
rect 6289 33212 6585 33232
rect 6345 33210 6369 33212
rect 6425 33210 6449 33212
rect 6505 33210 6529 33212
rect 6367 33158 6369 33210
rect 6431 33158 6443 33210
rect 6505 33158 6507 33210
rect 6345 33156 6369 33158
rect 6425 33156 6449 33158
rect 6505 33156 6529 33158
rect 6289 33136 6585 33156
rect 6184 32904 6236 32910
rect 6184 32846 6236 32852
rect 6368 32904 6420 32910
rect 6368 32846 6420 32852
rect 6196 32570 6224 32846
rect 6184 32564 6236 32570
rect 6184 32506 6236 32512
rect 6090 32192 6146 32201
rect 6090 32127 6146 32136
rect 6000 29028 6052 29034
rect 6000 28970 6052 28976
rect 6012 27010 6040 28970
rect 6104 28778 6132 32127
rect 6196 32026 6224 32506
rect 6380 32502 6408 32846
rect 6368 32496 6420 32502
rect 6368 32438 6420 32444
rect 6289 32124 6585 32144
rect 6345 32122 6369 32124
rect 6425 32122 6449 32124
rect 6505 32122 6529 32124
rect 6367 32070 6369 32122
rect 6431 32070 6443 32122
rect 6505 32070 6507 32122
rect 6345 32068 6369 32070
rect 6425 32068 6449 32070
rect 6505 32068 6529 32070
rect 6289 32048 6585 32068
rect 6656 32026 6684 33623
rect 6736 33448 6788 33454
rect 6736 33390 6788 33396
rect 6748 33289 6776 33390
rect 6828 33312 6880 33318
rect 6734 33280 6790 33289
rect 6828 33254 6880 33260
rect 6734 33215 6790 33224
rect 6840 32910 6868 33254
rect 6828 32904 6880 32910
rect 6828 32846 6880 32852
rect 6184 32020 6236 32026
rect 6184 31962 6236 31968
rect 6644 32020 6696 32026
rect 6644 31962 6696 31968
rect 6656 31142 6684 31962
rect 6828 31952 6880 31958
rect 6828 31894 6880 31900
rect 6840 31414 6868 31894
rect 6932 31482 6960 33798
rect 6920 31476 6972 31482
rect 6920 31418 6972 31424
rect 6828 31408 6880 31414
rect 6828 31350 6880 31356
rect 6644 31136 6696 31142
rect 6644 31078 6696 31084
rect 6289 31036 6585 31056
rect 6345 31034 6369 31036
rect 6425 31034 6449 31036
rect 6505 31034 6529 31036
rect 6367 30982 6369 31034
rect 6431 30982 6443 31034
rect 6505 30982 6507 31034
rect 6345 30980 6369 30982
rect 6425 30980 6449 30982
rect 6505 30980 6529 30982
rect 6289 30960 6585 30980
rect 6184 30796 6236 30802
rect 6184 30738 6236 30744
rect 6196 30161 6224 30738
rect 6182 30152 6238 30161
rect 6182 30087 6184 30096
rect 6236 30087 6238 30096
rect 6184 30058 6236 30064
rect 6289 29948 6585 29968
rect 6345 29946 6369 29948
rect 6425 29946 6449 29948
rect 6505 29946 6529 29948
rect 6367 29894 6369 29946
rect 6431 29894 6443 29946
rect 6505 29894 6507 29946
rect 6345 29892 6369 29894
rect 6425 29892 6449 29894
rect 6505 29892 6529 29894
rect 6289 29872 6585 29892
rect 6289 28860 6585 28880
rect 6345 28858 6369 28860
rect 6425 28858 6449 28860
rect 6505 28858 6529 28860
rect 6367 28806 6369 28858
rect 6431 28806 6443 28858
rect 6505 28806 6507 28858
rect 6345 28804 6369 28806
rect 6425 28804 6449 28806
rect 6505 28804 6529 28806
rect 6289 28784 6585 28804
rect 6104 28750 6224 28778
rect 6092 28688 6144 28694
rect 6092 28630 6144 28636
rect 6104 27878 6132 28630
rect 6196 27985 6224 28750
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6182 27976 6238 27985
rect 6564 27946 6592 28494
rect 6182 27911 6238 27920
rect 6552 27940 6604 27946
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 6104 27130 6132 27814
rect 6196 27554 6224 27911
rect 6552 27882 6604 27888
rect 6289 27772 6585 27792
rect 6345 27770 6369 27772
rect 6425 27770 6449 27772
rect 6505 27770 6529 27772
rect 6367 27718 6369 27770
rect 6431 27718 6443 27770
rect 6505 27718 6507 27770
rect 6345 27716 6369 27718
rect 6425 27716 6449 27718
rect 6505 27716 6529 27718
rect 6289 27696 6585 27716
rect 6196 27526 6408 27554
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6184 27056 6236 27062
rect 6012 26982 6132 27010
rect 6184 26998 6236 27004
rect 6000 26852 6052 26858
rect 6000 26794 6052 26800
rect 5828 17326 5948 17354
rect 5828 14929 5856 17326
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5814 14920 5870 14929
rect 5814 14855 5870 14864
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5460 10198 5488 10610
rect 5552 10266 5580 11154
rect 5736 11150 5764 12922
rect 5828 12918 5856 13398
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5632 11144 5684 11150
rect 5632 11086 5684 11092
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5644 10742 5672 11086
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5644 10198 5672 10678
rect 5828 10470 5856 12718
rect 5920 10538 5948 17206
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 6012 9382 6040 26794
rect 6104 17270 6132 26982
rect 6196 26586 6224 26998
rect 6380 26858 6408 27526
rect 6368 26852 6420 26858
rect 6368 26794 6420 26800
rect 6289 26684 6585 26704
rect 6345 26682 6369 26684
rect 6425 26682 6449 26684
rect 6505 26682 6529 26684
rect 6367 26630 6369 26682
rect 6431 26630 6443 26682
rect 6505 26630 6507 26682
rect 6345 26628 6369 26630
rect 6425 26628 6449 26630
rect 6505 26628 6529 26630
rect 6289 26608 6585 26628
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6289 25596 6585 25616
rect 6345 25594 6369 25596
rect 6425 25594 6449 25596
rect 6505 25594 6529 25596
rect 6367 25542 6369 25594
rect 6431 25542 6443 25594
rect 6505 25542 6507 25594
rect 6345 25540 6369 25542
rect 6425 25540 6449 25542
rect 6505 25540 6529 25542
rect 6289 25520 6585 25540
rect 6289 24508 6585 24528
rect 6345 24506 6369 24508
rect 6425 24506 6449 24508
rect 6505 24506 6529 24508
rect 6367 24454 6369 24506
rect 6431 24454 6443 24506
rect 6505 24454 6507 24506
rect 6345 24452 6369 24454
rect 6425 24452 6449 24454
rect 6505 24452 6529 24454
rect 6289 24432 6585 24452
rect 6289 23420 6585 23440
rect 6345 23418 6369 23420
rect 6425 23418 6449 23420
rect 6505 23418 6529 23420
rect 6367 23366 6369 23418
rect 6431 23366 6443 23418
rect 6505 23366 6507 23418
rect 6345 23364 6369 23366
rect 6425 23364 6449 23366
rect 6505 23364 6529 23366
rect 6289 23344 6585 23364
rect 6184 22500 6236 22506
rect 6184 22442 6236 22448
rect 6196 22234 6224 22442
rect 6289 22332 6585 22352
rect 6345 22330 6369 22332
rect 6425 22330 6449 22332
rect 6505 22330 6529 22332
rect 6367 22278 6369 22330
rect 6431 22278 6443 22330
rect 6505 22278 6507 22330
rect 6345 22276 6369 22278
rect 6425 22276 6449 22278
rect 6505 22276 6529 22278
rect 6289 22256 6585 22276
rect 6184 22228 6236 22234
rect 6184 22170 6236 22176
rect 6656 21593 6684 31078
rect 6826 30968 6882 30977
rect 6748 30912 6826 30920
rect 6748 30892 6828 30912
rect 6748 29850 6776 30892
rect 6880 30903 6882 30912
rect 6828 30874 6880 30880
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 6840 30394 6868 30670
rect 6920 30592 6972 30598
rect 6920 30534 6972 30540
rect 6828 30388 6880 30394
rect 6828 30330 6880 30336
rect 6932 30258 6960 30534
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 6748 23905 6776 29786
rect 6840 29714 6868 29990
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6840 29306 6868 29650
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 7024 29034 7052 34496
rect 7380 34478 7432 34484
rect 7392 33930 7420 34478
rect 7380 33924 7432 33930
rect 7380 33866 7432 33872
rect 7564 33856 7616 33862
rect 7564 33798 7616 33804
rect 7576 33561 7604 33798
rect 7562 33552 7618 33561
rect 7562 33487 7618 33496
rect 7104 33380 7156 33386
rect 7104 33322 7156 33328
rect 7116 33046 7144 33322
rect 7472 33312 7524 33318
rect 7472 33254 7524 33260
rect 7380 33108 7432 33114
rect 7380 33050 7432 33056
rect 7104 33040 7156 33046
rect 7104 32982 7156 32988
rect 7116 31822 7144 32982
rect 7288 32904 7340 32910
rect 7288 32846 7340 32852
rect 7300 32366 7328 32846
rect 7392 32570 7420 33050
rect 7380 32564 7432 32570
rect 7380 32506 7432 32512
rect 7288 32360 7340 32366
rect 7286 32328 7288 32337
rect 7340 32328 7342 32337
rect 7286 32263 7342 32272
rect 7196 31952 7248 31958
rect 7194 31920 7196 31929
rect 7248 31920 7250 31929
rect 7194 31855 7250 31864
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7116 30802 7144 31758
rect 7380 31748 7432 31754
rect 7380 31690 7432 31696
rect 7392 31142 7420 31690
rect 7288 31136 7340 31142
rect 7288 31078 7340 31084
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 7300 30666 7328 31078
rect 7288 30660 7340 30666
rect 7288 30602 7340 30608
rect 7196 30048 7248 30054
rect 7194 30016 7196 30025
rect 7248 30016 7250 30025
rect 7194 29951 7250 29960
rect 7300 29850 7328 30602
rect 7484 30258 7512 33254
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7576 30938 7604 31282
rect 7564 30932 7616 30938
rect 7564 30874 7616 30880
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7484 29782 7512 30194
rect 7472 29776 7524 29782
rect 7472 29718 7524 29724
rect 7288 29096 7340 29102
rect 7286 29064 7288 29073
rect 7340 29064 7342 29073
rect 7012 29028 7064 29034
rect 7286 28999 7342 29008
rect 7012 28970 7064 28976
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6840 27713 6868 27814
rect 6826 27704 6882 27713
rect 6826 27639 6882 27648
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6840 26042 6868 26862
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 6734 23896 6790 23905
rect 6734 23831 6790 23840
rect 6736 23792 6788 23798
rect 6736 23734 6788 23740
rect 6642 21584 6698 21593
rect 6642 21519 6698 21528
rect 6289 21244 6585 21264
rect 6345 21242 6369 21244
rect 6425 21242 6449 21244
rect 6505 21242 6529 21244
rect 6367 21190 6369 21242
rect 6431 21190 6443 21242
rect 6505 21190 6507 21242
rect 6345 21188 6369 21190
rect 6425 21188 6449 21190
rect 6505 21188 6529 21190
rect 6289 21168 6585 21188
rect 6644 20528 6696 20534
rect 6644 20470 6696 20476
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6196 17082 6224 20198
rect 6289 20156 6585 20176
rect 6345 20154 6369 20156
rect 6425 20154 6449 20156
rect 6505 20154 6529 20156
rect 6367 20102 6369 20154
rect 6431 20102 6443 20154
rect 6505 20102 6507 20154
rect 6345 20100 6369 20102
rect 6425 20100 6449 20102
rect 6505 20100 6529 20102
rect 6289 20080 6585 20100
rect 6656 19990 6684 20470
rect 6644 19984 6696 19990
rect 6644 19926 6696 19932
rect 6656 19514 6684 19926
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6289 19068 6585 19088
rect 6345 19066 6369 19068
rect 6425 19066 6449 19068
rect 6505 19066 6529 19068
rect 6367 19014 6369 19066
rect 6431 19014 6443 19066
rect 6505 19014 6507 19066
rect 6345 19012 6369 19014
rect 6425 19012 6449 19014
rect 6505 19012 6529 19014
rect 6289 18992 6585 19012
rect 6276 18624 6328 18630
rect 6276 18566 6328 18572
rect 6288 18290 6316 18566
rect 6276 18284 6328 18290
rect 6276 18226 6328 18232
rect 6289 17980 6585 18000
rect 6345 17978 6369 17980
rect 6425 17978 6449 17980
rect 6505 17978 6529 17980
rect 6367 17926 6369 17978
rect 6431 17926 6443 17978
rect 6505 17926 6507 17978
rect 6345 17924 6369 17926
rect 6425 17924 6449 17926
rect 6505 17924 6529 17926
rect 6289 17904 6585 17924
rect 6104 17054 6224 17082
rect 6104 13954 6132 17054
rect 6644 16992 6696 16998
rect 6644 16934 6696 16940
rect 6289 16892 6585 16912
rect 6345 16890 6369 16892
rect 6425 16890 6449 16892
rect 6505 16890 6529 16892
rect 6367 16838 6369 16890
rect 6431 16838 6443 16890
rect 6505 16838 6507 16890
rect 6345 16836 6369 16838
rect 6425 16836 6449 16838
rect 6505 16836 6529 16838
rect 6289 16816 6585 16836
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6196 16046 6224 16594
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6288 16046 6316 16526
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6196 15366 6224 15982
rect 6289 15804 6585 15824
rect 6345 15802 6369 15804
rect 6425 15802 6449 15804
rect 6505 15802 6529 15804
rect 6367 15750 6369 15802
rect 6431 15750 6443 15802
rect 6505 15750 6507 15802
rect 6345 15748 6369 15750
rect 6425 15748 6449 15750
rect 6505 15748 6529 15750
rect 6289 15728 6585 15748
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6196 14822 6224 15302
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6196 14074 6224 14758
rect 6289 14716 6585 14736
rect 6345 14714 6369 14716
rect 6425 14714 6449 14716
rect 6505 14714 6529 14716
rect 6367 14662 6369 14714
rect 6431 14662 6443 14714
rect 6505 14662 6507 14714
rect 6345 14660 6369 14662
rect 6425 14660 6449 14662
rect 6505 14660 6529 14662
rect 6289 14640 6585 14660
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6104 13926 6224 13954
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6104 12442 6132 13466
rect 6196 12850 6224 13926
rect 6289 13628 6585 13648
rect 6345 13626 6369 13628
rect 6425 13626 6449 13628
rect 6505 13626 6529 13628
rect 6367 13574 6369 13626
rect 6431 13574 6443 13626
rect 6505 13574 6507 13626
rect 6345 13572 6369 13574
rect 6425 13572 6449 13574
rect 6505 13572 6529 13574
rect 6289 13552 6585 13572
rect 6656 13462 6684 16934
rect 6748 14074 6776 23734
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 23338 6960 23462
rect 6840 23310 6960 23338
rect 6840 22574 6868 23310
rect 6920 23044 6972 23050
rect 6920 22986 6972 22992
rect 6932 22574 6960 22986
rect 6828 22568 6880 22574
rect 6828 22510 6880 22516
rect 6920 22568 6972 22574
rect 6920 22510 6972 22516
rect 7024 21010 7052 28970
rect 7288 28620 7340 28626
rect 7288 28562 7340 28568
rect 7300 28218 7328 28562
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 7300 27674 7328 28154
rect 7288 27668 7340 27674
rect 7288 27610 7340 27616
rect 7484 27033 7512 29718
rect 7668 27441 7696 34682
rect 7760 34649 7788 39520
rect 8220 35714 8248 39520
rect 8128 35686 8248 35714
rect 7932 34944 7984 34950
rect 7932 34886 7984 34892
rect 7746 34640 7802 34649
rect 7746 34575 7802 34584
rect 7944 34542 7972 34886
rect 7932 34536 7984 34542
rect 7932 34478 7984 34484
rect 7840 33924 7892 33930
rect 7840 33866 7892 33872
rect 7852 33454 7880 33866
rect 7840 33448 7892 33454
rect 7840 33390 7892 33396
rect 7746 33144 7802 33153
rect 7746 33079 7802 33088
rect 7760 32910 7788 33079
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7852 32366 7880 33390
rect 7944 32570 7972 34478
rect 8024 33108 8076 33114
rect 8024 33050 8076 33056
rect 8036 33017 8064 33050
rect 8022 33008 8078 33017
rect 8022 32943 8078 32952
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 7840 32360 7892 32366
rect 7840 32302 7892 32308
rect 8024 32360 8076 32366
rect 8024 32302 8076 32308
rect 7852 31686 7880 32302
rect 7932 31816 7984 31822
rect 7932 31758 7984 31764
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7748 31136 7800 31142
rect 7748 31078 7800 31084
rect 7852 31090 7880 31622
rect 7944 31482 7972 31758
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 8036 31385 8064 32302
rect 8022 31376 8078 31385
rect 8022 31311 8078 31320
rect 7654 27432 7710 27441
rect 7654 27367 7710 27376
rect 7470 27024 7526 27033
rect 7470 26959 7526 26968
rect 7196 26852 7248 26858
rect 7196 26794 7248 26800
rect 7208 26586 7236 26794
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 7484 25906 7512 26959
rect 7472 25900 7524 25906
rect 7472 25842 7524 25848
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 7300 25498 7328 25638
rect 7288 25492 7340 25498
rect 7288 25434 7340 25440
rect 7196 24064 7248 24070
rect 7196 24006 7248 24012
rect 7208 23322 7236 24006
rect 7196 23316 7248 23322
rect 7196 23258 7248 23264
rect 7300 22681 7328 25434
rect 7668 24750 7696 27367
rect 7760 26586 7788 31078
rect 7852 31062 7972 31090
rect 7840 29096 7892 29102
rect 7840 29038 7892 29044
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7656 24744 7708 24750
rect 7562 24712 7618 24721
rect 7656 24686 7708 24692
rect 7562 24647 7618 24656
rect 7576 24342 7604 24647
rect 7852 24596 7880 29038
rect 7944 27946 7972 31062
rect 8036 29850 8064 31311
rect 8128 30190 8156 35686
rect 8588 34066 8616 39520
rect 8956 37210 8984 39520
rect 8680 37182 8984 37210
rect 8484 34060 8536 34066
rect 8484 34002 8536 34008
rect 8576 34060 8628 34066
rect 8576 34002 8628 34008
rect 8300 32768 8352 32774
rect 8300 32710 8352 32716
rect 8312 32366 8340 32710
rect 8392 32564 8444 32570
rect 8392 32506 8444 32512
rect 8300 32360 8352 32366
rect 8300 32302 8352 32308
rect 8404 32212 8432 32506
rect 8220 32184 8432 32212
rect 8220 31346 8248 32184
rect 8496 32042 8524 34002
rect 8680 32473 8708 37182
rect 8956 37020 9252 37040
rect 9012 37018 9036 37020
rect 9092 37018 9116 37020
rect 9172 37018 9196 37020
rect 9034 36966 9036 37018
rect 9098 36966 9110 37018
rect 9172 36966 9174 37018
rect 9012 36964 9036 36966
rect 9092 36964 9116 36966
rect 9172 36964 9196 36966
rect 8956 36944 9252 36964
rect 8956 35932 9252 35952
rect 9012 35930 9036 35932
rect 9092 35930 9116 35932
rect 9172 35930 9196 35932
rect 9034 35878 9036 35930
rect 9098 35878 9110 35930
rect 9172 35878 9174 35930
rect 9012 35876 9036 35878
rect 9092 35876 9116 35878
rect 9172 35876 9196 35878
rect 8956 35856 9252 35876
rect 8760 35148 8812 35154
rect 8760 35090 8812 35096
rect 8772 34542 8800 35090
rect 8956 34844 9252 34864
rect 9012 34842 9036 34844
rect 9092 34842 9116 34844
rect 9172 34842 9196 34844
rect 9034 34790 9036 34842
rect 9098 34790 9110 34842
rect 9172 34790 9174 34842
rect 9012 34788 9036 34790
rect 9092 34788 9116 34790
rect 9172 34788 9196 34790
rect 8956 34768 9252 34788
rect 8760 34536 8812 34542
rect 8760 34478 8812 34484
rect 8666 32464 8722 32473
rect 8666 32399 8722 32408
rect 8312 32014 8524 32042
rect 8312 31482 8340 32014
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8576 31340 8628 31346
rect 8576 31282 8628 31288
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8116 30184 8168 30190
rect 8116 30126 8168 30132
rect 8024 29844 8076 29850
rect 8024 29786 8076 29792
rect 8024 29708 8076 29714
rect 8024 29650 8076 29656
rect 8036 29034 8064 29650
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8116 29232 8168 29238
rect 8116 29174 8168 29180
rect 8024 29028 8076 29034
rect 8024 28970 8076 28976
rect 7932 27940 7984 27946
rect 7932 27882 7984 27888
rect 7932 27464 7984 27470
rect 7932 27406 7984 27412
rect 7944 26926 7972 27406
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 7932 26920 7984 26926
rect 7930 26888 7932 26897
rect 7984 26888 7986 26897
rect 7930 26823 7986 26832
rect 8036 26586 8064 27270
rect 8024 26580 8076 26586
rect 8024 26522 8076 26528
rect 8128 26518 8156 29174
rect 8220 27860 8248 29582
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8404 28014 8432 28426
rect 8392 28008 8444 28014
rect 8392 27950 8444 27956
rect 8300 27872 8352 27878
rect 8220 27832 8300 27860
rect 8116 26512 8168 26518
rect 8116 26454 8168 26460
rect 7932 26376 7984 26382
rect 7932 26318 7984 26324
rect 7944 26042 7972 26318
rect 7932 26036 7984 26042
rect 7932 25978 7984 25984
rect 8128 25922 8156 26454
rect 8220 26382 8248 27832
rect 8300 27814 8352 27820
rect 8404 27674 8432 27950
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8298 27568 8354 27577
rect 8298 27503 8300 27512
rect 8352 27503 8354 27512
rect 8300 27474 8352 27480
rect 8312 27334 8340 27474
rect 8496 27418 8524 31078
rect 8588 30938 8616 31282
rect 8576 30932 8628 30938
rect 8576 30874 8628 30880
rect 8576 29028 8628 29034
rect 8680 29016 8708 32399
rect 8628 28988 8708 29016
rect 8576 28970 8628 28976
rect 8588 28422 8616 28970
rect 8576 28416 8628 28422
rect 8576 28358 8628 28364
rect 8404 27390 8524 27418
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8312 26042 8340 26522
rect 8300 26036 8352 26042
rect 8300 25978 8352 25984
rect 8128 25906 8340 25922
rect 8128 25900 8352 25906
rect 8128 25894 8300 25900
rect 8300 25842 8352 25848
rect 8208 25152 8260 25158
rect 8208 25094 8260 25100
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 7668 24568 7880 24596
rect 7932 24608 7984 24614
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7576 23798 7604 24278
rect 7564 23792 7616 23798
rect 7564 23734 7616 23740
rect 7472 23112 7524 23118
rect 7472 23054 7524 23060
rect 7286 22672 7342 22681
rect 7286 22607 7342 22616
rect 7104 22568 7156 22574
rect 7104 22510 7156 22516
rect 7116 21894 7144 22510
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 7116 21078 7144 21830
rect 7104 21072 7156 21078
rect 7104 21014 7156 21020
rect 7012 21004 7064 21010
rect 7012 20946 7064 20952
rect 7196 21004 7248 21010
rect 7196 20946 7248 20952
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20262 6868 20878
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6932 20398 6960 20810
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 7116 20466 7144 20742
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6932 19514 6960 20334
rect 7012 20324 7064 20330
rect 7012 20266 7064 20272
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7024 19310 7052 20266
rect 7208 20262 7236 20946
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 18970 7052 19246
rect 7104 19168 7156 19174
rect 7104 19110 7156 19116
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7116 18170 7144 19110
rect 7024 18142 7144 18170
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17202 6960 17478
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6932 16810 6960 17138
rect 6840 16782 6960 16810
rect 6840 16250 6868 16782
rect 6828 16244 6880 16250
rect 6828 16186 6880 16192
rect 6828 16040 6880 16046
rect 6828 15982 6880 15988
rect 6920 16040 6972 16046
rect 6920 15982 6972 15988
rect 6840 14958 6868 15982
rect 6932 15706 6960 15982
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 14952 6880 14958
rect 6828 14894 6880 14900
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 6736 14068 6788 14074
rect 6736 14010 6788 14016
rect 6748 13870 6776 14010
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13530 6868 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6472 12986 6500 13262
rect 6932 13190 6960 14418
rect 7024 13546 7052 18142
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 7116 14822 7144 15506
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7116 13682 7144 14758
rect 7208 13818 7236 20198
rect 7300 16726 7328 22607
rect 7484 22234 7512 23054
rect 7472 22228 7524 22234
rect 7472 22170 7524 22176
rect 7668 21350 7696 24568
rect 7932 24550 7984 24556
rect 7944 24410 7972 24550
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 7944 23866 7972 24142
rect 7932 23860 7984 23866
rect 7932 23802 7984 23808
rect 7944 23338 7972 23802
rect 8036 23662 8064 24754
rect 8220 24614 8248 25094
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 7852 23310 7972 23338
rect 7852 21962 7880 23310
rect 8036 23254 8064 23598
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8024 23248 8076 23254
rect 8076 23208 8156 23236
rect 8024 23190 8076 23196
rect 8022 23080 8078 23089
rect 8022 23015 8078 23024
rect 7932 22092 7984 22098
rect 7932 22034 7984 22040
rect 7840 21956 7892 21962
rect 7840 21898 7892 21904
rect 7852 21690 7880 21898
rect 7840 21684 7892 21690
rect 7840 21626 7892 21632
rect 7656 21344 7708 21350
rect 7656 21286 7708 21292
rect 7748 21072 7800 21078
rect 7562 21040 7618 21049
rect 7748 21014 7800 21020
rect 7562 20975 7618 20984
rect 7576 20942 7604 20975
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7760 20466 7788 21014
rect 7852 20942 7880 21626
rect 7944 21622 7972 22034
rect 8036 22030 8064 23015
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 7932 21616 7984 21622
rect 7932 21558 7984 21564
rect 8128 21554 8156 23208
rect 8220 22794 8248 23462
rect 8220 22778 8340 22794
rect 8220 22772 8352 22778
rect 8220 22766 8300 22772
rect 8300 22714 8352 22720
rect 8404 22658 8432 27390
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8496 26314 8524 27270
rect 8588 26353 8616 28358
rect 8772 27690 8800 34478
rect 8852 34400 8904 34406
rect 8852 34342 8904 34348
rect 8864 33998 8892 34342
rect 8852 33992 8904 33998
rect 8852 33934 8904 33940
rect 8864 33658 8892 33934
rect 8956 33756 9252 33776
rect 9012 33754 9036 33756
rect 9092 33754 9116 33756
rect 9172 33754 9196 33756
rect 9034 33702 9036 33754
rect 9098 33702 9110 33754
rect 9172 33702 9174 33754
rect 9012 33700 9036 33702
rect 9092 33700 9116 33702
rect 9172 33700 9196 33702
rect 8956 33680 9252 33700
rect 8852 33652 8904 33658
rect 8852 33594 8904 33600
rect 9310 33280 9366 33289
rect 9310 33215 9366 33224
rect 8956 32668 9252 32688
rect 9012 32666 9036 32668
rect 9092 32666 9116 32668
rect 9172 32666 9196 32668
rect 9034 32614 9036 32666
rect 9098 32614 9110 32666
rect 9172 32614 9174 32666
rect 9012 32612 9036 32614
rect 9092 32612 9116 32614
rect 9172 32612 9196 32614
rect 8956 32592 9252 32612
rect 8852 32020 8904 32026
rect 8852 31962 8904 31968
rect 8864 31278 8892 31962
rect 8956 31580 9252 31600
rect 9012 31578 9036 31580
rect 9092 31578 9116 31580
rect 9172 31578 9196 31580
rect 9034 31526 9036 31578
rect 9098 31526 9110 31578
rect 9172 31526 9174 31578
rect 9012 31524 9036 31526
rect 9092 31524 9116 31526
rect 9172 31524 9196 31526
rect 8956 31504 9252 31524
rect 8852 31272 8904 31278
rect 8852 31214 8904 31220
rect 8956 30492 9252 30512
rect 9012 30490 9036 30492
rect 9092 30490 9116 30492
rect 9172 30490 9196 30492
rect 9034 30438 9036 30490
rect 9098 30438 9110 30490
rect 9172 30438 9174 30490
rect 9012 30436 9036 30438
rect 9092 30436 9116 30438
rect 9172 30436 9196 30438
rect 8956 30416 9252 30436
rect 8852 30116 8904 30122
rect 8852 30058 8904 30064
rect 8680 27662 8800 27690
rect 8574 26344 8630 26353
rect 8484 26308 8536 26314
rect 8574 26279 8630 26288
rect 8484 26250 8536 26256
rect 8484 24608 8536 24614
rect 8484 24550 8536 24556
rect 8220 22630 8432 22658
rect 8220 22012 8248 22630
rect 8220 21984 8340 22012
rect 8116 21548 8168 21554
rect 8116 21490 8168 21496
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7852 20534 7880 20878
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7760 20058 7788 20402
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7852 19378 7880 20470
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7654 19272 7710 19281
rect 7654 19207 7710 19216
rect 7668 19174 7696 19207
rect 7656 19168 7708 19174
rect 7656 19110 7708 19116
rect 7852 18970 7880 19314
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7944 18850 7972 21286
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8128 19145 8156 19178
rect 8114 19136 8170 19145
rect 8114 19071 8170 19080
rect 7852 18822 7972 18850
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7760 17785 7788 17818
rect 7746 17776 7802 17785
rect 7746 17711 7802 17720
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 7392 16998 7420 17478
rect 7656 17196 7708 17202
rect 7656 17138 7708 17144
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7286 16552 7342 16561
rect 7286 16487 7342 16496
rect 7300 16114 7328 16487
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7392 15706 7420 16934
rect 7668 16794 7696 17138
rect 7852 16969 7880 18822
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8036 17882 8064 18566
rect 8128 18222 8156 19071
rect 8116 18216 8168 18222
rect 8116 18158 8168 18164
rect 8024 17876 8076 17882
rect 8024 17818 8076 17824
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7944 17338 7972 17614
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7838 16960 7894 16969
rect 7838 16895 7894 16904
rect 7656 16788 7708 16794
rect 7656 16730 7708 16736
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7576 15434 7604 16050
rect 7564 15428 7616 15434
rect 7564 15370 7616 15376
rect 7286 14920 7342 14929
rect 7286 14855 7342 14864
rect 7300 14550 7328 14855
rect 7378 14648 7434 14657
rect 7378 14583 7434 14592
rect 7288 14544 7340 14550
rect 7288 14486 7340 14492
rect 7392 14482 7420 14583
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7576 14414 7604 15370
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7300 13938 7328 14282
rect 7564 14272 7616 14278
rect 7668 14226 7696 16730
rect 7748 16040 7800 16046
rect 7746 16008 7748 16017
rect 7800 16008 7802 16017
rect 7746 15943 7802 15952
rect 7852 15502 7880 16895
rect 8036 16794 8064 17818
rect 8116 17740 8168 17746
rect 8116 17682 8168 17688
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7748 14816 7800 14822
rect 7852 14804 7880 15438
rect 7800 14776 7880 14804
rect 7748 14758 7800 14764
rect 7616 14220 7696 14226
rect 7564 14214 7696 14220
rect 7576 14198 7696 14214
rect 7576 13938 7604 14198
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7208 13790 7328 13818
rect 7116 13654 7236 13682
rect 7024 13518 7144 13546
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6184 12844 6236 12850
rect 6184 12786 6236 12792
rect 6182 12744 6238 12753
rect 6182 12679 6238 12688
rect 6196 12442 6224 12679
rect 6289 12540 6585 12560
rect 6345 12538 6369 12540
rect 6425 12538 6449 12540
rect 6505 12538 6529 12540
rect 6367 12486 6369 12538
rect 6431 12486 6443 12538
rect 6505 12486 6507 12538
rect 6345 12484 6369 12486
rect 6425 12484 6449 12486
rect 6505 12484 6529 12486
rect 6289 12464 6585 12484
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6656 12238 6684 13126
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6840 12442 6868 12922
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6184 11620 6236 11626
rect 6184 11562 6236 11568
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10674 6132 11086
rect 6092 10668 6144 10674
rect 6092 10610 6144 10616
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5540 7744 5592 7750
rect 5540 7686 5592 7692
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5460 6662 5488 7346
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5552 6338 5580 7686
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5644 7002 5672 7142
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5736 6458 5764 6802
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5460 6322 5580 6338
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5448 6316 5580 6322
rect 5500 6310 5580 6316
rect 5448 6258 5500 6264
rect 5460 5710 5488 6258
rect 5644 5710 5672 6326
rect 5736 5914 5764 6394
rect 6012 6186 6040 9318
rect 6104 7206 6132 10610
rect 6196 9518 6224 11562
rect 6289 11452 6585 11472
rect 6345 11450 6369 11452
rect 6425 11450 6449 11452
rect 6505 11450 6529 11452
rect 6367 11398 6369 11450
rect 6431 11398 6443 11450
rect 6505 11398 6507 11450
rect 6345 11396 6369 11398
rect 6425 11396 6449 11398
rect 6505 11396 6529 11398
rect 6289 11376 6585 11396
rect 6656 11354 6684 12174
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6748 11150 6776 11494
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6289 10364 6585 10384
rect 6345 10362 6369 10364
rect 6425 10362 6449 10364
rect 6505 10362 6529 10364
rect 6367 10310 6369 10362
rect 6431 10310 6443 10362
rect 6505 10310 6507 10362
rect 6345 10308 6369 10310
rect 6425 10308 6449 10310
rect 6505 10308 6529 10310
rect 6289 10288 6585 10308
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6840 9518 6868 10066
rect 6184 9512 6236 9518
rect 6184 9454 6236 9460
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 6289 9276 6585 9296
rect 6345 9274 6369 9276
rect 6425 9274 6449 9276
rect 6505 9274 6529 9276
rect 6367 9222 6369 9274
rect 6431 9222 6443 9274
rect 6505 9222 6507 9274
rect 6345 9220 6369 9222
rect 6425 9220 6449 9222
rect 6505 9220 6529 9222
rect 6289 9200 6585 9220
rect 6932 8480 6960 13126
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7024 9654 7052 12310
rect 7116 10418 7144 13518
rect 7208 12374 7236 13654
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7196 12232 7248 12238
rect 7300 12209 7328 13790
rect 7380 13456 7432 13462
rect 7380 13398 7432 13404
rect 7392 12986 7420 13398
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7484 12782 7512 13126
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7196 12174 7248 12180
rect 7286 12200 7342 12209
rect 7208 11898 7236 12174
rect 7286 12135 7342 12144
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7392 11694 7420 12038
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7380 10532 7432 10538
rect 7380 10474 7432 10480
rect 7288 10464 7340 10470
rect 7116 10390 7236 10418
rect 7392 10441 7420 10474
rect 7288 10406 7340 10412
rect 7378 10432 7434 10441
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7116 9722 7144 10202
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6932 8452 7144 8480
rect 6552 8424 6604 8430
rect 6550 8392 6552 8401
rect 6604 8392 6606 8401
rect 6550 8327 6606 8336
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6289 8188 6585 8208
rect 6345 8186 6369 8188
rect 6425 8186 6449 8188
rect 6505 8186 6529 8188
rect 6367 8134 6369 8186
rect 6431 8134 6443 8186
rect 6505 8134 6507 8186
rect 6345 8132 6369 8134
rect 6425 8132 6449 8134
rect 6505 8132 6529 8134
rect 6289 8112 6585 8132
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 7410 6592 7686
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6840 7206 6868 7822
rect 6932 7342 6960 8298
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6104 6390 6132 7142
rect 6289 7100 6585 7120
rect 6345 7098 6369 7100
rect 6425 7098 6449 7100
rect 6505 7098 6529 7100
rect 6367 7046 6369 7098
rect 6431 7046 6443 7098
rect 6505 7046 6507 7098
rect 6345 7044 6369 7046
rect 6425 7044 6449 7046
rect 6505 7044 6529 7046
rect 6289 7024 6585 7044
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6000 6180 6052 6186
rect 6000 6122 6052 6128
rect 6736 6112 6788 6118
rect 5814 6080 5870 6089
rect 6736 6054 6788 6060
rect 5814 6015 5870 6024
rect 5724 5908 5776 5914
rect 5724 5850 5776 5856
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5356 5160 5408 5166
rect 5276 5108 5356 5114
rect 5276 5102 5408 5108
rect 5276 5086 5396 5102
rect 5172 3664 5224 3670
rect 5172 3606 5224 3612
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4804 3528 4856 3534
rect 4526 3496 4582 3505
rect 4804 3470 4856 3476
rect 4526 3431 4582 3440
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4540 480 4568 3431
rect 4816 2990 4844 3470
rect 4988 3460 5040 3466
rect 4988 3402 5040 3408
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4816 2514 4844 2926
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5000 480 5028 3402
rect 5092 2922 5120 3538
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 5092 2009 5120 2858
rect 5276 2650 5304 5086
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5460 4826 5488 5646
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 4826 5580 5510
rect 5644 5370 5672 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5446 4584 5502 4593
rect 5828 4554 5856 6015
rect 6289 6012 6585 6032
rect 6345 6010 6369 6012
rect 6425 6010 6449 6012
rect 6505 6010 6529 6012
rect 6367 5958 6369 6010
rect 6431 5958 6443 6010
rect 6505 5958 6507 6010
rect 6345 5956 6369 5958
rect 6425 5956 6449 5958
rect 6505 5956 6529 5958
rect 6289 5936 6585 5956
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6012 4758 6040 5782
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6000 4752 6052 4758
rect 6000 4694 6052 4700
rect 5446 4519 5502 4528
rect 5816 4548 5868 4554
rect 5460 4078 5488 4519
rect 5816 4490 5868 4496
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5644 4146 5672 4422
rect 6012 4214 6040 4694
rect 6000 4208 6052 4214
rect 6000 4150 6052 4156
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 4004 5408 4010
rect 5356 3946 5408 3952
rect 5368 3738 5396 3946
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5354 2816 5410 2825
rect 5354 2751 5410 2760
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5170 2544 5226 2553
rect 5170 2479 5172 2488
rect 5224 2479 5226 2488
rect 5172 2450 5224 2456
rect 5078 2000 5134 2009
rect 5078 1935 5134 1944
rect 5368 480 5396 2751
rect 5460 2378 5488 4014
rect 5644 3194 5672 4082
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 5736 480 5764 4082
rect 6104 1442 6132 4966
rect 6289 4924 6585 4944
rect 6345 4922 6369 4924
rect 6425 4922 6449 4924
rect 6505 4922 6529 4924
rect 6367 4870 6369 4922
rect 6431 4870 6443 4922
rect 6505 4870 6507 4922
rect 6345 4868 6369 4870
rect 6425 4868 6449 4870
rect 6505 4868 6529 4870
rect 6289 4848 6585 4868
rect 6656 4622 6684 5850
rect 6644 4616 6696 4622
rect 6644 4558 6696 4564
rect 6656 4282 6684 4558
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6552 4208 6604 4214
rect 6552 4150 6604 4156
rect 6564 4010 6592 4150
rect 6748 4128 6776 6054
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6840 4282 6868 4762
rect 6932 4758 6960 7142
rect 7024 5846 7052 7686
rect 7012 5840 7064 5846
rect 7116 5817 7144 8452
rect 7012 5782 7064 5788
rect 7102 5808 7158 5817
rect 7102 5743 7158 5752
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6828 4276 6880 4282
rect 6828 4218 6880 4224
rect 7024 4214 7052 4966
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 6920 4140 6972 4146
rect 6748 4100 6920 4128
rect 6920 4082 6972 4088
rect 6642 4040 6698 4049
rect 6552 4004 6604 4010
rect 6642 3975 6698 3984
rect 6552 3946 6604 3952
rect 6289 3836 6585 3856
rect 6345 3834 6369 3836
rect 6425 3834 6449 3836
rect 6505 3834 6529 3836
rect 6367 3782 6369 3834
rect 6431 3782 6443 3834
rect 6505 3782 6507 3834
rect 6345 3780 6369 3782
rect 6425 3780 6449 3782
rect 6505 3780 6529 3782
rect 6289 3760 6585 3780
rect 6656 3602 6684 3975
rect 6932 3738 6960 4082
rect 7116 4078 7144 5510
rect 7208 5370 7236 10390
rect 7300 8072 7328 10406
rect 7378 10367 7434 10376
rect 7378 10160 7434 10169
rect 7378 10095 7380 10104
rect 7432 10095 7434 10104
rect 7380 10066 7432 10072
rect 7380 9036 7432 9042
rect 7380 8978 7432 8984
rect 7392 8362 7420 8978
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7300 8044 7420 8072
rect 7392 7993 7420 8044
rect 7378 7984 7434 7993
rect 7288 7948 7340 7954
rect 7378 7919 7434 7928
rect 7288 7890 7340 7896
rect 7300 7274 7328 7890
rect 7288 7268 7340 7274
rect 7288 7210 7340 7216
rect 7300 7002 7328 7210
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7208 5166 7236 5306
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6920 3732 6972 3738
rect 6920 3674 6972 3680
rect 6644 3596 6696 3602
rect 6644 3538 6696 3544
rect 6656 3194 6684 3538
rect 7116 3194 7144 4014
rect 7300 3602 7328 6938
rect 7484 6458 7512 12582
rect 7576 11286 7604 13874
rect 7654 13832 7710 13841
rect 7654 13767 7710 13776
rect 7668 12646 7696 13767
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7668 11694 7696 12378
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7668 11354 7696 11630
rect 7656 11348 7708 11354
rect 7656 11290 7708 11296
rect 7564 11280 7616 11286
rect 7564 11222 7616 11228
rect 7576 10674 7604 11222
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7576 10198 7604 10610
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7576 9722 7604 10134
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7760 9489 7788 14758
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7852 14074 7880 14486
rect 7840 14068 7892 14074
rect 7840 14010 7892 14016
rect 7852 13977 7880 14010
rect 7838 13968 7894 13977
rect 7838 13903 7894 13912
rect 7838 13696 7894 13705
rect 7838 13631 7894 13640
rect 7852 12714 7880 13631
rect 7840 12708 7892 12714
rect 7840 12650 7892 12656
rect 7746 9480 7802 9489
rect 7564 9444 7616 9450
rect 7746 9415 7802 9424
rect 7564 9386 7616 9392
rect 7576 8838 7604 9386
rect 7760 9042 7788 9415
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 7852 8922 7880 12650
rect 7760 8894 7880 8922
rect 7564 8832 7616 8838
rect 7564 8774 7616 8780
rect 7576 8362 7604 8774
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7380 5636 7432 5642
rect 7380 5578 7432 5584
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 6642 3088 6698 3097
rect 6642 3023 6698 3032
rect 6918 3088 6974 3097
rect 6918 3023 6974 3032
rect 6289 2748 6585 2768
rect 6345 2746 6369 2748
rect 6425 2746 6449 2748
rect 6505 2746 6529 2748
rect 6367 2694 6369 2746
rect 6431 2694 6443 2746
rect 6505 2694 6507 2746
rect 6345 2692 6369 2694
rect 6425 2692 6449 2694
rect 6505 2692 6529 2694
rect 6289 2672 6585 2692
rect 6104 1414 6224 1442
rect 6196 480 6224 1414
rect 6656 1034 6684 3023
rect 6564 1006 6684 1034
rect 6564 480 6592 1006
rect 6932 480 6960 3023
rect 7102 2952 7158 2961
rect 7102 2887 7158 2896
rect 7116 2650 7144 2887
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7392 480 7420 5578
rect 7484 2825 7512 6122
rect 7576 5556 7604 8298
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 7410 7696 7686
rect 7760 7546 7788 8894
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 7852 8498 7880 8774
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7656 7404 7708 7410
rect 7656 7346 7708 7352
rect 7760 6202 7788 7482
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 7002 7880 7278
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7760 6174 7880 6202
rect 7656 6112 7708 6118
rect 7708 6072 7788 6100
rect 7656 6054 7708 6060
rect 7656 5568 7708 5574
rect 7576 5528 7656 5556
rect 7656 5510 7708 5516
rect 7668 5302 7696 5510
rect 7656 5296 7708 5302
rect 7562 5264 7618 5273
rect 7656 5238 7708 5244
rect 7562 5199 7618 5208
rect 7576 2938 7604 5199
rect 7654 3632 7710 3641
rect 7654 3567 7710 3576
rect 7668 3534 7696 3567
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3058 7696 3470
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7576 2910 7696 2938
rect 7470 2816 7526 2825
rect 7470 2751 7526 2760
rect 7470 2680 7526 2689
rect 7668 2650 7696 2910
rect 7470 2615 7472 2624
rect 7524 2615 7526 2624
rect 7656 2644 7708 2650
rect 7472 2586 7524 2592
rect 7656 2586 7708 2592
rect 7760 480 7788 6072
rect 7852 4049 7880 6174
rect 7838 4040 7894 4049
rect 7838 3975 7894 3984
rect 7944 3516 7972 16662
rect 8024 16584 8076 16590
rect 8024 16526 8076 16532
rect 8036 15570 8064 16526
rect 8128 15910 8156 17682
rect 8220 16658 8248 19246
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8024 15564 8076 15570
rect 8024 15506 8076 15512
rect 8116 14884 8168 14890
rect 8116 14826 8168 14832
rect 8024 14816 8076 14822
rect 8024 14758 8076 14764
rect 8036 14618 8064 14758
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8128 14278 8156 14826
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8036 13530 8064 13738
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8128 13326 8156 14214
rect 8208 13728 8260 13734
rect 8208 13670 8260 13676
rect 8116 13320 8168 13326
rect 8116 13262 8168 13268
rect 8128 12850 8156 13262
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 12442 8156 12786
rect 8116 12436 8168 12442
rect 8116 12378 8168 12384
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8401 8064 8774
rect 8022 8392 8078 8401
rect 8022 8327 8078 8336
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 8036 6186 8064 8230
rect 8220 7857 8248 13670
rect 8312 8106 8340 21984
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 20806 8432 21286
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8404 19310 8432 20742
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8404 18834 8432 19110
rect 8496 18850 8524 24550
rect 8588 21350 8616 26279
rect 8680 25838 8708 27662
rect 8760 27600 8812 27606
rect 8760 27542 8812 27548
rect 8772 26926 8800 27542
rect 8864 27402 8892 30058
rect 8956 29404 9252 29424
rect 9012 29402 9036 29404
rect 9092 29402 9116 29404
rect 9172 29402 9196 29404
rect 9034 29350 9036 29402
rect 9098 29350 9110 29402
rect 9172 29350 9174 29402
rect 9012 29348 9036 29350
rect 9092 29348 9116 29350
rect 9172 29348 9196 29350
rect 8956 29328 9252 29348
rect 9036 29164 9088 29170
rect 9036 29106 9088 29112
rect 9048 28966 9076 29106
rect 9036 28960 9088 28966
rect 9036 28902 9088 28908
rect 9048 28490 9076 28902
rect 9036 28484 9088 28490
rect 9036 28426 9088 28432
rect 8956 28316 9252 28336
rect 9012 28314 9036 28316
rect 9092 28314 9116 28316
rect 9172 28314 9196 28316
rect 9034 28262 9036 28314
rect 9098 28262 9110 28314
rect 9172 28262 9174 28314
rect 9012 28260 9036 28262
rect 9092 28260 9116 28262
rect 9172 28260 9196 28262
rect 8956 28240 9252 28260
rect 9034 27704 9090 27713
rect 9034 27639 9090 27648
rect 9048 27606 9076 27639
rect 9036 27600 9088 27606
rect 9036 27542 9088 27548
rect 8852 27396 8904 27402
rect 8852 27338 8904 27344
rect 8760 26920 8812 26926
rect 8760 26862 8812 26868
rect 8864 26489 8892 27338
rect 8956 27228 9252 27248
rect 9012 27226 9036 27228
rect 9092 27226 9116 27228
rect 9172 27226 9196 27228
rect 9034 27174 9036 27226
rect 9098 27174 9110 27226
rect 9172 27174 9174 27226
rect 9012 27172 9036 27174
rect 9092 27172 9116 27174
rect 9172 27172 9196 27174
rect 8956 27152 9252 27172
rect 8942 27024 8998 27033
rect 8942 26959 8944 26968
rect 8996 26959 8998 26968
rect 8944 26930 8996 26936
rect 8956 26586 8984 26930
rect 8944 26580 8996 26586
rect 8944 26522 8996 26528
rect 8850 26480 8906 26489
rect 8850 26415 8906 26424
rect 8956 26140 9252 26160
rect 9012 26138 9036 26140
rect 9092 26138 9116 26140
rect 9172 26138 9196 26140
rect 9034 26086 9036 26138
rect 9098 26086 9110 26138
rect 9172 26086 9174 26138
rect 9012 26084 9036 26086
rect 9092 26084 9116 26086
rect 9172 26084 9196 26086
rect 8956 26064 9252 26084
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8576 21344 8628 21350
rect 8576 21286 8628 21292
rect 8680 18986 8708 25774
rect 8956 25052 9252 25072
rect 9012 25050 9036 25052
rect 9092 25050 9116 25052
rect 9172 25050 9196 25052
rect 9034 24998 9036 25050
rect 9098 24998 9110 25050
rect 9172 24998 9174 25050
rect 9012 24996 9036 24998
rect 9092 24996 9116 24998
rect 9172 24996 9196 24998
rect 8956 24976 9252 24996
rect 9324 24818 9352 33215
rect 9416 33017 9444 39520
rect 9588 35488 9640 35494
rect 9588 35430 9640 35436
rect 9496 35148 9548 35154
rect 9496 35090 9548 35096
rect 9508 34406 9536 35090
rect 9496 34400 9548 34406
rect 9496 34342 9548 34348
rect 9508 34202 9536 34342
rect 9496 34196 9548 34202
rect 9496 34138 9548 34144
rect 9402 33008 9458 33017
rect 9402 32943 9458 32952
rect 9416 32201 9444 32943
rect 9402 32192 9458 32201
rect 9402 32127 9458 32136
rect 9600 31822 9628 35430
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9692 34746 9720 35022
rect 9680 34740 9732 34746
rect 9680 34682 9732 34688
rect 9678 34640 9734 34649
rect 9678 34575 9734 34584
rect 9692 33590 9720 34575
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 9588 31816 9640 31822
rect 9588 31758 9640 31764
rect 9588 31680 9640 31686
rect 9588 31622 9640 31628
rect 9692 31634 9720 31826
rect 9784 31754 9812 39520
rect 9864 35760 9916 35766
rect 9862 35728 9864 35737
rect 9916 35728 9918 35737
rect 9862 35663 9918 35672
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9876 34202 9904 34546
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 9862 33416 9918 33425
rect 9862 33351 9918 33360
rect 9876 32842 9904 33351
rect 9956 33108 10008 33114
rect 9956 33050 10008 33056
rect 9864 32836 9916 32842
rect 9864 32778 9916 32784
rect 9968 32722 9996 33050
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 9876 32694 9996 32722
rect 9876 31929 9904 32694
rect 10060 32026 10088 32846
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 9862 31920 9918 31929
rect 9862 31855 9918 31864
rect 9772 31748 9824 31754
rect 9772 31690 9824 31696
rect 9600 31498 9628 31622
rect 9692 31606 9812 31634
rect 9600 31482 9720 31498
rect 9600 31476 9732 31482
rect 9600 31470 9680 31476
rect 9600 29594 9628 31470
rect 9680 31418 9732 31424
rect 9784 31142 9812 31606
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9772 30592 9824 30598
rect 9772 30534 9824 30540
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9385 29566 9628 29594
rect 9385 28801 9413 29566
rect 9588 29504 9640 29510
rect 9588 29446 9640 29452
rect 9600 29050 9628 29446
rect 9692 29170 9720 29990
rect 9680 29164 9732 29170
rect 9680 29106 9732 29112
rect 9600 29022 9720 29050
rect 9588 28960 9640 28966
rect 9588 28902 9640 28908
rect 9385 28792 9458 28801
rect 9385 28750 9402 28792
rect 9402 28727 9458 28736
rect 9494 27568 9550 27577
rect 9494 27503 9550 27512
rect 9508 27130 9536 27503
rect 9496 27124 9548 27130
rect 9496 27066 9548 27072
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9508 26058 9536 26250
rect 9600 26217 9628 28902
rect 9692 28218 9720 29022
rect 9680 28212 9732 28218
rect 9680 28154 9732 28160
rect 9784 27334 9812 30534
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9772 27056 9824 27062
rect 9772 26998 9824 27004
rect 9586 26208 9642 26217
rect 9586 26143 9642 26152
rect 9508 26030 9720 26058
rect 9586 25936 9642 25945
rect 9586 25871 9642 25880
rect 9600 25702 9628 25871
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9508 25294 9536 25638
rect 9692 25378 9720 26030
rect 9600 25350 9720 25378
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9508 24954 9536 25230
rect 9600 25106 9628 25350
rect 9678 25256 9734 25265
rect 9678 25191 9680 25200
rect 9732 25191 9734 25200
rect 9680 25162 9732 25168
rect 9600 25078 9720 25106
rect 9496 24948 9548 24954
rect 9496 24890 9548 24896
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8852 24744 8904 24750
rect 8852 24686 8904 24692
rect 8772 19174 8800 24686
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8680 18958 8800 18986
rect 8392 18828 8444 18834
rect 8496 18822 8708 18850
rect 8392 18770 8444 18776
rect 8404 17338 8432 18770
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8496 17610 8524 18702
rect 8588 18222 8616 18702
rect 8576 18216 8628 18222
rect 8576 18158 8628 18164
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 17678 8616 18022
rect 8576 17672 8628 17678
rect 8576 17614 8628 17620
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8588 17202 8616 17478
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8484 16108 8536 16114
rect 8484 16050 8536 16056
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 14074 8432 15846
rect 8496 14958 8524 16050
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8588 14890 8616 17138
rect 8576 14884 8628 14890
rect 8576 14826 8628 14832
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8680 13530 8708 18822
rect 8772 14482 8800 18958
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8864 14362 8892 24686
rect 9692 24274 9720 25078
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9680 24064 9732 24070
rect 9680 24006 9732 24012
rect 8956 23964 9252 23984
rect 9012 23962 9036 23964
rect 9092 23962 9116 23964
rect 9172 23962 9196 23964
rect 9034 23910 9036 23962
rect 9098 23910 9110 23962
rect 9172 23910 9174 23962
rect 9012 23908 9036 23910
rect 9092 23908 9116 23910
rect 9172 23908 9196 23910
rect 8956 23888 9252 23908
rect 9586 23216 9642 23225
rect 9586 23151 9588 23160
rect 9640 23151 9642 23160
rect 9588 23122 9640 23128
rect 9692 23089 9720 24006
rect 9678 23080 9734 23089
rect 9678 23015 9734 23024
rect 8956 22876 9252 22896
rect 9012 22874 9036 22876
rect 9092 22874 9116 22876
rect 9172 22874 9196 22876
rect 9034 22822 9036 22874
rect 9098 22822 9110 22874
rect 9172 22822 9174 22874
rect 9012 22820 9036 22822
rect 9092 22820 9116 22822
rect 9172 22820 9196 22822
rect 8956 22800 9252 22820
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 8956 21788 9252 21808
rect 9012 21786 9036 21788
rect 9092 21786 9116 21788
rect 9172 21786 9196 21788
rect 9034 21734 9036 21786
rect 9098 21734 9110 21786
rect 9172 21734 9174 21786
rect 9012 21732 9036 21734
rect 9092 21732 9116 21734
rect 9172 21732 9196 21734
rect 8956 21712 9252 21732
rect 9692 21457 9720 21830
rect 9678 21448 9734 21457
rect 9312 21412 9364 21418
rect 9678 21383 9734 21392
rect 9312 21354 9364 21360
rect 8956 20700 9252 20720
rect 9012 20698 9036 20700
rect 9092 20698 9116 20700
rect 9172 20698 9196 20700
rect 9034 20646 9036 20698
rect 9098 20646 9110 20698
rect 9172 20646 9174 20698
rect 9012 20644 9036 20646
rect 9092 20644 9116 20646
rect 9172 20644 9196 20646
rect 8956 20624 9252 20644
rect 9324 20602 9352 21354
rect 9404 20800 9456 20806
rect 9404 20742 9456 20748
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 9416 20534 9444 20742
rect 9586 20632 9642 20641
rect 9586 20567 9642 20576
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9416 20398 9444 20470
rect 9600 20466 9628 20567
rect 9588 20460 9640 20466
rect 9588 20402 9640 20408
rect 9404 20392 9456 20398
rect 9404 20334 9456 20340
rect 9586 20360 9642 20369
rect 9586 20295 9642 20304
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9508 20058 9536 20198
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 8956 19612 9252 19632
rect 9012 19610 9036 19612
rect 9092 19610 9116 19612
rect 9172 19610 9196 19612
rect 9034 19558 9036 19610
rect 9098 19558 9110 19610
rect 9172 19558 9174 19610
rect 9012 19556 9036 19558
rect 9092 19556 9116 19558
rect 9172 19556 9196 19558
rect 8956 19536 9252 19556
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 19145 9168 19246
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 9126 19136 9182 19145
rect 9126 19071 9182 19080
rect 9324 18630 9352 19178
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 8956 18524 9252 18544
rect 9012 18522 9036 18524
rect 9092 18522 9116 18524
rect 9172 18522 9196 18524
rect 9034 18470 9036 18522
rect 9098 18470 9110 18522
rect 9172 18470 9174 18522
rect 9012 18468 9036 18470
rect 9092 18468 9116 18470
rect 9172 18468 9196 18470
rect 8956 18448 9252 18468
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9232 17898 9260 18090
rect 9324 18086 9352 18566
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9232 17870 9352 17898
rect 8956 17436 9252 17456
rect 9012 17434 9036 17436
rect 9092 17434 9116 17436
rect 9172 17434 9196 17436
rect 9034 17382 9036 17434
rect 9098 17382 9110 17434
rect 9172 17382 9174 17434
rect 9012 17380 9036 17382
rect 9092 17380 9116 17382
rect 9172 17380 9196 17382
rect 8956 17360 9252 17380
rect 8942 17232 8998 17241
rect 8942 17167 8998 17176
rect 9128 17196 9180 17202
rect 8956 16998 8984 17167
rect 9128 17138 9180 17144
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 8956 16726 8984 16934
rect 8944 16720 8996 16726
rect 8944 16662 8996 16668
rect 9048 16658 9076 16934
rect 9140 16658 9168 17138
rect 9036 16652 9088 16658
rect 9036 16594 9088 16600
rect 9128 16652 9180 16658
rect 9128 16594 9180 16600
rect 8956 16348 9252 16368
rect 9012 16346 9036 16348
rect 9092 16346 9116 16348
rect 9172 16346 9196 16348
rect 9034 16294 9036 16346
rect 9098 16294 9110 16346
rect 9172 16294 9174 16346
rect 9012 16292 9036 16294
rect 9092 16292 9116 16294
rect 9172 16292 9196 16294
rect 8956 16272 9252 16292
rect 8956 15260 9252 15280
rect 9012 15258 9036 15260
rect 9092 15258 9116 15260
rect 9172 15258 9196 15260
rect 9034 15206 9036 15258
rect 9098 15206 9110 15258
rect 9172 15206 9174 15258
rect 9012 15204 9036 15206
rect 9092 15204 9116 15206
rect 9172 15204 9196 15206
rect 8956 15184 9252 15204
rect 9324 14822 9352 17870
rect 9508 17377 9536 19110
rect 9494 17368 9550 17377
rect 9494 17303 9550 17312
rect 9600 17252 9628 20295
rect 9784 17898 9812 26998
rect 9876 26926 9904 31855
rect 9956 31748 10008 31754
rect 9956 31690 10008 31696
rect 9968 31385 9996 31690
rect 9954 31376 10010 31385
rect 9954 31311 10010 31320
rect 10060 30938 10088 31962
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 9956 30184 10008 30190
rect 9956 30126 10008 30132
rect 9968 27538 9996 30126
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 10060 28762 10088 29106
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 10046 27976 10102 27985
rect 10046 27911 10048 27920
rect 10100 27911 10102 27920
rect 10048 27882 10100 27888
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9954 27432 10010 27441
rect 9954 27367 10010 27376
rect 9968 27130 9996 27367
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 9864 26920 9916 26926
rect 9864 26862 9916 26868
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 26376 9916 26382
rect 9862 26344 9864 26353
rect 9916 26344 9918 26353
rect 9862 26279 9918 26288
rect 9862 26208 9918 26217
rect 9862 26143 9918 26152
rect 9876 24410 9904 26143
rect 9968 25838 9996 26726
rect 9956 25832 10008 25838
rect 9956 25774 10008 25780
rect 9968 25498 9996 25774
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 10060 25378 10088 27270
rect 10152 27130 10180 39520
rect 10232 34060 10284 34066
rect 10232 34002 10284 34008
rect 10244 33114 10272 34002
rect 10324 33992 10376 33998
rect 10612 33946 10640 39520
rect 10692 35488 10744 35494
rect 10692 35430 10744 35436
rect 10324 33934 10376 33940
rect 10336 33590 10364 33934
rect 10428 33918 10640 33946
rect 10324 33584 10376 33590
rect 10322 33552 10324 33561
rect 10376 33552 10378 33561
rect 10322 33487 10378 33496
rect 10232 33108 10284 33114
rect 10232 33050 10284 33056
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 10336 32502 10364 32846
rect 10324 32496 10376 32502
rect 10324 32438 10376 32444
rect 10230 32328 10286 32337
rect 10230 32263 10286 32272
rect 10244 32026 10272 32263
rect 10322 32192 10378 32201
rect 10322 32127 10378 32136
rect 10336 32026 10364 32127
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10244 29850 10272 30194
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10244 29170 10272 29446
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10244 28626 10272 29106
rect 10232 28620 10284 28626
rect 10232 28562 10284 28568
rect 10244 27674 10272 28562
rect 10232 27668 10284 27674
rect 10232 27610 10284 27616
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10336 26976 10364 31962
rect 10428 27062 10456 33918
rect 10508 33856 10560 33862
rect 10508 33798 10560 33804
rect 10520 33386 10548 33798
rect 10598 33416 10654 33425
rect 10508 33380 10560 33386
rect 10598 33351 10654 33360
rect 10508 33322 10560 33328
rect 10520 33114 10548 33322
rect 10612 33318 10640 33351
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10600 33108 10652 33114
rect 10600 33050 10652 33056
rect 10612 32570 10640 33050
rect 10600 32564 10652 32570
rect 10600 32506 10652 32512
rect 10704 32230 10732 35430
rect 10784 34944 10836 34950
rect 10784 34886 10836 34892
rect 10796 34474 10824 34886
rect 10784 34468 10836 34474
rect 10784 34410 10836 34416
rect 10796 33998 10824 34410
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 33658 10824 33934
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10796 33153 10824 33254
rect 10782 33144 10838 33153
rect 10782 33079 10838 33088
rect 10782 32872 10838 32881
rect 10782 32807 10838 32816
rect 10796 32570 10824 32807
rect 10784 32564 10836 32570
rect 10784 32506 10836 32512
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10796 32026 10824 32370
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10600 31748 10652 31754
rect 10600 31690 10652 31696
rect 10506 31376 10562 31385
rect 10612 31346 10640 31690
rect 10692 31680 10744 31686
rect 10692 31622 10744 31628
rect 10506 31311 10562 31320
rect 10600 31340 10652 31346
rect 10520 31142 10548 31311
rect 10600 31282 10652 31288
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10520 30598 10548 31078
rect 10612 30938 10640 31282
rect 10600 30932 10652 30938
rect 10600 30874 10652 30880
rect 10508 30592 10560 30598
rect 10508 30534 10560 30540
rect 10704 28506 10732 31622
rect 10980 30977 11008 39520
rect 11244 34400 11296 34406
rect 11244 34342 11296 34348
rect 11256 34134 11284 34342
rect 11244 34128 11296 34134
rect 11244 34070 11296 34076
rect 11060 34060 11112 34066
rect 11060 34002 11112 34008
rect 10966 30968 11022 30977
rect 10966 30903 11022 30912
rect 11072 30802 11100 34002
rect 11256 33522 11284 34070
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 11152 33448 11204 33454
rect 11152 33390 11204 33396
rect 11164 32842 11192 33390
rect 11152 32836 11204 32842
rect 11152 32778 11204 32784
rect 11256 32774 11284 33458
rect 11244 32768 11296 32774
rect 11244 32710 11296 32716
rect 11152 32224 11204 32230
rect 11152 32166 11204 32172
rect 11060 30796 11112 30802
rect 11060 30738 11112 30744
rect 11072 29866 11100 30738
rect 10980 29838 11100 29866
rect 10980 29782 11008 29838
rect 10968 29776 11020 29782
rect 10968 29718 11020 29724
rect 10980 29306 11008 29718
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 10968 29300 11020 29306
rect 10968 29242 11020 29248
rect 10980 28558 11008 29242
rect 11072 28966 11100 29650
rect 11164 29102 11192 32166
rect 11256 32026 11284 32710
rect 11244 32020 11296 32026
rect 11244 31962 11296 31968
rect 11242 30016 11298 30025
rect 11242 29951 11298 29960
rect 11152 29096 11204 29102
rect 11152 29038 11204 29044
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 10612 28478 10732 28506
rect 10968 28552 11020 28558
rect 10968 28494 11020 28500
rect 10506 28112 10562 28121
rect 10506 28047 10562 28056
rect 10520 27878 10548 28047
rect 10508 27872 10560 27878
rect 10508 27814 10560 27820
rect 10520 27674 10548 27814
rect 10508 27668 10560 27674
rect 10508 27610 10560 27616
rect 10416 27056 10468 27062
rect 10416 26998 10468 27004
rect 10244 26948 10364 26976
rect 10138 26752 10194 26761
rect 10138 26687 10194 26696
rect 9968 25350 10088 25378
rect 9864 24404 9916 24410
rect 9864 24346 9916 24352
rect 9876 23866 9904 24346
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9864 22500 9916 22506
rect 9864 22442 9916 22448
rect 9876 21962 9904 22442
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9876 21554 9904 21898
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9876 21010 9904 21490
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9968 20040 9996 25350
rect 10152 24614 10180 26687
rect 10244 25158 10272 26948
rect 10416 26920 10468 26926
rect 10322 26888 10378 26897
rect 10416 26862 10468 26868
rect 10322 26823 10378 26832
rect 10336 26586 10364 26823
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10324 25288 10376 25294
rect 10324 25230 10376 25236
rect 10232 25152 10284 25158
rect 10232 25094 10284 25100
rect 10336 24993 10364 25230
rect 10322 24984 10378 24993
rect 10322 24919 10324 24928
rect 10376 24919 10378 24928
rect 10324 24890 10376 24896
rect 10336 24859 10364 24890
rect 10232 24812 10284 24818
rect 10232 24754 10284 24760
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10244 24206 10272 24754
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10232 24200 10284 24206
rect 10232 24142 10284 24148
rect 10244 23866 10272 24142
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10232 23860 10284 23866
rect 10232 23802 10284 23808
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 10060 21350 10088 21966
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 21146 10088 21286
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 10048 20052 10100 20058
rect 9968 20012 10048 20040
rect 10048 19994 10100 20000
rect 9956 19916 10008 19922
rect 9956 19858 10008 19864
rect 9968 18766 9996 19858
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9784 17870 9904 17898
rect 9772 17740 9824 17746
rect 9772 17682 9824 17688
rect 9416 17224 9628 17252
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 8772 14334 8892 14362
rect 8772 13818 8800 14334
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8864 13938 8892 14214
rect 8956 14172 9252 14192
rect 9012 14170 9036 14172
rect 9092 14170 9116 14172
rect 9172 14170 9196 14172
rect 9034 14118 9036 14170
rect 9098 14118 9110 14170
rect 9172 14118 9174 14170
rect 9012 14116 9036 14118
rect 9092 14116 9116 14118
rect 9172 14116 9196 14118
rect 8956 14096 9252 14116
rect 9324 14006 9352 14758
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8772 13790 8892 13818
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 8680 12986 8708 13466
rect 8772 13462 8800 13670
rect 8760 13456 8812 13462
rect 8760 13398 8812 13404
rect 8864 13394 8892 13790
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8864 13138 8892 13330
rect 8772 13110 8892 13138
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8772 12850 8800 13110
rect 8956 13084 9252 13104
rect 9012 13082 9036 13084
rect 9092 13082 9116 13084
rect 9172 13082 9196 13084
rect 9034 13030 9036 13082
rect 9098 13030 9110 13082
rect 9172 13030 9174 13082
rect 9012 13028 9036 13030
rect 9092 13028 9116 13030
rect 9172 13028 9196 13030
rect 8956 13008 9252 13028
rect 8852 12980 8904 12986
rect 8852 12922 8904 12928
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8760 12844 8812 12850
rect 8760 12786 8812 12792
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8404 12442 8432 12718
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10266 8432 10406
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8496 9081 8524 12786
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8482 9072 8538 9081
rect 8482 9007 8538 9016
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8496 8498 8524 8910
rect 8680 8634 8708 9318
rect 8864 9178 8892 12922
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 12170 8984 12718
rect 9324 12714 9352 13126
rect 9312 12708 9364 12714
rect 9312 12650 9364 12656
rect 9324 12238 9352 12650
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8956 11996 9252 12016
rect 9012 11994 9036 11996
rect 9092 11994 9116 11996
rect 9172 11994 9196 11996
rect 9034 11942 9036 11994
rect 9098 11942 9110 11994
rect 9172 11942 9174 11994
rect 9012 11940 9036 11942
rect 9092 11940 9116 11942
rect 9172 11940 9196 11942
rect 8956 11920 9252 11940
rect 9324 11898 9352 12174
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 8956 10908 9252 10928
rect 9012 10906 9036 10908
rect 9092 10906 9116 10908
rect 9172 10906 9196 10908
rect 9034 10854 9036 10906
rect 9098 10854 9110 10906
rect 9172 10854 9174 10906
rect 9012 10852 9036 10854
rect 9092 10852 9116 10854
rect 9172 10852 9196 10854
rect 8956 10832 9252 10852
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8956 9820 9252 9840
rect 9012 9818 9036 9820
rect 9092 9818 9116 9820
rect 9172 9818 9196 9820
rect 9034 9766 9036 9818
rect 9098 9766 9110 9818
rect 9172 9766 9174 9818
rect 9012 9764 9036 9766
rect 9092 9764 9116 9766
rect 9172 9764 9196 9766
rect 8956 9744 9252 9764
rect 9324 9586 9352 9862
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8758 9072 8814 9081
rect 8758 9007 8814 9016
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8312 8078 8524 8106
rect 8300 7880 8352 7886
rect 8206 7848 8262 7857
rect 8300 7822 8352 7828
rect 8206 7783 8262 7792
rect 8312 7002 8340 7822
rect 8496 7002 8524 8078
rect 8680 8022 8708 8366
rect 8772 8090 8800 9007
rect 8864 8634 8892 9114
rect 9232 8945 9260 9318
rect 9218 8936 9274 8945
rect 9218 8871 9274 8880
rect 8956 8732 9252 8752
rect 9012 8730 9036 8732
rect 9092 8730 9116 8732
rect 9172 8730 9196 8732
rect 9034 8678 9036 8730
rect 9098 8678 9110 8730
rect 9172 8678 9174 8730
rect 9012 8676 9036 8678
rect 9092 8676 9116 8678
rect 9172 8676 9196 8678
rect 8956 8656 9252 8676
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8496 6458 8524 6938
rect 8484 6452 8536 6458
rect 8536 6412 8616 6440
rect 8484 6394 8536 6400
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8036 5370 8064 5714
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8128 5234 8156 5646
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8128 5001 8156 5170
rect 8114 4992 8170 5001
rect 8114 4927 8170 4936
rect 8208 4820 8260 4826
rect 8312 4808 8340 6054
rect 8392 5092 8444 5098
rect 8496 5080 8524 6258
rect 8588 5778 8616 6412
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8576 5568 8628 5574
rect 8680 5556 8708 6054
rect 8628 5528 8708 5556
rect 8576 5510 8628 5516
rect 8444 5052 8524 5080
rect 8392 5034 8444 5040
rect 8260 4780 8340 4808
rect 8208 4762 8260 4768
rect 8024 4684 8076 4690
rect 8024 4626 8076 4632
rect 8036 4282 8064 4626
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8024 4276 8076 4282
rect 8024 4218 8076 4224
rect 8128 3670 8156 4422
rect 8220 3738 8248 4762
rect 8404 4554 8432 5034
rect 8772 4826 8800 8026
rect 8864 6866 8892 8570
rect 8956 7644 9252 7664
rect 9012 7642 9036 7644
rect 9092 7642 9116 7644
rect 9172 7642 9196 7644
rect 9034 7590 9036 7642
rect 9098 7590 9110 7642
rect 9172 7590 9174 7642
rect 9012 7588 9036 7590
rect 9092 7588 9116 7590
rect 9172 7588 9196 7590
rect 8956 7568 9252 7588
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 8956 6905 8984 7142
rect 8942 6896 8998 6905
rect 8852 6860 8904 6866
rect 8942 6831 8998 6840
rect 8852 6802 8904 6808
rect 9140 6798 9168 7346
rect 9416 6905 9444 17224
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9692 17082 9720 17138
rect 9508 17054 9720 17082
rect 9508 15978 9536 17054
rect 9680 16992 9732 16998
rect 9678 16960 9680 16969
rect 9732 16960 9734 16969
rect 9784 16946 9812 17682
rect 9734 16918 9812 16946
rect 9678 16895 9734 16904
rect 9588 16720 9640 16726
rect 9588 16662 9640 16668
rect 9680 16720 9732 16726
rect 9680 16662 9732 16668
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15706 9536 15914
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9600 15586 9628 16662
rect 9692 16250 9720 16662
rect 9876 16266 9904 17870
rect 9968 17066 9996 18702
rect 10152 17762 10180 23802
rect 10336 23526 10364 24210
rect 10324 23520 10376 23526
rect 10324 23462 10376 23468
rect 10232 23180 10284 23186
rect 10232 23122 10284 23128
rect 10244 22030 10272 23122
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 10244 21690 10272 21966
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10232 20256 10284 20262
rect 10232 20198 10284 20204
rect 10060 17734 10180 17762
rect 10060 17270 10088 17734
rect 10140 17672 10192 17678
rect 10244 17649 10272 20198
rect 10140 17614 10192 17620
rect 10230 17640 10286 17649
rect 10152 17338 10180 17614
rect 10230 17575 10286 17584
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10048 17264 10100 17270
rect 10048 17206 10100 17212
rect 10060 17134 10088 17206
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16238 9904 16266
rect 9508 15558 9628 15586
rect 9680 15564 9732 15570
rect 9508 8514 9536 15558
rect 9680 15506 9732 15512
rect 9692 15450 9720 15506
rect 9600 15422 9720 15450
rect 9600 14618 9628 15422
rect 9784 14657 9812 16238
rect 9862 16144 9918 16153
rect 9862 16079 9918 16088
rect 9876 15706 9904 16079
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9770 14648 9826 14657
rect 9588 14612 9640 14618
rect 9770 14583 9826 14592
rect 9588 14554 9640 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 11121 9628 14418
rect 9968 13394 9996 17002
rect 10060 16561 10088 17070
rect 10152 16794 10180 17274
rect 10336 17066 10364 23462
rect 10428 19990 10456 26862
rect 10508 26784 10560 26790
rect 10612 26761 10640 28478
rect 10692 28416 10744 28422
rect 10692 28358 10744 28364
rect 10704 28082 10732 28358
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10980 28014 11008 28494
rect 10968 28008 11020 28014
rect 10968 27950 11020 27956
rect 10980 27470 11008 27950
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 10784 27124 10836 27130
rect 10784 27066 10836 27072
rect 10690 27024 10746 27033
rect 10690 26959 10746 26968
rect 10508 26726 10560 26732
rect 10598 26752 10654 26761
rect 10520 26382 10548 26726
rect 10598 26687 10654 26696
rect 10704 26602 10732 26959
rect 10612 26586 10732 26602
rect 10612 26580 10744 26586
rect 10612 26574 10692 26580
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10612 26042 10640 26574
rect 10692 26522 10744 26528
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10704 26042 10732 26386
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10612 25294 10640 25978
rect 10796 25922 10824 27066
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26382 10916 26930
rect 10980 26790 11008 27406
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 10876 26376 10928 26382
rect 10876 26318 10928 26324
rect 10704 25894 10824 25922
rect 10600 25288 10652 25294
rect 10600 25230 10652 25236
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10520 21146 10548 25094
rect 10704 22556 10732 25894
rect 10888 25498 10916 26318
rect 10980 25770 11008 26726
rect 10968 25764 11020 25770
rect 10968 25706 11020 25712
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10796 22658 10824 25230
rect 10888 24818 10916 25434
rect 10876 24812 10928 24818
rect 10876 24754 10928 24760
rect 10888 24410 10916 24754
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10980 24206 11008 25706
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 11072 24818 11100 25298
rect 11060 24812 11112 24818
rect 11060 24754 11112 24760
rect 10968 24200 11020 24206
rect 10968 24142 11020 24148
rect 10980 23526 11008 24142
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10980 23254 11008 23462
rect 11072 23322 11100 23802
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10968 23248 11020 23254
rect 10968 23190 11020 23196
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 10888 22778 10916 23122
rect 10876 22772 10928 22778
rect 10876 22714 10928 22720
rect 10796 22630 10916 22658
rect 10704 22528 10824 22556
rect 10796 22030 10824 22528
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10520 19854 10548 20266
rect 10416 19848 10468 19854
rect 10416 19790 10468 19796
rect 10508 19848 10560 19854
rect 10508 19790 10560 19796
rect 10428 18630 10456 19790
rect 10520 19514 10548 19790
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10416 18624 10468 18630
rect 10416 18566 10468 18572
rect 10428 17105 10456 18566
rect 10414 17096 10470 17105
rect 10324 17060 10376 17066
rect 10414 17031 10470 17040
rect 10324 17002 10376 17008
rect 10140 16788 10192 16794
rect 10336 16776 10364 17002
rect 10140 16730 10192 16736
rect 10244 16748 10364 16776
rect 10046 16552 10102 16561
rect 10102 16510 10180 16538
rect 10046 16487 10102 16496
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 10060 16250 10088 16390
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10046 16008 10102 16017
rect 10046 15943 10102 15952
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12442 9996 13330
rect 9956 12436 10008 12442
rect 9956 12378 10008 12384
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 9968 11898 9996 12106
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 9586 11112 9642 11121
rect 9586 11047 9642 11056
rect 9968 10266 9996 11834
rect 9956 10260 10008 10266
rect 9876 10220 9956 10248
rect 9876 9722 9904 10220
rect 9956 10202 10008 10208
rect 10060 10146 10088 15943
rect 9968 10118 10088 10146
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9680 9580 9732 9586
rect 9680 9522 9732 9528
rect 9692 9178 9720 9522
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9876 9110 9904 9658
rect 9864 9104 9916 9110
rect 9968 9081 9996 10118
rect 10046 10024 10102 10033
rect 10046 9959 10102 9968
rect 9864 9046 9916 9052
rect 9954 9072 10010 9081
rect 9954 9007 9956 9016
rect 10008 9007 10010 9016
rect 9956 8978 10008 8984
rect 9968 8566 9996 8978
rect 9956 8560 10008 8566
rect 9508 8486 9628 8514
rect 9956 8502 10008 8508
rect 9600 8430 9628 8486
rect 9588 8424 9640 8430
rect 9640 8372 9812 8378
rect 9588 8366 9812 8372
rect 9600 8350 9812 8366
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9402 6896 9458 6905
rect 9312 6860 9364 6866
rect 9402 6831 9458 6840
rect 9312 6802 9364 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6322 8892 6598
rect 8956 6556 9252 6576
rect 9012 6554 9036 6556
rect 9092 6554 9116 6556
rect 9172 6554 9196 6556
rect 9034 6502 9036 6554
rect 9098 6502 9110 6554
rect 9172 6502 9174 6554
rect 9012 6500 9036 6502
rect 9092 6500 9116 6502
rect 9172 6500 9196 6502
rect 8956 6480 9252 6500
rect 9324 6458 9352 6802
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 9310 6216 9366 6225
rect 9310 6151 9366 6160
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8208 3732 8260 3738
rect 8208 3674 8260 3680
rect 8116 3664 8168 3670
rect 8116 3606 8168 3612
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7852 3488 7972 3516
rect 7852 2310 7880 3488
rect 7930 3224 7986 3233
rect 7930 3159 7986 3168
rect 7944 2990 7972 3159
rect 8036 3058 8064 3538
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7944 2553 7972 2926
rect 7930 2544 7986 2553
rect 7930 2479 7986 2488
rect 8404 2428 8432 4218
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8666 3904 8722 3913
rect 8588 2446 8616 3878
rect 8666 3839 8722 3848
rect 8220 2400 8432 2428
rect 8576 2440 8628 2446
rect 7840 2304 7892 2310
rect 7840 2246 7892 2252
rect 8220 480 8248 2400
rect 8576 2382 8628 2388
rect 8680 1034 8708 3839
rect 8772 3738 8800 4762
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 8772 3369 8800 3470
rect 8758 3360 8814 3369
rect 8758 3295 8814 3304
rect 8864 1442 8892 6054
rect 8956 5468 9252 5488
rect 9012 5466 9036 5468
rect 9092 5466 9116 5468
rect 9172 5466 9196 5468
rect 9034 5414 9036 5466
rect 9098 5414 9110 5466
rect 9172 5414 9174 5466
rect 9012 5412 9036 5414
rect 9092 5412 9116 5414
rect 9172 5412 9196 5414
rect 8956 5392 9252 5412
rect 9324 5098 9352 6151
rect 9508 5370 9536 6734
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9312 5092 9364 5098
rect 9312 5034 9364 5040
rect 8956 4380 9252 4400
rect 9012 4378 9036 4380
rect 9092 4378 9116 4380
rect 9172 4378 9196 4380
rect 9034 4326 9036 4378
rect 9098 4326 9110 4378
rect 9172 4326 9174 4378
rect 9012 4324 9036 4326
rect 9092 4324 9116 4326
rect 9172 4324 9196 4326
rect 8956 4304 9252 4324
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9140 3670 9168 4082
rect 9128 3664 9180 3670
rect 9128 3606 9180 3612
rect 8956 3292 9252 3312
rect 9012 3290 9036 3292
rect 9092 3290 9116 3292
rect 9172 3290 9196 3292
rect 9034 3238 9036 3290
rect 9098 3238 9110 3290
rect 9172 3238 9174 3290
rect 9012 3236 9036 3238
rect 9092 3236 9116 3238
rect 9172 3236 9196 3238
rect 8956 3216 9252 3236
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 9048 2446 9076 2858
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8956 2204 9252 2224
rect 9012 2202 9036 2204
rect 9092 2202 9116 2204
rect 9172 2202 9196 2204
rect 9034 2150 9036 2202
rect 9098 2150 9110 2202
rect 9172 2150 9174 2202
rect 9012 2148 9036 2150
rect 9092 2148 9116 2150
rect 9172 2148 9196 2150
rect 8956 2128 9252 2148
rect 8864 1414 8984 1442
rect 8588 1006 8708 1034
rect 8588 480 8616 1006
rect 8956 480 8984 1414
rect 9324 1034 9352 5034
rect 9600 4978 9628 8026
rect 9680 6180 9732 6186
rect 9680 6122 9732 6128
rect 9692 5846 9720 6122
rect 9680 5840 9732 5846
rect 9678 5808 9680 5817
rect 9732 5808 9734 5817
rect 9678 5743 9734 5752
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9508 4950 9628 4978
rect 9508 4690 9536 4950
rect 9692 4842 9720 5578
rect 9600 4814 9720 4842
rect 9600 4758 9628 4814
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9496 4684 9548 4690
rect 9496 4626 9548 4632
rect 9494 4176 9550 4185
rect 9494 4111 9550 4120
rect 9404 3936 9456 3942
rect 9508 3924 9536 4111
rect 9600 4078 9628 4694
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4072 9640 4078
rect 9588 4014 9640 4020
rect 9456 3896 9536 3924
rect 9404 3878 9456 3884
rect 9508 3738 9536 3896
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9416 2582 9444 3606
rect 9496 2848 9548 2854
rect 9496 2790 9548 2796
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9508 2514 9536 2790
rect 9600 2650 9628 3674
rect 9692 3194 9720 4558
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9324 1006 9444 1034
rect 9416 480 9444 1006
rect 9784 480 9812 8350
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 3641 9904 6054
rect 9968 3777 9996 6598
rect 10060 4162 10088 9959
rect 10152 9178 10180 16510
rect 10244 16017 10272 16748
rect 10230 16008 10286 16017
rect 10230 15943 10286 15952
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10336 15162 10364 15438
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10244 14074 10272 14894
rect 10336 14618 10364 15098
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10428 14498 10456 17031
rect 10506 16688 10562 16697
rect 10506 16623 10508 16632
rect 10560 16623 10562 16632
rect 10508 16594 10560 16600
rect 10520 15706 10548 16594
rect 10508 15700 10560 15706
rect 10612 15688 10640 21966
rect 10784 21888 10836 21894
rect 10782 21856 10784 21865
rect 10836 21856 10838 21865
rect 10782 21791 10838 21800
rect 10796 21486 10824 21791
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10796 20398 10824 21082
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10704 19281 10732 19994
rect 10796 19417 10824 20334
rect 10782 19408 10838 19417
rect 10782 19343 10784 19352
rect 10836 19343 10838 19352
rect 10784 19314 10836 19320
rect 10690 19272 10746 19281
rect 10690 19207 10746 19216
rect 10782 17640 10838 17649
rect 10782 17575 10838 17584
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17202 10732 17478
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10704 16794 10732 17138
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10612 15660 10732 15688
rect 10508 15642 10560 15648
rect 10520 15502 10548 15642
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10520 15094 10548 15438
rect 10508 15088 10560 15094
rect 10508 15030 10560 15036
rect 10704 14521 10732 15660
rect 10796 14958 10824 17575
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10336 14470 10456 14498
rect 10690 14512 10746 14521
rect 10600 14476 10652 14482
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10244 13870 10272 14010
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10244 9178 10272 13806
rect 10336 13326 10364 14470
rect 10690 14447 10746 14456
rect 10600 14418 10652 14424
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10428 14074 10456 14350
rect 10416 14068 10468 14074
rect 10416 14010 10468 14016
rect 10506 13968 10562 13977
rect 10506 13903 10562 13912
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12628 10364 13262
rect 10416 12640 10468 12646
rect 10336 12600 10416 12628
rect 10416 12582 10468 12588
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10152 8537 10180 9114
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10138 8528 10194 8537
rect 10138 8463 10194 8472
rect 10152 8090 10180 8463
rect 10244 8090 10272 8842
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10230 7848 10286 7857
rect 10230 7783 10286 7792
rect 10244 7206 10272 7783
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10336 6769 10364 12378
rect 10428 7313 10456 12582
rect 10414 7304 10470 7313
rect 10414 7239 10470 7248
rect 10322 6760 10378 6769
rect 10322 6695 10378 6704
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10152 4570 10180 6054
rect 10336 5250 10364 6695
rect 10244 5222 10364 5250
rect 10244 4690 10272 5222
rect 10324 5160 10376 5166
rect 10322 5128 10324 5137
rect 10376 5128 10378 5137
rect 10322 5063 10378 5072
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10428 4622 10456 7239
rect 10520 6186 10548 13903
rect 10612 13530 10640 14418
rect 10600 13524 10652 13530
rect 10600 13466 10652 13472
rect 10704 13410 10732 14447
rect 10796 14414 10824 14758
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10796 14278 10824 14350
rect 10784 14272 10836 14278
rect 10784 14214 10836 14220
rect 10796 14006 10824 14214
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10888 13818 10916 22630
rect 10980 19854 11008 23190
rect 11164 21049 11192 27610
rect 11256 22148 11284 29951
rect 11348 27878 11376 39520
rect 11808 37754 11836 39520
rect 11440 37726 11836 37754
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 11336 27600 11388 27606
rect 11336 27542 11388 27548
rect 11348 27130 11376 27542
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11440 22148 11468 37726
rect 11622 37564 11918 37584
rect 11678 37562 11702 37564
rect 11758 37562 11782 37564
rect 11838 37562 11862 37564
rect 11700 37510 11702 37562
rect 11764 37510 11776 37562
rect 11838 37510 11840 37562
rect 11678 37508 11702 37510
rect 11758 37508 11782 37510
rect 11838 37508 11862 37510
rect 11622 37488 11918 37508
rect 11622 36476 11918 36496
rect 11678 36474 11702 36476
rect 11758 36474 11782 36476
rect 11838 36474 11862 36476
rect 11700 36422 11702 36474
rect 11764 36422 11776 36474
rect 11838 36422 11840 36474
rect 11678 36420 11702 36422
rect 11758 36420 11782 36422
rect 11838 36420 11862 36422
rect 11622 36400 11918 36420
rect 11622 35388 11918 35408
rect 11678 35386 11702 35388
rect 11758 35386 11782 35388
rect 11838 35386 11862 35388
rect 11700 35334 11702 35386
rect 11764 35334 11776 35386
rect 11838 35334 11840 35386
rect 11678 35332 11702 35334
rect 11758 35332 11782 35334
rect 11838 35332 11862 35334
rect 11622 35312 11918 35332
rect 12072 34604 12124 34610
rect 12072 34546 12124 34552
rect 11622 34300 11918 34320
rect 11678 34298 11702 34300
rect 11758 34298 11782 34300
rect 11838 34298 11862 34300
rect 11700 34246 11702 34298
rect 11764 34246 11776 34298
rect 11838 34246 11840 34298
rect 11678 34244 11702 34246
rect 11758 34244 11782 34246
rect 11838 34244 11862 34246
rect 11622 34224 11918 34244
rect 12084 34134 12112 34546
rect 12072 34128 12124 34134
rect 12072 34070 12124 34076
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 11808 33658 11836 34002
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 11622 33212 11918 33232
rect 11678 33210 11702 33212
rect 11758 33210 11782 33212
rect 11838 33210 11862 33212
rect 11700 33158 11702 33210
rect 11764 33158 11776 33210
rect 11838 33158 11840 33210
rect 11678 33156 11702 33158
rect 11758 33156 11782 33158
rect 11838 33156 11862 33158
rect 11622 33136 11918 33156
rect 11520 33040 11572 33046
rect 11520 32982 11572 32988
rect 11532 32026 11560 32982
rect 12072 32836 12124 32842
rect 12072 32778 12124 32784
rect 11796 32768 11848 32774
rect 11796 32710 11848 32716
rect 11808 32570 11836 32710
rect 12084 32570 12112 32778
rect 11796 32564 11848 32570
rect 11796 32506 11848 32512
rect 12072 32564 12124 32570
rect 12072 32506 12124 32512
rect 11622 32124 11918 32144
rect 11678 32122 11702 32124
rect 11758 32122 11782 32124
rect 11838 32122 11862 32124
rect 11700 32070 11702 32122
rect 11764 32070 11776 32122
rect 11838 32070 11840 32122
rect 11678 32068 11702 32070
rect 11758 32068 11782 32070
rect 11838 32068 11862 32070
rect 11622 32048 11918 32068
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 12072 31680 12124 31686
rect 12072 31622 12124 31628
rect 11622 31036 11918 31056
rect 11678 31034 11702 31036
rect 11758 31034 11782 31036
rect 11838 31034 11862 31036
rect 11700 30982 11702 31034
rect 11764 30982 11776 31034
rect 11838 30982 11840 31034
rect 11678 30980 11702 30982
rect 11758 30980 11782 30982
rect 11838 30980 11862 30982
rect 11622 30960 11918 30980
rect 12084 30870 12112 31622
rect 12072 30864 12124 30870
rect 12072 30806 12124 30812
rect 11612 30796 11664 30802
rect 11612 30738 11664 30744
rect 11624 30394 11652 30738
rect 12084 30394 12112 30806
rect 11612 30388 11664 30394
rect 11612 30330 11664 30336
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 11622 29948 11918 29968
rect 11678 29946 11702 29948
rect 11758 29946 11782 29948
rect 11838 29946 11862 29948
rect 11700 29894 11702 29946
rect 11764 29894 11776 29946
rect 11838 29894 11840 29946
rect 11678 29892 11702 29894
rect 11758 29892 11782 29894
rect 11838 29892 11862 29894
rect 11622 29872 11918 29892
rect 11980 29028 12032 29034
rect 11980 28970 12032 28976
rect 11992 28914 12020 28970
rect 11992 28886 12112 28914
rect 11622 28860 11918 28880
rect 11678 28858 11702 28860
rect 11758 28858 11782 28860
rect 11838 28858 11862 28860
rect 11700 28806 11702 28858
rect 11764 28806 11776 28858
rect 11838 28806 11840 28858
rect 11678 28804 11702 28806
rect 11758 28804 11782 28806
rect 11838 28804 11862 28806
rect 11622 28784 11918 28804
rect 11622 27772 11918 27792
rect 11678 27770 11702 27772
rect 11758 27770 11782 27772
rect 11838 27770 11862 27772
rect 11700 27718 11702 27770
rect 11764 27718 11776 27770
rect 11838 27718 11840 27770
rect 11678 27716 11702 27718
rect 11758 27716 11782 27718
rect 11838 27716 11862 27718
rect 11622 27696 11918 27716
rect 12084 27713 12112 28886
rect 12070 27704 12126 27713
rect 12176 27674 12204 39520
rect 12348 35080 12400 35086
rect 12348 35022 12400 35028
rect 12360 34746 12388 35022
rect 12348 34740 12400 34746
rect 12348 34682 12400 34688
rect 12360 34542 12388 34682
rect 12348 34536 12400 34542
rect 12348 34478 12400 34484
rect 12440 34400 12492 34406
rect 12440 34342 12492 34348
rect 12452 33454 12480 34342
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12348 33312 12400 33318
rect 12348 33254 12400 33260
rect 12360 33046 12388 33254
rect 12348 33040 12400 33046
rect 12348 32982 12400 32988
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12256 32564 12308 32570
rect 12256 32506 12308 32512
rect 12268 32230 12296 32506
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12070 27639 12126 27648
rect 12164 27668 12216 27674
rect 12164 27610 12216 27616
rect 12070 27568 12126 27577
rect 12070 27503 12126 27512
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 26586 11560 26726
rect 11622 26684 11918 26704
rect 11678 26682 11702 26684
rect 11758 26682 11782 26684
rect 11838 26682 11862 26684
rect 11700 26630 11702 26682
rect 11764 26630 11776 26682
rect 11838 26630 11840 26682
rect 11678 26628 11702 26630
rect 11758 26628 11782 26630
rect 11838 26628 11862 26630
rect 11622 26608 11918 26628
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11532 24886 11560 26522
rect 11888 26376 11940 26382
rect 11888 26318 11940 26324
rect 11900 25838 11928 26318
rect 11888 25832 11940 25838
rect 11888 25774 11940 25780
rect 12084 25650 12112 27503
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 12176 26994 12204 27270
rect 12164 26988 12216 26994
rect 12164 26930 12216 26936
rect 12176 26790 12204 26930
rect 12164 26784 12216 26790
rect 12164 26726 12216 26732
rect 12176 26450 12204 26726
rect 12164 26444 12216 26450
rect 12164 26386 12216 26392
rect 12176 25974 12204 26386
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 12084 25622 12204 25650
rect 11622 25596 11918 25616
rect 11678 25594 11702 25596
rect 11758 25594 11782 25596
rect 11838 25594 11862 25596
rect 11700 25542 11702 25594
rect 11764 25542 11776 25594
rect 11838 25542 11840 25594
rect 11678 25540 11702 25542
rect 11758 25540 11782 25542
rect 11838 25540 11862 25542
rect 11622 25520 11918 25540
rect 12070 24984 12126 24993
rect 12070 24919 12126 24928
rect 11520 24880 11572 24886
rect 11520 24822 11572 24828
rect 11622 24508 11918 24528
rect 11678 24506 11702 24508
rect 11758 24506 11782 24508
rect 11838 24506 11862 24508
rect 11700 24454 11702 24506
rect 11764 24454 11776 24506
rect 11838 24454 11840 24506
rect 11678 24452 11702 24454
rect 11758 24452 11782 24454
rect 11838 24452 11862 24454
rect 11622 24432 11918 24452
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11532 23526 11560 24210
rect 11520 23520 11572 23526
rect 11520 23462 11572 23468
rect 11622 23420 11918 23440
rect 11678 23418 11702 23420
rect 11758 23418 11782 23420
rect 11838 23418 11862 23420
rect 11700 23366 11702 23418
rect 11764 23366 11776 23418
rect 11838 23366 11840 23418
rect 11678 23364 11702 23366
rect 11758 23364 11782 23366
rect 11838 23364 11862 23366
rect 11622 23344 11918 23364
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11808 22710 11836 23054
rect 11796 22704 11848 22710
rect 11794 22672 11796 22681
rect 11848 22672 11850 22681
rect 11794 22607 11850 22616
rect 11622 22332 11918 22352
rect 11678 22330 11702 22332
rect 11758 22330 11782 22332
rect 11838 22330 11862 22332
rect 11700 22278 11702 22330
rect 11764 22278 11776 22330
rect 11838 22278 11840 22330
rect 11678 22276 11702 22278
rect 11758 22276 11782 22278
rect 11838 22276 11862 22278
rect 11622 22256 11918 22276
rect 11247 22120 11284 22148
rect 11431 22120 11468 22148
rect 11247 22012 11275 22120
rect 11336 22024 11388 22030
rect 11247 21984 11284 22012
rect 11256 21486 11284 21984
rect 11431 22012 11459 22120
rect 11431 21984 11468 22012
rect 11336 21966 11388 21972
rect 11348 21690 11376 21966
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11440 21078 11468 21984
rect 11520 21344 11572 21350
rect 11520 21286 11572 21292
rect 11532 21146 11560 21286
rect 11622 21244 11918 21264
rect 11678 21242 11702 21244
rect 11758 21242 11782 21244
rect 11838 21242 11862 21244
rect 11700 21190 11702 21242
rect 11764 21190 11776 21242
rect 11838 21190 11840 21242
rect 11678 21188 11702 21190
rect 11758 21188 11782 21190
rect 11838 21188 11862 21190
rect 11622 21168 11918 21188
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11428 21072 11480 21078
rect 11150 21040 11206 21049
rect 11428 21014 11480 21020
rect 11150 20975 11206 20984
rect 11440 20058 11468 21014
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11532 20913 11560 20946
rect 11612 20936 11664 20942
rect 11518 20904 11574 20913
rect 11612 20878 11664 20884
rect 11518 20839 11574 20848
rect 11532 20262 11560 20839
rect 11624 20466 11652 20878
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 10968 19848 11020 19854
rect 11164 19825 11192 19994
rect 11428 19848 11480 19854
rect 10968 19790 11020 19796
rect 11150 19816 11206 19825
rect 11428 19790 11480 19796
rect 11150 19751 11206 19760
rect 11440 19378 11468 19790
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11428 19372 11480 19378
rect 11428 19314 11480 19320
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 15156 11020 15162
rect 11072 15144 11100 15574
rect 11020 15116 11100 15144
rect 10968 15098 11020 15104
rect 10796 13790 10916 13818
rect 10796 13705 10824 13790
rect 10876 13728 10928 13734
rect 10782 13696 10838 13705
rect 10876 13670 10928 13676
rect 10782 13631 10838 13640
rect 10704 13382 10824 13410
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10704 12986 10732 13262
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10704 12764 10732 12922
rect 10612 12736 10732 12764
rect 10612 12306 10640 12736
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10612 11898 10640 12242
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10796 10282 10824 13382
rect 10888 13258 10916 13670
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 11164 12918 11192 19314
rect 11440 19145 11468 19314
rect 11426 19136 11482 19145
rect 11426 19071 11482 19080
rect 11440 17746 11468 19071
rect 11428 17740 11480 17746
rect 11428 17682 11480 17688
rect 11440 17338 11468 17682
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11440 16726 11468 17274
rect 11428 16720 11480 16726
rect 11428 16662 11480 16668
rect 11440 16250 11468 16662
rect 11428 16244 11480 16250
rect 11428 16186 11480 16192
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11348 13734 11376 14758
rect 11440 14482 11468 16186
rect 11532 15065 11560 20198
rect 11622 20156 11918 20176
rect 11678 20154 11702 20156
rect 11758 20154 11782 20156
rect 11838 20154 11862 20156
rect 11700 20102 11702 20154
rect 11764 20102 11776 20154
rect 11838 20102 11840 20154
rect 11678 20100 11702 20102
rect 11758 20100 11782 20102
rect 11838 20100 11862 20102
rect 11622 20080 11918 20100
rect 12084 20097 12112 24919
rect 12176 23100 12204 25622
rect 12268 23254 12296 32166
rect 12360 30954 12388 32846
rect 12440 32768 12492 32774
rect 12440 32710 12492 32716
rect 12452 32570 12480 32710
rect 12440 32564 12492 32570
rect 12440 32506 12492 32512
rect 12544 32366 12572 39520
rect 12900 34944 12952 34950
rect 12900 34886 12952 34892
rect 12912 34610 12940 34886
rect 12900 34604 12952 34610
rect 12900 34546 12952 34552
rect 12900 33856 12952 33862
rect 12900 33798 12952 33804
rect 12912 33522 12940 33798
rect 12900 33516 12952 33522
rect 12900 33458 12952 33464
rect 12714 33416 12770 33425
rect 12912 33402 12940 33458
rect 12714 33351 12770 33360
rect 12820 33374 12940 33402
rect 12728 33114 12756 33351
rect 12716 33108 12768 33114
rect 12716 33050 12768 33056
rect 12624 32972 12676 32978
rect 12624 32914 12676 32920
rect 12636 32881 12664 32914
rect 12622 32872 12678 32881
rect 12622 32807 12678 32816
rect 12636 32570 12664 32807
rect 12624 32564 12676 32570
rect 12624 32506 12676 32512
rect 12728 32502 12756 33050
rect 12820 32910 12848 33374
rect 12900 33312 12952 33318
rect 12900 33254 12952 33260
rect 12808 32904 12860 32910
rect 12808 32846 12860 32852
rect 12716 32496 12768 32502
rect 12716 32438 12768 32444
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 12544 32026 12572 32302
rect 12532 32020 12584 32026
rect 12532 31962 12584 31968
rect 12820 31822 12848 32846
rect 12912 32774 12940 33254
rect 12900 32768 12952 32774
rect 12900 32710 12952 32716
rect 12808 31816 12860 31822
rect 12808 31758 12860 31764
rect 12360 30938 12480 30954
rect 12360 30932 12492 30938
rect 12360 30926 12440 30932
rect 12360 28694 12388 30926
rect 12440 30874 12492 30880
rect 12532 28960 12584 28966
rect 12532 28902 12584 28908
rect 12348 28688 12400 28694
rect 12348 28630 12400 28636
rect 12360 28218 12388 28630
rect 12544 28490 12572 28902
rect 12532 28484 12584 28490
rect 12532 28426 12584 28432
rect 12348 28212 12400 28218
rect 12348 28154 12400 28160
rect 12808 27328 12860 27334
rect 12808 27270 12860 27276
rect 12820 26897 12848 27270
rect 13004 27033 13032 39520
rect 13372 35714 13400 39520
rect 13096 35686 13400 35714
rect 12990 27024 13046 27033
rect 12990 26959 13046 26968
rect 12806 26888 12862 26897
rect 12806 26823 12808 26832
rect 12860 26823 12862 26832
rect 12808 26794 12860 26800
rect 12440 26784 12492 26790
rect 12820 26763 12848 26794
rect 12900 26784 12952 26790
rect 12440 26726 12492 26732
rect 12900 26726 12952 26732
rect 12452 24970 12480 26726
rect 12912 26586 12940 26726
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12360 24942 12480 24970
rect 12360 24818 12388 24942
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12256 23248 12308 23254
rect 12256 23190 12308 23196
rect 12360 23186 12388 23462
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12176 23072 12296 23100
rect 12164 22976 12216 22982
rect 12164 22918 12216 22924
rect 12176 22166 12204 22918
rect 12164 22160 12216 22166
rect 12164 22102 12216 22108
rect 12176 21146 12204 22102
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12070 20088 12126 20097
rect 12070 20023 12126 20032
rect 12070 19952 12126 19961
rect 11796 19916 11848 19922
rect 12070 19887 12126 19896
rect 11796 19858 11848 19864
rect 11808 19514 11836 19858
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 12084 19378 12112 19887
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11622 19068 11918 19088
rect 11678 19066 11702 19068
rect 11758 19066 11782 19068
rect 11838 19066 11862 19068
rect 11700 19014 11702 19066
rect 11764 19014 11776 19066
rect 11838 19014 11840 19066
rect 11678 19012 11702 19014
rect 11758 19012 11782 19014
rect 11838 19012 11862 19014
rect 11622 18992 11918 19012
rect 11622 17980 11918 18000
rect 11678 17978 11702 17980
rect 11758 17978 11782 17980
rect 11838 17978 11862 17980
rect 11700 17926 11702 17978
rect 11764 17926 11776 17978
rect 11838 17926 11840 17978
rect 11678 17924 11702 17926
rect 11758 17924 11782 17926
rect 11838 17924 11862 17926
rect 11622 17904 11918 17924
rect 11622 16892 11918 16912
rect 11678 16890 11702 16892
rect 11758 16890 11782 16892
rect 11838 16890 11862 16892
rect 11700 16838 11702 16890
rect 11764 16838 11776 16890
rect 11838 16838 11840 16890
rect 11678 16836 11702 16838
rect 11758 16836 11782 16838
rect 11838 16836 11862 16838
rect 11622 16816 11918 16836
rect 11622 15804 11918 15824
rect 11678 15802 11702 15804
rect 11758 15802 11782 15804
rect 11838 15802 11862 15804
rect 11700 15750 11702 15802
rect 11764 15750 11776 15802
rect 11838 15750 11840 15802
rect 11678 15748 11702 15750
rect 11758 15748 11782 15750
rect 11838 15748 11862 15750
rect 11622 15728 11918 15748
rect 11992 15722 12020 19314
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 16998 12204 17682
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 11992 15694 12112 15722
rect 11980 15632 12032 15638
rect 11980 15574 12032 15580
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11518 15056 11574 15065
rect 11518 14991 11574 15000
rect 11428 14476 11480 14482
rect 11428 14418 11480 14424
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11440 13002 11468 14418
rect 11348 12974 11468 13002
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11348 12374 11376 12974
rect 11428 12912 11480 12918
rect 11428 12854 11480 12860
rect 11336 12368 11388 12374
rect 11336 12310 11388 12316
rect 11242 10432 11298 10441
rect 11242 10367 11298 10376
rect 10612 10254 10824 10282
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10416 4616 10468 4622
rect 10152 4542 10272 4570
rect 10416 4558 10468 4564
rect 10244 4486 10272 4542
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10060 4134 10180 4162
rect 10152 4078 10180 4134
rect 10140 4072 10192 4078
rect 10046 4040 10102 4049
rect 10140 4014 10192 4020
rect 10046 3975 10102 3984
rect 10060 3942 10088 3975
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9954 3768 10010 3777
rect 9954 3703 10010 3712
rect 9862 3632 9918 3641
rect 9862 3567 9918 3576
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9876 3097 9904 3334
rect 9862 3088 9918 3097
rect 9862 3023 9918 3032
rect 10152 480 10180 4014
rect 10244 3942 10272 4422
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3534 10272 3878
rect 10336 3738 10364 3946
rect 10428 3913 10456 4558
rect 10414 3904 10470 3913
rect 10414 3839 10470 3848
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10520 3618 10548 6122
rect 10612 6118 10640 10254
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10704 9586 10732 10134
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10704 8906 10732 9522
rect 10888 9518 10916 9862
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10876 9512 10928 9518
rect 10782 9480 10838 9489
rect 10876 9454 10928 9460
rect 10782 9415 10838 9424
rect 10796 9382 10824 9415
rect 10784 9376 10836 9382
rect 10980 9330 11008 9522
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10784 9318 10836 9324
rect 10888 9302 11008 9330
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10692 8900 10744 8906
rect 10692 8842 10744 8848
rect 10704 8634 10732 8842
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10704 7478 10732 8570
rect 10796 8514 10824 9114
rect 10888 8838 10916 9302
rect 11072 8906 11100 9386
rect 11150 8936 11206 8945
rect 11060 8900 11112 8906
rect 11150 8871 11206 8880
rect 11060 8842 11112 8848
rect 10876 8832 10928 8838
rect 10874 8800 10876 8809
rect 10928 8800 10930 8809
rect 10874 8735 10930 8744
rect 10796 8486 10916 8514
rect 10782 8392 10838 8401
rect 10782 8327 10838 8336
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10704 6934 10732 7414
rect 10796 7410 10824 8327
rect 10784 7404 10836 7410
rect 10784 7346 10836 7352
rect 10796 7002 10824 7346
rect 10784 6996 10836 7002
rect 10784 6938 10836 6944
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10612 5370 10640 5714
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10704 4826 10732 5646
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10796 4758 10824 5646
rect 10888 5302 10916 8486
rect 11072 8090 11100 8842
rect 11164 8090 11192 8871
rect 11256 8430 11284 10367
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7546 11100 7890
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7002 11192 8026
rect 11348 7886 11376 8570
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11348 7478 11376 7822
rect 11336 7472 11388 7478
rect 11336 7414 11388 7420
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10888 5098 10916 5238
rect 10876 5092 10928 5098
rect 10876 5034 10928 5040
rect 11164 5001 11192 5306
rect 11348 5234 11376 5714
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11150 4992 11206 5001
rect 11150 4927 11206 4936
rect 10784 4752 10836 4758
rect 10690 4720 10746 4729
rect 10784 4694 10836 4700
rect 10690 4655 10746 4664
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10612 3738 10640 4082
rect 10600 3732 10652 3738
rect 10600 3674 10652 3680
rect 10520 3590 10640 3618
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10612 480 10640 3590
rect 10704 3074 10732 4655
rect 10796 3738 10824 4694
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10888 4282 10916 4558
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11164 3602 11192 4927
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11256 4078 11284 4626
rect 11348 4622 11376 5170
rect 11440 5166 11468 12854
rect 11428 5160 11480 5166
rect 11428 5102 11480 5108
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11348 4146 11376 4558
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11256 3738 11284 3878
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11256 3602 11284 3674
rect 10784 3596 10836 3602
rect 10784 3538 10836 3544
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10796 3233 10824 3538
rect 10782 3224 10838 3233
rect 10782 3159 10784 3168
rect 10836 3159 10838 3168
rect 10784 3130 10836 3136
rect 10704 3046 10916 3074
rect 10888 2666 10916 3046
rect 10888 2638 11008 2666
rect 11164 2650 11192 3538
rect 11426 3496 11482 3505
rect 11426 3431 11482 3440
rect 11440 3194 11468 3431
rect 11428 3188 11480 3194
rect 11428 3130 11480 3136
rect 11334 2816 11390 2825
rect 11334 2751 11390 2760
rect 10980 480 11008 2638
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11348 480 11376 2751
rect 11532 1442 11560 14991
rect 11716 14890 11744 15438
rect 11704 14884 11756 14890
rect 11704 14826 11756 14832
rect 11622 14716 11918 14736
rect 11678 14714 11702 14716
rect 11758 14714 11782 14716
rect 11838 14714 11862 14716
rect 11700 14662 11702 14714
rect 11764 14662 11776 14714
rect 11838 14662 11840 14714
rect 11678 14660 11702 14662
rect 11758 14660 11782 14662
rect 11838 14660 11862 14662
rect 11622 14640 11918 14660
rect 11992 14618 12020 15574
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11888 14476 11940 14482
rect 11888 14418 11940 14424
rect 11808 14074 11836 14418
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11900 13938 11928 14418
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11992 13841 12020 14010
rect 11978 13832 12034 13841
rect 11978 13767 12034 13776
rect 11622 13628 11918 13648
rect 11678 13626 11702 13628
rect 11758 13626 11782 13628
rect 11838 13626 11862 13628
rect 11700 13574 11702 13626
rect 11764 13574 11776 13626
rect 11838 13574 11840 13626
rect 11678 13572 11702 13574
rect 11758 13572 11782 13574
rect 11838 13572 11862 13574
rect 11622 13552 11918 13572
rect 12084 13530 12112 15694
rect 12176 15502 12204 16934
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12176 14822 12204 14962
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 12176 14550 12204 14758
rect 12164 14544 12216 14550
rect 12164 14486 12216 14492
rect 12164 13932 12216 13938
rect 12164 13874 12216 13880
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11992 12918 12020 13330
rect 12084 12986 12112 13466
rect 12176 13326 12204 13874
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12986 12204 13262
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11622 12540 11918 12560
rect 11678 12538 11702 12540
rect 11758 12538 11782 12540
rect 11838 12538 11862 12540
rect 11700 12486 11702 12538
rect 11764 12486 11776 12538
rect 11838 12486 11840 12538
rect 11678 12484 11702 12486
rect 11758 12484 11782 12486
rect 11838 12484 11862 12486
rect 11622 12464 11918 12484
rect 12176 12442 12204 12922
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11622 11452 11918 11472
rect 11678 11450 11702 11452
rect 11758 11450 11782 11452
rect 11838 11450 11862 11452
rect 11700 11398 11702 11450
rect 11764 11398 11776 11450
rect 11838 11398 11840 11450
rect 11678 11396 11702 11398
rect 11758 11396 11782 11398
rect 11838 11396 11862 11398
rect 11622 11376 11918 11396
rect 12070 11112 12126 11121
rect 12070 11047 12126 11056
rect 11622 10364 11918 10384
rect 11678 10362 11702 10364
rect 11758 10362 11782 10364
rect 11838 10362 11862 10364
rect 11700 10310 11702 10362
rect 11764 10310 11776 10362
rect 11838 10310 11840 10362
rect 11678 10308 11702 10310
rect 11758 10308 11782 10310
rect 11838 10308 11862 10310
rect 11622 10288 11918 10308
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11622 9276 11918 9296
rect 11678 9274 11702 9276
rect 11758 9274 11782 9276
rect 11838 9274 11862 9276
rect 11700 9222 11702 9274
rect 11764 9222 11776 9274
rect 11838 9222 11840 9274
rect 11678 9220 11702 9222
rect 11758 9220 11782 9222
rect 11838 9220 11862 9222
rect 11622 9200 11918 9220
rect 11992 9110 12020 9862
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11716 8566 11744 8978
rect 11992 8634 12020 9046
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11622 8188 11918 8208
rect 11678 8186 11702 8188
rect 11758 8186 11782 8188
rect 11838 8186 11862 8188
rect 11700 8134 11702 8186
rect 11764 8134 11776 8186
rect 11838 8134 11840 8186
rect 11678 8132 11702 8134
rect 11758 8132 11782 8134
rect 11838 8132 11862 8134
rect 11622 8112 11918 8132
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11622 7100 11918 7120
rect 11678 7098 11702 7100
rect 11758 7098 11782 7100
rect 11838 7098 11862 7100
rect 11700 7046 11702 7098
rect 11764 7046 11776 7098
rect 11838 7046 11840 7098
rect 11678 7044 11702 7046
rect 11758 7044 11782 7046
rect 11838 7044 11862 7046
rect 11622 7024 11918 7044
rect 11622 6012 11918 6032
rect 11678 6010 11702 6012
rect 11758 6010 11782 6012
rect 11838 6010 11862 6012
rect 11700 5958 11702 6010
rect 11764 5958 11776 6010
rect 11838 5958 11840 6010
rect 11678 5956 11702 5958
rect 11758 5956 11782 5958
rect 11838 5956 11862 5958
rect 11622 5936 11918 5956
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11808 5370 11836 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11622 4924 11918 4944
rect 11678 4922 11702 4924
rect 11758 4922 11782 4924
rect 11838 4922 11862 4924
rect 11700 4870 11702 4922
rect 11764 4870 11776 4922
rect 11838 4870 11840 4922
rect 11678 4868 11702 4870
rect 11758 4868 11782 4870
rect 11838 4868 11862 4870
rect 11622 4848 11918 4868
rect 11622 3836 11918 3856
rect 11678 3834 11702 3836
rect 11758 3834 11782 3836
rect 11838 3834 11862 3836
rect 11700 3782 11702 3834
rect 11764 3782 11776 3834
rect 11838 3782 11840 3834
rect 11678 3780 11702 3782
rect 11758 3780 11782 3782
rect 11838 3780 11862 3782
rect 11622 3760 11918 3780
rect 11992 3074 12020 7142
rect 12084 3194 12112 11047
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12176 6769 12204 6802
rect 12162 6760 12218 6769
rect 12162 6695 12218 6704
rect 12176 6458 12204 6695
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12176 5574 12204 6394
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12176 4185 12204 4422
rect 12162 4176 12218 4185
rect 12162 4111 12218 4120
rect 12268 3754 12296 23072
rect 12452 22522 12480 24006
rect 13096 23322 13124 35686
rect 13174 34640 13230 34649
rect 13174 34575 13230 34584
rect 13634 34640 13690 34649
rect 13634 34575 13690 34584
rect 13188 34542 13216 34575
rect 13176 34536 13228 34542
rect 13176 34478 13228 34484
rect 13542 33416 13598 33425
rect 13542 33351 13598 33360
rect 13176 32360 13228 32366
rect 13176 32302 13228 32308
rect 12624 23316 12676 23322
rect 12624 23258 12676 23264
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12636 23118 12664 23258
rect 12716 23248 12768 23254
rect 12716 23190 12768 23196
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12360 22494 12480 22522
rect 12360 22030 12388 22494
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 22098 12480 22374
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12348 22024 12400 22030
rect 12348 21966 12400 21972
rect 12544 21894 12572 22578
rect 12728 22574 12756 23190
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12532 21888 12584 21894
rect 12438 21856 12494 21865
rect 12532 21830 12584 21836
rect 12438 21791 12494 21800
rect 12452 21690 12480 21791
rect 12440 21684 12492 21690
rect 12440 21626 12492 21632
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12360 14074 12388 15506
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14618 12480 14758
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12544 14006 12572 21830
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12636 20806 12664 21490
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12636 20641 12664 20742
rect 12622 20632 12678 20641
rect 12622 20567 12678 20576
rect 12636 20058 12664 20567
rect 12624 20052 12676 20058
rect 12624 19994 12676 20000
rect 12728 14890 12756 22510
rect 12808 22500 12860 22506
rect 12808 22442 12860 22448
rect 12820 22234 12848 22442
rect 12808 22228 12860 22234
rect 12808 22170 12860 22176
rect 13004 21554 13032 22578
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13084 21480 13136 21486
rect 13084 21422 13136 21428
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 16697 13032 17478
rect 12990 16688 13046 16697
rect 12990 16623 13046 16632
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12716 14884 12768 14890
rect 12716 14826 12768 14832
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12544 13870 12572 13942
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12636 13530 12664 13670
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12356 12572 12854
rect 12544 12328 12664 12356
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9586 12572 9862
rect 12636 9602 12664 12328
rect 12912 10146 12940 14894
rect 12912 10118 13032 10146
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12532 9580 12584 9586
rect 12636 9574 12756 9602
rect 12532 9522 12584 9528
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12452 8634 12480 9318
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12636 6458 12664 6802
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12348 5840 12400 5846
rect 12348 5782 12400 5788
rect 12360 5370 12388 5782
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12728 4826 12756 9574
rect 12820 9518 12848 9862
rect 12912 9722 12940 9998
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12912 8838 12940 9658
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 8498 12940 8774
rect 12900 8492 12952 8498
rect 12820 8452 12900 8480
rect 12820 8022 12848 8452
rect 12900 8434 12952 8440
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12912 8090 12940 8230
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 8016 12860 8022
rect 12912 7993 12940 8026
rect 12808 7958 12860 7964
rect 12898 7984 12954 7993
rect 12898 7919 12954 7928
rect 13004 5114 13032 10118
rect 13096 8922 13124 21422
rect 13188 15706 13216 32302
rect 13556 31482 13584 33351
rect 13544 31476 13596 31482
rect 13544 31418 13596 31424
rect 13452 31272 13504 31278
rect 13452 31214 13504 31220
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13280 24993 13308 26250
rect 13266 24984 13322 24993
rect 13266 24919 13322 24928
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22642 13308 22918
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13464 19378 13492 31214
rect 13648 22574 13676 34575
rect 13740 31385 13768 39520
rect 14108 39494 14228 39520
rect 13726 31376 13782 31385
rect 13726 31311 13782 31320
rect 14108 24857 14136 39494
rect 14568 37210 14596 39520
rect 14936 39494 15056 39520
rect 14568 37182 14688 37210
rect 14289 37020 14585 37040
rect 14345 37018 14369 37020
rect 14425 37018 14449 37020
rect 14505 37018 14529 37020
rect 14367 36966 14369 37018
rect 14431 36966 14443 37018
rect 14505 36966 14507 37018
rect 14345 36964 14369 36966
rect 14425 36964 14449 36966
rect 14505 36964 14529 36966
rect 14289 36944 14585 36964
rect 14289 35932 14585 35952
rect 14345 35930 14369 35932
rect 14425 35930 14449 35932
rect 14505 35930 14529 35932
rect 14367 35878 14369 35930
rect 14431 35878 14443 35930
rect 14505 35878 14507 35930
rect 14345 35876 14369 35878
rect 14425 35876 14449 35878
rect 14505 35876 14529 35878
rect 14289 35856 14585 35876
rect 14289 34844 14585 34864
rect 14345 34842 14369 34844
rect 14425 34842 14449 34844
rect 14505 34842 14529 34844
rect 14367 34790 14369 34842
rect 14431 34790 14443 34842
rect 14505 34790 14507 34842
rect 14345 34788 14369 34790
rect 14425 34788 14449 34790
rect 14505 34788 14529 34790
rect 14289 34768 14585 34788
rect 14289 33756 14585 33776
rect 14345 33754 14369 33756
rect 14425 33754 14449 33756
rect 14505 33754 14529 33756
rect 14367 33702 14369 33754
rect 14431 33702 14443 33754
rect 14505 33702 14507 33754
rect 14345 33700 14369 33702
rect 14425 33700 14449 33702
rect 14505 33700 14529 33702
rect 14289 33680 14585 33700
rect 14289 32668 14585 32688
rect 14345 32666 14369 32668
rect 14425 32666 14449 32668
rect 14505 32666 14529 32668
rect 14367 32614 14369 32666
rect 14431 32614 14443 32666
rect 14505 32614 14507 32666
rect 14345 32612 14369 32614
rect 14425 32612 14449 32614
rect 14505 32612 14529 32614
rect 14289 32592 14585 32612
rect 14289 31580 14585 31600
rect 14345 31578 14369 31580
rect 14425 31578 14449 31580
rect 14505 31578 14529 31580
rect 14367 31526 14369 31578
rect 14431 31526 14443 31578
rect 14505 31526 14507 31578
rect 14345 31524 14369 31526
rect 14425 31524 14449 31526
rect 14505 31524 14529 31526
rect 14289 31504 14585 31524
rect 14289 30492 14585 30512
rect 14345 30490 14369 30492
rect 14425 30490 14449 30492
rect 14505 30490 14529 30492
rect 14367 30438 14369 30490
rect 14431 30438 14443 30490
rect 14505 30438 14507 30490
rect 14345 30436 14369 30438
rect 14425 30436 14449 30438
rect 14505 30436 14529 30438
rect 14289 30416 14585 30436
rect 14660 29753 14688 37182
rect 14646 29744 14702 29753
rect 14646 29679 14702 29688
rect 14289 29404 14585 29424
rect 14345 29402 14369 29404
rect 14425 29402 14449 29404
rect 14505 29402 14529 29404
rect 14367 29350 14369 29402
rect 14431 29350 14443 29402
rect 14505 29350 14507 29402
rect 14345 29348 14369 29350
rect 14425 29348 14449 29350
rect 14505 29348 14529 29350
rect 14289 29328 14585 29348
rect 14289 28316 14585 28336
rect 14345 28314 14369 28316
rect 14425 28314 14449 28316
rect 14505 28314 14529 28316
rect 14367 28262 14369 28314
rect 14431 28262 14443 28314
rect 14505 28262 14507 28314
rect 14345 28260 14369 28262
rect 14425 28260 14449 28262
rect 14505 28260 14529 28262
rect 14289 28240 14585 28260
rect 15028 27577 15056 39494
rect 15396 32337 15424 39520
rect 15764 34649 15792 39520
rect 15750 34640 15806 34649
rect 15750 34575 15806 34584
rect 15382 32328 15438 32337
rect 15382 32263 15438 32272
rect 15014 27568 15070 27577
rect 15014 27503 15070 27512
rect 14289 27228 14585 27248
rect 14345 27226 14369 27228
rect 14425 27226 14449 27228
rect 14505 27226 14529 27228
rect 14367 27174 14369 27226
rect 14431 27174 14443 27226
rect 14505 27174 14507 27226
rect 14345 27172 14369 27174
rect 14425 27172 14449 27174
rect 14505 27172 14529 27174
rect 14289 27152 14585 27172
rect 14289 26140 14585 26160
rect 14345 26138 14369 26140
rect 14425 26138 14449 26140
rect 14505 26138 14529 26140
rect 14367 26086 14369 26138
rect 14431 26086 14443 26138
rect 14505 26086 14507 26138
rect 14345 26084 14369 26086
rect 14425 26084 14449 26086
rect 14505 26084 14529 26086
rect 14289 26064 14585 26084
rect 14289 25052 14585 25072
rect 14345 25050 14369 25052
rect 14425 25050 14449 25052
rect 14505 25050 14529 25052
rect 14367 24998 14369 25050
rect 14431 24998 14443 25050
rect 14505 24998 14507 25050
rect 14345 24996 14369 24998
rect 14425 24996 14449 24998
rect 14505 24996 14529 24998
rect 14289 24976 14585 24996
rect 14094 24848 14150 24857
rect 14094 24783 14150 24792
rect 14289 23964 14585 23984
rect 14345 23962 14369 23964
rect 14425 23962 14449 23964
rect 14505 23962 14529 23964
rect 14367 23910 14369 23962
rect 14431 23910 14443 23962
rect 14505 23910 14507 23962
rect 14345 23908 14369 23910
rect 14425 23908 14449 23910
rect 14505 23908 14529 23910
rect 14289 23888 14585 23908
rect 14289 22876 14585 22896
rect 14345 22874 14369 22876
rect 14425 22874 14449 22876
rect 14505 22874 14529 22876
rect 14367 22822 14369 22874
rect 14431 22822 14443 22874
rect 14505 22822 14507 22874
rect 14345 22820 14369 22822
rect 14425 22820 14449 22822
rect 14505 22820 14529 22822
rect 14289 22800 14585 22820
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 14289 21788 14585 21808
rect 14345 21786 14369 21788
rect 14425 21786 14449 21788
rect 14505 21786 14529 21788
rect 14367 21734 14369 21786
rect 14431 21734 14443 21786
rect 14505 21734 14507 21786
rect 14345 21732 14369 21734
rect 14425 21732 14449 21734
rect 14505 21732 14529 21734
rect 14289 21712 14585 21732
rect 14289 20700 14585 20720
rect 14345 20698 14369 20700
rect 14425 20698 14449 20700
rect 14505 20698 14529 20700
rect 14367 20646 14369 20698
rect 14431 20646 14443 20698
rect 14505 20646 14507 20698
rect 14345 20644 14369 20646
rect 14425 20644 14449 20646
rect 14505 20644 14529 20646
rect 14289 20624 14585 20644
rect 14289 19612 14585 19632
rect 14345 19610 14369 19612
rect 14425 19610 14449 19612
rect 14505 19610 14529 19612
rect 14367 19558 14369 19610
rect 14431 19558 14443 19610
rect 14505 19558 14507 19610
rect 14345 19556 14369 19558
rect 14425 19556 14449 19558
rect 14505 19556 14529 19558
rect 14289 19536 14585 19556
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13188 14958 13216 15642
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13372 10554 13400 19314
rect 14289 18524 14585 18544
rect 14345 18522 14369 18524
rect 14425 18522 14449 18524
rect 14505 18522 14529 18524
rect 14367 18470 14369 18522
rect 14431 18470 14443 18522
rect 14505 18470 14507 18522
rect 14345 18468 14369 18470
rect 14425 18468 14449 18470
rect 14505 18468 14529 18470
rect 14289 18448 14585 18468
rect 14289 17436 14585 17456
rect 14345 17434 14369 17436
rect 14425 17434 14449 17436
rect 14505 17434 14529 17436
rect 14367 17382 14369 17434
rect 14431 17382 14443 17434
rect 14505 17382 14507 17434
rect 14345 17380 14369 17382
rect 14425 17380 14449 17382
rect 14505 17380 14529 17382
rect 14289 17360 14585 17380
rect 14289 16348 14585 16368
rect 14345 16346 14369 16348
rect 14425 16346 14449 16348
rect 14505 16346 14529 16348
rect 14367 16294 14369 16346
rect 14431 16294 14443 16346
rect 14505 16294 14507 16346
rect 14345 16292 14369 16294
rect 14425 16292 14449 16294
rect 14505 16292 14529 16294
rect 14289 16272 14585 16292
rect 14289 15260 14585 15280
rect 14345 15258 14369 15260
rect 14425 15258 14449 15260
rect 14505 15258 14529 15260
rect 14367 15206 14369 15258
rect 14431 15206 14443 15258
rect 14505 15206 14507 15258
rect 14345 15204 14369 15206
rect 14425 15204 14449 15206
rect 14505 15204 14529 15206
rect 14289 15184 14585 15204
rect 14004 14884 14056 14890
rect 14004 14826 14056 14832
rect 13726 12200 13782 12209
rect 13726 12135 13782 12144
rect 13280 10526 13400 10554
rect 13280 9489 13308 10526
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13372 10266 13400 10406
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 13372 9722 13400 10202
rect 13450 10160 13506 10169
rect 13450 10095 13452 10104
rect 13504 10095 13506 10104
rect 13452 10066 13504 10072
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13464 9654 13492 10066
rect 13452 9648 13504 9654
rect 13452 9590 13504 9596
rect 13266 9480 13322 9489
rect 13266 9415 13322 9424
rect 13096 8894 13400 8922
rect 13084 8832 13136 8838
rect 13082 8800 13084 8809
rect 13136 8800 13138 8809
rect 13082 8735 13138 8744
rect 13096 6866 13124 8735
rect 13174 8392 13230 8401
rect 13174 8327 13176 8336
rect 13228 8327 13230 8336
rect 13176 8298 13228 8304
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12912 5086 13032 5114
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12544 4282 12572 4762
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12636 4282 12664 4558
rect 12532 4276 12584 4282
rect 12452 4236 12532 4264
rect 12452 3924 12480 4236
rect 12532 4218 12584 4224
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12636 4162 12664 4218
rect 12544 4134 12664 4162
rect 12716 4140 12768 4146
rect 12544 4049 12572 4134
rect 12716 4082 12768 4088
rect 12624 4072 12676 4078
rect 12530 4040 12586 4049
rect 12624 4014 12676 4020
rect 12530 3975 12586 3984
rect 12452 3896 12572 3924
rect 12268 3726 12480 3754
rect 12452 3233 12480 3726
rect 12438 3224 12494 3233
rect 12072 3188 12124 3194
rect 12438 3159 12494 3168
rect 12072 3130 12124 3136
rect 11992 3046 12112 3074
rect 11622 2748 11918 2768
rect 11678 2746 11702 2748
rect 11758 2746 11782 2748
rect 11838 2746 11862 2748
rect 11700 2694 11702 2746
rect 11764 2694 11776 2746
rect 11838 2694 11840 2746
rect 11678 2692 11702 2694
rect 11758 2692 11782 2694
rect 11838 2692 11862 2694
rect 11622 2672 11918 2692
rect 12084 2666 12112 3046
rect 12084 2638 12204 2666
rect 12452 2650 12480 3159
rect 11532 1414 11836 1442
rect 11808 480 11836 1414
rect 12176 480 12204 2638
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12544 480 12572 3896
rect 12636 2650 12664 4014
rect 12728 3670 12756 4082
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12728 3466 12756 3606
rect 12716 3460 12768 3466
rect 12716 3402 12768 3408
rect 12912 2922 12940 5086
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12898 2544 12954 2553
rect 13004 2514 13032 4966
rect 13188 4758 13216 5510
rect 13176 4752 13228 4758
rect 13228 4712 13308 4740
rect 13176 4694 13228 4700
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4078 13216 4422
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13084 3936 13136 3942
rect 13084 3878 13136 3884
rect 13096 3398 13124 3878
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3194 13124 3334
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 13280 3058 13308 4712
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12898 2479 12954 2488
rect 12992 2508 13044 2514
rect 12912 2394 12940 2479
rect 12992 2450 13044 2456
rect 13280 2446 13308 2994
rect 13268 2440 13320 2446
rect 12912 2366 13032 2394
rect 13268 2382 13320 2388
rect 13004 480 13032 2366
rect 13372 480 13400 8894
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 5846 13492 6598
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13740 480 13768 12135
rect 14016 7546 14044 14826
rect 14289 14172 14585 14192
rect 14345 14170 14369 14172
rect 14425 14170 14449 14172
rect 14505 14170 14529 14172
rect 14367 14118 14369 14170
rect 14431 14118 14443 14170
rect 14505 14118 14507 14170
rect 14345 14116 14369 14118
rect 14425 14116 14449 14118
rect 14505 14116 14529 14118
rect 14289 14096 14585 14116
rect 14289 13084 14585 13104
rect 14345 13082 14369 13084
rect 14425 13082 14449 13084
rect 14505 13082 14529 13084
rect 14367 13030 14369 13082
rect 14431 13030 14443 13082
rect 14505 13030 14507 13082
rect 14345 13028 14369 13030
rect 14425 13028 14449 13030
rect 14505 13028 14529 13030
rect 14289 13008 14585 13028
rect 14289 11996 14585 12016
rect 14345 11994 14369 11996
rect 14425 11994 14449 11996
rect 14505 11994 14529 11996
rect 14367 11942 14369 11994
rect 14431 11942 14443 11994
rect 14505 11942 14507 11994
rect 14345 11940 14369 11942
rect 14425 11940 14449 11942
rect 14505 11940 14529 11942
rect 14289 11920 14585 11940
rect 14289 10908 14585 10928
rect 14345 10906 14369 10908
rect 14425 10906 14449 10908
rect 14505 10906 14529 10908
rect 14367 10854 14369 10906
rect 14431 10854 14443 10906
rect 14505 10854 14507 10906
rect 14345 10852 14369 10854
rect 14425 10852 14449 10854
rect 14505 10852 14529 10854
rect 14289 10832 14585 10852
rect 14289 9820 14585 9840
rect 14345 9818 14369 9820
rect 14425 9818 14449 9820
rect 14505 9818 14529 9820
rect 14367 9766 14369 9818
rect 14431 9766 14443 9818
rect 14505 9766 14507 9818
rect 14345 9764 14369 9766
rect 14425 9764 14449 9766
rect 14505 9764 14529 9766
rect 14289 9744 14585 9764
rect 14289 8732 14585 8752
rect 14345 8730 14369 8732
rect 14425 8730 14449 8732
rect 14505 8730 14529 8732
rect 14367 8678 14369 8730
rect 14431 8678 14443 8730
rect 14505 8678 14507 8730
rect 14345 8676 14369 8678
rect 14425 8676 14449 8678
rect 14505 8676 14529 8678
rect 14289 8656 14585 8676
rect 14646 8392 14702 8401
rect 14646 8327 14702 8336
rect 14289 7644 14585 7664
rect 14345 7642 14369 7644
rect 14425 7642 14449 7644
rect 14505 7642 14529 7644
rect 14367 7590 14369 7642
rect 14431 7590 14443 7642
rect 14505 7590 14507 7642
rect 14345 7588 14369 7590
rect 14425 7588 14449 7590
rect 14505 7588 14529 7590
rect 14289 7568 14585 7588
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14289 6556 14585 6576
rect 14345 6554 14369 6556
rect 14425 6554 14449 6556
rect 14505 6554 14529 6556
rect 14367 6502 14369 6554
rect 14431 6502 14443 6554
rect 14505 6502 14507 6554
rect 14345 6500 14369 6502
rect 14425 6500 14449 6502
rect 14505 6500 14529 6502
rect 14289 6480 14585 6500
rect 14289 5468 14585 5488
rect 14345 5466 14369 5468
rect 14425 5466 14449 5468
rect 14505 5466 14529 5468
rect 14367 5414 14369 5466
rect 14431 5414 14443 5466
rect 14505 5414 14507 5466
rect 14345 5412 14369 5414
rect 14425 5412 14449 5414
rect 14505 5412 14529 5414
rect 14289 5392 14585 5412
rect 14289 4380 14585 4400
rect 14345 4378 14369 4380
rect 14425 4378 14449 4380
rect 14505 4378 14529 4380
rect 14367 4326 14369 4378
rect 14431 4326 14443 4378
rect 14505 4326 14507 4378
rect 14345 4324 14369 4326
rect 14425 4324 14449 4326
rect 14505 4324 14529 4326
rect 14289 4304 14585 4324
rect 14289 3292 14585 3312
rect 14345 3290 14369 3292
rect 14425 3290 14449 3292
rect 14505 3290 14529 3292
rect 14367 3238 14369 3290
rect 14431 3238 14443 3290
rect 14505 3238 14507 3290
rect 14345 3236 14369 3238
rect 14425 3236 14449 3238
rect 14505 3236 14529 3238
rect 14289 3216 14585 3236
rect 14289 2204 14585 2224
rect 14345 2202 14369 2204
rect 14425 2202 14449 2204
rect 14505 2202 14529 2204
rect 14367 2150 14369 2202
rect 14431 2150 14443 2202
rect 14505 2150 14507 2202
rect 14345 2148 14369 2150
rect 14425 2148 14449 2150
rect 14505 2148 14529 2150
rect 14289 2128 14585 2148
rect 14186 2000 14242 2009
rect 14186 1935 14242 1944
rect 14200 480 14228 1935
rect 14660 1442 14688 8327
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15382 6896 15438 6905
rect 15382 6831 15438 6840
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14568 1414 14688 1442
rect 14568 480 14596 1414
rect 14936 480 14964 2790
rect 15396 480 15424 6831
rect 15764 480 15792 7482
rect 202 0 258 480
rect 570 0 626 480
rect 938 0 994 480
rect 1398 0 1454 480
rect 1766 0 1822 480
rect 2134 0 2190 480
rect 2594 0 2650 480
rect 2962 0 3018 480
rect 3330 0 3386 480
rect 3790 0 3846 480
rect 4158 0 4214 480
rect 4526 0 4582 480
rect 4986 0 5042 480
rect 5354 0 5410 480
rect 5722 0 5778 480
rect 6182 0 6238 480
rect 6550 0 6606 480
rect 6918 0 6974 480
rect 7378 0 7434 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8574 0 8630 480
rect 8942 0 8998 480
rect 9402 0 9458 480
rect 9770 0 9826 480
rect 10138 0 10194 480
rect 10598 0 10654 480
rect 10966 0 11022 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12162 0 12218 480
rect 12530 0 12586 480
rect 12990 0 13046 480
rect 13358 0 13414 480
rect 13726 0 13782 480
rect 14186 0 14242 480
rect 14554 0 14610 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15750 0 15806 480
<< via2 >>
rect 570 35808 626 35864
rect 1490 36352 1546 36408
rect 2686 38664 2742 38720
rect 2594 35264 2650 35320
rect 1766 35128 1822 35184
rect 1582 34040 1638 34096
rect 1398 33496 1454 33552
rect 1582 31592 1638 31648
rect 1582 29300 1638 29336
rect 1582 29280 1584 29300
rect 1584 29280 1636 29300
rect 1636 29280 1638 29300
rect 1950 33380 2006 33416
rect 1950 33360 1952 33380
rect 1952 33360 2004 33380
rect 2004 33360 2006 33380
rect 2410 30232 2466 30288
rect 2318 29028 2374 29064
rect 2318 29008 2320 29028
rect 2320 29008 2372 29028
rect 2372 29008 2374 29028
rect 1582 26968 1638 27024
rect 2226 26832 2282 26888
rect 1582 24520 1638 24576
rect 3622 37018 3678 37020
rect 3702 37018 3758 37020
rect 3782 37018 3838 37020
rect 3862 37018 3918 37020
rect 3622 36966 3648 37018
rect 3648 36966 3678 37018
rect 3702 36966 3712 37018
rect 3712 36966 3758 37018
rect 3782 36966 3828 37018
rect 3828 36966 3838 37018
rect 3862 36966 3892 37018
rect 3892 36966 3918 37018
rect 3622 36964 3678 36966
rect 3702 36964 3758 36966
rect 3782 36964 3838 36966
rect 3862 36964 3918 36966
rect 3622 35930 3678 35932
rect 3702 35930 3758 35932
rect 3782 35930 3838 35932
rect 3862 35930 3918 35932
rect 3622 35878 3648 35930
rect 3648 35878 3678 35930
rect 3702 35878 3712 35930
rect 3712 35878 3758 35930
rect 3782 35878 3828 35930
rect 3828 35878 3838 35930
rect 3862 35878 3892 35930
rect 3892 35878 3918 35930
rect 3622 35876 3678 35878
rect 3702 35876 3758 35878
rect 3782 35876 3838 35878
rect 3862 35876 3918 35878
rect 3422 35828 3478 35864
rect 3422 35808 3424 35828
rect 3424 35808 3476 35828
rect 3476 35808 3478 35828
rect 2594 32272 2650 32328
rect 2594 28872 2650 28928
rect 2502 25200 2558 25256
rect 2778 27532 2834 27568
rect 2778 27512 2780 27532
rect 2780 27512 2832 27532
rect 2832 27512 2834 27532
rect 1674 22228 1730 22264
rect 1674 22208 1676 22228
rect 1676 22208 1728 22228
rect 1728 22208 1730 22228
rect 1582 21936 1638 21992
rect 1950 21412 2006 21448
rect 1950 21392 1952 21412
rect 1952 21392 2004 21412
rect 2004 21392 2006 21412
rect 1582 19896 1638 19952
rect 1950 17720 2006 17776
rect 1582 17584 1638 17640
rect 2410 16788 2466 16824
rect 2410 16768 2412 16788
rect 2412 16768 2464 16788
rect 2464 16768 2466 16788
rect 1398 16088 1454 16144
rect 1490 15136 1546 15192
rect 3622 34842 3678 34844
rect 3702 34842 3758 34844
rect 3782 34842 3838 34844
rect 3862 34842 3918 34844
rect 3622 34790 3648 34842
rect 3648 34790 3678 34842
rect 3702 34790 3712 34842
rect 3712 34790 3758 34842
rect 3782 34790 3828 34842
rect 3828 34790 3838 34842
rect 3862 34790 3892 34842
rect 3892 34790 3918 34842
rect 3622 34788 3678 34790
rect 3702 34788 3758 34790
rect 3782 34788 3838 34790
rect 3862 34788 3918 34790
rect 3622 33754 3678 33756
rect 3702 33754 3758 33756
rect 3782 33754 3838 33756
rect 3862 33754 3918 33756
rect 3622 33702 3648 33754
rect 3648 33702 3678 33754
rect 3702 33702 3712 33754
rect 3712 33702 3758 33754
rect 3782 33702 3828 33754
rect 3828 33702 3838 33754
rect 3862 33702 3892 33754
rect 3892 33702 3918 33754
rect 3622 33700 3678 33702
rect 3702 33700 3758 33702
rect 3782 33700 3838 33702
rect 3862 33700 3918 33702
rect 3622 32666 3678 32668
rect 3702 32666 3758 32668
rect 3782 32666 3838 32668
rect 3862 32666 3918 32668
rect 3622 32614 3648 32666
rect 3648 32614 3678 32666
rect 3702 32614 3712 32666
rect 3712 32614 3758 32666
rect 3782 32614 3828 32666
rect 3828 32614 3838 32666
rect 3862 32614 3892 32666
rect 3892 32614 3918 32666
rect 3622 32612 3678 32614
rect 3702 32612 3758 32614
rect 3782 32612 3838 32614
rect 3862 32612 3918 32614
rect 3698 32408 3754 32464
rect 3606 32172 3608 32192
rect 3608 32172 3660 32192
rect 3660 32172 3662 32192
rect 3606 32136 3662 32172
rect 3622 31578 3678 31580
rect 3702 31578 3758 31580
rect 3782 31578 3838 31580
rect 3862 31578 3918 31580
rect 3622 31526 3648 31578
rect 3648 31526 3678 31578
rect 3702 31526 3712 31578
rect 3712 31526 3758 31578
rect 3782 31526 3828 31578
rect 3828 31526 3838 31578
rect 3862 31526 3892 31578
rect 3892 31526 3918 31578
rect 3622 31524 3678 31526
rect 3702 31524 3758 31526
rect 3782 31524 3838 31526
rect 3862 31524 3918 31526
rect 3622 30490 3678 30492
rect 3702 30490 3758 30492
rect 3782 30490 3838 30492
rect 3862 30490 3918 30492
rect 3622 30438 3648 30490
rect 3648 30438 3678 30490
rect 3702 30438 3712 30490
rect 3712 30438 3758 30490
rect 3782 30438 3828 30490
rect 3828 30438 3838 30490
rect 3862 30438 3892 30490
rect 3892 30438 3918 30490
rect 3622 30436 3678 30438
rect 3702 30436 3758 30438
rect 3782 30436 3838 30438
rect 3862 30436 3918 30438
rect 4066 33632 4122 33688
rect 4526 35672 4582 35728
rect 3622 29402 3678 29404
rect 3702 29402 3758 29404
rect 3782 29402 3838 29404
rect 3862 29402 3918 29404
rect 3622 29350 3648 29402
rect 3648 29350 3678 29402
rect 3702 29350 3712 29402
rect 3712 29350 3758 29402
rect 3782 29350 3828 29402
rect 3828 29350 3838 29402
rect 3862 29350 3892 29402
rect 3892 29350 3918 29402
rect 3622 29348 3678 29350
rect 3702 29348 3758 29350
rect 3782 29348 3838 29350
rect 3862 29348 3918 29350
rect 4342 30096 4398 30152
rect 3622 28314 3678 28316
rect 3702 28314 3758 28316
rect 3782 28314 3838 28316
rect 3862 28314 3918 28316
rect 3622 28262 3648 28314
rect 3648 28262 3678 28314
rect 3702 28262 3712 28314
rect 3712 28262 3758 28314
rect 3782 28262 3828 28314
rect 3828 28262 3838 28314
rect 3862 28262 3892 28314
rect 3892 28262 3918 28314
rect 3622 28260 3678 28262
rect 3702 28260 3758 28262
rect 3782 28260 3838 28262
rect 3862 28260 3918 28262
rect 4250 28056 4306 28112
rect 3622 27226 3678 27228
rect 3702 27226 3758 27228
rect 3782 27226 3838 27228
rect 3862 27226 3918 27228
rect 3622 27174 3648 27226
rect 3648 27174 3678 27226
rect 3702 27174 3712 27226
rect 3712 27174 3758 27226
rect 3782 27174 3828 27226
rect 3828 27174 3838 27226
rect 3862 27174 3892 27226
rect 3892 27174 3918 27226
rect 3622 27172 3678 27174
rect 3702 27172 3758 27174
rect 3782 27172 3838 27174
rect 3862 27172 3918 27174
rect 3622 26138 3678 26140
rect 3702 26138 3758 26140
rect 3782 26138 3838 26140
rect 3862 26138 3918 26140
rect 3622 26086 3648 26138
rect 3648 26086 3678 26138
rect 3702 26086 3712 26138
rect 3712 26086 3758 26138
rect 3782 26086 3828 26138
rect 3828 26086 3838 26138
rect 3862 26086 3892 26138
rect 3892 26086 3918 26138
rect 3622 26084 3678 26086
rect 3702 26084 3758 26086
rect 3782 26084 3838 26086
rect 3862 26084 3918 26086
rect 3622 25050 3678 25052
rect 3702 25050 3758 25052
rect 3782 25050 3838 25052
rect 3862 25050 3918 25052
rect 3622 24998 3648 25050
rect 3648 24998 3678 25050
rect 3702 24998 3712 25050
rect 3712 24998 3758 25050
rect 3782 24998 3828 25050
rect 3828 24998 3838 25050
rect 3862 24998 3892 25050
rect 3892 24998 3918 25050
rect 3622 24996 3678 24998
rect 3702 24996 3758 24998
rect 3782 24996 3838 24998
rect 3862 24996 3918 24998
rect 3622 23962 3678 23964
rect 3702 23962 3758 23964
rect 3782 23962 3838 23964
rect 3862 23962 3918 23964
rect 3622 23910 3648 23962
rect 3648 23910 3678 23962
rect 3702 23910 3712 23962
rect 3712 23910 3758 23962
rect 3782 23910 3828 23962
rect 3828 23910 3838 23962
rect 3862 23910 3892 23962
rect 3892 23910 3918 23962
rect 3622 23908 3678 23910
rect 3702 23908 3758 23910
rect 3782 23908 3838 23910
rect 3862 23908 3918 23910
rect 3146 17584 3202 17640
rect 3622 22874 3678 22876
rect 3702 22874 3758 22876
rect 3782 22874 3838 22876
rect 3862 22874 3918 22876
rect 3622 22822 3648 22874
rect 3648 22822 3678 22874
rect 3702 22822 3712 22874
rect 3712 22822 3758 22874
rect 3782 22822 3828 22874
rect 3828 22822 3838 22874
rect 3862 22822 3892 22874
rect 3892 22822 3918 22874
rect 3622 22820 3678 22822
rect 3702 22820 3758 22822
rect 3782 22820 3838 22822
rect 3862 22820 3918 22822
rect 3622 21786 3678 21788
rect 3702 21786 3758 21788
rect 3782 21786 3838 21788
rect 3862 21786 3918 21788
rect 3622 21734 3648 21786
rect 3648 21734 3678 21786
rect 3702 21734 3712 21786
rect 3712 21734 3758 21786
rect 3782 21734 3828 21786
rect 3828 21734 3838 21786
rect 3862 21734 3892 21786
rect 3892 21734 3918 21786
rect 3622 21732 3678 21734
rect 3702 21732 3758 21734
rect 3782 21732 3838 21734
rect 3862 21732 3918 21734
rect 3622 20698 3678 20700
rect 3702 20698 3758 20700
rect 3782 20698 3838 20700
rect 3862 20698 3918 20700
rect 3622 20646 3648 20698
rect 3648 20646 3678 20698
rect 3702 20646 3712 20698
rect 3712 20646 3758 20698
rect 3782 20646 3828 20698
rect 3828 20646 3838 20698
rect 3862 20646 3892 20698
rect 3892 20646 3918 20698
rect 3622 20644 3678 20646
rect 3702 20644 3758 20646
rect 3782 20644 3838 20646
rect 3862 20644 3918 20646
rect 3422 19352 3478 19408
rect 3622 19610 3678 19612
rect 3702 19610 3758 19612
rect 3782 19610 3838 19612
rect 3862 19610 3918 19612
rect 3622 19558 3648 19610
rect 3648 19558 3678 19610
rect 3702 19558 3712 19610
rect 3712 19558 3758 19610
rect 3782 19558 3828 19610
rect 3828 19558 3838 19610
rect 3862 19558 3892 19610
rect 3892 19558 3918 19610
rect 3622 19556 3678 19558
rect 3702 19556 3758 19558
rect 3782 19556 3838 19558
rect 3862 19556 3918 19558
rect 3622 18522 3678 18524
rect 3702 18522 3758 18524
rect 3782 18522 3838 18524
rect 3862 18522 3918 18524
rect 3622 18470 3648 18522
rect 3648 18470 3678 18522
rect 3702 18470 3712 18522
rect 3712 18470 3758 18522
rect 3782 18470 3828 18522
rect 3828 18470 3838 18522
rect 3862 18470 3892 18522
rect 3892 18470 3918 18522
rect 3622 18468 3678 18470
rect 3702 18468 3758 18470
rect 3782 18468 3838 18470
rect 3862 18468 3918 18470
rect 3622 17434 3678 17436
rect 3702 17434 3758 17436
rect 3782 17434 3838 17436
rect 3862 17434 3918 17436
rect 3622 17382 3648 17434
rect 3648 17382 3678 17434
rect 3702 17382 3712 17434
rect 3712 17382 3758 17434
rect 3782 17382 3828 17434
rect 3828 17382 3838 17434
rect 3862 17382 3892 17434
rect 3892 17382 3918 17434
rect 3622 17380 3678 17382
rect 3702 17380 3758 17382
rect 3782 17380 3838 17382
rect 3862 17380 3918 17382
rect 3622 16346 3678 16348
rect 3702 16346 3758 16348
rect 3782 16346 3838 16348
rect 3862 16346 3918 16348
rect 3622 16294 3648 16346
rect 3648 16294 3678 16346
rect 3702 16294 3712 16346
rect 3712 16294 3758 16346
rect 3782 16294 3828 16346
rect 3828 16294 3838 16346
rect 3862 16294 3892 16346
rect 3892 16294 3918 16346
rect 3622 16292 3678 16294
rect 3702 16292 3758 16294
rect 3782 16292 3838 16294
rect 3862 16292 3918 16294
rect 3622 15258 3678 15260
rect 3702 15258 3758 15260
rect 3782 15258 3838 15260
rect 3862 15258 3918 15260
rect 3622 15206 3648 15258
rect 3648 15206 3678 15258
rect 3702 15206 3712 15258
rect 3712 15206 3758 15258
rect 3782 15206 3828 15258
rect 3828 15206 3838 15258
rect 3862 15206 3892 15258
rect 3892 15206 3918 15258
rect 3622 15204 3678 15206
rect 3702 15204 3758 15206
rect 3782 15204 3838 15206
rect 3862 15204 3918 15206
rect 3330 14592 3386 14648
rect 3622 14170 3678 14172
rect 3702 14170 3758 14172
rect 3782 14170 3838 14172
rect 3862 14170 3918 14172
rect 3622 14118 3648 14170
rect 3648 14118 3678 14170
rect 3702 14118 3712 14170
rect 3712 14118 3758 14170
rect 3782 14118 3828 14170
rect 3828 14118 3838 14170
rect 3862 14118 3892 14170
rect 3892 14118 3918 14170
rect 3622 14116 3678 14118
rect 3702 14116 3758 14118
rect 3782 14116 3838 14118
rect 3862 14116 3918 14118
rect 1582 12824 1638 12880
rect 3622 13082 3678 13084
rect 3702 13082 3758 13084
rect 3782 13082 3838 13084
rect 3862 13082 3918 13084
rect 3622 13030 3648 13082
rect 3648 13030 3678 13082
rect 3702 13030 3712 13082
rect 3712 13030 3758 13082
rect 3782 13030 3828 13082
rect 3828 13030 3838 13082
rect 3862 13030 3892 13082
rect 3892 13030 3918 13082
rect 3622 13028 3678 13030
rect 3702 13028 3758 13030
rect 3782 13028 3838 13030
rect 3862 13028 3918 13030
rect 1674 12708 1730 12744
rect 1674 12688 1676 12708
rect 1676 12688 1728 12708
rect 1728 12688 1730 12708
rect 3622 11994 3678 11996
rect 3702 11994 3758 11996
rect 3782 11994 3838 11996
rect 3862 11994 3918 11996
rect 3622 11942 3648 11994
rect 3648 11942 3678 11994
rect 3702 11942 3712 11994
rect 3712 11942 3758 11994
rect 3782 11942 3828 11994
rect 3828 11942 3838 11994
rect 3862 11942 3892 11994
rect 3892 11942 3918 11994
rect 3622 11940 3678 11942
rect 3702 11940 3758 11942
rect 3782 11940 3838 11942
rect 3862 11940 3918 11942
rect 1582 10512 1638 10568
rect 3622 10906 3678 10908
rect 3702 10906 3758 10908
rect 3782 10906 3838 10908
rect 3862 10906 3918 10908
rect 3622 10854 3648 10906
rect 3648 10854 3678 10906
rect 3702 10854 3712 10906
rect 3712 10854 3758 10906
rect 3782 10854 3828 10906
rect 3828 10854 3838 10906
rect 3862 10854 3892 10906
rect 3892 10854 3918 10906
rect 3622 10852 3678 10854
rect 3702 10852 3758 10854
rect 3782 10852 3838 10854
rect 3862 10852 3918 10854
rect 3146 8336 3202 8392
rect 2778 8064 2834 8120
rect 570 4120 626 4176
rect 2134 5616 2190 5672
rect 1950 4564 1952 4584
rect 1952 4564 2004 4584
rect 2004 4564 2006 4584
rect 1582 3440 1638 3496
rect 1950 4528 2006 4564
rect 2410 5208 2466 5264
rect 2410 5092 2466 5128
rect 2410 5072 2412 5092
rect 2412 5072 2464 5092
rect 2464 5072 2466 5092
rect 3054 6060 3056 6080
rect 3056 6060 3108 6080
rect 3108 6060 3110 6080
rect 3054 6024 3110 6060
rect 2686 5752 2742 5808
rect 1858 3712 1914 3768
rect 1766 3440 1822 3496
rect 1674 2488 1730 2544
rect 1950 2760 2006 2816
rect 1490 1128 1546 1184
rect 2226 3068 2228 3088
rect 2228 3068 2280 3088
rect 2280 3068 2282 3088
rect 2226 3032 2282 3068
rect 3054 4120 3110 4176
rect 2870 3596 2926 3632
rect 2870 3576 2872 3596
rect 2872 3576 2924 3596
rect 2924 3576 2926 3596
rect 5078 35284 5134 35320
rect 5078 35264 5080 35284
rect 5080 35264 5132 35284
rect 5132 35264 5134 35284
rect 4986 30232 5042 30288
rect 5078 29688 5134 29744
rect 4894 29008 4950 29064
rect 4894 24812 4950 24848
rect 4894 24792 4896 24812
rect 4896 24792 4948 24812
rect 4948 24792 4950 24812
rect 4802 23840 4858 23896
rect 4618 20848 4674 20904
rect 4710 19796 4712 19816
rect 4712 19796 4764 19816
rect 4764 19796 4766 19816
rect 4710 19760 4766 19796
rect 4250 17620 4252 17640
rect 4252 17620 4304 17640
rect 4304 17620 4306 17640
rect 4250 17584 4306 17620
rect 4526 16788 4582 16824
rect 4526 16768 4528 16788
rect 4528 16768 4580 16788
rect 4580 16768 4582 16788
rect 4434 15000 4490 15056
rect 4618 13776 4674 13832
rect 3622 9818 3678 9820
rect 3702 9818 3758 9820
rect 3782 9818 3838 9820
rect 3862 9818 3918 9820
rect 3622 9766 3648 9818
rect 3648 9766 3678 9818
rect 3702 9766 3712 9818
rect 3712 9766 3758 9818
rect 3782 9766 3828 9818
rect 3828 9766 3838 9818
rect 3862 9766 3892 9818
rect 3892 9766 3918 9818
rect 3622 9764 3678 9766
rect 3702 9764 3758 9766
rect 3782 9764 3838 9766
rect 3862 9764 3918 9766
rect 3330 9460 3332 9480
rect 3332 9460 3384 9480
rect 3384 9460 3386 9480
rect 3330 9424 3386 9460
rect 3622 8730 3678 8732
rect 3702 8730 3758 8732
rect 3782 8730 3838 8732
rect 3862 8730 3918 8732
rect 3622 8678 3648 8730
rect 3648 8678 3678 8730
rect 3702 8678 3712 8730
rect 3712 8678 3758 8730
rect 3782 8678 3828 8730
rect 3828 8678 3838 8730
rect 3862 8678 3892 8730
rect 3892 8678 3918 8730
rect 3622 8676 3678 8678
rect 3702 8676 3758 8678
rect 3782 8676 3838 8678
rect 3862 8676 3918 8678
rect 3790 8492 3846 8528
rect 3790 8472 3792 8492
rect 3792 8472 3844 8492
rect 3844 8472 3846 8492
rect 3622 7642 3678 7644
rect 3702 7642 3758 7644
rect 3782 7642 3838 7644
rect 3862 7642 3918 7644
rect 3622 7590 3648 7642
rect 3648 7590 3678 7642
rect 3702 7590 3712 7642
rect 3712 7590 3758 7642
rect 3782 7590 3828 7642
rect 3828 7590 3838 7642
rect 3862 7590 3892 7642
rect 3892 7590 3918 7642
rect 3622 7588 3678 7590
rect 3702 7588 3758 7590
rect 3782 7588 3838 7590
rect 3862 7588 3918 7590
rect 3622 6554 3678 6556
rect 3702 6554 3758 6556
rect 3782 6554 3838 6556
rect 3862 6554 3918 6556
rect 3622 6502 3648 6554
rect 3648 6502 3678 6554
rect 3702 6502 3712 6554
rect 3712 6502 3758 6554
rect 3782 6502 3828 6554
rect 3828 6502 3838 6554
rect 3862 6502 3892 6554
rect 3892 6502 3918 6554
rect 3622 6500 3678 6502
rect 3702 6500 3758 6502
rect 3782 6500 3838 6502
rect 3862 6500 3918 6502
rect 3622 5466 3678 5468
rect 3702 5466 3758 5468
rect 3782 5466 3838 5468
rect 3862 5466 3918 5468
rect 3622 5414 3648 5466
rect 3648 5414 3678 5466
rect 3702 5414 3712 5466
rect 3712 5414 3758 5466
rect 3782 5414 3828 5466
rect 3828 5414 3838 5466
rect 3862 5414 3892 5466
rect 3892 5414 3918 5466
rect 3622 5412 3678 5414
rect 3702 5412 3758 5414
rect 3782 5412 3838 5414
rect 3862 5412 3918 5414
rect 3622 4378 3678 4380
rect 3702 4378 3758 4380
rect 3782 4378 3838 4380
rect 3862 4378 3918 4380
rect 3622 4326 3648 4378
rect 3648 4326 3678 4378
rect 3702 4326 3712 4378
rect 3712 4326 3758 4378
rect 3782 4326 3828 4378
rect 3828 4326 3838 4378
rect 3862 4326 3892 4378
rect 3892 4326 3918 4378
rect 3622 4324 3678 4326
rect 3702 4324 3758 4326
rect 3782 4324 3838 4326
rect 3862 4324 3918 4326
rect 6289 37562 6345 37564
rect 6369 37562 6425 37564
rect 6449 37562 6505 37564
rect 6529 37562 6585 37564
rect 6289 37510 6315 37562
rect 6315 37510 6345 37562
rect 6369 37510 6379 37562
rect 6379 37510 6425 37562
rect 6449 37510 6495 37562
rect 6495 37510 6505 37562
rect 6529 37510 6559 37562
rect 6559 37510 6585 37562
rect 6289 37508 6345 37510
rect 6369 37508 6425 37510
rect 6449 37508 6505 37510
rect 6529 37508 6585 37510
rect 6289 36474 6345 36476
rect 6369 36474 6425 36476
rect 6449 36474 6505 36476
rect 6529 36474 6585 36476
rect 6289 36422 6315 36474
rect 6315 36422 6345 36474
rect 6369 36422 6379 36474
rect 6379 36422 6425 36474
rect 6449 36422 6495 36474
rect 6495 36422 6505 36474
rect 6529 36422 6559 36474
rect 6559 36422 6585 36474
rect 6289 36420 6345 36422
rect 6369 36420 6425 36422
rect 6449 36420 6505 36422
rect 6529 36420 6585 36422
rect 5722 29144 5778 29200
rect 5722 24928 5778 24984
rect 5630 24656 5686 24712
rect 5170 23160 5226 23216
rect 5170 22208 5226 22264
rect 5354 21528 5410 21584
rect 4894 13776 4950 13832
rect 5170 19352 5226 19408
rect 5078 14612 5134 14648
rect 5078 14592 5080 14612
rect 5080 14592 5132 14612
rect 5132 14592 5134 14612
rect 4986 11600 5042 11656
rect 5722 21256 5778 21312
rect 5446 17176 5502 17232
rect 5354 17076 5356 17096
rect 5356 17076 5408 17096
rect 5408 17076 5410 17096
rect 5354 17040 5410 17076
rect 5354 14492 5356 14512
rect 5356 14492 5408 14512
rect 5408 14492 5410 14512
rect 5354 14456 5410 14492
rect 5170 9968 5226 10024
rect 4986 6180 5042 6216
rect 4986 6160 4988 6180
rect 4988 6160 5040 6180
rect 5040 6160 5042 6180
rect 4894 4664 4950 4720
rect 3622 3290 3678 3292
rect 3702 3290 3758 3292
rect 3782 3290 3838 3292
rect 3862 3290 3918 3292
rect 3622 3238 3648 3290
rect 3648 3238 3678 3290
rect 3702 3238 3712 3290
rect 3712 3238 3758 3290
rect 3782 3238 3828 3290
rect 3828 3238 3838 3290
rect 3862 3238 3892 3290
rect 3892 3238 3918 3290
rect 3622 3236 3678 3238
rect 3702 3236 3758 3238
rect 3782 3236 3838 3238
rect 3862 3236 3918 3238
rect 4158 2896 4214 2952
rect 3622 2202 3678 2204
rect 3702 2202 3758 2204
rect 3782 2202 3838 2204
rect 3862 2202 3918 2204
rect 3622 2150 3648 2202
rect 3648 2150 3678 2202
rect 3702 2150 3712 2202
rect 3712 2150 3758 2202
rect 3782 2150 3828 2202
rect 3828 2150 3838 2202
rect 3862 2150 3892 2202
rect 3892 2150 3918 2202
rect 3622 2148 3678 2150
rect 3702 2148 3758 2150
rect 3782 2148 3838 2150
rect 3862 2148 3918 2150
rect 4618 3576 4674 3632
rect 5262 7268 5318 7304
rect 5262 7248 5264 7268
rect 5264 7248 5316 7268
rect 5316 7248 5318 7268
rect 5262 6704 5318 6760
rect 6289 35386 6345 35388
rect 6369 35386 6425 35388
rect 6449 35386 6505 35388
rect 6529 35386 6585 35388
rect 6289 35334 6315 35386
rect 6315 35334 6345 35386
rect 6369 35334 6379 35386
rect 6379 35334 6425 35386
rect 6449 35334 6495 35386
rect 6495 35334 6505 35386
rect 6529 35334 6559 35386
rect 6559 35334 6585 35386
rect 6289 35332 6345 35334
rect 6369 35332 6425 35334
rect 6449 35332 6505 35334
rect 6529 35332 6585 35334
rect 7562 35128 7618 35184
rect 6289 34298 6345 34300
rect 6369 34298 6425 34300
rect 6449 34298 6505 34300
rect 6529 34298 6585 34300
rect 6289 34246 6315 34298
rect 6315 34246 6345 34298
rect 6369 34246 6379 34298
rect 6379 34246 6425 34298
rect 6449 34246 6495 34298
rect 6495 34246 6505 34298
rect 6529 34246 6559 34298
rect 6559 34246 6585 34298
rect 6289 34244 6345 34246
rect 6369 34244 6425 34246
rect 6449 34244 6505 34246
rect 6529 34244 6585 34246
rect 6642 33632 6698 33688
rect 6289 33210 6345 33212
rect 6369 33210 6425 33212
rect 6449 33210 6505 33212
rect 6529 33210 6585 33212
rect 6289 33158 6315 33210
rect 6315 33158 6345 33210
rect 6369 33158 6379 33210
rect 6379 33158 6425 33210
rect 6449 33158 6495 33210
rect 6495 33158 6505 33210
rect 6529 33158 6559 33210
rect 6559 33158 6585 33210
rect 6289 33156 6345 33158
rect 6369 33156 6425 33158
rect 6449 33156 6505 33158
rect 6529 33156 6585 33158
rect 6090 32136 6146 32192
rect 6289 32122 6345 32124
rect 6369 32122 6425 32124
rect 6449 32122 6505 32124
rect 6529 32122 6585 32124
rect 6289 32070 6315 32122
rect 6315 32070 6345 32122
rect 6369 32070 6379 32122
rect 6379 32070 6425 32122
rect 6449 32070 6495 32122
rect 6495 32070 6505 32122
rect 6529 32070 6559 32122
rect 6559 32070 6585 32122
rect 6289 32068 6345 32070
rect 6369 32068 6425 32070
rect 6449 32068 6505 32070
rect 6529 32068 6585 32070
rect 6734 33224 6790 33280
rect 6289 31034 6345 31036
rect 6369 31034 6425 31036
rect 6449 31034 6505 31036
rect 6529 31034 6585 31036
rect 6289 30982 6315 31034
rect 6315 30982 6345 31034
rect 6369 30982 6379 31034
rect 6379 30982 6425 31034
rect 6449 30982 6495 31034
rect 6495 30982 6505 31034
rect 6529 30982 6559 31034
rect 6559 30982 6585 31034
rect 6289 30980 6345 30982
rect 6369 30980 6425 30982
rect 6449 30980 6505 30982
rect 6529 30980 6585 30982
rect 6182 30116 6238 30152
rect 6182 30096 6184 30116
rect 6184 30096 6236 30116
rect 6236 30096 6238 30116
rect 6289 29946 6345 29948
rect 6369 29946 6425 29948
rect 6449 29946 6505 29948
rect 6529 29946 6585 29948
rect 6289 29894 6315 29946
rect 6315 29894 6345 29946
rect 6369 29894 6379 29946
rect 6379 29894 6425 29946
rect 6449 29894 6495 29946
rect 6495 29894 6505 29946
rect 6529 29894 6559 29946
rect 6559 29894 6585 29946
rect 6289 29892 6345 29894
rect 6369 29892 6425 29894
rect 6449 29892 6505 29894
rect 6529 29892 6585 29894
rect 6289 28858 6345 28860
rect 6369 28858 6425 28860
rect 6449 28858 6505 28860
rect 6529 28858 6585 28860
rect 6289 28806 6315 28858
rect 6315 28806 6345 28858
rect 6369 28806 6379 28858
rect 6379 28806 6425 28858
rect 6449 28806 6495 28858
rect 6495 28806 6505 28858
rect 6529 28806 6559 28858
rect 6559 28806 6585 28858
rect 6289 28804 6345 28806
rect 6369 28804 6425 28806
rect 6449 28804 6505 28806
rect 6529 28804 6585 28806
rect 6182 27920 6238 27976
rect 6289 27770 6345 27772
rect 6369 27770 6425 27772
rect 6449 27770 6505 27772
rect 6529 27770 6585 27772
rect 6289 27718 6315 27770
rect 6315 27718 6345 27770
rect 6369 27718 6379 27770
rect 6379 27718 6425 27770
rect 6449 27718 6495 27770
rect 6495 27718 6505 27770
rect 6529 27718 6559 27770
rect 6559 27718 6585 27770
rect 6289 27716 6345 27718
rect 6369 27716 6425 27718
rect 6449 27716 6505 27718
rect 6529 27716 6585 27718
rect 5814 14864 5870 14920
rect 6289 26682 6345 26684
rect 6369 26682 6425 26684
rect 6449 26682 6505 26684
rect 6529 26682 6585 26684
rect 6289 26630 6315 26682
rect 6315 26630 6345 26682
rect 6369 26630 6379 26682
rect 6379 26630 6425 26682
rect 6449 26630 6495 26682
rect 6495 26630 6505 26682
rect 6529 26630 6559 26682
rect 6559 26630 6585 26682
rect 6289 26628 6345 26630
rect 6369 26628 6425 26630
rect 6449 26628 6505 26630
rect 6529 26628 6585 26630
rect 6289 25594 6345 25596
rect 6369 25594 6425 25596
rect 6449 25594 6505 25596
rect 6529 25594 6585 25596
rect 6289 25542 6315 25594
rect 6315 25542 6345 25594
rect 6369 25542 6379 25594
rect 6379 25542 6425 25594
rect 6449 25542 6495 25594
rect 6495 25542 6505 25594
rect 6529 25542 6559 25594
rect 6559 25542 6585 25594
rect 6289 25540 6345 25542
rect 6369 25540 6425 25542
rect 6449 25540 6505 25542
rect 6529 25540 6585 25542
rect 6289 24506 6345 24508
rect 6369 24506 6425 24508
rect 6449 24506 6505 24508
rect 6529 24506 6585 24508
rect 6289 24454 6315 24506
rect 6315 24454 6345 24506
rect 6369 24454 6379 24506
rect 6379 24454 6425 24506
rect 6449 24454 6495 24506
rect 6495 24454 6505 24506
rect 6529 24454 6559 24506
rect 6559 24454 6585 24506
rect 6289 24452 6345 24454
rect 6369 24452 6425 24454
rect 6449 24452 6505 24454
rect 6529 24452 6585 24454
rect 6289 23418 6345 23420
rect 6369 23418 6425 23420
rect 6449 23418 6505 23420
rect 6529 23418 6585 23420
rect 6289 23366 6315 23418
rect 6315 23366 6345 23418
rect 6369 23366 6379 23418
rect 6379 23366 6425 23418
rect 6449 23366 6495 23418
rect 6495 23366 6505 23418
rect 6529 23366 6559 23418
rect 6559 23366 6585 23418
rect 6289 23364 6345 23366
rect 6369 23364 6425 23366
rect 6449 23364 6505 23366
rect 6529 23364 6585 23366
rect 6289 22330 6345 22332
rect 6369 22330 6425 22332
rect 6449 22330 6505 22332
rect 6529 22330 6585 22332
rect 6289 22278 6315 22330
rect 6315 22278 6345 22330
rect 6369 22278 6379 22330
rect 6379 22278 6425 22330
rect 6449 22278 6495 22330
rect 6495 22278 6505 22330
rect 6529 22278 6559 22330
rect 6559 22278 6585 22330
rect 6289 22276 6345 22278
rect 6369 22276 6425 22278
rect 6449 22276 6505 22278
rect 6529 22276 6585 22278
rect 6826 30932 6882 30968
rect 6826 30912 6828 30932
rect 6828 30912 6880 30932
rect 6880 30912 6882 30932
rect 7562 33496 7618 33552
rect 7286 32308 7288 32328
rect 7288 32308 7340 32328
rect 7340 32308 7342 32328
rect 7286 32272 7342 32308
rect 7194 31900 7196 31920
rect 7196 31900 7248 31920
rect 7248 31900 7250 31920
rect 7194 31864 7250 31900
rect 7194 29996 7196 30016
rect 7196 29996 7248 30016
rect 7248 29996 7250 30016
rect 7194 29960 7250 29996
rect 7286 29044 7288 29064
rect 7288 29044 7340 29064
rect 7340 29044 7342 29064
rect 7286 29008 7342 29044
rect 6826 27648 6882 27704
rect 6734 23840 6790 23896
rect 6642 21528 6698 21584
rect 6289 21242 6345 21244
rect 6369 21242 6425 21244
rect 6449 21242 6505 21244
rect 6529 21242 6585 21244
rect 6289 21190 6315 21242
rect 6315 21190 6345 21242
rect 6369 21190 6379 21242
rect 6379 21190 6425 21242
rect 6449 21190 6495 21242
rect 6495 21190 6505 21242
rect 6529 21190 6559 21242
rect 6559 21190 6585 21242
rect 6289 21188 6345 21190
rect 6369 21188 6425 21190
rect 6449 21188 6505 21190
rect 6529 21188 6585 21190
rect 6289 20154 6345 20156
rect 6369 20154 6425 20156
rect 6449 20154 6505 20156
rect 6529 20154 6585 20156
rect 6289 20102 6315 20154
rect 6315 20102 6345 20154
rect 6369 20102 6379 20154
rect 6379 20102 6425 20154
rect 6449 20102 6495 20154
rect 6495 20102 6505 20154
rect 6529 20102 6559 20154
rect 6559 20102 6585 20154
rect 6289 20100 6345 20102
rect 6369 20100 6425 20102
rect 6449 20100 6505 20102
rect 6529 20100 6585 20102
rect 6289 19066 6345 19068
rect 6369 19066 6425 19068
rect 6449 19066 6505 19068
rect 6529 19066 6585 19068
rect 6289 19014 6315 19066
rect 6315 19014 6345 19066
rect 6369 19014 6379 19066
rect 6379 19014 6425 19066
rect 6449 19014 6495 19066
rect 6495 19014 6505 19066
rect 6529 19014 6559 19066
rect 6559 19014 6585 19066
rect 6289 19012 6345 19014
rect 6369 19012 6425 19014
rect 6449 19012 6505 19014
rect 6529 19012 6585 19014
rect 6289 17978 6345 17980
rect 6369 17978 6425 17980
rect 6449 17978 6505 17980
rect 6529 17978 6585 17980
rect 6289 17926 6315 17978
rect 6315 17926 6345 17978
rect 6369 17926 6379 17978
rect 6379 17926 6425 17978
rect 6449 17926 6495 17978
rect 6495 17926 6505 17978
rect 6529 17926 6559 17978
rect 6559 17926 6585 17978
rect 6289 17924 6345 17926
rect 6369 17924 6425 17926
rect 6449 17924 6505 17926
rect 6529 17924 6585 17926
rect 6289 16890 6345 16892
rect 6369 16890 6425 16892
rect 6449 16890 6505 16892
rect 6529 16890 6585 16892
rect 6289 16838 6315 16890
rect 6315 16838 6345 16890
rect 6369 16838 6379 16890
rect 6379 16838 6425 16890
rect 6449 16838 6495 16890
rect 6495 16838 6505 16890
rect 6529 16838 6559 16890
rect 6559 16838 6585 16890
rect 6289 16836 6345 16838
rect 6369 16836 6425 16838
rect 6449 16836 6505 16838
rect 6529 16836 6585 16838
rect 6289 15802 6345 15804
rect 6369 15802 6425 15804
rect 6449 15802 6505 15804
rect 6529 15802 6585 15804
rect 6289 15750 6315 15802
rect 6315 15750 6345 15802
rect 6369 15750 6379 15802
rect 6379 15750 6425 15802
rect 6449 15750 6495 15802
rect 6495 15750 6505 15802
rect 6529 15750 6559 15802
rect 6559 15750 6585 15802
rect 6289 15748 6345 15750
rect 6369 15748 6425 15750
rect 6449 15748 6505 15750
rect 6529 15748 6585 15750
rect 6289 14714 6345 14716
rect 6369 14714 6425 14716
rect 6449 14714 6505 14716
rect 6529 14714 6585 14716
rect 6289 14662 6315 14714
rect 6315 14662 6345 14714
rect 6369 14662 6379 14714
rect 6379 14662 6425 14714
rect 6449 14662 6495 14714
rect 6495 14662 6505 14714
rect 6529 14662 6559 14714
rect 6559 14662 6585 14714
rect 6289 14660 6345 14662
rect 6369 14660 6425 14662
rect 6449 14660 6505 14662
rect 6529 14660 6585 14662
rect 6289 13626 6345 13628
rect 6369 13626 6425 13628
rect 6449 13626 6505 13628
rect 6529 13626 6585 13628
rect 6289 13574 6315 13626
rect 6315 13574 6345 13626
rect 6369 13574 6379 13626
rect 6379 13574 6425 13626
rect 6449 13574 6495 13626
rect 6495 13574 6505 13626
rect 6529 13574 6559 13626
rect 6559 13574 6585 13626
rect 6289 13572 6345 13574
rect 6369 13572 6425 13574
rect 6449 13572 6505 13574
rect 6529 13572 6585 13574
rect 7746 34584 7802 34640
rect 7746 33088 7802 33144
rect 8022 32952 8078 33008
rect 8022 31320 8078 31376
rect 7654 27376 7710 27432
rect 7470 26968 7526 27024
rect 7562 24656 7618 24712
rect 8956 37018 9012 37020
rect 9036 37018 9092 37020
rect 9116 37018 9172 37020
rect 9196 37018 9252 37020
rect 8956 36966 8982 37018
rect 8982 36966 9012 37018
rect 9036 36966 9046 37018
rect 9046 36966 9092 37018
rect 9116 36966 9162 37018
rect 9162 36966 9172 37018
rect 9196 36966 9226 37018
rect 9226 36966 9252 37018
rect 8956 36964 9012 36966
rect 9036 36964 9092 36966
rect 9116 36964 9172 36966
rect 9196 36964 9252 36966
rect 8956 35930 9012 35932
rect 9036 35930 9092 35932
rect 9116 35930 9172 35932
rect 9196 35930 9252 35932
rect 8956 35878 8982 35930
rect 8982 35878 9012 35930
rect 9036 35878 9046 35930
rect 9046 35878 9092 35930
rect 9116 35878 9162 35930
rect 9162 35878 9172 35930
rect 9196 35878 9226 35930
rect 9226 35878 9252 35930
rect 8956 35876 9012 35878
rect 9036 35876 9092 35878
rect 9116 35876 9172 35878
rect 9196 35876 9252 35878
rect 8956 34842 9012 34844
rect 9036 34842 9092 34844
rect 9116 34842 9172 34844
rect 9196 34842 9252 34844
rect 8956 34790 8982 34842
rect 8982 34790 9012 34842
rect 9036 34790 9046 34842
rect 9046 34790 9092 34842
rect 9116 34790 9162 34842
rect 9162 34790 9172 34842
rect 9196 34790 9226 34842
rect 9226 34790 9252 34842
rect 8956 34788 9012 34790
rect 9036 34788 9092 34790
rect 9116 34788 9172 34790
rect 9196 34788 9252 34790
rect 8666 32408 8722 32464
rect 7930 26868 7932 26888
rect 7932 26868 7984 26888
rect 7984 26868 7986 26888
rect 7930 26832 7986 26868
rect 8298 27532 8354 27568
rect 8298 27512 8300 27532
rect 8300 27512 8352 27532
rect 8352 27512 8354 27532
rect 7286 22616 7342 22672
rect 8022 23024 8078 23080
rect 7562 20984 7618 21040
rect 8956 33754 9012 33756
rect 9036 33754 9092 33756
rect 9116 33754 9172 33756
rect 9196 33754 9252 33756
rect 8956 33702 8982 33754
rect 8982 33702 9012 33754
rect 9036 33702 9046 33754
rect 9046 33702 9092 33754
rect 9116 33702 9162 33754
rect 9162 33702 9172 33754
rect 9196 33702 9226 33754
rect 9226 33702 9252 33754
rect 8956 33700 9012 33702
rect 9036 33700 9092 33702
rect 9116 33700 9172 33702
rect 9196 33700 9252 33702
rect 9310 33224 9366 33280
rect 8956 32666 9012 32668
rect 9036 32666 9092 32668
rect 9116 32666 9172 32668
rect 9196 32666 9252 32668
rect 8956 32614 8982 32666
rect 8982 32614 9012 32666
rect 9036 32614 9046 32666
rect 9046 32614 9092 32666
rect 9116 32614 9162 32666
rect 9162 32614 9172 32666
rect 9196 32614 9226 32666
rect 9226 32614 9252 32666
rect 8956 32612 9012 32614
rect 9036 32612 9092 32614
rect 9116 32612 9172 32614
rect 9196 32612 9252 32614
rect 8956 31578 9012 31580
rect 9036 31578 9092 31580
rect 9116 31578 9172 31580
rect 9196 31578 9252 31580
rect 8956 31526 8982 31578
rect 8982 31526 9012 31578
rect 9036 31526 9046 31578
rect 9046 31526 9092 31578
rect 9116 31526 9162 31578
rect 9162 31526 9172 31578
rect 9196 31526 9226 31578
rect 9226 31526 9252 31578
rect 8956 31524 9012 31526
rect 9036 31524 9092 31526
rect 9116 31524 9172 31526
rect 9196 31524 9252 31526
rect 8956 30490 9012 30492
rect 9036 30490 9092 30492
rect 9116 30490 9172 30492
rect 9196 30490 9252 30492
rect 8956 30438 8982 30490
rect 8982 30438 9012 30490
rect 9036 30438 9046 30490
rect 9046 30438 9092 30490
rect 9116 30438 9162 30490
rect 9162 30438 9172 30490
rect 9196 30438 9226 30490
rect 9226 30438 9252 30490
rect 8956 30436 9012 30438
rect 9036 30436 9092 30438
rect 9116 30436 9172 30438
rect 9196 30436 9252 30438
rect 8574 26288 8630 26344
rect 7654 19216 7710 19272
rect 8114 19080 8170 19136
rect 7746 17720 7802 17776
rect 7286 16496 7342 16552
rect 7838 16904 7894 16960
rect 7286 14864 7342 14920
rect 7378 14592 7434 14648
rect 7746 15988 7748 16008
rect 7748 15988 7800 16008
rect 7800 15988 7802 16008
rect 7746 15952 7802 15988
rect 6182 12688 6238 12744
rect 6289 12538 6345 12540
rect 6369 12538 6425 12540
rect 6449 12538 6505 12540
rect 6529 12538 6585 12540
rect 6289 12486 6315 12538
rect 6315 12486 6345 12538
rect 6369 12486 6379 12538
rect 6379 12486 6425 12538
rect 6449 12486 6495 12538
rect 6495 12486 6505 12538
rect 6529 12486 6559 12538
rect 6559 12486 6585 12538
rect 6289 12484 6345 12486
rect 6369 12484 6425 12486
rect 6449 12484 6505 12486
rect 6529 12484 6585 12486
rect 6289 11450 6345 11452
rect 6369 11450 6425 11452
rect 6449 11450 6505 11452
rect 6529 11450 6585 11452
rect 6289 11398 6315 11450
rect 6315 11398 6345 11450
rect 6369 11398 6379 11450
rect 6379 11398 6425 11450
rect 6449 11398 6495 11450
rect 6495 11398 6505 11450
rect 6529 11398 6559 11450
rect 6559 11398 6585 11450
rect 6289 11396 6345 11398
rect 6369 11396 6425 11398
rect 6449 11396 6505 11398
rect 6529 11396 6585 11398
rect 6289 10362 6345 10364
rect 6369 10362 6425 10364
rect 6449 10362 6505 10364
rect 6529 10362 6585 10364
rect 6289 10310 6315 10362
rect 6315 10310 6345 10362
rect 6369 10310 6379 10362
rect 6379 10310 6425 10362
rect 6449 10310 6495 10362
rect 6495 10310 6505 10362
rect 6529 10310 6559 10362
rect 6559 10310 6585 10362
rect 6289 10308 6345 10310
rect 6369 10308 6425 10310
rect 6449 10308 6505 10310
rect 6529 10308 6585 10310
rect 6289 9274 6345 9276
rect 6369 9274 6425 9276
rect 6449 9274 6505 9276
rect 6529 9274 6585 9276
rect 6289 9222 6315 9274
rect 6315 9222 6345 9274
rect 6369 9222 6379 9274
rect 6379 9222 6425 9274
rect 6449 9222 6495 9274
rect 6495 9222 6505 9274
rect 6529 9222 6559 9274
rect 6559 9222 6585 9274
rect 6289 9220 6345 9222
rect 6369 9220 6425 9222
rect 6449 9220 6505 9222
rect 6529 9220 6585 9222
rect 7286 12144 7342 12200
rect 6550 8372 6552 8392
rect 6552 8372 6604 8392
rect 6604 8372 6606 8392
rect 6550 8336 6606 8372
rect 6289 8186 6345 8188
rect 6369 8186 6425 8188
rect 6449 8186 6505 8188
rect 6529 8186 6585 8188
rect 6289 8134 6315 8186
rect 6315 8134 6345 8186
rect 6369 8134 6379 8186
rect 6379 8134 6425 8186
rect 6449 8134 6495 8186
rect 6495 8134 6505 8186
rect 6529 8134 6559 8186
rect 6559 8134 6585 8186
rect 6289 8132 6345 8134
rect 6369 8132 6425 8134
rect 6449 8132 6505 8134
rect 6529 8132 6585 8134
rect 6289 7098 6345 7100
rect 6369 7098 6425 7100
rect 6449 7098 6505 7100
rect 6529 7098 6585 7100
rect 6289 7046 6315 7098
rect 6315 7046 6345 7098
rect 6369 7046 6379 7098
rect 6379 7046 6425 7098
rect 6449 7046 6495 7098
rect 6495 7046 6505 7098
rect 6529 7046 6559 7098
rect 6559 7046 6585 7098
rect 6289 7044 6345 7046
rect 6369 7044 6425 7046
rect 6449 7044 6505 7046
rect 6529 7044 6585 7046
rect 5814 6024 5870 6080
rect 4526 3440 4582 3496
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5446 4528 5502 4584
rect 6289 6010 6345 6012
rect 6369 6010 6425 6012
rect 6449 6010 6505 6012
rect 6529 6010 6585 6012
rect 6289 5958 6315 6010
rect 6315 5958 6345 6010
rect 6369 5958 6379 6010
rect 6379 5958 6425 6010
rect 6449 5958 6495 6010
rect 6495 5958 6505 6010
rect 6529 5958 6559 6010
rect 6559 5958 6585 6010
rect 6289 5956 6345 5958
rect 6369 5956 6425 5958
rect 6449 5956 6505 5958
rect 6529 5956 6585 5958
rect 5354 2760 5410 2816
rect 5170 2508 5226 2544
rect 5170 2488 5172 2508
rect 5172 2488 5224 2508
rect 5224 2488 5226 2508
rect 5078 1944 5134 2000
rect 6289 4922 6345 4924
rect 6369 4922 6425 4924
rect 6449 4922 6505 4924
rect 6529 4922 6585 4924
rect 6289 4870 6315 4922
rect 6315 4870 6345 4922
rect 6369 4870 6379 4922
rect 6379 4870 6425 4922
rect 6449 4870 6495 4922
rect 6495 4870 6505 4922
rect 6529 4870 6559 4922
rect 6559 4870 6585 4922
rect 6289 4868 6345 4870
rect 6369 4868 6425 4870
rect 6449 4868 6505 4870
rect 6529 4868 6585 4870
rect 7102 5752 7158 5808
rect 6642 3984 6698 4040
rect 6289 3834 6345 3836
rect 6369 3834 6425 3836
rect 6449 3834 6505 3836
rect 6529 3834 6585 3836
rect 6289 3782 6315 3834
rect 6315 3782 6345 3834
rect 6369 3782 6379 3834
rect 6379 3782 6425 3834
rect 6449 3782 6495 3834
rect 6495 3782 6505 3834
rect 6529 3782 6559 3834
rect 6559 3782 6585 3834
rect 6289 3780 6345 3782
rect 6369 3780 6425 3782
rect 6449 3780 6505 3782
rect 6529 3780 6585 3782
rect 7378 10376 7434 10432
rect 7378 10124 7434 10160
rect 7378 10104 7380 10124
rect 7380 10104 7432 10124
rect 7432 10104 7434 10124
rect 7378 7928 7434 7984
rect 7654 13776 7710 13832
rect 7838 13912 7894 13968
rect 7838 13640 7894 13696
rect 7746 9424 7802 9480
rect 6642 3032 6698 3088
rect 6918 3032 6974 3088
rect 6289 2746 6345 2748
rect 6369 2746 6425 2748
rect 6449 2746 6505 2748
rect 6529 2746 6585 2748
rect 6289 2694 6315 2746
rect 6315 2694 6345 2746
rect 6369 2694 6379 2746
rect 6379 2694 6425 2746
rect 6449 2694 6495 2746
rect 6495 2694 6505 2746
rect 6529 2694 6559 2746
rect 6559 2694 6585 2746
rect 6289 2692 6345 2694
rect 6369 2692 6425 2694
rect 6449 2692 6505 2694
rect 6529 2692 6585 2694
rect 7102 2896 7158 2952
rect 7562 5208 7618 5264
rect 7654 3576 7710 3632
rect 7470 2760 7526 2816
rect 7470 2644 7526 2680
rect 7470 2624 7472 2644
rect 7472 2624 7524 2644
rect 7524 2624 7526 2644
rect 7838 3984 7894 4040
rect 8022 8336 8078 8392
rect 8956 29402 9012 29404
rect 9036 29402 9092 29404
rect 9116 29402 9172 29404
rect 9196 29402 9252 29404
rect 8956 29350 8982 29402
rect 8982 29350 9012 29402
rect 9036 29350 9046 29402
rect 9046 29350 9092 29402
rect 9116 29350 9162 29402
rect 9162 29350 9172 29402
rect 9196 29350 9226 29402
rect 9226 29350 9252 29402
rect 8956 29348 9012 29350
rect 9036 29348 9092 29350
rect 9116 29348 9172 29350
rect 9196 29348 9252 29350
rect 8956 28314 9012 28316
rect 9036 28314 9092 28316
rect 9116 28314 9172 28316
rect 9196 28314 9252 28316
rect 8956 28262 8982 28314
rect 8982 28262 9012 28314
rect 9036 28262 9046 28314
rect 9046 28262 9092 28314
rect 9116 28262 9162 28314
rect 9162 28262 9172 28314
rect 9196 28262 9226 28314
rect 9226 28262 9252 28314
rect 8956 28260 9012 28262
rect 9036 28260 9092 28262
rect 9116 28260 9172 28262
rect 9196 28260 9252 28262
rect 9034 27648 9090 27704
rect 8956 27226 9012 27228
rect 9036 27226 9092 27228
rect 9116 27226 9172 27228
rect 9196 27226 9252 27228
rect 8956 27174 8982 27226
rect 8982 27174 9012 27226
rect 9036 27174 9046 27226
rect 9046 27174 9092 27226
rect 9116 27174 9162 27226
rect 9162 27174 9172 27226
rect 9196 27174 9226 27226
rect 9226 27174 9252 27226
rect 8956 27172 9012 27174
rect 9036 27172 9092 27174
rect 9116 27172 9172 27174
rect 9196 27172 9252 27174
rect 8942 26988 8998 27024
rect 8942 26968 8944 26988
rect 8944 26968 8996 26988
rect 8996 26968 8998 26988
rect 8850 26424 8906 26480
rect 8956 26138 9012 26140
rect 9036 26138 9092 26140
rect 9116 26138 9172 26140
rect 9196 26138 9252 26140
rect 8956 26086 8982 26138
rect 8982 26086 9012 26138
rect 9036 26086 9046 26138
rect 9046 26086 9092 26138
rect 9116 26086 9162 26138
rect 9162 26086 9172 26138
rect 9196 26086 9226 26138
rect 9226 26086 9252 26138
rect 8956 26084 9012 26086
rect 9036 26084 9092 26086
rect 9116 26084 9172 26086
rect 9196 26084 9252 26086
rect 8956 25050 9012 25052
rect 9036 25050 9092 25052
rect 9116 25050 9172 25052
rect 9196 25050 9252 25052
rect 8956 24998 8982 25050
rect 8982 24998 9012 25050
rect 9036 24998 9046 25050
rect 9046 24998 9092 25050
rect 9116 24998 9162 25050
rect 9162 24998 9172 25050
rect 9196 24998 9226 25050
rect 9226 24998 9252 25050
rect 8956 24996 9012 24998
rect 9036 24996 9092 24998
rect 9116 24996 9172 24998
rect 9196 24996 9252 24998
rect 9402 32952 9458 33008
rect 9402 32136 9458 32192
rect 9678 34584 9734 34640
rect 9862 35708 9864 35728
rect 9864 35708 9916 35728
rect 9916 35708 9918 35728
rect 9862 35672 9918 35708
rect 9862 33360 9918 33416
rect 9862 31864 9918 31920
rect 9402 28736 9458 28792
rect 9494 27512 9550 27568
rect 9586 26152 9642 26208
rect 9586 25880 9642 25936
rect 9678 25220 9734 25256
rect 9678 25200 9680 25220
rect 9680 25200 9732 25220
rect 9732 25200 9734 25220
rect 8956 23962 9012 23964
rect 9036 23962 9092 23964
rect 9116 23962 9172 23964
rect 9196 23962 9252 23964
rect 8956 23910 8982 23962
rect 8982 23910 9012 23962
rect 9036 23910 9046 23962
rect 9046 23910 9092 23962
rect 9116 23910 9162 23962
rect 9162 23910 9172 23962
rect 9196 23910 9226 23962
rect 9226 23910 9252 23962
rect 8956 23908 9012 23910
rect 9036 23908 9092 23910
rect 9116 23908 9172 23910
rect 9196 23908 9252 23910
rect 9586 23180 9642 23216
rect 9586 23160 9588 23180
rect 9588 23160 9640 23180
rect 9640 23160 9642 23180
rect 9678 23024 9734 23080
rect 8956 22874 9012 22876
rect 9036 22874 9092 22876
rect 9116 22874 9172 22876
rect 9196 22874 9252 22876
rect 8956 22822 8982 22874
rect 8982 22822 9012 22874
rect 9036 22822 9046 22874
rect 9046 22822 9092 22874
rect 9116 22822 9162 22874
rect 9162 22822 9172 22874
rect 9196 22822 9226 22874
rect 9226 22822 9252 22874
rect 8956 22820 9012 22822
rect 9036 22820 9092 22822
rect 9116 22820 9172 22822
rect 9196 22820 9252 22822
rect 8956 21786 9012 21788
rect 9036 21786 9092 21788
rect 9116 21786 9172 21788
rect 9196 21786 9252 21788
rect 8956 21734 8982 21786
rect 8982 21734 9012 21786
rect 9036 21734 9046 21786
rect 9046 21734 9092 21786
rect 9116 21734 9162 21786
rect 9162 21734 9172 21786
rect 9196 21734 9226 21786
rect 9226 21734 9252 21786
rect 8956 21732 9012 21734
rect 9036 21732 9092 21734
rect 9116 21732 9172 21734
rect 9196 21732 9252 21734
rect 9678 21392 9734 21448
rect 8956 20698 9012 20700
rect 9036 20698 9092 20700
rect 9116 20698 9172 20700
rect 9196 20698 9252 20700
rect 8956 20646 8982 20698
rect 8982 20646 9012 20698
rect 9036 20646 9046 20698
rect 9046 20646 9092 20698
rect 9116 20646 9162 20698
rect 9162 20646 9172 20698
rect 9196 20646 9226 20698
rect 9226 20646 9252 20698
rect 8956 20644 9012 20646
rect 9036 20644 9092 20646
rect 9116 20644 9172 20646
rect 9196 20644 9252 20646
rect 9586 20576 9642 20632
rect 9586 20304 9642 20360
rect 8956 19610 9012 19612
rect 9036 19610 9092 19612
rect 9116 19610 9172 19612
rect 9196 19610 9252 19612
rect 8956 19558 8982 19610
rect 8982 19558 9012 19610
rect 9036 19558 9046 19610
rect 9046 19558 9092 19610
rect 9116 19558 9162 19610
rect 9162 19558 9172 19610
rect 9196 19558 9226 19610
rect 9226 19558 9252 19610
rect 8956 19556 9012 19558
rect 9036 19556 9092 19558
rect 9116 19556 9172 19558
rect 9196 19556 9252 19558
rect 9126 19080 9182 19136
rect 8956 18522 9012 18524
rect 9036 18522 9092 18524
rect 9116 18522 9172 18524
rect 9196 18522 9252 18524
rect 8956 18470 8982 18522
rect 8982 18470 9012 18522
rect 9036 18470 9046 18522
rect 9046 18470 9092 18522
rect 9116 18470 9162 18522
rect 9162 18470 9172 18522
rect 9196 18470 9226 18522
rect 9226 18470 9252 18522
rect 8956 18468 9012 18470
rect 9036 18468 9092 18470
rect 9116 18468 9172 18470
rect 9196 18468 9252 18470
rect 8956 17434 9012 17436
rect 9036 17434 9092 17436
rect 9116 17434 9172 17436
rect 9196 17434 9252 17436
rect 8956 17382 8982 17434
rect 8982 17382 9012 17434
rect 9036 17382 9046 17434
rect 9046 17382 9092 17434
rect 9116 17382 9162 17434
rect 9162 17382 9172 17434
rect 9196 17382 9226 17434
rect 9226 17382 9252 17434
rect 8956 17380 9012 17382
rect 9036 17380 9092 17382
rect 9116 17380 9172 17382
rect 9196 17380 9252 17382
rect 8942 17176 8998 17232
rect 8956 16346 9012 16348
rect 9036 16346 9092 16348
rect 9116 16346 9172 16348
rect 9196 16346 9252 16348
rect 8956 16294 8982 16346
rect 8982 16294 9012 16346
rect 9036 16294 9046 16346
rect 9046 16294 9092 16346
rect 9116 16294 9162 16346
rect 9162 16294 9172 16346
rect 9196 16294 9226 16346
rect 9226 16294 9252 16346
rect 8956 16292 9012 16294
rect 9036 16292 9092 16294
rect 9116 16292 9172 16294
rect 9196 16292 9252 16294
rect 8956 15258 9012 15260
rect 9036 15258 9092 15260
rect 9116 15258 9172 15260
rect 9196 15258 9252 15260
rect 8956 15206 8982 15258
rect 8982 15206 9012 15258
rect 9036 15206 9046 15258
rect 9046 15206 9092 15258
rect 9116 15206 9162 15258
rect 9162 15206 9172 15258
rect 9196 15206 9226 15258
rect 9226 15206 9252 15258
rect 8956 15204 9012 15206
rect 9036 15204 9092 15206
rect 9116 15204 9172 15206
rect 9196 15204 9252 15206
rect 9494 17312 9550 17368
rect 9954 31320 10010 31376
rect 10046 27940 10102 27976
rect 10046 27920 10048 27940
rect 10048 27920 10100 27940
rect 10100 27920 10102 27940
rect 9954 27376 10010 27432
rect 9862 26324 9864 26344
rect 9864 26324 9916 26344
rect 9916 26324 9918 26344
rect 9862 26288 9918 26324
rect 9862 26152 9918 26208
rect 10322 33532 10324 33552
rect 10324 33532 10376 33552
rect 10376 33532 10378 33552
rect 10322 33496 10378 33532
rect 10230 32272 10286 32328
rect 10322 32136 10378 32192
rect 10598 33360 10654 33416
rect 10782 33088 10838 33144
rect 10782 32816 10838 32872
rect 10506 31320 10562 31376
rect 10966 30912 11022 30968
rect 11242 29960 11298 30016
rect 10506 28056 10562 28112
rect 10138 26696 10194 26752
rect 10322 26832 10378 26888
rect 10322 24948 10378 24984
rect 10322 24928 10324 24948
rect 10324 24928 10376 24948
rect 10376 24928 10378 24948
rect 8956 14170 9012 14172
rect 9036 14170 9092 14172
rect 9116 14170 9172 14172
rect 9196 14170 9252 14172
rect 8956 14118 8982 14170
rect 8982 14118 9012 14170
rect 9036 14118 9046 14170
rect 9046 14118 9092 14170
rect 9116 14118 9162 14170
rect 9162 14118 9172 14170
rect 9196 14118 9226 14170
rect 9226 14118 9252 14170
rect 8956 14116 9012 14118
rect 9036 14116 9092 14118
rect 9116 14116 9172 14118
rect 9196 14116 9252 14118
rect 8956 13082 9012 13084
rect 9036 13082 9092 13084
rect 9116 13082 9172 13084
rect 9196 13082 9252 13084
rect 8956 13030 8982 13082
rect 8982 13030 9012 13082
rect 9036 13030 9046 13082
rect 9046 13030 9092 13082
rect 9116 13030 9162 13082
rect 9162 13030 9172 13082
rect 9196 13030 9226 13082
rect 9226 13030 9252 13082
rect 8956 13028 9012 13030
rect 9036 13028 9092 13030
rect 9116 13028 9172 13030
rect 9196 13028 9252 13030
rect 8482 9016 8538 9072
rect 8956 11994 9012 11996
rect 9036 11994 9092 11996
rect 9116 11994 9172 11996
rect 9196 11994 9252 11996
rect 8956 11942 8982 11994
rect 8982 11942 9012 11994
rect 9036 11942 9046 11994
rect 9046 11942 9092 11994
rect 9116 11942 9162 11994
rect 9162 11942 9172 11994
rect 9196 11942 9226 11994
rect 9226 11942 9252 11994
rect 8956 11940 9012 11942
rect 9036 11940 9092 11942
rect 9116 11940 9172 11942
rect 9196 11940 9252 11942
rect 8956 10906 9012 10908
rect 9036 10906 9092 10908
rect 9116 10906 9172 10908
rect 9196 10906 9252 10908
rect 8956 10854 8982 10906
rect 8982 10854 9012 10906
rect 9036 10854 9046 10906
rect 9046 10854 9092 10906
rect 9116 10854 9162 10906
rect 9162 10854 9172 10906
rect 9196 10854 9226 10906
rect 9226 10854 9252 10906
rect 8956 10852 9012 10854
rect 9036 10852 9092 10854
rect 9116 10852 9172 10854
rect 9196 10852 9252 10854
rect 8956 9818 9012 9820
rect 9036 9818 9092 9820
rect 9116 9818 9172 9820
rect 9196 9818 9252 9820
rect 8956 9766 8982 9818
rect 8982 9766 9012 9818
rect 9036 9766 9046 9818
rect 9046 9766 9092 9818
rect 9116 9766 9162 9818
rect 9162 9766 9172 9818
rect 9196 9766 9226 9818
rect 9226 9766 9252 9818
rect 8956 9764 9012 9766
rect 9036 9764 9092 9766
rect 9116 9764 9172 9766
rect 9196 9764 9252 9766
rect 8758 9016 8814 9072
rect 8206 7792 8262 7848
rect 9218 8880 9274 8936
rect 8956 8730 9012 8732
rect 9036 8730 9092 8732
rect 9116 8730 9172 8732
rect 9196 8730 9252 8732
rect 8956 8678 8982 8730
rect 8982 8678 9012 8730
rect 9036 8678 9046 8730
rect 9046 8678 9092 8730
rect 9116 8678 9162 8730
rect 9162 8678 9172 8730
rect 9196 8678 9226 8730
rect 9226 8678 9252 8730
rect 8956 8676 9012 8678
rect 9036 8676 9092 8678
rect 9116 8676 9172 8678
rect 9196 8676 9252 8678
rect 8114 4936 8170 4992
rect 8956 7642 9012 7644
rect 9036 7642 9092 7644
rect 9116 7642 9172 7644
rect 9196 7642 9252 7644
rect 8956 7590 8982 7642
rect 8982 7590 9012 7642
rect 9036 7590 9046 7642
rect 9046 7590 9092 7642
rect 9116 7590 9162 7642
rect 9162 7590 9172 7642
rect 9196 7590 9226 7642
rect 9226 7590 9252 7642
rect 8956 7588 9012 7590
rect 9036 7588 9092 7590
rect 9116 7588 9172 7590
rect 9196 7588 9252 7590
rect 8942 6840 8998 6896
rect 9678 16940 9680 16960
rect 9680 16940 9732 16960
rect 9732 16940 9734 16960
rect 9678 16904 9734 16940
rect 10230 17584 10286 17640
rect 9862 16088 9918 16144
rect 9770 14592 9826 14648
rect 10690 26968 10746 27024
rect 10598 26696 10654 26752
rect 10414 17040 10470 17096
rect 10046 16496 10102 16552
rect 10046 15952 10102 16008
rect 9586 11056 9642 11112
rect 10046 9968 10102 10024
rect 9954 9036 10010 9072
rect 9954 9016 9956 9036
rect 9956 9016 10008 9036
rect 10008 9016 10010 9036
rect 9402 6840 9458 6896
rect 8956 6554 9012 6556
rect 9036 6554 9092 6556
rect 9116 6554 9172 6556
rect 9196 6554 9252 6556
rect 8956 6502 8982 6554
rect 8982 6502 9012 6554
rect 9036 6502 9046 6554
rect 9046 6502 9092 6554
rect 9116 6502 9162 6554
rect 9162 6502 9172 6554
rect 9196 6502 9226 6554
rect 9226 6502 9252 6554
rect 8956 6500 9012 6502
rect 9036 6500 9092 6502
rect 9116 6500 9172 6502
rect 9196 6500 9252 6502
rect 9310 6160 9366 6216
rect 7930 3168 7986 3224
rect 7930 2488 7986 2544
rect 8666 3848 8722 3904
rect 8758 3304 8814 3360
rect 8956 5466 9012 5468
rect 9036 5466 9092 5468
rect 9116 5466 9172 5468
rect 9196 5466 9252 5468
rect 8956 5414 8982 5466
rect 8982 5414 9012 5466
rect 9036 5414 9046 5466
rect 9046 5414 9092 5466
rect 9116 5414 9162 5466
rect 9162 5414 9172 5466
rect 9196 5414 9226 5466
rect 9226 5414 9252 5466
rect 8956 5412 9012 5414
rect 9036 5412 9092 5414
rect 9116 5412 9172 5414
rect 9196 5412 9252 5414
rect 8956 4378 9012 4380
rect 9036 4378 9092 4380
rect 9116 4378 9172 4380
rect 9196 4378 9252 4380
rect 8956 4326 8982 4378
rect 8982 4326 9012 4378
rect 9036 4326 9046 4378
rect 9046 4326 9092 4378
rect 9116 4326 9162 4378
rect 9162 4326 9172 4378
rect 9196 4326 9226 4378
rect 9226 4326 9252 4378
rect 8956 4324 9012 4326
rect 9036 4324 9092 4326
rect 9116 4324 9172 4326
rect 9196 4324 9252 4326
rect 8956 3290 9012 3292
rect 9036 3290 9092 3292
rect 9116 3290 9172 3292
rect 9196 3290 9252 3292
rect 8956 3238 8982 3290
rect 8982 3238 9012 3290
rect 9036 3238 9046 3290
rect 9046 3238 9092 3290
rect 9116 3238 9162 3290
rect 9162 3238 9172 3290
rect 9196 3238 9226 3290
rect 9226 3238 9252 3290
rect 8956 3236 9012 3238
rect 9036 3236 9092 3238
rect 9116 3236 9172 3238
rect 9196 3236 9252 3238
rect 8956 2202 9012 2204
rect 9036 2202 9092 2204
rect 9116 2202 9172 2204
rect 9196 2202 9252 2204
rect 8956 2150 8982 2202
rect 8982 2150 9012 2202
rect 9036 2150 9046 2202
rect 9046 2150 9092 2202
rect 9116 2150 9162 2202
rect 9162 2150 9172 2202
rect 9196 2150 9226 2202
rect 9226 2150 9252 2202
rect 8956 2148 9012 2150
rect 9036 2148 9092 2150
rect 9116 2148 9172 2150
rect 9196 2148 9252 2150
rect 9678 5788 9680 5808
rect 9680 5788 9732 5808
rect 9732 5788 9734 5808
rect 9678 5752 9734 5788
rect 9494 4120 9550 4176
rect 10230 15952 10286 16008
rect 10506 16652 10562 16688
rect 10506 16632 10508 16652
rect 10508 16632 10560 16652
rect 10560 16632 10562 16652
rect 10782 21836 10784 21856
rect 10784 21836 10836 21856
rect 10836 21836 10838 21856
rect 10782 21800 10838 21836
rect 10782 19372 10838 19408
rect 10782 19352 10784 19372
rect 10784 19352 10836 19372
rect 10836 19352 10838 19372
rect 10690 19216 10746 19272
rect 10782 17584 10838 17640
rect 10690 14456 10746 14512
rect 10506 13912 10562 13968
rect 10138 8472 10194 8528
rect 10230 7792 10286 7848
rect 10414 7248 10470 7304
rect 10322 6704 10378 6760
rect 10322 5108 10324 5128
rect 10324 5108 10376 5128
rect 10376 5108 10378 5128
rect 10322 5072 10378 5108
rect 11622 37562 11678 37564
rect 11702 37562 11758 37564
rect 11782 37562 11838 37564
rect 11862 37562 11918 37564
rect 11622 37510 11648 37562
rect 11648 37510 11678 37562
rect 11702 37510 11712 37562
rect 11712 37510 11758 37562
rect 11782 37510 11828 37562
rect 11828 37510 11838 37562
rect 11862 37510 11892 37562
rect 11892 37510 11918 37562
rect 11622 37508 11678 37510
rect 11702 37508 11758 37510
rect 11782 37508 11838 37510
rect 11862 37508 11918 37510
rect 11622 36474 11678 36476
rect 11702 36474 11758 36476
rect 11782 36474 11838 36476
rect 11862 36474 11918 36476
rect 11622 36422 11648 36474
rect 11648 36422 11678 36474
rect 11702 36422 11712 36474
rect 11712 36422 11758 36474
rect 11782 36422 11828 36474
rect 11828 36422 11838 36474
rect 11862 36422 11892 36474
rect 11892 36422 11918 36474
rect 11622 36420 11678 36422
rect 11702 36420 11758 36422
rect 11782 36420 11838 36422
rect 11862 36420 11918 36422
rect 11622 35386 11678 35388
rect 11702 35386 11758 35388
rect 11782 35386 11838 35388
rect 11862 35386 11918 35388
rect 11622 35334 11648 35386
rect 11648 35334 11678 35386
rect 11702 35334 11712 35386
rect 11712 35334 11758 35386
rect 11782 35334 11828 35386
rect 11828 35334 11838 35386
rect 11862 35334 11892 35386
rect 11892 35334 11918 35386
rect 11622 35332 11678 35334
rect 11702 35332 11758 35334
rect 11782 35332 11838 35334
rect 11862 35332 11918 35334
rect 11622 34298 11678 34300
rect 11702 34298 11758 34300
rect 11782 34298 11838 34300
rect 11862 34298 11918 34300
rect 11622 34246 11648 34298
rect 11648 34246 11678 34298
rect 11702 34246 11712 34298
rect 11712 34246 11758 34298
rect 11782 34246 11828 34298
rect 11828 34246 11838 34298
rect 11862 34246 11892 34298
rect 11892 34246 11918 34298
rect 11622 34244 11678 34246
rect 11702 34244 11758 34246
rect 11782 34244 11838 34246
rect 11862 34244 11918 34246
rect 11622 33210 11678 33212
rect 11702 33210 11758 33212
rect 11782 33210 11838 33212
rect 11862 33210 11918 33212
rect 11622 33158 11648 33210
rect 11648 33158 11678 33210
rect 11702 33158 11712 33210
rect 11712 33158 11758 33210
rect 11782 33158 11828 33210
rect 11828 33158 11838 33210
rect 11862 33158 11892 33210
rect 11892 33158 11918 33210
rect 11622 33156 11678 33158
rect 11702 33156 11758 33158
rect 11782 33156 11838 33158
rect 11862 33156 11918 33158
rect 11622 32122 11678 32124
rect 11702 32122 11758 32124
rect 11782 32122 11838 32124
rect 11862 32122 11918 32124
rect 11622 32070 11648 32122
rect 11648 32070 11678 32122
rect 11702 32070 11712 32122
rect 11712 32070 11758 32122
rect 11782 32070 11828 32122
rect 11828 32070 11838 32122
rect 11862 32070 11892 32122
rect 11892 32070 11918 32122
rect 11622 32068 11678 32070
rect 11702 32068 11758 32070
rect 11782 32068 11838 32070
rect 11862 32068 11918 32070
rect 11622 31034 11678 31036
rect 11702 31034 11758 31036
rect 11782 31034 11838 31036
rect 11862 31034 11918 31036
rect 11622 30982 11648 31034
rect 11648 30982 11678 31034
rect 11702 30982 11712 31034
rect 11712 30982 11758 31034
rect 11782 30982 11828 31034
rect 11828 30982 11838 31034
rect 11862 30982 11892 31034
rect 11892 30982 11918 31034
rect 11622 30980 11678 30982
rect 11702 30980 11758 30982
rect 11782 30980 11838 30982
rect 11862 30980 11918 30982
rect 11622 29946 11678 29948
rect 11702 29946 11758 29948
rect 11782 29946 11838 29948
rect 11862 29946 11918 29948
rect 11622 29894 11648 29946
rect 11648 29894 11678 29946
rect 11702 29894 11712 29946
rect 11712 29894 11758 29946
rect 11782 29894 11828 29946
rect 11828 29894 11838 29946
rect 11862 29894 11892 29946
rect 11892 29894 11918 29946
rect 11622 29892 11678 29894
rect 11702 29892 11758 29894
rect 11782 29892 11838 29894
rect 11862 29892 11918 29894
rect 11622 28858 11678 28860
rect 11702 28858 11758 28860
rect 11782 28858 11838 28860
rect 11862 28858 11918 28860
rect 11622 28806 11648 28858
rect 11648 28806 11678 28858
rect 11702 28806 11712 28858
rect 11712 28806 11758 28858
rect 11782 28806 11828 28858
rect 11828 28806 11838 28858
rect 11862 28806 11892 28858
rect 11892 28806 11918 28858
rect 11622 28804 11678 28806
rect 11702 28804 11758 28806
rect 11782 28804 11838 28806
rect 11862 28804 11918 28806
rect 11622 27770 11678 27772
rect 11702 27770 11758 27772
rect 11782 27770 11838 27772
rect 11862 27770 11918 27772
rect 11622 27718 11648 27770
rect 11648 27718 11678 27770
rect 11702 27718 11712 27770
rect 11712 27718 11758 27770
rect 11782 27718 11828 27770
rect 11828 27718 11838 27770
rect 11862 27718 11892 27770
rect 11892 27718 11918 27770
rect 11622 27716 11678 27718
rect 11702 27716 11758 27718
rect 11782 27716 11838 27718
rect 11862 27716 11918 27718
rect 12070 27648 12126 27704
rect 12070 27512 12126 27568
rect 11622 26682 11678 26684
rect 11702 26682 11758 26684
rect 11782 26682 11838 26684
rect 11862 26682 11918 26684
rect 11622 26630 11648 26682
rect 11648 26630 11678 26682
rect 11702 26630 11712 26682
rect 11712 26630 11758 26682
rect 11782 26630 11828 26682
rect 11828 26630 11838 26682
rect 11862 26630 11892 26682
rect 11892 26630 11918 26682
rect 11622 26628 11678 26630
rect 11702 26628 11758 26630
rect 11782 26628 11838 26630
rect 11862 26628 11918 26630
rect 11622 25594 11678 25596
rect 11702 25594 11758 25596
rect 11782 25594 11838 25596
rect 11862 25594 11918 25596
rect 11622 25542 11648 25594
rect 11648 25542 11678 25594
rect 11702 25542 11712 25594
rect 11712 25542 11758 25594
rect 11782 25542 11828 25594
rect 11828 25542 11838 25594
rect 11862 25542 11892 25594
rect 11892 25542 11918 25594
rect 11622 25540 11678 25542
rect 11702 25540 11758 25542
rect 11782 25540 11838 25542
rect 11862 25540 11918 25542
rect 12070 24928 12126 24984
rect 11622 24506 11678 24508
rect 11702 24506 11758 24508
rect 11782 24506 11838 24508
rect 11862 24506 11918 24508
rect 11622 24454 11648 24506
rect 11648 24454 11678 24506
rect 11702 24454 11712 24506
rect 11712 24454 11758 24506
rect 11782 24454 11828 24506
rect 11828 24454 11838 24506
rect 11862 24454 11892 24506
rect 11892 24454 11918 24506
rect 11622 24452 11678 24454
rect 11702 24452 11758 24454
rect 11782 24452 11838 24454
rect 11862 24452 11918 24454
rect 11622 23418 11678 23420
rect 11702 23418 11758 23420
rect 11782 23418 11838 23420
rect 11862 23418 11918 23420
rect 11622 23366 11648 23418
rect 11648 23366 11678 23418
rect 11702 23366 11712 23418
rect 11712 23366 11758 23418
rect 11782 23366 11828 23418
rect 11828 23366 11838 23418
rect 11862 23366 11892 23418
rect 11892 23366 11918 23418
rect 11622 23364 11678 23366
rect 11702 23364 11758 23366
rect 11782 23364 11838 23366
rect 11862 23364 11918 23366
rect 11794 22652 11796 22672
rect 11796 22652 11848 22672
rect 11848 22652 11850 22672
rect 11794 22616 11850 22652
rect 11622 22330 11678 22332
rect 11702 22330 11758 22332
rect 11782 22330 11838 22332
rect 11862 22330 11918 22332
rect 11622 22278 11648 22330
rect 11648 22278 11678 22330
rect 11702 22278 11712 22330
rect 11712 22278 11758 22330
rect 11782 22278 11828 22330
rect 11828 22278 11838 22330
rect 11862 22278 11892 22330
rect 11892 22278 11918 22330
rect 11622 22276 11678 22278
rect 11702 22276 11758 22278
rect 11782 22276 11838 22278
rect 11862 22276 11918 22278
rect 11622 21242 11678 21244
rect 11702 21242 11758 21244
rect 11782 21242 11838 21244
rect 11862 21242 11918 21244
rect 11622 21190 11648 21242
rect 11648 21190 11678 21242
rect 11702 21190 11712 21242
rect 11712 21190 11758 21242
rect 11782 21190 11828 21242
rect 11828 21190 11838 21242
rect 11862 21190 11892 21242
rect 11892 21190 11918 21242
rect 11622 21188 11678 21190
rect 11702 21188 11758 21190
rect 11782 21188 11838 21190
rect 11862 21188 11918 21190
rect 11150 20984 11206 21040
rect 11518 20848 11574 20904
rect 11150 19760 11206 19816
rect 10782 13640 10838 13696
rect 11426 19080 11482 19136
rect 11622 20154 11678 20156
rect 11702 20154 11758 20156
rect 11782 20154 11838 20156
rect 11862 20154 11918 20156
rect 11622 20102 11648 20154
rect 11648 20102 11678 20154
rect 11702 20102 11712 20154
rect 11712 20102 11758 20154
rect 11782 20102 11828 20154
rect 11828 20102 11838 20154
rect 11862 20102 11892 20154
rect 11892 20102 11918 20154
rect 11622 20100 11678 20102
rect 11702 20100 11758 20102
rect 11782 20100 11838 20102
rect 11862 20100 11918 20102
rect 12714 33360 12770 33416
rect 12622 32816 12678 32872
rect 12990 26968 13046 27024
rect 12806 26852 12862 26888
rect 12806 26832 12808 26852
rect 12808 26832 12860 26852
rect 12860 26832 12862 26852
rect 12070 20032 12126 20088
rect 12070 19896 12126 19952
rect 11622 19066 11678 19068
rect 11702 19066 11758 19068
rect 11782 19066 11838 19068
rect 11862 19066 11918 19068
rect 11622 19014 11648 19066
rect 11648 19014 11678 19066
rect 11702 19014 11712 19066
rect 11712 19014 11758 19066
rect 11782 19014 11828 19066
rect 11828 19014 11838 19066
rect 11862 19014 11892 19066
rect 11892 19014 11918 19066
rect 11622 19012 11678 19014
rect 11702 19012 11758 19014
rect 11782 19012 11838 19014
rect 11862 19012 11918 19014
rect 11622 17978 11678 17980
rect 11702 17978 11758 17980
rect 11782 17978 11838 17980
rect 11862 17978 11918 17980
rect 11622 17926 11648 17978
rect 11648 17926 11678 17978
rect 11702 17926 11712 17978
rect 11712 17926 11758 17978
rect 11782 17926 11828 17978
rect 11828 17926 11838 17978
rect 11862 17926 11892 17978
rect 11892 17926 11918 17978
rect 11622 17924 11678 17926
rect 11702 17924 11758 17926
rect 11782 17924 11838 17926
rect 11862 17924 11918 17926
rect 11622 16890 11678 16892
rect 11702 16890 11758 16892
rect 11782 16890 11838 16892
rect 11862 16890 11918 16892
rect 11622 16838 11648 16890
rect 11648 16838 11678 16890
rect 11702 16838 11712 16890
rect 11712 16838 11758 16890
rect 11782 16838 11828 16890
rect 11828 16838 11838 16890
rect 11862 16838 11892 16890
rect 11892 16838 11918 16890
rect 11622 16836 11678 16838
rect 11702 16836 11758 16838
rect 11782 16836 11838 16838
rect 11862 16836 11918 16838
rect 11622 15802 11678 15804
rect 11702 15802 11758 15804
rect 11782 15802 11838 15804
rect 11862 15802 11918 15804
rect 11622 15750 11648 15802
rect 11648 15750 11678 15802
rect 11702 15750 11712 15802
rect 11712 15750 11758 15802
rect 11782 15750 11828 15802
rect 11828 15750 11838 15802
rect 11862 15750 11892 15802
rect 11892 15750 11918 15802
rect 11622 15748 11678 15750
rect 11702 15748 11758 15750
rect 11782 15748 11838 15750
rect 11862 15748 11918 15750
rect 11518 15000 11574 15056
rect 11242 10376 11298 10432
rect 10046 3984 10102 4040
rect 9954 3712 10010 3768
rect 9862 3576 9918 3632
rect 9862 3032 9918 3088
rect 10414 3848 10470 3904
rect 10782 9424 10838 9480
rect 11150 8880 11206 8936
rect 10874 8780 10876 8800
rect 10876 8780 10928 8800
rect 10928 8780 10930 8800
rect 10874 8744 10930 8780
rect 10782 8336 10838 8392
rect 11150 4936 11206 4992
rect 10690 4664 10746 4720
rect 10782 3188 10838 3224
rect 10782 3168 10784 3188
rect 10784 3168 10836 3188
rect 10836 3168 10838 3188
rect 11426 3440 11482 3496
rect 11334 2760 11390 2816
rect 11622 14714 11678 14716
rect 11702 14714 11758 14716
rect 11782 14714 11838 14716
rect 11862 14714 11918 14716
rect 11622 14662 11648 14714
rect 11648 14662 11678 14714
rect 11702 14662 11712 14714
rect 11712 14662 11758 14714
rect 11782 14662 11828 14714
rect 11828 14662 11838 14714
rect 11862 14662 11892 14714
rect 11892 14662 11918 14714
rect 11622 14660 11678 14662
rect 11702 14660 11758 14662
rect 11782 14660 11838 14662
rect 11862 14660 11918 14662
rect 11978 13776 12034 13832
rect 11622 13626 11678 13628
rect 11702 13626 11758 13628
rect 11782 13626 11838 13628
rect 11862 13626 11918 13628
rect 11622 13574 11648 13626
rect 11648 13574 11678 13626
rect 11702 13574 11712 13626
rect 11712 13574 11758 13626
rect 11782 13574 11828 13626
rect 11828 13574 11838 13626
rect 11862 13574 11892 13626
rect 11892 13574 11918 13626
rect 11622 13572 11678 13574
rect 11702 13572 11758 13574
rect 11782 13572 11838 13574
rect 11862 13572 11918 13574
rect 11622 12538 11678 12540
rect 11702 12538 11758 12540
rect 11782 12538 11838 12540
rect 11862 12538 11918 12540
rect 11622 12486 11648 12538
rect 11648 12486 11678 12538
rect 11702 12486 11712 12538
rect 11712 12486 11758 12538
rect 11782 12486 11828 12538
rect 11828 12486 11838 12538
rect 11862 12486 11892 12538
rect 11892 12486 11918 12538
rect 11622 12484 11678 12486
rect 11702 12484 11758 12486
rect 11782 12484 11838 12486
rect 11862 12484 11918 12486
rect 11622 11450 11678 11452
rect 11702 11450 11758 11452
rect 11782 11450 11838 11452
rect 11862 11450 11918 11452
rect 11622 11398 11648 11450
rect 11648 11398 11678 11450
rect 11702 11398 11712 11450
rect 11712 11398 11758 11450
rect 11782 11398 11828 11450
rect 11828 11398 11838 11450
rect 11862 11398 11892 11450
rect 11892 11398 11918 11450
rect 11622 11396 11678 11398
rect 11702 11396 11758 11398
rect 11782 11396 11838 11398
rect 11862 11396 11918 11398
rect 12070 11056 12126 11112
rect 11622 10362 11678 10364
rect 11702 10362 11758 10364
rect 11782 10362 11838 10364
rect 11862 10362 11918 10364
rect 11622 10310 11648 10362
rect 11648 10310 11678 10362
rect 11702 10310 11712 10362
rect 11712 10310 11758 10362
rect 11782 10310 11828 10362
rect 11828 10310 11838 10362
rect 11862 10310 11892 10362
rect 11892 10310 11918 10362
rect 11622 10308 11678 10310
rect 11702 10308 11758 10310
rect 11782 10308 11838 10310
rect 11862 10308 11918 10310
rect 11622 9274 11678 9276
rect 11702 9274 11758 9276
rect 11782 9274 11838 9276
rect 11862 9274 11918 9276
rect 11622 9222 11648 9274
rect 11648 9222 11678 9274
rect 11702 9222 11712 9274
rect 11712 9222 11758 9274
rect 11782 9222 11828 9274
rect 11828 9222 11838 9274
rect 11862 9222 11892 9274
rect 11892 9222 11918 9274
rect 11622 9220 11678 9222
rect 11702 9220 11758 9222
rect 11782 9220 11838 9222
rect 11862 9220 11918 9222
rect 11622 8186 11678 8188
rect 11702 8186 11758 8188
rect 11782 8186 11838 8188
rect 11862 8186 11918 8188
rect 11622 8134 11648 8186
rect 11648 8134 11678 8186
rect 11702 8134 11712 8186
rect 11712 8134 11758 8186
rect 11782 8134 11828 8186
rect 11828 8134 11838 8186
rect 11862 8134 11892 8186
rect 11892 8134 11918 8186
rect 11622 8132 11678 8134
rect 11702 8132 11758 8134
rect 11782 8132 11838 8134
rect 11862 8132 11918 8134
rect 11622 7098 11678 7100
rect 11702 7098 11758 7100
rect 11782 7098 11838 7100
rect 11862 7098 11918 7100
rect 11622 7046 11648 7098
rect 11648 7046 11678 7098
rect 11702 7046 11712 7098
rect 11712 7046 11758 7098
rect 11782 7046 11828 7098
rect 11828 7046 11838 7098
rect 11862 7046 11892 7098
rect 11892 7046 11918 7098
rect 11622 7044 11678 7046
rect 11702 7044 11758 7046
rect 11782 7044 11838 7046
rect 11862 7044 11918 7046
rect 11622 6010 11678 6012
rect 11702 6010 11758 6012
rect 11782 6010 11838 6012
rect 11862 6010 11918 6012
rect 11622 5958 11648 6010
rect 11648 5958 11678 6010
rect 11702 5958 11712 6010
rect 11712 5958 11758 6010
rect 11782 5958 11828 6010
rect 11828 5958 11838 6010
rect 11862 5958 11892 6010
rect 11892 5958 11918 6010
rect 11622 5956 11678 5958
rect 11702 5956 11758 5958
rect 11782 5956 11838 5958
rect 11862 5956 11918 5958
rect 11622 4922 11678 4924
rect 11702 4922 11758 4924
rect 11782 4922 11838 4924
rect 11862 4922 11918 4924
rect 11622 4870 11648 4922
rect 11648 4870 11678 4922
rect 11702 4870 11712 4922
rect 11712 4870 11758 4922
rect 11782 4870 11828 4922
rect 11828 4870 11838 4922
rect 11862 4870 11892 4922
rect 11892 4870 11918 4922
rect 11622 4868 11678 4870
rect 11702 4868 11758 4870
rect 11782 4868 11838 4870
rect 11862 4868 11918 4870
rect 11622 3834 11678 3836
rect 11702 3834 11758 3836
rect 11782 3834 11838 3836
rect 11862 3834 11918 3836
rect 11622 3782 11648 3834
rect 11648 3782 11678 3834
rect 11702 3782 11712 3834
rect 11712 3782 11758 3834
rect 11782 3782 11828 3834
rect 11828 3782 11838 3834
rect 11862 3782 11892 3834
rect 11892 3782 11918 3834
rect 11622 3780 11678 3782
rect 11702 3780 11758 3782
rect 11782 3780 11838 3782
rect 11862 3780 11918 3782
rect 12162 6704 12218 6760
rect 12162 4120 12218 4176
rect 13174 34584 13230 34640
rect 13634 34584 13690 34640
rect 13542 33360 13598 33416
rect 12438 21800 12494 21856
rect 12622 20576 12678 20632
rect 12990 16632 13046 16688
rect 12898 7928 12954 7984
rect 13266 24928 13322 24984
rect 13726 31320 13782 31376
rect 14289 37018 14345 37020
rect 14369 37018 14425 37020
rect 14449 37018 14505 37020
rect 14529 37018 14585 37020
rect 14289 36966 14315 37018
rect 14315 36966 14345 37018
rect 14369 36966 14379 37018
rect 14379 36966 14425 37018
rect 14449 36966 14495 37018
rect 14495 36966 14505 37018
rect 14529 36966 14559 37018
rect 14559 36966 14585 37018
rect 14289 36964 14345 36966
rect 14369 36964 14425 36966
rect 14449 36964 14505 36966
rect 14529 36964 14585 36966
rect 14289 35930 14345 35932
rect 14369 35930 14425 35932
rect 14449 35930 14505 35932
rect 14529 35930 14585 35932
rect 14289 35878 14315 35930
rect 14315 35878 14345 35930
rect 14369 35878 14379 35930
rect 14379 35878 14425 35930
rect 14449 35878 14495 35930
rect 14495 35878 14505 35930
rect 14529 35878 14559 35930
rect 14559 35878 14585 35930
rect 14289 35876 14345 35878
rect 14369 35876 14425 35878
rect 14449 35876 14505 35878
rect 14529 35876 14585 35878
rect 14289 34842 14345 34844
rect 14369 34842 14425 34844
rect 14449 34842 14505 34844
rect 14529 34842 14585 34844
rect 14289 34790 14315 34842
rect 14315 34790 14345 34842
rect 14369 34790 14379 34842
rect 14379 34790 14425 34842
rect 14449 34790 14495 34842
rect 14495 34790 14505 34842
rect 14529 34790 14559 34842
rect 14559 34790 14585 34842
rect 14289 34788 14345 34790
rect 14369 34788 14425 34790
rect 14449 34788 14505 34790
rect 14529 34788 14585 34790
rect 14289 33754 14345 33756
rect 14369 33754 14425 33756
rect 14449 33754 14505 33756
rect 14529 33754 14585 33756
rect 14289 33702 14315 33754
rect 14315 33702 14345 33754
rect 14369 33702 14379 33754
rect 14379 33702 14425 33754
rect 14449 33702 14495 33754
rect 14495 33702 14505 33754
rect 14529 33702 14559 33754
rect 14559 33702 14585 33754
rect 14289 33700 14345 33702
rect 14369 33700 14425 33702
rect 14449 33700 14505 33702
rect 14529 33700 14585 33702
rect 14289 32666 14345 32668
rect 14369 32666 14425 32668
rect 14449 32666 14505 32668
rect 14529 32666 14585 32668
rect 14289 32614 14315 32666
rect 14315 32614 14345 32666
rect 14369 32614 14379 32666
rect 14379 32614 14425 32666
rect 14449 32614 14495 32666
rect 14495 32614 14505 32666
rect 14529 32614 14559 32666
rect 14559 32614 14585 32666
rect 14289 32612 14345 32614
rect 14369 32612 14425 32614
rect 14449 32612 14505 32614
rect 14529 32612 14585 32614
rect 14289 31578 14345 31580
rect 14369 31578 14425 31580
rect 14449 31578 14505 31580
rect 14529 31578 14585 31580
rect 14289 31526 14315 31578
rect 14315 31526 14345 31578
rect 14369 31526 14379 31578
rect 14379 31526 14425 31578
rect 14449 31526 14495 31578
rect 14495 31526 14505 31578
rect 14529 31526 14559 31578
rect 14559 31526 14585 31578
rect 14289 31524 14345 31526
rect 14369 31524 14425 31526
rect 14449 31524 14505 31526
rect 14529 31524 14585 31526
rect 14289 30490 14345 30492
rect 14369 30490 14425 30492
rect 14449 30490 14505 30492
rect 14529 30490 14585 30492
rect 14289 30438 14315 30490
rect 14315 30438 14345 30490
rect 14369 30438 14379 30490
rect 14379 30438 14425 30490
rect 14449 30438 14495 30490
rect 14495 30438 14505 30490
rect 14529 30438 14559 30490
rect 14559 30438 14585 30490
rect 14289 30436 14345 30438
rect 14369 30436 14425 30438
rect 14449 30436 14505 30438
rect 14529 30436 14585 30438
rect 14646 29688 14702 29744
rect 14289 29402 14345 29404
rect 14369 29402 14425 29404
rect 14449 29402 14505 29404
rect 14529 29402 14585 29404
rect 14289 29350 14315 29402
rect 14315 29350 14345 29402
rect 14369 29350 14379 29402
rect 14379 29350 14425 29402
rect 14449 29350 14495 29402
rect 14495 29350 14505 29402
rect 14529 29350 14559 29402
rect 14559 29350 14585 29402
rect 14289 29348 14345 29350
rect 14369 29348 14425 29350
rect 14449 29348 14505 29350
rect 14529 29348 14585 29350
rect 14289 28314 14345 28316
rect 14369 28314 14425 28316
rect 14449 28314 14505 28316
rect 14529 28314 14585 28316
rect 14289 28262 14315 28314
rect 14315 28262 14345 28314
rect 14369 28262 14379 28314
rect 14379 28262 14425 28314
rect 14449 28262 14495 28314
rect 14495 28262 14505 28314
rect 14529 28262 14559 28314
rect 14559 28262 14585 28314
rect 14289 28260 14345 28262
rect 14369 28260 14425 28262
rect 14449 28260 14505 28262
rect 14529 28260 14585 28262
rect 15750 34584 15806 34640
rect 15382 32272 15438 32328
rect 15014 27512 15070 27568
rect 14289 27226 14345 27228
rect 14369 27226 14425 27228
rect 14449 27226 14505 27228
rect 14529 27226 14585 27228
rect 14289 27174 14315 27226
rect 14315 27174 14345 27226
rect 14369 27174 14379 27226
rect 14379 27174 14425 27226
rect 14449 27174 14495 27226
rect 14495 27174 14505 27226
rect 14529 27174 14559 27226
rect 14559 27174 14585 27226
rect 14289 27172 14345 27174
rect 14369 27172 14425 27174
rect 14449 27172 14505 27174
rect 14529 27172 14585 27174
rect 14289 26138 14345 26140
rect 14369 26138 14425 26140
rect 14449 26138 14505 26140
rect 14529 26138 14585 26140
rect 14289 26086 14315 26138
rect 14315 26086 14345 26138
rect 14369 26086 14379 26138
rect 14379 26086 14425 26138
rect 14449 26086 14495 26138
rect 14495 26086 14505 26138
rect 14529 26086 14559 26138
rect 14559 26086 14585 26138
rect 14289 26084 14345 26086
rect 14369 26084 14425 26086
rect 14449 26084 14505 26086
rect 14529 26084 14585 26086
rect 14289 25050 14345 25052
rect 14369 25050 14425 25052
rect 14449 25050 14505 25052
rect 14529 25050 14585 25052
rect 14289 24998 14315 25050
rect 14315 24998 14345 25050
rect 14369 24998 14379 25050
rect 14379 24998 14425 25050
rect 14449 24998 14495 25050
rect 14495 24998 14505 25050
rect 14529 24998 14559 25050
rect 14559 24998 14585 25050
rect 14289 24996 14345 24998
rect 14369 24996 14425 24998
rect 14449 24996 14505 24998
rect 14529 24996 14585 24998
rect 14094 24792 14150 24848
rect 14289 23962 14345 23964
rect 14369 23962 14425 23964
rect 14449 23962 14505 23964
rect 14529 23962 14585 23964
rect 14289 23910 14315 23962
rect 14315 23910 14345 23962
rect 14369 23910 14379 23962
rect 14379 23910 14425 23962
rect 14449 23910 14495 23962
rect 14495 23910 14505 23962
rect 14529 23910 14559 23962
rect 14559 23910 14585 23962
rect 14289 23908 14345 23910
rect 14369 23908 14425 23910
rect 14449 23908 14505 23910
rect 14529 23908 14585 23910
rect 14289 22874 14345 22876
rect 14369 22874 14425 22876
rect 14449 22874 14505 22876
rect 14529 22874 14585 22876
rect 14289 22822 14315 22874
rect 14315 22822 14345 22874
rect 14369 22822 14379 22874
rect 14379 22822 14425 22874
rect 14449 22822 14495 22874
rect 14495 22822 14505 22874
rect 14529 22822 14559 22874
rect 14559 22822 14585 22874
rect 14289 22820 14345 22822
rect 14369 22820 14425 22822
rect 14449 22820 14505 22822
rect 14529 22820 14585 22822
rect 14289 21786 14345 21788
rect 14369 21786 14425 21788
rect 14449 21786 14505 21788
rect 14529 21786 14585 21788
rect 14289 21734 14315 21786
rect 14315 21734 14345 21786
rect 14369 21734 14379 21786
rect 14379 21734 14425 21786
rect 14449 21734 14495 21786
rect 14495 21734 14505 21786
rect 14529 21734 14559 21786
rect 14559 21734 14585 21786
rect 14289 21732 14345 21734
rect 14369 21732 14425 21734
rect 14449 21732 14505 21734
rect 14529 21732 14585 21734
rect 14289 20698 14345 20700
rect 14369 20698 14425 20700
rect 14449 20698 14505 20700
rect 14529 20698 14585 20700
rect 14289 20646 14315 20698
rect 14315 20646 14345 20698
rect 14369 20646 14379 20698
rect 14379 20646 14425 20698
rect 14449 20646 14495 20698
rect 14495 20646 14505 20698
rect 14529 20646 14559 20698
rect 14559 20646 14585 20698
rect 14289 20644 14345 20646
rect 14369 20644 14425 20646
rect 14449 20644 14505 20646
rect 14529 20644 14585 20646
rect 14289 19610 14345 19612
rect 14369 19610 14425 19612
rect 14449 19610 14505 19612
rect 14529 19610 14585 19612
rect 14289 19558 14315 19610
rect 14315 19558 14345 19610
rect 14369 19558 14379 19610
rect 14379 19558 14425 19610
rect 14449 19558 14495 19610
rect 14495 19558 14505 19610
rect 14529 19558 14559 19610
rect 14559 19558 14585 19610
rect 14289 19556 14345 19558
rect 14369 19556 14425 19558
rect 14449 19556 14505 19558
rect 14529 19556 14585 19558
rect 14289 18522 14345 18524
rect 14369 18522 14425 18524
rect 14449 18522 14505 18524
rect 14529 18522 14585 18524
rect 14289 18470 14315 18522
rect 14315 18470 14345 18522
rect 14369 18470 14379 18522
rect 14379 18470 14425 18522
rect 14449 18470 14495 18522
rect 14495 18470 14505 18522
rect 14529 18470 14559 18522
rect 14559 18470 14585 18522
rect 14289 18468 14345 18470
rect 14369 18468 14425 18470
rect 14449 18468 14505 18470
rect 14529 18468 14585 18470
rect 14289 17434 14345 17436
rect 14369 17434 14425 17436
rect 14449 17434 14505 17436
rect 14529 17434 14585 17436
rect 14289 17382 14315 17434
rect 14315 17382 14345 17434
rect 14369 17382 14379 17434
rect 14379 17382 14425 17434
rect 14449 17382 14495 17434
rect 14495 17382 14505 17434
rect 14529 17382 14559 17434
rect 14559 17382 14585 17434
rect 14289 17380 14345 17382
rect 14369 17380 14425 17382
rect 14449 17380 14505 17382
rect 14529 17380 14585 17382
rect 14289 16346 14345 16348
rect 14369 16346 14425 16348
rect 14449 16346 14505 16348
rect 14529 16346 14585 16348
rect 14289 16294 14315 16346
rect 14315 16294 14345 16346
rect 14369 16294 14379 16346
rect 14379 16294 14425 16346
rect 14449 16294 14495 16346
rect 14495 16294 14505 16346
rect 14529 16294 14559 16346
rect 14559 16294 14585 16346
rect 14289 16292 14345 16294
rect 14369 16292 14425 16294
rect 14449 16292 14505 16294
rect 14529 16292 14585 16294
rect 14289 15258 14345 15260
rect 14369 15258 14425 15260
rect 14449 15258 14505 15260
rect 14529 15258 14585 15260
rect 14289 15206 14315 15258
rect 14315 15206 14345 15258
rect 14369 15206 14379 15258
rect 14379 15206 14425 15258
rect 14449 15206 14495 15258
rect 14495 15206 14505 15258
rect 14529 15206 14559 15258
rect 14559 15206 14585 15258
rect 14289 15204 14345 15206
rect 14369 15204 14425 15206
rect 14449 15204 14505 15206
rect 14529 15204 14585 15206
rect 13726 12144 13782 12200
rect 13450 10124 13506 10160
rect 13450 10104 13452 10124
rect 13452 10104 13504 10124
rect 13504 10104 13506 10124
rect 13266 9424 13322 9480
rect 13082 8780 13084 8800
rect 13084 8780 13136 8800
rect 13136 8780 13138 8800
rect 13082 8744 13138 8780
rect 13174 8356 13230 8392
rect 13174 8336 13176 8356
rect 13176 8336 13228 8356
rect 13228 8336 13230 8356
rect 12530 3984 12586 4040
rect 12438 3168 12494 3224
rect 11622 2746 11678 2748
rect 11702 2746 11758 2748
rect 11782 2746 11838 2748
rect 11862 2746 11918 2748
rect 11622 2694 11648 2746
rect 11648 2694 11678 2746
rect 11702 2694 11712 2746
rect 11712 2694 11758 2746
rect 11782 2694 11828 2746
rect 11828 2694 11838 2746
rect 11862 2694 11892 2746
rect 11892 2694 11918 2746
rect 11622 2692 11678 2694
rect 11702 2692 11758 2694
rect 11782 2692 11838 2694
rect 11862 2692 11918 2694
rect 12898 2488 12954 2544
rect 14289 14170 14345 14172
rect 14369 14170 14425 14172
rect 14449 14170 14505 14172
rect 14529 14170 14585 14172
rect 14289 14118 14315 14170
rect 14315 14118 14345 14170
rect 14369 14118 14379 14170
rect 14379 14118 14425 14170
rect 14449 14118 14495 14170
rect 14495 14118 14505 14170
rect 14529 14118 14559 14170
rect 14559 14118 14585 14170
rect 14289 14116 14345 14118
rect 14369 14116 14425 14118
rect 14449 14116 14505 14118
rect 14529 14116 14585 14118
rect 14289 13082 14345 13084
rect 14369 13082 14425 13084
rect 14449 13082 14505 13084
rect 14529 13082 14585 13084
rect 14289 13030 14315 13082
rect 14315 13030 14345 13082
rect 14369 13030 14379 13082
rect 14379 13030 14425 13082
rect 14449 13030 14495 13082
rect 14495 13030 14505 13082
rect 14529 13030 14559 13082
rect 14559 13030 14585 13082
rect 14289 13028 14345 13030
rect 14369 13028 14425 13030
rect 14449 13028 14505 13030
rect 14529 13028 14585 13030
rect 14289 11994 14345 11996
rect 14369 11994 14425 11996
rect 14449 11994 14505 11996
rect 14529 11994 14585 11996
rect 14289 11942 14315 11994
rect 14315 11942 14345 11994
rect 14369 11942 14379 11994
rect 14379 11942 14425 11994
rect 14449 11942 14495 11994
rect 14495 11942 14505 11994
rect 14529 11942 14559 11994
rect 14559 11942 14585 11994
rect 14289 11940 14345 11942
rect 14369 11940 14425 11942
rect 14449 11940 14505 11942
rect 14529 11940 14585 11942
rect 14289 10906 14345 10908
rect 14369 10906 14425 10908
rect 14449 10906 14505 10908
rect 14529 10906 14585 10908
rect 14289 10854 14315 10906
rect 14315 10854 14345 10906
rect 14369 10854 14379 10906
rect 14379 10854 14425 10906
rect 14449 10854 14495 10906
rect 14495 10854 14505 10906
rect 14529 10854 14559 10906
rect 14559 10854 14585 10906
rect 14289 10852 14345 10854
rect 14369 10852 14425 10854
rect 14449 10852 14505 10854
rect 14529 10852 14585 10854
rect 14289 9818 14345 9820
rect 14369 9818 14425 9820
rect 14449 9818 14505 9820
rect 14529 9818 14585 9820
rect 14289 9766 14315 9818
rect 14315 9766 14345 9818
rect 14369 9766 14379 9818
rect 14379 9766 14425 9818
rect 14449 9766 14495 9818
rect 14495 9766 14505 9818
rect 14529 9766 14559 9818
rect 14559 9766 14585 9818
rect 14289 9764 14345 9766
rect 14369 9764 14425 9766
rect 14449 9764 14505 9766
rect 14529 9764 14585 9766
rect 14289 8730 14345 8732
rect 14369 8730 14425 8732
rect 14449 8730 14505 8732
rect 14529 8730 14585 8732
rect 14289 8678 14315 8730
rect 14315 8678 14345 8730
rect 14369 8678 14379 8730
rect 14379 8678 14425 8730
rect 14449 8678 14495 8730
rect 14495 8678 14505 8730
rect 14529 8678 14559 8730
rect 14559 8678 14585 8730
rect 14289 8676 14345 8678
rect 14369 8676 14425 8678
rect 14449 8676 14505 8678
rect 14529 8676 14585 8678
rect 14646 8336 14702 8392
rect 14289 7642 14345 7644
rect 14369 7642 14425 7644
rect 14449 7642 14505 7644
rect 14529 7642 14585 7644
rect 14289 7590 14315 7642
rect 14315 7590 14345 7642
rect 14369 7590 14379 7642
rect 14379 7590 14425 7642
rect 14449 7590 14495 7642
rect 14495 7590 14505 7642
rect 14529 7590 14559 7642
rect 14559 7590 14585 7642
rect 14289 7588 14345 7590
rect 14369 7588 14425 7590
rect 14449 7588 14505 7590
rect 14529 7588 14585 7590
rect 14289 6554 14345 6556
rect 14369 6554 14425 6556
rect 14449 6554 14505 6556
rect 14529 6554 14585 6556
rect 14289 6502 14315 6554
rect 14315 6502 14345 6554
rect 14369 6502 14379 6554
rect 14379 6502 14425 6554
rect 14449 6502 14495 6554
rect 14495 6502 14505 6554
rect 14529 6502 14559 6554
rect 14559 6502 14585 6554
rect 14289 6500 14345 6502
rect 14369 6500 14425 6502
rect 14449 6500 14505 6502
rect 14529 6500 14585 6502
rect 14289 5466 14345 5468
rect 14369 5466 14425 5468
rect 14449 5466 14505 5468
rect 14529 5466 14585 5468
rect 14289 5414 14315 5466
rect 14315 5414 14345 5466
rect 14369 5414 14379 5466
rect 14379 5414 14425 5466
rect 14449 5414 14495 5466
rect 14495 5414 14505 5466
rect 14529 5414 14559 5466
rect 14559 5414 14585 5466
rect 14289 5412 14345 5414
rect 14369 5412 14425 5414
rect 14449 5412 14505 5414
rect 14529 5412 14585 5414
rect 14289 4378 14345 4380
rect 14369 4378 14425 4380
rect 14449 4378 14505 4380
rect 14529 4378 14585 4380
rect 14289 4326 14315 4378
rect 14315 4326 14345 4378
rect 14369 4326 14379 4378
rect 14379 4326 14425 4378
rect 14449 4326 14495 4378
rect 14495 4326 14505 4378
rect 14529 4326 14559 4378
rect 14559 4326 14585 4378
rect 14289 4324 14345 4326
rect 14369 4324 14425 4326
rect 14449 4324 14505 4326
rect 14529 4324 14585 4326
rect 14289 3290 14345 3292
rect 14369 3290 14425 3292
rect 14449 3290 14505 3292
rect 14529 3290 14585 3292
rect 14289 3238 14315 3290
rect 14315 3238 14345 3290
rect 14369 3238 14379 3290
rect 14379 3238 14425 3290
rect 14449 3238 14495 3290
rect 14495 3238 14505 3290
rect 14529 3238 14559 3290
rect 14559 3238 14585 3290
rect 14289 3236 14345 3238
rect 14369 3236 14425 3238
rect 14449 3236 14505 3238
rect 14529 3236 14585 3238
rect 14289 2202 14345 2204
rect 14369 2202 14425 2204
rect 14449 2202 14505 2204
rect 14529 2202 14585 2204
rect 14289 2150 14315 2202
rect 14315 2150 14345 2202
rect 14369 2150 14379 2202
rect 14379 2150 14425 2202
rect 14449 2150 14495 2202
rect 14495 2150 14505 2202
rect 14529 2150 14559 2202
rect 14559 2150 14585 2202
rect 14289 2148 14345 2150
rect 14369 2148 14425 2150
rect 14449 2148 14505 2150
rect 14529 2148 14585 2150
rect 14186 1944 14242 2000
rect 15382 6840 15438 6896
<< metal3 >>
rect 0 38722 480 38752
rect 2681 38722 2747 38725
rect 0 38720 2747 38722
rect 0 38664 2686 38720
rect 2742 38664 2747 38720
rect 0 38662 2747 38664
rect 0 38632 480 38662
rect 2681 38659 2747 38662
rect 6277 37568 6597 37569
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 37503 6597 37504
rect 11610 37568 11930 37569
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 37503 11930 37504
rect 3610 37024 3930 37025
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3930 37024
rect 3610 36959 3930 36960
rect 8944 37024 9264 37025
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 36959 9264 36960
rect 14277 37024 14597 37025
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 36959 14597 36960
rect 6277 36480 6597 36481
rect 0 36410 480 36440
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 36415 6597 36416
rect 11610 36480 11930 36481
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 36415 11930 36416
rect 1485 36410 1551 36413
rect 0 36408 1551 36410
rect 0 36352 1490 36408
rect 1546 36352 1551 36408
rect 0 36350 1551 36352
rect 0 36320 480 36350
rect 1485 36347 1551 36350
rect 3610 35936 3930 35937
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3930 35936
rect 3610 35871 3930 35872
rect 8944 35936 9264 35937
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 35871 9264 35872
rect 14277 35936 14597 35937
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 35871 14597 35872
rect 565 35866 631 35869
rect 3417 35866 3483 35869
rect 565 35864 3483 35866
rect 565 35808 570 35864
rect 626 35808 3422 35864
rect 3478 35808 3483 35864
rect 565 35806 3483 35808
rect 565 35803 631 35806
rect 3417 35803 3483 35806
rect 4521 35730 4587 35733
rect 9857 35730 9923 35733
rect 4521 35728 9923 35730
rect 4521 35672 4526 35728
rect 4582 35672 9862 35728
rect 9918 35672 9923 35728
rect 4521 35670 9923 35672
rect 4521 35667 4587 35670
rect 9857 35667 9923 35670
rect 6277 35392 6597 35393
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 35327 6597 35328
rect 11610 35392 11930 35393
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 35327 11930 35328
rect 2589 35322 2655 35325
rect 5073 35322 5139 35325
rect 2589 35320 5139 35322
rect 2589 35264 2594 35320
rect 2650 35264 5078 35320
rect 5134 35264 5139 35320
rect 2589 35262 5139 35264
rect 2589 35259 2655 35262
rect 5073 35259 5139 35262
rect 1761 35186 1827 35189
rect 7557 35186 7623 35189
rect 1761 35184 7623 35186
rect 1761 35128 1766 35184
rect 1822 35128 7562 35184
rect 7618 35128 7623 35184
rect 1761 35126 7623 35128
rect 1761 35123 1827 35126
rect 7557 35123 7623 35126
rect 3610 34848 3930 34849
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3930 34848
rect 3610 34783 3930 34784
rect 8944 34848 9264 34849
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 34783 9264 34784
rect 14277 34848 14597 34849
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 34783 14597 34784
rect 7741 34642 7807 34645
rect 9673 34642 9739 34645
rect 7741 34640 9739 34642
rect 7741 34584 7746 34640
rect 7802 34584 9678 34640
rect 9734 34584 9739 34640
rect 7741 34582 9739 34584
rect 7741 34579 7807 34582
rect 9673 34579 9739 34582
rect 13169 34642 13235 34645
rect 13629 34642 13695 34645
rect 15745 34642 15811 34645
rect 13169 34640 15811 34642
rect 13169 34584 13174 34640
rect 13230 34584 13634 34640
rect 13690 34584 15750 34640
rect 15806 34584 15811 34640
rect 13169 34582 15811 34584
rect 13169 34579 13235 34582
rect 13629 34579 13695 34582
rect 15745 34579 15811 34582
rect 6277 34304 6597 34305
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 34239 6597 34240
rect 11610 34304 11930 34305
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 34239 11930 34240
rect 0 34098 480 34128
rect 1577 34098 1643 34101
rect 0 34096 1643 34098
rect 0 34040 1582 34096
rect 1638 34040 1643 34096
rect 0 34038 1643 34040
rect 0 34008 480 34038
rect 1577 34035 1643 34038
rect 3610 33760 3930 33761
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3930 33760
rect 3610 33695 3930 33696
rect 8944 33760 9264 33761
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 33695 9264 33696
rect 14277 33760 14597 33761
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 33695 14597 33696
rect 4061 33690 4127 33693
rect 6637 33690 6703 33693
rect 4061 33688 7850 33690
rect 4061 33632 4066 33688
rect 4122 33632 6642 33688
rect 6698 33632 7850 33688
rect 4061 33630 7850 33632
rect 4061 33627 4127 33630
rect 6637 33627 6703 33630
rect 1393 33554 1459 33557
rect 7557 33554 7623 33557
rect 1393 33552 7623 33554
rect 1393 33496 1398 33552
rect 1454 33496 7562 33552
rect 7618 33496 7623 33552
rect 1393 33494 7623 33496
rect 7790 33554 7850 33630
rect 10317 33554 10383 33557
rect 7790 33552 10383 33554
rect 7790 33496 10322 33552
rect 10378 33496 10383 33552
rect 7790 33494 10383 33496
rect 1393 33491 1459 33494
rect 7557 33491 7623 33494
rect 10317 33491 10383 33494
rect 1945 33418 2011 33421
rect 9857 33418 9923 33421
rect 1945 33416 9923 33418
rect 1945 33360 1950 33416
rect 2006 33360 9862 33416
rect 9918 33360 9923 33416
rect 1945 33358 9923 33360
rect 1945 33355 2011 33358
rect 9857 33355 9923 33358
rect 10593 33418 10659 33421
rect 12709 33418 12775 33421
rect 10593 33416 12775 33418
rect 10593 33360 10598 33416
rect 10654 33360 12714 33416
rect 12770 33360 12775 33416
rect 10593 33358 12775 33360
rect 10593 33355 10659 33358
rect 12709 33355 12775 33358
rect 13537 33418 13603 33421
rect 15520 33418 16000 33448
rect 13537 33416 16000 33418
rect 13537 33360 13542 33416
rect 13598 33360 16000 33416
rect 13537 33358 16000 33360
rect 13537 33355 13603 33358
rect 15520 33328 16000 33358
rect 6729 33282 6795 33285
rect 9305 33282 9371 33285
rect 6729 33280 9371 33282
rect 6729 33224 6734 33280
rect 6790 33224 9310 33280
rect 9366 33224 9371 33280
rect 6729 33222 9371 33224
rect 6729 33219 6795 33222
rect 9305 33219 9371 33222
rect 6277 33216 6597 33217
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 33151 6597 33152
rect 11610 33216 11930 33217
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 33151 11930 33152
rect 7741 33146 7807 33149
rect 10777 33146 10843 33149
rect 7741 33144 10843 33146
rect 7741 33088 7746 33144
rect 7802 33088 10782 33144
rect 10838 33088 10843 33144
rect 7741 33086 10843 33088
rect 7741 33083 7807 33086
rect 10777 33083 10843 33086
rect 8017 33010 8083 33013
rect 9397 33010 9463 33013
rect 8017 33008 9463 33010
rect 8017 32952 8022 33008
rect 8078 32952 9402 33008
rect 9458 32952 9463 33008
rect 8017 32950 9463 32952
rect 8017 32947 8083 32950
rect 9397 32947 9463 32950
rect 10777 32874 10843 32877
rect 12617 32874 12683 32877
rect 10777 32872 12683 32874
rect 10777 32816 10782 32872
rect 10838 32816 12622 32872
rect 12678 32816 12683 32872
rect 10777 32814 12683 32816
rect 10777 32811 10843 32814
rect 12617 32811 12683 32814
rect 3610 32672 3930 32673
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3930 32672
rect 3610 32607 3930 32608
rect 8944 32672 9264 32673
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 32607 9264 32608
rect 14277 32672 14597 32673
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 32607 14597 32608
rect 3693 32466 3759 32469
rect 8661 32466 8727 32469
rect 3693 32464 8727 32466
rect 3693 32408 3698 32464
rect 3754 32408 8666 32464
rect 8722 32408 8727 32464
rect 3693 32406 8727 32408
rect 3693 32403 3759 32406
rect 8661 32403 8727 32406
rect 2589 32330 2655 32333
rect 7281 32330 7347 32333
rect 2589 32328 7347 32330
rect 2589 32272 2594 32328
rect 2650 32272 7286 32328
rect 7342 32272 7347 32328
rect 2589 32270 7347 32272
rect 2589 32267 2655 32270
rect 7281 32267 7347 32270
rect 10225 32330 10291 32333
rect 15377 32330 15443 32333
rect 10225 32328 15443 32330
rect 10225 32272 10230 32328
rect 10286 32272 15382 32328
rect 15438 32272 15443 32328
rect 10225 32270 15443 32272
rect 10225 32267 10291 32270
rect 15377 32267 15443 32270
rect 3601 32194 3667 32197
rect 6085 32194 6151 32197
rect 3601 32192 6151 32194
rect 3601 32136 3606 32192
rect 3662 32136 6090 32192
rect 6146 32136 6151 32192
rect 3601 32134 6151 32136
rect 3601 32131 3667 32134
rect 6085 32131 6151 32134
rect 9397 32194 9463 32197
rect 10317 32194 10383 32197
rect 9397 32192 10383 32194
rect 9397 32136 9402 32192
rect 9458 32136 10322 32192
rect 10378 32136 10383 32192
rect 9397 32134 10383 32136
rect 9397 32131 9463 32134
rect 10317 32131 10383 32134
rect 6277 32128 6597 32129
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 32063 6597 32064
rect 11610 32128 11930 32129
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 32063 11930 32064
rect 7189 31922 7255 31925
rect 9857 31922 9923 31925
rect 7189 31920 9923 31922
rect 7189 31864 7194 31920
rect 7250 31864 9862 31920
rect 9918 31864 9923 31920
rect 7189 31862 9923 31864
rect 7189 31859 7255 31862
rect 9857 31859 9923 31862
rect 0 31650 480 31680
rect 1577 31650 1643 31653
rect 0 31648 1643 31650
rect 0 31592 1582 31648
rect 1638 31592 1643 31648
rect 0 31590 1643 31592
rect 0 31560 480 31590
rect 1577 31587 1643 31590
rect 3610 31584 3930 31585
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3930 31584
rect 3610 31519 3930 31520
rect 8944 31584 9264 31585
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 31519 9264 31520
rect 14277 31584 14597 31585
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 31519 14597 31520
rect 8017 31378 8083 31381
rect 9949 31378 10015 31381
rect 8017 31376 10015 31378
rect 8017 31320 8022 31376
rect 8078 31320 9954 31376
rect 10010 31320 10015 31376
rect 8017 31318 10015 31320
rect 8017 31315 8083 31318
rect 9949 31315 10015 31318
rect 10501 31378 10567 31381
rect 13721 31378 13787 31381
rect 10501 31376 13787 31378
rect 10501 31320 10506 31376
rect 10562 31320 13726 31376
rect 13782 31320 13787 31376
rect 10501 31318 13787 31320
rect 10501 31315 10567 31318
rect 13721 31315 13787 31318
rect 6277 31040 6597 31041
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 30975 6597 30976
rect 11610 31040 11930 31041
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 30975 11930 30976
rect 6821 30970 6887 30973
rect 10961 30970 11027 30973
rect 6821 30968 11027 30970
rect 6821 30912 6826 30968
rect 6882 30912 10966 30968
rect 11022 30912 11027 30968
rect 6821 30910 11027 30912
rect 6821 30907 6887 30910
rect 10961 30907 11027 30910
rect 3610 30496 3930 30497
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3930 30496
rect 3610 30431 3930 30432
rect 8944 30496 9264 30497
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 30431 9264 30432
rect 14277 30496 14597 30497
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 30431 14597 30432
rect 2405 30290 2471 30293
rect 4981 30290 5047 30293
rect 2405 30288 5047 30290
rect 2405 30232 2410 30288
rect 2466 30232 4986 30288
rect 5042 30232 5047 30288
rect 2405 30230 5047 30232
rect 2405 30227 2471 30230
rect 4981 30227 5047 30230
rect 4337 30154 4403 30157
rect 6177 30154 6243 30157
rect 4337 30152 6243 30154
rect 4337 30096 4342 30152
rect 4398 30096 6182 30152
rect 6238 30096 6243 30152
rect 4337 30094 6243 30096
rect 4337 30091 4403 30094
rect 6177 30091 6243 30094
rect 7189 30018 7255 30021
rect 11237 30018 11303 30021
rect 7189 30016 11303 30018
rect 7189 29960 7194 30016
rect 7250 29960 11242 30016
rect 11298 29960 11303 30016
rect 7189 29958 11303 29960
rect 7189 29955 7255 29958
rect 11237 29955 11303 29958
rect 6277 29952 6597 29953
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 29887 6597 29888
rect 11610 29952 11930 29953
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 29887 11930 29888
rect 5073 29746 5139 29749
rect 14641 29746 14707 29749
rect 5073 29744 14707 29746
rect 5073 29688 5078 29744
rect 5134 29688 14646 29744
rect 14702 29688 14707 29744
rect 5073 29686 14707 29688
rect 5073 29683 5139 29686
rect 3610 29408 3930 29409
rect 0 29338 480 29368
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3930 29408
rect 3610 29343 3930 29344
rect 1577 29338 1643 29341
rect 0 29336 1643 29338
rect 0 29280 1582 29336
rect 1638 29280 1643 29336
rect 0 29278 1643 29280
rect 0 29248 480 29278
rect 1577 29275 1643 29278
rect 5766 29205 5826 29686
rect 14641 29683 14707 29686
rect 8944 29408 9264 29409
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 29343 9264 29344
rect 14277 29408 14597 29409
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 29343 14597 29344
rect 5717 29200 5826 29205
rect 5717 29144 5722 29200
rect 5778 29144 5826 29200
rect 5717 29142 5826 29144
rect 5717 29139 5783 29142
rect 2313 29066 2379 29069
rect 4889 29066 4955 29069
rect 7281 29066 7347 29069
rect 2313 29064 4955 29066
rect 2313 29008 2318 29064
rect 2374 29008 4894 29064
rect 4950 29008 4955 29064
rect 2313 29006 4955 29008
rect 2313 29003 2379 29006
rect 4889 29003 4955 29006
rect 6134 29064 7347 29066
rect 6134 29008 7286 29064
rect 7342 29008 7347 29064
rect 6134 29006 7347 29008
rect 2589 28930 2655 28933
rect 6134 28930 6194 29006
rect 7281 29003 7347 29006
rect 2589 28928 6194 28930
rect 2589 28872 2594 28928
rect 2650 28872 6194 28928
rect 2589 28870 6194 28872
rect 2589 28867 2655 28870
rect 6277 28864 6597 28865
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 28799 6597 28800
rect 11610 28864 11930 28865
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 11610 28799 11930 28800
rect 9397 28796 9463 28797
rect 9397 28794 9444 28796
rect 9352 28792 9444 28794
rect 9352 28736 9402 28792
rect 9352 28734 9444 28736
rect 9397 28732 9444 28734
rect 9508 28732 9514 28796
rect 9397 28731 9463 28732
rect 3610 28320 3930 28321
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3930 28320
rect 3610 28255 3930 28256
rect 8944 28320 9264 28321
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 28255 9264 28256
rect 14277 28320 14597 28321
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 14277 28255 14597 28256
rect 4245 28114 4311 28117
rect 10501 28114 10567 28117
rect 4245 28112 10567 28114
rect 4245 28056 4250 28112
rect 4306 28056 10506 28112
rect 10562 28056 10567 28112
rect 4245 28054 10567 28056
rect 4245 28051 4311 28054
rect 10501 28051 10567 28054
rect 6177 27978 6243 27981
rect 10041 27978 10107 27981
rect 6177 27976 10107 27978
rect 6177 27920 6182 27976
rect 6238 27920 10046 27976
rect 10102 27920 10107 27976
rect 6177 27918 10107 27920
rect 6177 27915 6243 27918
rect 10041 27915 10107 27918
rect 6277 27776 6597 27777
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 27711 6597 27712
rect 11610 27776 11930 27777
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 27711 11930 27712
rect 6821 27706 6887 27709
rect 9029 27706 9095 27709
rect 12065 27708 12131 27709
rect 6821 27704 9095 27706
rect 6821 27648 6826 27704
rect 6882 27648 9034 27704
rect 9090 27648 9095 27704
rect 6821 27646 9095 27648
rect 6821 27643 6887 27646
rect 9029 27643 9095 27646
rect 12014 27644 12020 27708
rect 12084 27706 12131 27708
rect 12084 27704 12176 27706
rect 12126 27648 12176 27704
rect 12084 27646 12176 27648
rect 12084 27644 12131 27646
rect 12065 27643 12131 27644
rect 2773 27570 2839 27573
rect 8293 27570 8359 27573
rect 2773 27568 8359 27570
rect 2773 27512 2778 27568
rect 2834 27512 8298 27568
rect 8354 27512 8359 27568
rect 2773 27510 8359 27512
rect 2773 27507 2839 27510
rect 8293 27507 8359 27510
rect 9489 27570 9555 27573
rect 12065 27570 12131 27573
rect 15009 27570 15075 27573
rect 9489 27568 15075 27570
rect 9489 27512 9494 27568
rect 9550 27512 12070 27568
rect 12126 27512 15014 27568
rect 15070 27512 15075 27568
rect 9489 27510 15075 27512
rect 9489 27507 9555 27510
rect 12065 27507 12131 27510
rect 15009 27507 15075 27510
rect 7649 27434 7715 27437
rect 9949 27434 10015 27437
rect 7649 27432 10015 27434
rect 7649 27376 7654 27432
rect 7710 27376 9954 27432
rect 10010 27376 10015 27432
rect 7649 27374 10015 27376
rect 7649 27371 7715 27374
rect 9949 27371 10015 27374
rect 3610 27232 3930 27233
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3930 27232
rect 3610 27167 3930 27168
rect 8944 27232 9264 27233
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 27167 9264 27168
rect 14277 27232 14597 27233
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 27167 14597 27168
rect 0 27026 480 27056
rect 1577 27026 1643 27029
rect 0 27024 1643 27026
rect 0 26968 1582 27024
rect 1638 26968 1643 27024
rect 0 26966 1643 26968
rect 0 26936 480 26966
rect 1577 26963 1643 26966
rect 7465 27026 7531 27029
rect 8937 27026 9003 27029
rect 7465 27024 9003 27026
rect 7465 26968 7470 27024
rect 7526 26968 8942 27024
rect 8998 26968 9003 27024
rect 7465 26966 9003 26968
rect 7465 26963 7531 26966
rect 8937 26963 9003 26966
rect 10685 27026 10751 27029
rect 12985 27026 13051 27029
rect 10685 27024 13051 27026
rect 10685 26968 10690 27024
rect 10746 26968 12990 27024
rect 13046 26968 13051 27024
rect 10685 26966 13051 26968
rect 10685 26963 10751 26966
rect 12985 26963 13051 26966
rect 2221 26890 2287 26893
rect 7925 26890 7991 26893
rect 2221 26888 7991 26890
rect 2221 26832 2226 26888
rect 2282 26832 7930 26888
rect 7986 26832 7991 26888
rect 2221 26830 7991 26832
rect 2221 26827 2287 26830
rect 7925 26827 7991 26830
rect 10317 26890 10383 26893
rect 12801 26890 12867 26893
rect 10317 26888 12867 26890
rect 10317 26832 10322 26888
rect 10378 26832 12806 26888
rect 12862 26832 12867 26888
rect 10317 26830 12867 26832
rect 10317 26827 10383 26830
rect 12801 26827 12867 26830
rect 10133 26754 10199 26757
rect 10593 26754 10659 26757
rect 10133 26752 10659 26754
rect 10133 26696 10138 26752
rect 10194 26696 10598 26752
rect 10654 26696 10659 26752
rect 10133 26694 10659 26696
rect 10133 26691 10199 26694
rect 10593 26691 10659 26694
rect 6277 26688 6597 26689
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 26623 6597 26624
rect 11610 26688 11930 26689
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 26623 11930 26624
rect 8845 26482 8911 26485
rect 8845 26480 10058 26482
rect 8845 26424 8850 26480
rect 8906 26424 10058 26480
rect 8845 26422 10058 26424
rect 8845 26419 8911 26422
rect 8569 26346 8635 26349
rect 9857 26346 9923 26349
rect 8569 26344 9923 26346
rect 8569 26288 8574 26344
rect 8630 26288 9862 26344
rect 9918 26288 9923 26344
rect 8569 26286 9923 26288
rect 8569 26283 8635 26286
rect 9857 26283 9923 26286
rect 9581 26210 9647 26213
rect 9857 26210 9923 26213
rect 9998 26210 10058 26422
rect 9581 26208 9690 26210
rect 9581 26152 9586 26208
rect 9642 26152 9690 26208
rect 9581 26147 9690 26152
rect 9857 26208 10058 26210
rect 9857 26152 9862 26208
rect 9918 26152 10058 26208
rect 9857 26150 10058 26152
rect 9857 26147 9923 26150
rect 3610 26144 3930 26145
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3930 26144
rect 3610 26079 3930 26080
rect 8944 26144 9264 26145
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 26079 9264 26080
rect 9630 25941 9690 26147
rect 14277 26144 14597 26145
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 26079 14597 26080
rect 9581 25936 9690 25941
rect 9581 25880 9586 25936
rect 9642 25880 9690 25936
rect 9581 25878 9690 25880
rect 9581 25875 9647 25878
rect 6277 25600 6597 25601
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 6277 25535 6597 25536
rect 11610 25600 11930 25601
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 25535 11930 25536
rect 2497 25258 2563 25261
rect 9673 25258 9739 25261
rect 2497 25256 9739 25258
rect 2497 25200 2502 25256
rect 2558 25200 9678 25256
rect 9734 25200 9739 25256
rect 2497 25198 9739 25200
rect 2497 25195 2563 25198
rect 9673 25195 9739 25198
rect 3610 25056 3930 25057
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3930 25056
rect 3610 24991 3930 24992
rect 8944 25056 9264 25057
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 24991 9264 24992
rect 14277 25056 14597 25057
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 24991 14597 24992
rect 5717 24988 5783 24989
rect 5717 24984 5764 24988
rect 5828 24986 5834 24988
rect 10317 24986 10383 24989
rect 12065 24986 12131 24989
rect 13261 24986 13327 24989
rect 5717 24928 5722 24984
rect 5717 24924 5764 24928
rect 5828 24926 5874 24986
rect 10317 24984 13327 24986
rect 10317 24928 10322 24984
rect 10378 24928 12070 24984
rect 12126 24928 13266 24984
rect 13322 24928 13327 24984
rect 10317 24926 13327 24928
rect 5828 24924 5834 24926
rect 5717 24923 5783 24924
rect 10317 24923 10383 24926
rect 12065 24923 12131 24926
rect 13261 24923 13327 24926
rect 4889 24850 4955 24853
rect 14089 24850 14155 24853
rect 4889 24848 14155 24850
rect 4889 24792 4894 24848
rect 4950 24792 14094 24848
rect 14150 24792 14155 24848
rect 4889 24790 14155 24792
rect 4889 24787 4955 24790
rect 14089 24787 14155 24790
rect 5625 24714 5691 24717
rect 7557 24714 7623 24717
rect 5625 24712 7623 24714
rect 5625 24656 5630 24712
rect 5686 24656 7562 24712
rect 7618 24656 7623 24712
rect 5625 24654 7623 24656
rect 5625 24651 5691 24654
rect 7557 24651 7623 24654
rect 0 24578 480 24608
rect 1577 24578 1643 24581
rect 0 24576 1643 24578
rect 0 24520 1582 24576
rect 1638 24520 1643 24576
rect 0 24518 1643 24520
rect 0 24488 480 24518
rect 1577 24515 1643 24518
rect 6277 24512 6597 24513
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 24447 6597 24448
rect 11610 24512 11930 24513
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 24447 11930 24448
rect 3610 23968 3930 23969
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3930 23968
rect 3610 23903 3930 23904
rect 8944 23968 9264 23969
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 23903 9264 23904
rect 14277 23968 14597 23969
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 23903 14597 23904
rect 4797 23898 4863 23901
rect 6729 23898 6795 23901
rect 4797 23896 6795 23898
rect 4797 23840 4802 23896
rect 4858 23840 6734 23896
rect 6790 23840 6795 23896
rect 4797 23838 6795 23840
rect 4797 23835 4863 23838
rect 6729 23835 6795 23838
rect 6277 23424 6597 23425
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 23359 6597 23360
rect 11610 23424 11930 23425
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 23359 11930 23360
rect 5165 23218 5231 23221
rect 9581 23218 9647 23221
rect 5165 23216 9647 23218
rect 5165 23160 5170 23216
rect 5226 23160 9586 23216
rect 9642 23160 9647 23216
rect 5165 23158 9647 23160
rect 5165 23155 5231 23158
rect 9581 23155 9647 23158
rect 8017 23082 8083 23085
rect 9673 23082 9739 23085
rect 8017 23080 9739 23082
rect 8017 23024 8022 23080
rect 8078 23024 9678 23080
rect 9734 23024 9739 23080
rect 8017 23022 9739 23024
rect 8017 23019 8083 23022
rect 9673 23019 9739 23022
rect 3610 22880 3930 22881
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3930 22880
rect 3610 22815 3930 22816
rect 8944 22880 9264 22881
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 22815 9264 22816
rect 14277 22880 14597 22881
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 22815 14597 22816
rect 7281 22674 7347 22677
rect 11789 22674 11855 22677
rect 7281 22672 11855 22674
rect 7281 22616 7286 22672
rect 7342 22616 11794 22672
rect 11850 22616 11855 22672
rect 7281 22614 11855 22616
rect 7281 22611 7347 22614
rect 11789 22611 11855 22614
rect 6277 22336 6597 22337
rect 0 22266 480 22296
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 6277 22271 6597 22272
rect 11610 22336 11930 22337
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 22271 11930 22272
rect 1669 22266 1735 22269
rect 5165 22266 5231 22269
rect 0 22206 1594 22266
rect 0 22176 480 22206
rect 1534 21997 1594 22206
rect 1669 22264 5231 22266
rect 1669 22208 1674 22264
rect 1730 22208 5170 22264
rect 5226 22208 5231 22264
rect 1669 22206 5231 22208
rect 1669 22203 1735 22206
rect 5165 22203 5231 22206
rect 1534 21992 1643 21997
rect 1534 21936 1582 21992
rect 1638 21936 1643 21992
rect 1534 21934 1643 21936
rect 1577 21931 1643 21934
rect 10777 21858 10843 21861
rect 12433 21858 12499 21861
rect 10777 21856 12499 21858
rect 10777 21800 10782 21856
rect 10838 21800 12438 21856
rect 12494 21800 12499 21856
rect 10777 21798 12499 21800
rect 10777 21795 10843 21798
rect 12433 21795 12499 21798
rect 3610 21792 3930 21793
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3930 21792
rect 3610 21727 3930 21728
rect 8944 21792 9264 21793
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 21727 9264 21728
rect 14277 21792 14597 21793
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 21727 14597 21728
rect 5349 21586 5415 21589
rect 6637 21586 6703 21589
rect 5349 21584 6703 21586
rect 5349 21528 5354 21584
rect 5410 21528 6642 21584
rect 6698 21528 6703 21584
rect 5349 21526 6703 21528
rect 5349 21523 5415 21526
rect 6637 21523 6703 21526
rect 1945 21450 2011 21453
rect 9673 21450 9739 21453
rect 1945 21448 9739 21450
rect 1945 21392 1950 21448
rect 2006 21392 9678 21448
rect 9734 21392 9739 21448
rect 1945 21390 9739 21392
rect 1945 21387 2011 21390
rect 9673 21387 9739 21390
rect 5717 21316 5783 21317
rect 5717 21314 5764 21316
rect 5672 21312 5764 21314
rect 5672 21256 5722 21312
rect 5672 21254 5764 21256
rect 5717 21252 5764 21254
rect 5828 21252 5834 21316
rect 5717 21251 5783 21252
rect 6277 21248 6597 21249
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 21183 6597 21184
rect 11610 21248 11930 21249
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 11610 21183 11930 21184
rect 7557 21042 7623 21045
rect 11145 21042 11211 21045
rect 7557 21040 11211 21042
rect 7557 20984 7562 21040
rect 7618 20984 11150 21040
rect 11206 20984 11211 21040
rect 7557 20982 11211 20984
rect 7557 20979 7623 20982
rect 11145 20979 11211 20982
rect 4613 20906 4679 20909
rect 11513 20906 11579 20909
rect 4613 20904 11579 20906
rect 4613 20848 4618 20904
rect 4674 20848 11518 20904
rect 11574 20848 11579 20904
rect 4613 20846 11579 20848
rect 4613 20843 4679 20846
rect 11513 20843 11579 20846
rect 3610 20704 3930 20705
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3930 20704
rect 3610 20639 3930 20640
rect 8944 20704 9264 20705
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 20639 9264 20640
rect 14277 20704 14597 20705
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 14277 20639 14597 20640
rect 9581 20634 9647 20637
rect 12617 20634 12683 20637
rect 9581 20632 12683 20634
rect 9581 20576 9586 20632
rect 9642 20576 12622 20632
rect 12678 20576 12683 20632
rect 9581 20574 12683 20576
rect 9581 20571 9647 20574
rect 12617 20571 12683 20574
rect 9438 20300 9444 20364
rect 9508 20362 9514 20364
rect 9581 20362 9647 20365
rect 9508 20360 9647 20362
rect 9508 20304 9586 20360
rect 9642 20304 9647 20360
rect 9508 20302 9647 20304
rect 9508 20300 9514 20302
rect 9581 20299 9647 20302
rect 6277 20160 6597 20161
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 20095 6597 20096
rect 11610 20160 11930 20161
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 20095 11930 20096
rect 12065 20090 12131 20093
rect 15520 20090 16000 20120
rect 12065 20088 16000 20090
rect 12065 20032 12070 20088
rect 12126 20032 16000 20088
rect 12065 20030 16000 20032
rect 12065 20027 12131 20030
rect 15520 20000 16000 20030
rect 0 19954 480 19984
rect 1577 19954 1643 19957
rect 12065 19956 12131 19957
rect 0 19952 1643 19954
rect 0 19896 1582 19952
rect 1638 19896 1643 19952
rect 0 19894 1643 19896
rect 0 19864 480 19894
rect 1577 19891 1643 19894
rect 12014 19892 12020 19956
rect 12084 19954 12131 19956
rect 12084 19952 12176 19954
rect 12126 19896 12176 19952
rect 12084 19894 12176 19896
rect 12084 19892 12131 19894
rect 12065 19891 12131 19892
rect 4705 19818 4771 19821
rect 11145 19818 11211 19821
rect 4705 19816 11211 19818
rect 4705 19760 4710 19816
rect 4766 19760 11150 19816
rect 11206 19760 11211 19816
rect 4705 19758 11211 19760
rect 4705 19755 4771 19758
rect 11145 19755 11211 19758
rect 3610 19616 3930 19617
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3930 19616
rect 3610 19551 3930 19552
rect 8944 19616 9264 19617
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 19551 9264 19552
rect 14277 19616 14597 19617
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 19551 14597 19552
rect 3417 19410 3483 19413
rect 5165 19410 5231 19413
rect 10777 19410 10843 19413
rect 3417 19408 10843 19410
rect 3417 19352 3422 19408
rect 3478 19352 5170 19408
rect 5226 19352 10782 19408
rect 10838 19352 10843 19408
rect 3417 19350 10843 19352
rect 3417 19347 3483 19350
rect 5165 19347 5231 19350
rect 10777 19347 10843 19350
rect 7649 19274 7715 19277
rect 10685 19274 10751 19277
rect 7649 19272 10751 19274
rect 7649 19216 7654 19272
rect 7710 19216 10690 19272
rect 10746 19216 10751 19272
rect 7649 19214 10751 19216
rect 7649 19211 7715 19214
rect 10685 19211 10751 19214
rect 8109 19138 8175 19141
rect 9121 19138 9187 19141
rect 11421 19138 11487 19141
rect 8109 19136 11487 19138
rect 8109 19080 8114 19136
rect 8170 19080 9126 19136
rect 9182 19080 11426 19136
rect 11482 19080 11487 19136
rect 8109 19078 11487 19080
rect 8109 19075 8175 19078
rect 9121 19075 9187 19078
rect 11421 19075 11487 19078
rect 6277 19072 6597 19073
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 19007 6597 19008
rect 11610 19072 11930 19073
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 19007 11930 19008
rect 3610 18528 3930 18529
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3930 18528
rect 3610 18463 3930 18464
rect 8944 18528 9264 18529
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 18463 9264 18464
rect 14277 18528 14597 18529
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 18463 14597 18464
rect 6277 17984 6597 17985
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 6277 17919 6597 17920
rect 11610 17984 11930 17985
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 17919 11930 17920
rect 1945 17778 2011 17781
rect 7741 17778 7807 17781
rect 1945 17776 7807 17778
rect 1945 17720 1950 17776
rect 2006 17720 7746 17776
rect 7802 17720 7807 17776
rect 1945 17718 7807 17720
rect 1945 17715 2011 17718
rect 7741 17715 7807 17718
rect 0 17642 480 17672
rect 1577 17642 1643 17645
rect 0 17640 1643 17642
rect 0 17584 1582 17640
rect 1638 17584 1643 17640
rect 0 17582 1643 17584
rect 0 17552 480 17582
rect 1577 17579 1643 17582
rect 3141 17642 3207 17645
rect 4245 17642 4311 17645
rect 10225 17642 10291 17645
rect 10777 17642 10843 17645
rect 3141 17640 10843 17642
rect 3141 17584 3146 17640
rect 3202 17584 4250 17640
rect 4306 17584 10230 17640
rect 10286 17584 10782 17640
rect 10838 17584 10843 17640
rect 3141 17582 10843 17584
rect 3141 17579 3207 17582
rect 4245 17579 4311 17582
rect 10225 17579 10291 17582
rect 10777 17579 10843 17582
rect 3610 17440 3930 17441
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3930 17440
rect 3610 17375 3930 17376
rect 8944 17440 9264 17441
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 17375 9264 17376
rect 14277 17440 14597 17441
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 17375 14597 17376
rect 9489 17370 9555 17373
rect 9446 17368 9555 17370
rect 9446 17312 9494 17368
rect 9550 17312 9555 17368
rect 9446 17307 9555 17312
rect 5022 17172 5028 17236
rect 5092 17234 5098 17236
rect 5441 17234 5507 17237
rect 5092 17232 5507 17234
rect 5092 17176 5446 17232
rect 5502 17176 5507 17232
rect 5092 17174 5507 17176
rect 5092 17172 5098 17174
rect 5441 17171 5507 17174
rect 8937 17234 9003 17237
rect 9446 17234 9506 17307
rect 8937 17232 9506 17234
rect 8937 17176 8942 17232
rect 8998 17176 9506 17232
rect 8937 17174 9506 17176
rect 8937 17171 9003 17174
rect 5349 17098 5415 17101
rect 10409 17098 10475 17101
rect 5349 17096 10475 17098
rect 5349 17040 5354 17096
rect 5410 17040 10414 17096
rect 10470 17040 10475 17096
rect 5349 17038 10475 17040
rect 5349 17035 5415 17038
rect 10409 17035 10475 17038
rect 7833 16962 7899 16965
rect 9673 16962 9739 16965
rect 7833 16960 9739 16962
rect 7833 16904 7838 16960
rect 7894 16904 9678 16960
rect 9734 16904 9739 16960
rect 7833 16902 9739 16904
rect 7833 16899 7899 16902
rect 9673 16899 9739 16902
rect 6277 16896 6597 16897
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 16831 6597 16832
rect 11610 16896 11930 16897
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 16831 11930 16832
rect 2405 16826 2471 16829
rect 4521 16826 4587 16829
rect 2405 16824 4587 16826
rect 2405 16768 2410 16824
rect 2466 16768 4526 16824
rect 4582 16768 4587 16824
rect 2405 16766 4587 16768
rect 2405 16763 2471 16766
rect 4521 16763 4587 16766
rect 10501 16690 10567 16693
rect 12985 16690 13051 16693
rect 10501 16688 13051 16690
rect 10501 16632 10506 16688
rect 10562 16632 12990 16688
rect 13046 16632 13051 16688
rect 10501 16630 13051 16632
rect 10501 16627 10567 16630
rect 12985 16627 13051 16630
rect 7281 16554 7347 16557
rect 10041 16554 10107 16557
rect 7281 16552 10107 16554
rect 7281 16496 7286 16552
rect 7342 16496 10046 16552
rect 10102 16496 10107 16552
rect 7281 16494 10107 16496
rect 7281 16491 7347 16494
rect 10041 16491 10107 16494
rect 3610 16352 3930 16353
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3930 16352
rect 3610 16287 3930 16288
rect 8944 16352 9264 16353
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 16287 9264 16288
rect 14277 16352 14597 16353
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 16287 14597 16288
rect 1393 16146 1459 16149
rect 9857 16146 9923 16149
rect 1393 16144 9923 16146
rect 1393 16088 1398 16144
rect 1454 16088 9862 16144
rect 9918 16088 9923 16144
rect 1393 16086 9923 16088
rect 1393 16083 1459 16086
rect 9857 16083 9923 16086
rect 7741 16010 7807 16013
rect 10041 16010 10107 16013
rect 10225 16010 10291 16013
rect 7741 16008 10291 16010
rect 7741 15952 7746 16008
rect 7802 15952 10046 16008
rect 10102 15952 10230 16008
rect 10286 15952 10291 16008
rect 7741 15950 10291 15952
rect 7741 15947 7807 15950
rect 10041 15947 10107 15950
rect 10225 15947 10291 15950
rect 6277 15808 6597 15809
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 15743 6597 15744
rect 11610 15808 11930 15809
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 15743 11930 15744
rect 3610 15264 3930 15265
rect 0 15194 480 15224
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3930 15264
rect 3610 15199 3930 15200
rect 8944 15264 9264 15265
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 15199 9264 15200
rect 14277 15264 14597 15265
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 15199 14597 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 480 15134
rect 1485 15131 1551 15134
rect 4429 15058 4495 15061
rect 11513 15058 11579 15061
rect 4429 15056 11579 15058
rect 4429 15000 4434 15056
rect 4490 15000 11518 15056
rect 11574 15000 11579 15056
rect 4429 14998 11579 15000
rect 4429 14995 4495 14998
rect 11513 14995 11579 14998
rect 5809 14922 5875 14925
rect 7281 14922 7347 14925
rect 5809 14920 7347 14922
rect 5809 14864 5814 14920
rect 5870 14864 7286 14920
rect 7342 14864 7347 14920
rect 5809 14862 7347 14864
rect 5809 14859 5875 14862
rect 7281 14859 7347 14862
rect 6277 14720 6597 14721
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 14655 6597 14656
rect 11610 14720 11930 14721
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 14655 11930 14656
rect 3325 14650 3391 14653
rect 5073 14650 5139 14653
rect 3325 14648 5139 14650
rect 3325 14592 3330 14648
rect 3386 14592 5078 14648
rect 5134 14592 5139 14648
rect 3325 14590 5139 14592
rect 3325 14587 3391 14590
rect 5073 14587 5139 14590
rect 7373 14650 7439 14653
rect 9765 14650 9831 14653
rect 7373 14648 9831 14650
rect 7373 14592 7378 14648
rect 7434 14592 9770 14648
rect 9826 14592 9831 14648
rect 7373 14590 9831 14592
rect 7373 14587 7439 14590
rect 9765 14587 9831 14590
rect 5349 14514 5415 14517
rect 10685 14514 10751 14517
rect 5349 14512 10751 14514
rect 5349 14456 5354 14512
rect 5410 14456 10690 14512
rect 10746 14456 10751 14512
rect 5349 14454 10751 14456
rect 5349 14451 5415 14454
rect 10685 14451 10751 14454
rect 3610 14176 3930 14177
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3930 14176
rect 3610 14111 3930 14112
rect 8944 14176 9264 14177
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 14111 9264 14112
rect 14277 14176 14597 14177
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 14111 14597 14112
rect 7833 13970 7899 13973
rect 10501 13970 10567 13973
rect 7833 13968 10567 13970
rect 7833 13912 7838 13968
rect 7894 13912 10506 13968
rect 10562 13912 10567 13968
rect 7833 13910 10567 13912
rect 7833 13907 7899 13910
rect 10501 13907 10567 13910
rect 4613 13834 4679 13837
rect 4889 13834 4955 13837
rect 4613 13832 4955 13834
rect 4613 13776 4618 13832
rect 4674 13776 4894 13832
rect 4950 13776 4955 13832
rect 4613 13774 4955 13776
rect 4613 13771 4679 13774
rect 4889 13771 4955 13774
rect 7649 13834 7715 13837
rect 11973 13834 12039 13837
rect 7649 13832 12039 13834
rect 7649 13776 7654 13832
rect 7710 13776 11978 13832
rect 12034 13776 12039 13832
rect 7649 13774 12039 13776
rect 7649 13771 7715 13774
rect 11973 13771 12039 13774
rect 7833 13698 7899 13701
rect 10777 13698 10843 13701
rect 7833 13696 10843 13698
rect 7833 13640 7838 13696
rect 7894 13640 10782 13696
rect 10838 13640 10843 13696
rect 7833 13638 10843 13640
rect 7833 13635 7899 13638
rect 10777 13635 10843 13638
rect 6277 13632 6597 13633
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 13567 6597 13568
rect 11610 13632 11930 13633
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 13567 11930 13568
rect 3610 13088 3930 13089
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3930 13088
rect 3610 13023 3930 13024
rect 8944 13088 9264 13089
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 13023 9264 13024
rect 14277 13088 14597 13089
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 13023 14597 13024
rect 0 12882 480 12912
rect 1577 12882 1643 12885
rect 0 12880 1643 12882
rect 0 12824 1582 12880
rect 1638 12824 1643 12880
rect 0 12822 1643 12824
rect 0 12792 480 12822
rect 1577 12819 1643 12822
rect 1669 12746 1735 12749
rect 6177 12746 6243 12749
rect 1669 12744 6243 12746
rect 1669 12688 1674 12744
rect 1730 12688 6182 12744
rect 6238 12688 6243 12744
rect 1669 12686 6243 12688
rect 1669 12683 1735 12686
rect 6177 12683 6243 12686
rect 6277 12544 6597 12545
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 6277 12479 6597 12480
rect 11610 12544 11930 12545
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 12479 11930 12480
rect 7281 12202 7347 12205
rect 13721 12202 13787 12205
rect 7281 12200 13787 12202
rect 7281 12144 7286 12200
rect 7342 12144 13726 12200
rect 13782 12144 13787 12200
rect 7281 12142 13787 12144
rect 7281 12139 7347 12142
rect 13721 12139 13787 12142
rect 3610 12000 3930 12001
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3930 12000
rect 3610 11935 3930 11936
rect 8944 12000 9264 12001
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 11935 9264 11936
rect 14277 12000 14597 12001
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 11935 14597 11936
rect 4981 11660 5047 11661
rect 4981 11658 5028 11660
rect 4936 11656 5028 11658
rect 4936 11600 4986 11656
rect 4936 11598 5028 11600
rect 4981 11596 5028 11598
rect 5092 11596 5098 11660
rect 4981 11595 5047 11596
rect 6277 11456 6597 11457
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 11391 6597 11392
rect 11610 11456 11930 11457
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 11391 11930 11392
rect 9581 11114 9647 11117
rect 12065 11114 12131 11117
rect 9581 11112 12131 11114
rect 9581 11056 9586 11112
rect 9642 11056 12070 11112
rect 12126 11056 12131 11112
rect 9581 11054 12131 11056
rect 9581 11051 9647 11054
rect 12065 11051 12131 11054
rect 3610 10912 3930 10913
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3930 10912
rect 3610 10847 3930 10848
rect 8944 10912 9264 10913
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 10847 9264 10848
rect 14277 10912 14597 10913
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 10847 14597 10848
rect 0 10570 480 10600
rect 1577 10570 1643 10573
rect 0 10568 1643 10570
rect 0 10512 1582 10568
rect 1638 10512 1643 10568
rect 0 10510 1643 10512
rect 0 10480 480 10510
rect 1577 10507 1643 10510
rect 7373 10434 7439 10437
rect 11237 10434 11303 10437
rect 7373 10432 11303 10434
rect 7373 10376 7378 10432
rect 7434 10376 11242 10432
rect 11298 10376 11303 10432
rect 7373 10374 11303 10376
rect 7373 10371 7439 10374
rect 11237 10371 11303 10374
rect 6277 10368 6597 10369
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 10303 6597 10304
rect 11610 10368 11930 10369
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 10303 11930 10304
rect 7373 10162 7439 10165
rect 13445 10162 13511 10165
rect 7373 10160 13511 10162
rect 7373 10104 7378 10160
rect 7434 10104 13450 10160
rect 13506 10104 13511 10160
rect 7373 10102 13511 10104
rect 7373 10099 7439 10102
rect 13445 10099 13511 10102
rect 5165 10026 5231 10029
rect 10041 10026 10107 10029
rect 5165 10024 10107 10026
rect 5165 9968 5170 10024
rect 5226 9968 10046 10024
rect 10102 9968 10107 10024
rect 5165 9966 10107 9968
rect 5165 9963 5231 9966
rect 10041 9963 10107 9966
rect 3610 9824 3930 9825
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3930 9824
rect 3610 9759 3930 9760
rect 8944 9824 9264 9825
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 8944 9759 9264 9760
rect 14277 9824 14597 9825
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 9759 14597 9760
rect 3325 9482 3391 9485
rect 7741 9482 7807 9485
rect 3325 9480 7807 9482
rect 3325 9424 3330 9480
rect 3386 9424 7746 9480
rect 7802 9424 7807 9480
rect 3325 9422 7807 9424
rect 3325 9419 3391 9422
rect 7741 9419 7807 9422
rect 10777 9482 10843 9485
rect 13261 9482 13327 9485
rect 10777 9480 13327 9482
rect 10777 9424 10782 9480
rect 10838 9424 13266 9480
rect 13322 9424 13327 9480
rect 10777 9422 13327 9424
rect 10777 9419 10843 9422
rect 13261 9419 13327 9422
rect 6277 9280 6597 9281
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 9215 6597 9216
rect 11610 9280 11930 9281
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 9215 11930 9216
rect 7966 9012 7972 9076
rect 8036 9074 8042 9076
rect 8477 9074 8543 9077
rect 8036 9072 8543 9074
rect 8036 9016 8482 9072
rect 8538 9016 8543 9072
rect 8036 9014 8543 9016
rect 8036 9012 8042 9014
rect 8477 9011 8543 9014
rect 8753 9074 8819 9077
rect 9949 9074 10015 9077
rect 8753 9072 10015 9074
rect 8753 9016 8758 9072
rect 8814 9016 9954 9072
rect 10010 9016 10015 9072
rect 8753 9014 10015 9016
rect 8753 9011 8819 9014
rect 9949 9011 10015 9014
rect 9213 8938 9279 8941
rect 11145 8938 11211 8941
rect 9213 8936 11211 8938
rect 9213 8880 9218 8936
rect 9274 8880 11150 8936
rect 11206 8880 11211 8936
rect 9213 8878 11211 8880
rect 9213 8875 9279 8878
rect 11145 8875 11211 8878
rect 10869 8802 10935 8805
rect 13077 8802 13143 8805
rect 10869 8800 13143 8802
rect 10869 8744 10874 8800
rect 10930 8744 13082 8800
rect 13138 8744 13143 8800
rect 10869 8742 13143 8744
rect 10869 8739 10935 8742
rect 13077 8739 13143 8742
rect 3610 8736 3930 8737
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3930 8736
rect 3610 8671 3930 8672
rect 8944 8736 9264 8737
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 8671 9264 8672
rect 14277 8736 14597 8737
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 8671 14597 8672
rect 3785 8530 3851 8533
rect 10133 8530 10199 8533
rect 3785 8528 10199 8530
rect 3785 8472 3790 8528
rect 3846 8472 10138 8528
rect 10194 8472 10199 8528
rect 3785 8470 10199 8472
rect 3785 8467 3851 8470
rect 10133 8467 10199 8470
rect 3141 8394 3207 8397
rect 6545 8394 6611 8397
rect 3141 8392 6611 8394
rect 3141 8336 3146 8392
rect 3202 8336 6550 8392
rect 6606 8336 6611 8392
rect 3141 8334 6611 8336
rect 3141 8331 3207 8334
rect 6545 8331 6611 8334
rect 8017 8394 8083 8397
rect 10777 8394 10843 8397
rect 8017 8392 10843 8394
rect 8017 8336 8022 8392
rect 8078 8336 10782 8392
rect 10838 8336 10843 8392
rect 8017 8334 10843 8336
rect 8017 8331 8083 8334
rect 10777 8331 10843 8334
rect 13169 8394 13235 8397
rect 14641 8394 14707 8397
rect 13169 8392 14707 8394
rect 13169 8336 13174 8392
rect 13230 8336 14646 8392
rect 14702 8336 14707 8392
rect 13169 8334 14707 8336
rect 13169 8331 13235 8334
rect 14641 8331 14707 8334
rect 6277 8192 6597 8193
rect 0 8122 480 8152
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 8127 6597 8128
rect 11610 8192 11930 8193
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 8127 11930 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 480 8062
rect 2773 8059 2839 8062
rect 7373 7988 7439 7989
rect 7373 7986 7420 7988
rect 7292 7984 7420 7986
rect 7484 7986 7490 7988
rect 12893 7986 12959 7989
rect 7484 7984 12959 7986
rect 7292 7928 7378 7984
rect 7484 7928 12898 7984
rect 12954 7928 12959 7984
rect 7292 7926 7420 7928
rect 7373 7924 7420 7926
rect 7484 7926 12959 7928
rect 7484 7924 7490 7926
rect 7373 7923 7439 7924
rect 12893 7923 12959 7926
rect 8201 7850 8267 7853
rect 10225 7850 10291 7853
rect 8201 7848 10291 7850
rect 8201 7792 8206 7848
rect 8262 7792 10230 7848
rect 10286 7792 10291 7848
rect 8201 7790 10291 7792
rect 8201 7787 8267 7790
rect 10225 7787 10291 7790
rect 3610 7648 3930 7649
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3930 7648
rect 3610 7583 3930 7584
rect 8944 7648 9264 7649
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 7583 9264 7584
rect 14277 7648 14597 7649
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 7583 14597 7584
rect 5257 7306 5323 7309
rect 10409 7306 10475 7309
rect 5257 7304 10475 7306
rect 5257 7248 5262 7304
rect 5318 7248 10414 7304
rect 10470 7248 10475 7304
rect 5257 7246 10475 7248
rect 5257 7243 5323 7246
rect 10409 7243 10475 7246
rect 6277 7104 6597 7105
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 7039 6597 7040
rect 11610 7104 11930 7105
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 7039 11930 7040
rect 8937 6898 9003 6901
rect 9397 6898 9463 6901
rect 15377 6898 15443 6901
rect 8937 6896 15443 6898
rect 8937 6840 8942 6896
rect 8998 6840 9402 6896
rect 9458 6840 15382 6896
rect 15438 6840 15443 6896
rect 8937 6838 15443 6840
rect 8937 6835 9003 6838
rect 9397 6835 9463 6838
rect 15377 6835 15443 6838
rect 5257 6762 5323 6765
rect 10317 6762 10383 6765
rect 5257 6760 10383 6762
rect 5257 6704 5262 6760
rect 5318 6704 10322 6760
rect 10378 6704 10383 6760
rect 5257 6702 10383 6704
rect 5257 6699 5323 6702
rect 10317 6699 10383 6702
rect 12157 6762 12223 6765
rect 15520 6762 16000 6792
rect 12157 6760 16000 6762
rect 12157 6704 12162 6760
rect 12218 6704 16000 6760
rect 12157 6702 16000 6704
rect 12157 6699 12223 6702
rect 15520 6672 16000 6702
rect 3610 6560 3930 6561
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3930 6560
rect 3610 6495 3930 6496
rect 8944 6560 9264 6561
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 6495 9264 6496
rect 14277 6560 14597 6561
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 6495 14597 6496
rect 4981 6218 5047 6221
rect 9305 6218 9371 6221
rect 4981 6216 9371 6218
rect 4981 6160 4986 6216
rect 5042 6160 9310 6216
rect 9366 6160 9371 6216
rect 4981 6158 9371 6160
rect 4981 6155 5047 6158
rect 9305 6155 9371 6158
rect 3049 6082 3115 6085
rect 5809 6082 5875 6085
rect 3049 6080 5875 6082
rect 3049 6024 3054 6080
rect 3110 6024 5814 6080
rect 5870 6024 5875 6080
rect 3049 6022 5875 6024
rect 3049 6019 3115 6022
rect 5809 6019 5875 6022
rect 6277 6016 6597 6017
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 5951 6597 5952
rect 11610 6016 11930 6017
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 5951 11930 5952
rect 0 5810 480 5840
rect 2681 5810 2747 5813
rect 0 5808 2747 5810
rect 0 5752 2686 5808
rect 2742 5752 2747 5808
rect 0 5750 2747 5752
rect 0 5720 480 5750
rect 2681 5747 2747 5750
rect 7097 5810 7163 5813
rect 9673 5810 9739 5813
rect 7097 5808 9739 5810
rect 7097 5752 7102 5808
rect 7158 5752 9678 5808
rect 9734 5752 9739 5808
rect 7097 5750 9739 5752
rect 7097 5747 7163 5750
rect 9673 5747 9739 5750
rect 2129 5674 2195 5677
rect 7100 5674 7160 5747
rect 2129 5672 7160 5674
rect 2129 5616 2134 5672
rect 2190 5616 7160 5672
rect 2129 5614 7160 5616
rect 2129 5611 2195 5614
rect 3610 5472 3930 5473
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3930 5472
rect 3610 5407 3930 5408
rect 8944 5472 9264 5473
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 5407 9264 5408
rect 14277 5472 14597 5473
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 5407 14597 5408
rect 2405 5266 2471 5269
rect 7557 5266 7623 5269
rect 2405 5264 7623 5266
rect 2405 5208 2410 5264
rect 2466 5208 7562 5264
rect 7618 5208 7623 5264
rect 2405 5206 7623 5208
rect 2405 5203 2471 5206
rect 7557 5203 7623 5206
rect 2405 5130 2471 5133
rect 10317 5130 10383 5133
rect 2405 5128 10383 5130
rect 2405 5072 2410 5128
rect 2466 5072 10322 5128
rect 10378 5072 10383 5128
rect 2405 5070 10383 5072
rect 2405 5067 2471 5070
rect 5398 4997 5458 5070
rect 10317 5067 10383 5070
rect 5349 4992 5458 4997
rect 5349 4936 5354 4992
rect 5410 4936 5458 4992
rect 5349 4934 5458 4936
rect 8109 4994 8175 4997
rect 11145 4994 11211 4997
rect 8109 4992 11211 4994
rect 8109 4936 8114 4992
rect 8170 4936 11150 4992
rect 11206 4936 11211 4992
rect 8109 4934 11211 4936
rect 5349 4931 5415 4934
rect 8109 4931 8175 4934
rect 11145 4931 11211 4934
rect 6277 4928 6597 4929
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 4863 6597 4864
rect 11610 4928 11930 4929
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 4863 11930 4864
rect 4889 4722 4955 4725
rect 10685 4722 10751 4725
rect 4889 4720 10751 4722
rect 4889 4664 4894 4720
rect 4950 4664 10690 4720
rect 10746 4664 10751 4720
rect 4889 4662 10751 4664
rect 4889 4659 4955 4662
rect 10685 4659 10751 4662
rect 1945 4586 2011 4589
rect 5441 4586 5507 4589
rect 1945 4584 5507 4586
rect 1945 4528 1950 4584
rect 2006 4528 5446 4584
rect 5502 4528 5507 4584
rect 1945 4526 5507 4528
rect 1945 4523 2011 4526
rect 5441 4523 5507 4526
rect 3610 4384 3930 4385
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3930 4384
rect 3610 4319 3930 4320
rect 8944 4384 9264 4385
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 4319 9264 4320
rect 14277 4384 14597 4385
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 4319 14597 4320
rect 565 4178 631 4181
rect 3049 4178 3115 4181
rect 565 4176 3115 4178
rect 565 4120 570 4176
rect 626 4120 3054 4176
rect 3110 4120 3115 4176
rect 565 4118 3115 4120
rect 565 4115 631 4118
rect 3049 4115 3115 4118
rect 9489 4178 9555 4181
rect 12157 4178 12223 4181
rect 9489 4176 12223 4178
rect 9489 4120 9494 4176
rect 9550 4120 12162 4176
rect 12218 4120 12223 4176
rect 9489 4118 12223 4120
rect 9489 4115 9555 4118
rect 12157 4115 12223 4118
rect 6637 4042 6703 4045
rect 7833 4042 7899 4045
rect 6637 4040 7899 4042
rect 6637 3984 6642 4040
rect 6698 3984 7838 4040
rect 7894 3984 7899 4040
rect 6637 3982 7899 3984
rect 6637 3979 6703 3982
rect 7833 3979 7899 3982
rect 10041 4042 10107 4045
rect 12525 4042 12591 4045
rect 10041 4040 12591 4042
rect 10041 3984 10046 4040
rect 10102 3984 12530 4040
rect 12586 3984 12591 4040
rect 10041 3982 12591 3984
rect 10041 3979 10107 3982
rect 12525 3979 12591 3982
rect 8661 3906 8727 3909
rect 10409 3906 10475 3909
rect 8661 3904 10475 3906
rect 8661 3848 8666 3904
rect 8722 3848 10414 3904
rect 10470 3848 10475 3904
rect 8661 3846 10475 3848
rect 8661 3843 8727 3846
rect 10409 3843 10475 3846
rect 6277 3840 6597 3841
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 3775 6597 3776
rect 11610 3840 11930 3841
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 3775 11930 3776
rect 1853 3770 1919 3773
rect 9949 3770 10015 3773
rect 1853 3768 6194 3770
rect 1853 3712 1858 3768
rect 1914 3712 6194 3768
rect 1853 3710 6194 3712
rect 1853 3707 1919 3710
rect 2865 3634 2931 3637
rect 4613 3634 4679 3637
rect 2865 3632 4679 3634
rect 2865 3576 2870 3632
rect 2926 3576 4618 3632
rect 4674 3576 4679 3632
rect 2865 3574 4679 3576
rect 6134 3634 6194 3710
rect 6686 3768 10015 3770
rect 6686 3712 9954 3768
rect 10010 3712 10015 3768
rect 6686 3710 10015 3712
rect 6686 3634 6746 3710
rect 9949 3707 10015 3710
rect 6134 3574 6746 3634
rect 7649 3634 7715 3637
rect 9857 3634 9923 3637
rect 7649 3632 9923 3634
rect 7649 3576 7654 3632
rect 7710 3576 9862 3632
rect 9918 3576 9923 3632
rect 7649 3574 9923 3576
rect 2865 3571 2931 3574
rect 4613 3571 4679 3574
rect 7649 3571 7715 3574
rect 9857 3571 9923 3574
rect 0 3498 480 3528
rect 1577 3498 1643 3501
rect 0 3496 1643 3498
rect 0 3440 1582 3496
rect 1638 3440 1643 3496
rect 0 3438 1643 3440
rect 0 3408 480 3438
rect 1577 3435 1643 3438
rect 1761 3498 1827 3501
rect 4521 3498 4587 3501
rect 11421 3498 11487 3501
rect 1761 3496 4354 3498
rect 1761 3440 1766 3496
rect 1822 3440 4354 3496
rect 1761 3438 4354 3440
rect 1761 3435 1827 3438
rect 4294 3362 4354 3438
rect 4521 3496 11487 3498
rect 4521 3440 4526 3496
rect 4582 3440 11426 3496
rect 11482 3440 11487 3496
rect 4521 3438 11487 3440
rect 4521 3435 4587 3438
rect 11421 3435 11487 3438
rect 8753 3362 8819 3365
rect 4294 3360 8819 3362
rect 4294 3304 8758 3360
rect 8814 3304 8819 3360
rect 4294 3302 8819 3304
rect 8753 3299 8819 3302
rect 3610 3296 3930 3297
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3930 3296
rect 3610 3231 3930 3232
rect 8944 3296 9264 3297
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 8944 3231 9264 3232
rect 14277 3296 14597 3297
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 3231 14597 3232
rect 7925 3228 7991 3229
rect 7925 3226 7972 3228
rect 7880 3224 7972 3226
rect 7880 3168 7930 3224
rect 7880 3166 7972 3168
rect 7925 3164 7972 3166
rect 8036 3164 8042 3228
rect 10777 3226 10843 3229
rect 12433 3226 12499 3229
rect 10777 3224 12499 3226
rect 10777 3168 10782 3224
rect 10838 3168 12438 3224
rect 12494 3168 12499 3224
rect 10777 3166 12499 3168
rect 7925 3163 7991 3164
rect 10777 3163 10843 3166
rect 12433 3163 12499 3166
rect 2221 3090 2287 3093
rect 6637 3090 6703 3093
rect 2221 3088 6703 3090
rect 2221 3032 2226 3088
rect 2282 3032 6642 3088
rect 6698 3032 6703 3088
rect 2221 3030 6703 3032
rect 2221 3027 2287 3030
rect 6637 3027 6703 3030
rect 6913 3090 6979 3093
rect 9857 3090 9923 3093
rect 6913 3088 9923 3090
rect 6913 3032 6918 3088
rect 6974 3032 9862 3088
rect 9918 3032 9923 3088
rect 6913 3030 9923 3032
rect 6913 3027 6979 3030
rect 9857 3027 9923 3030
rect 4153 2954 4219 2957
rect 7097 2954 7163 2957
rect 4153 2952 7163 2954
rect 4153 2896 4158 2952
rect 4214 2896 7102 2952
rect 7158 2896 7163 2952
rect 4153 2894 7163 2896
rect 4153 2891 4219 2894
rect 7097 2891 7163 2894
rect 1945 2818 2011 2821
rect 5349 2818 5415 2821
rect 1945 2816 5415 2818
rect 1945 2760 1950 2816
rect 2006 2760 5354 2816
rect 5410 2760 5415 2816
rect 1945 2758 5415 2760
rect 1945 2755 2011 2758
rect 5349 2755 5415 2758
rect 7465 2818 7531 2821
rect 11329 2818 11395 2821
rect 7465 2816 11395 2818
rect 7465 2760 7470 2816
rect 7526 2760 11334 2816
rect 11390 2760 11395 2816
rect 7465 2758 11395 2760
rect 7465 2755 7531 2758
rect 11329 2755 11395 2758
rect 6277 2752 6597 2753
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2687 6597 2688
rect 11610 2752 11930 2753
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2687 11930 2688
rect 7465 2684 7531 2685
rect 7414 2620 7420 2684
rect 7484 2682 7531 2684
rect 7484 2680 7576 2682
rect 7526 2624 7576 2680
rect 7484 2622 7576 2624
rect 7484 2620 7531 2622
rect 7465 2619 7531 2620
rect 1669 2546 1735 2549
rect 5165 2546 5231 2549
rect 1669 2544 5231 2546
rect 1669 2488 1674 2544
rect 1730 2488 5170 2544
rect 5226 2488 5231 2544
rect 1669 2486 5231 2488
rect 1669 2483 1735 2486
rect 5165 2483 5231 2486
rect 7925 2546 7991 2549
rect 12893 2546 12959 2549
rect 7925 2544 12959 2546
rect 7925 2488 7930 2544
rect 7986 2488 12898 2544
rect 12954 2488 12959 2544
rect 7925 2486 12959 2488
rect 7925 2483 7991 2486
rect 12893 2483 12959 2486
rect 3610 2208 3930 2209
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3930 2208
rect 3610 2143 3930 2144
rect 8944 2208 9264 2209
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2143 9264 2144
rect 14277 2208 14597 2209
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2143 14597 2144
rect 5073 2002 5139 2005
rect 14181 2002 14247 2005
rect 5073 2000 14247 2002
rect 5073 1944 5078 2000
rect 5134 1944 14186 2000
rect 14242 1944 14247 2000
rect 5073 1942 14247 1944
rect 5073 1939 5139 1942
rect 14181 1939 14247 1942
rect 0 1186 480 1216
rect 1485 1186 1551 1189
rect 0 1184 1551 1186
rect 0 1128 1490 1184
rect 1546 1128 1551 1184
rect 0 1126 1551 1128
rect 0 1096 480 1126
rect 1485 1123 1551 1126
<< via3 >>
rect 6285 37564 6349 37568
rect 6285 37508 6289 37564
rect 6289 37508 6345 37564
rect 6345 37508 6349 37564
rect 6285 37504 6349 37508
rect 6365 37564 6429 37568
rect 6365 37508 6369 37564
rect 6369 37508 6425 37564
rect 6425 37508 6429 37564
rect 6365 37504 6429 37508
rect 6445 37564 6509 37568
rect 6445 37508 6449 37564
rect 6449 37508 6505 37564
rect 6505 37508 6509 37564
rect 6445 37504 6509 37508
rect 6525 37564 6589 37568
rect 6525 37508 6529 37564
rect 6529 37508 6585 37564
rect 6585 37508 6589 37564
rect 6525 37504 6589 37508
rect 11618 37564 11682 37568
rect 11618 37508 11622 37564
rect 11622 37508 11678 37564
rect 11678 37508 11682 37564
rect 11618 37504 11682 37508
rect 11698 37564 11762 37568
rect 11698 37508 11702 37564
rect 11702 37508 11758 37564
rect 11758 37508 11762 37564
rect 11698 37504 11762 37508
rect 11778 37564 11842 37568
rect 11778 37508 11782 37564
rect 11782 37508 11838 37564
rect 11838 37508 11842 37564
rect 11778 37504 11842 37508
rect 11858 37564 11922 37568
rect 11858 37508 11862 37564
rect 11862 37508 11918 37564
rect 11918 37508 11922 37564
rect 11858 37504 11922 37508
rect 3618 37020 3682 37024
rect 3618 36964 3622 37020
rect 3622 36964 3678 37020
rect 3678 36964 3682 37020
rect 3618 36960 3682 36964
rect 3698 37020 3762 37024
rect 3698 36964 3702 37020
rect 3702 36964 3758 37020
rect 3758 36964 3762 37020
rect 3698 36960 3762 36964
rect 3778 37020 3842 37024
rect 3778 36964 3782 37020
rect 3782 36964 3838 37020
rect 3838 36964 3842 37020
rect 3778 36960 3842 36964
rect 3858 37020 3922 37024
rect 3858 36964 3862 37020
rect 3862 36964 3918 37020
rect 3918 36964 3922 37020
rect 3858 36960 3922 36964
rect 8952 37020 9016 37024
rect 8952 36964 8956 37020
rect 8956 36964 9012 37020
rect 9012 36964 9016 37020
rect 8952 36960 9016 36964
rect 9032 37020 9096 37024
rect 9032 36964 9036 37020
rect 9036 36964 9092 37020
rect 9092 36964 9096 37020
rect 9032 36960 9096 36964
rect 9112 37020 9176 37024
rect 9112 36964 9116 37020
rect 9116 36964 9172 37020
rect 9172 36964 9176 37020
rect 9112 36960 9176 36964
rect 9192 37020 9256 37024
rect 9192 36964 9196 37020
rect 9196 36964 9252 37020
rect 9252 36964 9256 37020
rect 9192 36960 9256 36964
rect 14285 37020 14349 37024
rect 14285 36964 14289 37020
rect 14289 36964 14345 37020
rect 14345 36964 14349 37020
rect 14285 36960 14349 36964
rect 14365 37020 14429 37024
rect 14365 36964 14369 37020
rect 14369 36964 14425 37020
rect 14425 36964 14429 37020
rect 14365 36960 14429 36964
rect 14445 37020 14509 37024
rect 14445 36964 14449 37020
rect 14449 36964 14505 37020
rect 14505 36964 14509 37020
rect 14445 36960 14509 36964
rect 14525 37020 14589 37024
rect 14525 36964 14529 37020
rect 14529 36964 14585 37020
rect 14585 36964 14589 37020
rect 14525 36960 14589 36964
rect 6285 36476 6349 36480
rect 6285 36420 6289 36476
rect 6289 36420 6345 36476
rect 6345 36420 6349 36476
rect 6285 36416 6349 36420
rect 6365 36476 6429 36480
rect 6365 36420 6369 36476
rect 6369 36420 6425 36476
rect 6425 36420 6429 36476
rect 6365 36416 6429 36420
rect 6445 36476 6509 36480
rect 6445 36420 6449 36476
rect 6449 36420 6505 36476
rect 6505 36420 6509 36476
rect 6445 36416 6509 36420
rect 6525 36476 6589 36480
rect 6525 36420 6529 36476
rect 6529 36420 6585 36476
rect 6585 36420 6589 36476
rect 6525 36416 6589 36420
rect 11618 36476 11682 36480
rect 11618 36420 11622 36476
rect 11622 36420 11678 36476
rect 11678 36420 11682 36476
rect 11618 36416 11682 36420
rect 11698 36476 11762 36480
rect 11698 36420 11702 36476
rect 11702 36420 11758 36476
rect 11758 36420 11762 36476
rect 11698 36416 11762 36420
rect 11778 36476 11842 36480
rect 11778 36420 11782 36476
rect 11782 36420 11838 36476
rect 11838 36420 11842 36476
rect 11778 36416 11842 36420
rect 11858 36476 11922 36480
rect 11858 36420 11862 36476
rect 11862 36420 11918 36476
rect 11918 36420 11922 36476
rect 11858 36416 11922 36420
rect 3618 35932 3682 35936
rect 3618 35876 3622 35932
rect 3622 35876 3678 35932
rect 3678 35876 3682 35932
rect 3618 35872 3682 35876
rect 3698 35932 3762 35936
rect 3698 35876 3702 35932
rect 3702 35876 3758 35932
rect 3758 35876 3762 35932
rect 3698 35872 3762 35876
rect 3778 35932 3842 35936
rect 3778 35876 3782 35932
rect 3782 35876 3838 35932
rect 3838 35876 3842 35932
rect 3778 35872 3842 35876
rect 3858 35932 3922 35936
rect 3858 35876 3862 35932
rect 3862 35876 3918 35932
rect 3918 35876 3922 35932
rect 3858 35872 3922 35876
rect 8952 35932 9016 35936
rect 8952 35876 8956 35932
rect 8956 35876 9012 35932
rect 9012 35876 9016 35932
rect 8952 35872 9016 35876
rect 9032 35932 9096 35936
rect 9032 35876 9036 35932
rect 9036 35876 9092 35932
rect 9092 35876 9096 35932
rect 9032 35872 9096 35876
rect 9112 35932 9176 35936
rect 9112 35876 9116 35932
rect 9116 35876 9172 35932
rect 9172 35876 9176 35932
rect 9112 35872 9176 35876
rect 9192 35932 9256 35936
rect 9192 35876 9196 35932
rect 9196 35876 9252 35932
rect 9252 35876 9256 35932
rect 9192 35872 9256 35876
rect 14285 35932 14349 35936
rect 14285 35876 14289 35932
rect 14289 35876 14345 35932
rect 14345 35876 14349 35932
rect 14285 35872 14349 35876
rect 14365 35932 14429 35936
rect 14365 35876 14369 35932
rect 14369 35876 14425 35932
rect 14425 35876 14429 35932
rect 14365 35872 14429 35876
rect 14445 35932 14509 35936
rect 14445 35876 14449 35932
rect 14449 35876 14505 35932
rect 14505 35876 14509 35932
rect 14445 35872 14509 35876
rect 14525 35932 14589 35936
rect 14525 35876 14529 35932
rect 14529 35876 14585 35932
rect 14585 35876 14589 35932
rect 14525 35872 14589 35876
rect 6285 35388 6349 35392
rect 6285 35332 6289 35388
rect 6289 35332 6345 35388
rect 6345 35332 6349 35388
rect 6285 35328 6349 35332
rect 6365 35388 6429 35392
rect 6365 35332 6369 35388
rect 6369 35332 6425 35388
rect 6425 35332 6429 35388
rect 6365 35328 6429 35332
rect 6445 35388 6509 35392
rect 6445 35332 6449 35388
rect 6449 35332 6505 35388
rect 6505 35332 6509 35388
rect 6445 35328 6509 35332
rect 6525 35388 6589 35392
rect 6525 35332 6529 35388
rect 6529 35332 6585 35388
rect 6585 35332 6589 35388
rect 6525 35328 6589 35332
rect 11618 35388 11682 35392
rect 11618 35332 11622 35388
rect 11622 35332 11678 35388
rect 11678 35332 11682 35388
rect 11618 35328 11682 35332
rect 11698 35388 11762 35392
rect 11698 35332 11702 35388
rect 11702 35332 11758 35388
rect 11758 35332 11762 35388
rect 11698 35328 11762 35332
rect 11778 35388 11842 35392
rect 11778 35332 11782 35388
rect 11782 35332 11838 35388
rect 11838 35332 11842 35388
rect 11778 35328 11842 35332
rect 11858 35388 11922 35392
rect 11858 35332 11862 35388
rect 11862 35332 11918 35388
rect 11918 35332 11922 35388
rect 11858 35328 11922 35332
rect 3618 34844 3682 34848
rect 3618 34788 3622 34844
rect 3622 34788 3678 34844
rect 3678 34788 3682 34844
rect 3618 34784 3682 34788
rect 3698 34844 3762 34848
rect 3698 34788 3702 34844
rect 3702 34788 3758 34844
rect 3758 34788 3762 34844
rect 3698 34784 3762 34788
rect 3778 34844 3842 34848
rect 3778 34788 3782 34844
rect 3782 34788 3838 34844
rect 3838 34788 3842 34844
rect 3778 34784 3842 34788
rect 3858 34844 3922 34848
rect 3858 34788 3862 34844
rect 3862 34788 3918 34844
rect 3918 34788 3922 34844
rect 3858 34784 3922 34788
rect 8952 34844 9016 34848
rect 8952 34788 8956 34844
rect 8956 34788 9012 34844
rect 9012 34788 9016 34844
rect 8952 34784 9016 34788
rect 9032 34844 9096 34848
rect 9032 34788 9036 34844
rect 9036 34788 9092 34844
rect 9092 34788 9096 34844
rect 9032 34784 9096 34788
rect 9112 34844 9176 34848
rect 9112 34788 9116 34844
rect 9116 34788 9172 34844
rect 9172 34788 9176 34844
rect 9112 34784 9176 34788
rect 9192 34844 9256 34848
rect 9192 34788 9196 34844
rect 9196 34788 9252 34844
rect 9252 34788 9256 34844
rect 9192 34784 9256 34788
rect 14285 34844 14349 34848
rect 14285 34788 14289 34844
rect 14289 34788 14345 34844
rect 14345 34788 14349 34844
rect 14285 34784 14349 34788
rect 14365 34844 14429 34848
rect 14365 34788 14369 34844
rect 14369 34788 14425 34844
rect 14425 34788 14429 34844
rect 14365 34784 14429 34788
rect 14445 34844 14509 34848
rect 14445 34788 14449 34844
rect 14449 34788 14505 34844
rect 14505 34788 14509 34844
rect 14445 34784 14509 34788
rect 14525 34844 14589 34848
rect 14525 34788 14529 34844
rect 14529 34788 14585 34844
rect 14585 34788 14589 34844
rect 14525 34784 14589 34788
rect 6285 34300 6349 34304
rect 6285 34244 6289 34300
rect 6289 34244 6345 34300
rect 6345 34244 6349 34300
rect 6285 34240 6349 34244
rect 6365 34300 6429 34304
rect 6365 34244 6369 34300
rect 6369 34244 6425 34300
rect 6425 34244 6429 34300
rect 6365 34240 6429 34244
rect 6445 34300 6509 34304
rect 6445 34244 6449 34300
rect 6449 34244 6505 34300
rect 6505 34244 6509 34300
rect 6445 34240 6509 34244
rect 6525 34300 6589 34304
rect 6525 34244 6529 34300
rect 6529 34244 6585 34300
rect 6585 34244 6589 34300
rect 6525 34240 6589 34244
rect 11618 34300 11682 34304
rect 11618 34244 11622 34300
rect 11622 34244 11678 34300
rect 11678 34244 11682 34300
rect 11618 34240 11682 34244
rect 11698 34300 11762 34304
rect 11698 34244 11702 34300
rect 11702 34244 11758 34300
rect 11758 34244 11762 34300
rect 11698 34240 11762 34244
rect 11778 34300 11842 34304
rect 11778 34244 11782 34300
rect 11782 34244 11838 34300
rect 11838 34244 11842 34300
rect 11778 34240 11842 34244
rect 11858 34300 11922 34304
rect 11858 34244 11862 34300
rect 11862 34244 11918 34300
rect 11918 34244 11922 34300
rect 11858 34240 11922 34244
rect 3618 33756 3682 33760
rect 3618 33700 3622 33756
rect 3622 33700 3678 33756
rect 3678 33700 3682 33756
rect 3618 33696 3682 33700
rect 3698 33756 3762 33760
rect 3698 33700 3702 33756
rect 3702 33700 3758 33756
rect 3758 33700 3762 33756
rect 3698 33696 3762 33700
rect 3778 33756 3842 33760
rect 3778 33700 3782 33756
rect 3782 33700 3838 33756
rect 3838 33700 3842 33756
rect 3778 33696 3842 33700
rect 3858 33756 3922 33760
rect 3858 33700 3862 33756
rect 3862 33700 3918 33756
rect 3918 33700 3922 33756
rect 3858 33696 3922 33700
rect 8952 33756 9016 33760
rect 8952 33700 8956 33756
rect 8956 33700 9012 33756
rect 9012 33700 9016 33756
rect 8952 33696 9016 33700
rect 9032 33756 9096 33760
rect 9032 33700 9036 33756
rect 9036 33700 9092 33756
rect 9092 33700 9096 33756
rect 9032 33696 9096 33700
rect 9112 33756 9176 33760
rect 9112 33700 9116 33756
rect 9116 33700 9172 33756
rect 9172 33700 9176 33756
rect 9112 33696 9176 33700
rect 9192 33756 9256 33760
rect 9192 33700 9196 33756
rect 9196 33700 9252 33756
rect 9252 33700 9256 33756
rect 9192 33696 9256 33700
rect 14285 33756 14349 33760
rect 14285 33700 14289 33756
rect 14289 33700 14345 33756
rect 14345 33700 14349 33756
rect 14285 33696 14349 33700
rect 14365 33756 14429 33760
rect 14365 33700 14369 33756
rect 14369 33700 14425 33756
rect 14425 33700 14429 33756
rect 14365 33696 14429 33700
rect 14445 33756 14509 33760
rect 14445 33700 14449 33756
rect 14449 33700 14505 33756
rect 14505 33700 14509 33756
rect 14445 33696 14509 33700
rect 14525 33756 14589 33760
rect 14525 33700 14529 33756
rect 14529 33700 14585 33756
rect 14585 33700 14589 33756
rect 14525 33696 14589 33700
rect 6285 33212 6349 33216
rect 6285 33156 6289 33212
rect 6289 33156 6345 33212
rect 6345 33156 6349 33212
rect 6285 33152 6349 33156
rect 6365 33212 6429 33216
rect 6365 33156 6369 33212
rect 6369 33156 6425 33212
rect 6425 33156 6429 33212
rect 6365 33152 6429 33156
rect 6445 33212 6509 33216
rect 6445 33156 6449 33212
rect 6449 33156 6505 33212
rect 6505 33156 6509 33212
rect 6445 33152 6509 33156
rect 6525 33212 6589 33216
rect 6525 33156 6529 33212
rect 6529 33156 6585 33212
rect 6585 33156 6589 33212
rect 6525 33152 6589 33156
rect 11618 33212 11682 33216
rect 11618 33156 11622 33212
rect 11622 33156 11678 33212
rect 11678 33156 11682 33212
rect 11618 33152 11682 33156
rect 11698 33212 11762 33216
rect 11698 33156 11702 33212
rect 11702 33156 11758 33212
rect 11758 33156 11762 33212
rect 11698 33152 11762 33156
rect 11778 33212 11842 33216
rect 11778 33156 11782 33212
rect 11782 33156 11838 33212
rect 11838 33156 11842 33212
rect 11778 33152 11842 33156
rect 11858 33212 11922 33216
rect 11858 33156 11862 33212
rect 11862 33156 11918 33212
rect 11918 33156 11922 33212
rect 11858 33152 11922 33156
rect 3618 32668 3682 32672
rect 3618 32612 3622 32668
rect 3622 32612 3678 32668
rect 3678 32612 3682 32668
rect 3618 32608 3682 32612
rect 3698 32668 3762 32672
rect 3698 32612 3702 32668
rect 3702 32612 3758 32668
rect 3758 32612 3762 32668
rect 3698 32608 3762 32612
rect 3778 32668 3842 32672
rect 3778 32612 3782 32668
rect 3782 32612 3838 32668
rect 3838 32612 3842 32668
rect 3778 32608 3842 32612
rect 3858 32668 3922 32672
rect 3858 32612 3862 32668
rect 3862 32612 3918 32668
rect 3918 32612 3922 32668
rect 3858 32608 3922 32612
rect 8952 32668 9016 32672
rect 8952 32612 8956 32668
rect 8956 32612 9012 32668
rect 9012 32612 9016 32668
rect 8952 32608 9016 32612
rect 9032 32668 9096 32672
rect 9032 32612 9036 32668
rect 9036 32612 9092 32668
rect 9092 32612 9096 32668
rect 9032 32608 9096 32612
rect 9112 32668 9176 32672
rect 9112 32612 9116 32668
rect 9116 32612 9172 32668
rect 9172 32612 9176 32668
rect 9112 32608 9176 32612
rect 9192 32668 9256 32672
rect 9192 32612 9196 32668
rect 9196 32612 9252 32668
rect 9252 32612 9256 32668
rect 9192 32608 9256 32612
rect 14285 32668 14349 32672
rect 14285 32612 14289 32668
rect 14289 32612 14345 32668
rect 14345 32612 14349 32668
rect 14285 32608 14349 32612
rect 14365 32668 14429 32672
rect 14365 32612 14369 32668
rect 14369 32612 14425 32668
rect 14425 32612 14429 32668
rect 14365 32608 14429 32612
rect 14445 32668 14509 32672
rect 14445 32612 14449 32668
rect 14449 32612 14505 32668
rect 14505 32612 14509 32668
rect 14445 32608 14509 32612
rect 14525 32668 14589 32672
rect 14525 32612 14529 32668
rect 14529 32612 14585 32668
rect 14585 32612 14589 32668
rect 14525 32608 14589 32612
rect 6285 32124 6349 32128
rect 6285 32068 6289 32124
rect 6289 32068 6345 32124
rect 6345 32068 6349 32124
rect 6285 32064 6349 32068
rect 6365 32124 6429 32128
rect 6365 32068 6369 32124
rect 6369 32068 6425 32124
rect 6425 32068 6429 32124
rect 6365 32064 6429 32068
rect 6445 32124 6509 32128
rect 6445 32068 6449 32124
rect 6449 32068 6505 32124
rect 6505 32068 6509 32124
rect 6445 32064 6509 32068
rect 6525 32124 6589 32128
rect 6525 32068 6529 32124
rect 6529 32068 6585 32124
rect 6585 32068 6589 32124
rect 6525 32064 6589 32068
rect 11618 32124 11682 32128
rect 11618 32068 11622 32124
rect 11622 32068 11678 32124
rect 11678 32068 11682 32124
rect 11618 32064 11682 32068
rect 11698 32124 11762 32128
rect 11698 32068 11702 32124
rect 11702 32068 11758 32124
rect 11758 32068 11762 32124
rect 11698 32064 11762 32068
rect 11778 32124 11842 32128
rect 11778 32068 11782 32124
rect 11782 32068 11838 32124
rect 11838 32068 11842 32124
rect 11778 32064 11842 32068
rect 11858 32124 11922 32128
rect 11858 32068 11862 32124
rect 11862 32068 11918 32124
rect 11918 32068 11922 32124
rect 11858 32064 11922 32068
rect 3618 31580 3682 31584
rect 3618 31524 3622 31580
rect 3622 31524 3678 31580
rect 3678 31524 3682 31580
rect 3618 31520 3682 31524
rect 3698 31580 3762 31584
rect 3698 31524 3702 31580
rect 3702 31524 3758 31580
rect 3758 31524 3762 31580
rect 3698 31520 3762 31524
rect 3778 31580 3842 31584
rect 3778 31524 3782 31580
rect 3782 31524 3838 31580
rect 3838 31524 3842 31580
rect 3778 31520 3842 31524
rect 3858 31580 3922 31584
rect 3858 31524 3862 31580
rect 3862 31524 3918 31580
rect 3918 31524 3922 31580
rect 3858 31520 3922 31524
rect 8952 31580 9016 31584
rect 8952 31524 8956 31580
rect 8956 31524 9012 31580
rect 9012 31524 9016 31580
rect 8952 31520 9016 31524
rect 9032 31580 9096 31584
rect 9032 31524 9036 31580
rect 9036 31524 9092 31580
rect 9092 31524 9096 31580
rect 9032 31520 9096 31524
rect 9112 31580 9176 31584
rect 9112 31524 9116 31580
rect 9116 31524 9172 31580
rect 9172 31524 9176 31580
rect 9112 31520 9176 31524
rect 9192 31580 9256 31584
rect 9192 31524 9196 31580
rect 9196 31524 9252 31580
rect 9252 31524 9256 31580
rect 9192 31520 9256 31524
rect 14285 31580 14349 31584
rect 14285 31524 14289 31580
rect 14289 31524 14345 31580
rect 14345 31524 14349 31580
rect 14285 31520 14349 31524
rect 14365 31580 14429 31584
rect 14365 31524 14369 31580
rect 14369 31524 14425 31580
rect 14425 31524 14429 31580
rect 14365 31520 14429 31524
rect 14445 31580 14509 31584
rect 14445 31524 14449 31580
rect 14449 31524 14505 31580
rect 14505 31524 14509 31580
rect 14445 31520 14509 31524
rect 14525 31580 14589 31584
rect 14525 31524 14529 31580
rect 14529 31524 14585 31580
rect 14585 31524 14589 31580
rect 14525 31520 14589 31524
rect 6285 31036 6349 31040
rect 6285 30980 6289 31036
rect 6289 30980 6345 31036
rect 6345 30980 6349 31036
rect 6285 30976 6349 30980
rect 6365 31036 6429 31040
rect 6365 30980 6369 31036
rect 6369 30980 6425 31036
rect 6425 30980 6429 31036
rect 6365 30976 6429 30980
rect 6445 31036 6509 31040
rect 6445 30980 6449 31036
rect 6449 30980 6505 31036
rect 6505 30980 6509 31036
rect 6445 30976 6509 30980
rect 6525 31036 6589 31040
rect 6525 30980 6529 31036
rect 6529 30980 6585 31036
rect 6585 30980 6589 31036
rect 6525 30976 6589 30980
rect 11618 31036 11682 31040
rect 11618 30980 11622 31036
rect 11622 30980 11678 31036
rect 11678 30980 11682 31036
rect 11618 30976 11682 30980
rect 11698 31036 11762 31040
rect 11698 30980 11702 31036
rect 11702 30980 11758 31036
rect 11758 30980 11762 31036
rect 11698 30976 11762 30980
rect 11778 31036 11842 31040
rect 11778 30980 11782 31036
rect 11782 30980 11838 31036
rect 11838 30980 11842 31036
rect 11778 30976 11842 30980
rect 11858 31036 11922 31040
rect 11858 30980 11862 31036
rect 11862 30980 11918 31036
rect 11918 30980 11922 31036
rect 11858 30976 11922 30980
rect 3618 30492 3682 30496
rect 3618 30436 3622 30492
rect 3622 30436 3678 30492
rect 3678 30436 3682 30492
rect 3618 30432 3682 30436
rect 3698 30492 3762 30496
rect 3698 30436 3702 30492
rect 3702 30436 3758 30492
rect 3758 30436 3762 30492
rect 3698 30432 3762 30436
rect 3778 30492 3842 30496
rect 3778 30436 3782 30492
rect 3782 30436 3838 30492
rect 3838 30436 3842 30492
rect 3778 30432 3842 30436
rect 3858 30492 3922 30496
rect 3858 30436 3862 30492
rect 3862 30436 3918 30492
rect 3918 30436 3922 30492
rect 3858 30432 3922 30436
rect 8952 30492 9016 30496
rect 8952 30436 8956 30492
rect 8956 30436 9012 30492
rect 9012 30436 9016 30492
rect 8952 30432 9016 30436
rect 9032 30492 9096 30496
rect 9032 30436 9036 30492
rect 9036 30436 9092 30492
rect 9092 30436 9096 30492
rect 9032 30432 9096 30436
rect 9112 30492 9176 30496
rect 9112 30436 9116 30492
rect 9116 30436 9172 30492
rect 9172 30436 9176 30492
rect 9112 30432 9176 30436
rect 9192 30492 9256 30496
rect 9192 30436 9196 30492
rect 9196 30436 9252 30492
rect 9252 30436 9256 30492
rect 9192 30432 9256 30436
rect 14285 30492 14349 30496
rect 14285 30436 14289 30492
rect 14289 30436 14345 30492
rect 14345 30436 14349 30492
rect 14285 30432 14349 30436
rect 14365 30492 14429 30496
rect 14365 30436 14369 30492
rect 14369 30436 14425 30492
rect 14425 30436 14429 30492
rect 14365 30432 14429 30436
rect 14445 30492 14509 30496
rect 14445 30436 14449 30492
rect 14449 30436 14505 30492
rect 14505 30436 14509 30492
rect 14445 30432 14509 30436
rect 14525 30492 14589 30496
rect 14525 30436 14529 30492
rect 14529 30436 14585 30492
rect 14585 30436 14589 30492
rect 14525 30432 14589 30436
rect 6285 29948 6349 29952
rect 6285 29892 6289 29948
rect 6289 29892 6345 29948
rect 6345 29892 6349 29948
rect 6285 29888 6349 29892
rect 6365 29948 6429 29952
rect 6365 29892 6369 29948
rect 6369 29892 6425 29948
rect 6425 29892 6429 29948
rect 6365 29888 6429 29892
rect 6445 29948 6509 29952
rect 6445 29892 6449 29948
rect 6449 29892 6505 29948
rect 6505 29892 6509 29948
rect 6445 29888 6509 29892
rect 6525 29948 6589 29952
rect 6525 29892 6529 29948
rect 6529 29892 6585 29948
rect 6585 29892 6589 29948
rect 6525 29888 6589 29892
rect 11618 29948 11682 29952
rect 11618 29892 11622 29948
rect 11622 29892 11678 29948
rect 11678 29892 11682 29948
rect 11618 29888 11682 29892
rect 11698 29948 11762 29952
rect 11698 29892 11702 29948
rect 11702 29892 11758 29948
rect 11758 29892 11762 29948
rect 11698 29888 11762 29892
rect 11778 29948 11842 29952
rect 11778 29892 11782 29948
rect 11782 29892 11838 29948
rect 11838 29892 11842 29948
rect 11778 29888 11842 29892
rect 11858 29948 11922 29952
rect 11858 29892 11862 29948
rect 11862 29892 11918 29948
rect 11918 29892 11922 29948
rect 11858 29888 11922 29892
rect 3618 29404 3682 29408
rect 3618 29348 3622 29404
rect 3622 29348 3678 29404
rect 3678 29348 3682 29404
rect 3618 29344 3682 29348
rect 3698 29404 3762 29408
rect 3698 29348 3702 29404
rect 3702 29348 3758 29404
rect 3758 29348 3762 29404
rect 3698 29344 3762 29348
rect 3778 29404 3842 29408
rect 3778 29348 3782 29404
rect 3782 29348 3838 29404
rect 3838 29348 3842 29404
rect 3778 29344 3842 29348
rect 3858 29404 3922 29408
rect 3858 29348 3862 29404
rect 3862 29348 3918 29404
rect 3918 29348 3922 29404
rect 3858 29344 3922 29348
rect 8952 29404 9016 29408
rect 8952 29348 8956 29404
rect 8956 29348 9012 29404
rect 9012 29348 9016 29404
rect 8952 29344 9016 29348
rect 9032 29404 9096 29408
rect 9032 29348 9036 29404
rect 9036 29348 9092 29404
rect 9092 29348 9096 29404
rect 9032 29344 9096 29348
rect 9112 29404 9176 29408
rect 9112 29348 9116 29404
rect 9116 29348 9172 29404
rect 9172 29348 9176 29404
rect 9112 29344 9176 29348
rect 9192 29404 9256 29408
rect 9192 29348 9196 29404
rect 9196 29348 9252 29404
rect 9252 29348 9256 29404
rect 9192 29344 9256 29348
rect 14285 29404 14349 29408
rect 14285 29348 14289 29404
rect 14289 29348 14345 29404
rect 14345 29348 14349 29404
rect 14285 29344 14349 29348
rect 14365 29404 14429 29408
rect 14365 29348 14369 29404
rect 14369 29348 14425 29404
rect 14425 29348 14429 29404
rect 14365 29344 14429 29348
rect 14445 29404 14509 29408
rect 14445 29348 14449 29404
rect 14449 29348 14505 29404
rect 14505 29348 14509 29404
rect 14445 29344 14509 29348
rect 14525 29404 14589 29408
rect 14525 29348 14529 29404
rect 14529 29348 14585 29404
rect 14585 29348 14589 29404
rect 14525 29344 14589 29348
rect 6285 28860 6349 28864
rect 6285 28804 6289 28860
rect 6289 28804 6345 28860
rect 6345 28804 6349 28860
rect 6285 28800 6349 28804
rect 6365 28860 6429 28864
rect 6365 28804 6369 28860
rect 6369 28804 6425 28860
rect 6425 28804 6429 28860
rect 6365 28800 6429 28804
rect 6445 28860 6509 28864
rect 6445 28804 6449 28860
rect 6449 28804 6505 28860
rect 6505 28804 6509 28860
rect 6445 28800 6509 28804
rect 6525 28860 6589 28864
rect 6525 28804 6529 28860
rect 6529 28804 6585 28860
rect 6585 28804 6589 28860
rect 6525 28800 6589 28804
rect 11618 28860 11682 28864
rect 11618 28804 11622 28860
rect 11622 28804 11678 28860
rect 11678 28804 11682 28860
rect 11618 28800 11682 28804
rect 11698 28860 11762 28864
rect 11698 28804 11702 28860
rect 11702 28804 11758 28860
rect 11758 28804 11762 28860
rect 11698 28800 11762 28804
rect 11778 28860 11842 28864
rect 11778 28804 11782 28860
rect 11782 28804 11838 28860
rect 11838 28804 11842 28860
rect 11778 28800 11842 28804
rect 11858 28860 11922 28864
rect 11858 28804 11862 28860
rect 11862 28804 11918 28860
rect 11918 28804 11922 28860
rect 11858 28800 11922 28804
rect 9444 28792 9508 28796
rect 9444 28736 9458 28792
rect 9458 28736 9508 28792
rect 9444 28732 9508 28736
rect 3618 28316 3682 28320
rect 3618 28260 3622 28316
rect 3622 28260 3678 28316
rect 3678 28260 3682 28316
rect 3618 28256 3682 28260
rect 3698 28316 3762 28320
rect 3698 28260 3702 28316
rect 3702 28260 3758 28316
rect 3758 28260 3762 28316
rect 3698 28256 3762 28260
rect 3778 28316 3842 28320
rect 3778 28260 3782 28316
rect 3782 28260 3838 28316
rect 3838 28260 3842 28316
rect 3778 28256 3842 28260
rect 3858 28316 3922 28320
rect 3858 28260 3862 28316
rect 3862 28260 3918 28316
rect 3918 28260 3922 28316
rect 3858 28256 3922 28260
rect 8952 28316 9016 28320
rect 8952 28260 8956 28316
rect 8956 28260 9012 28316
rect 9012 28260 9016 28316
rect 8952 28256 9016 28260
rect 9032 28316 9096 28320
rect 9032 28260 9036 28316
rect 9036 28260 9092 28316
rect 9092 28260 9096 28316
rect 9032 28256 9096 28260
rect 9112 28316 9176 28320
rect 9112 28260 9116 28316
rect 9116 28260 9172 28316
rect 9172 28260 9176 28316
rect 9112 28256 9176 28260
rect 9192 28316 9256 28320
rect 9192 28260 9196 28316
rect 9196 28260 9252 28316
rect 9252 28260 9256 28316
rect 9192 28256 9256 28260
rect 14285 28316 14349 28320
rect 14285 28260 14289 28316
rect 14289 28260 14345 28316
rect 14345 28260 14349 28316
rect 14285 28256 14349 28260
rect 14365 28316 14429 28320
rect 14365 28260 14369 28316
rect 14369 28260 14425 28316
rect 14425 28260 14429 28316
rect 14365 28256 14429 28260
rect 14445 28316 14509 28320
rect 14445 28260 14449 28316
rect 14449 28260 14505 28316
rect 14505 28260 14509 28316
rect 14445 28256 14509 28260
rect 14525 28316 14589 28320
rect 14525 28260 14529 28316
rect 14529 28260 14585 28316
rect 14585 28260 14589 28316
rect 14525 28256 14589 28260
rect 6285 27772 6349 27776
rect 6285 27716 6289 27772
rect 6289 27716 6345 27772
rect 6345 27716 6349 27772
rect 6285 27712 6349 27716
rect 6365 27772 6429 27776
rect 6365 27716 6369 27772
rect 6369 27716 6425 27772
rect 6425 27716 6429 27772
rect 6365 27712 6429 27716
rect 6445 27772 6509 27776
rect 6445 27716 6449 27772
rect 6449 27716 6505 27772
rect 6505 27716 6509 27772
rect 6445 27712 6509 27716
rect 6525 27772 6589 27776
rect 6525 27716 6529 27772
rect 6529 27716 6585 27772
rect 6585 27716 6589 27772
rect 6525 27712 6589 27716
rect 11618 27772 11682 27776
rect 11618 27716 11622 27772
rect 11622 27716 11678 27772
rect 11678 27716 11682 27772
rect 11618 27712 11682 27716
rect 11698 27772 11762 27776
rect 11698 27716 11702 27772
rect 11702 27716 11758 27772
rect 11758 27716 11762 27772
rect 11698 27712 11762 27716
rect 11778 27772 11842 27776
rect 11778 27716 11782 27772
rect 11782 27716 11838 27772
rect 11838 27716 11842 27772
rect 11778 27712 11842 27716
rect 11858 27772 11922 27776
rect 11858 27716 11862 27772
rect 11862 27716 11918 27772
rect 11918 27716 11922 27772
rect 11858 27712 11922 27716
rect 12020 27704 12084 27708
rect 12020 27648 12070 27704
rect 12070 27648 12084 27704
rect 12020 27644 12084 27648
rect 3618 27228 3682 27232
rect 3618 27172 3622 27228
rect 3622 27172 3678 27228
rect 3678 27172 3682 27228
rect 3618 27168 3682 27172
rect 3698 27228 3762 27232
rect 3698 27172 3702 27228
rect 3702 27172 3758 27228
rect 3758 27172 3762 27228
rect 3698 27168 3762 27172
rect 3778 27228 3842 27232
rect 3778 27172 3782 27228
rect 3782 27172 3838 27228
rect 3838 27172 3842 27228
rect 3778 27168 3842 27172
rect 3858 27228 3922 27232
rect 3858 27172 3862 27228
rect 3862 27172 3918 27228
rect 3918 27172 3922 27228
rect 3858 27168 3922 27172
rect 8952 27228 9016 27232
rect 8952 27172 8956 27228
rect 8956 27172 9012 27228
rect 9012 27172 9016 27228
rect 8952 27168 9016 27172
rect 9032 27228 9096 27232
rect 9032 27172 9036 27228
rect 9036 27172 9092 27228
rect 9092 27172 9096 27228
rect 9032 27168 9096 27172
rect 9112 27228 9176 27232
rect 9112 27172 9116 27228
rect 9116 27172 9172 27228
rect 9172 27172 9176 27228
rect 9112 27168 9176 27172
rect 9192 27228 9256 27232
rect 9192 27172 9196 27228
rect 9196 27172 9252 27228
rect 9252 27172 9256 27228
rect 9192 27168 9256 27172
rect 14285 27228 14349 27232
rect 14285 27172 14289 27228
rect 14289 27172 14345 27228
rect 14345 27172 14349 27228
rect 14285 27168 14349 27172
rect 14365 27228 14429 27232
rect 14365 27172 14369 27228
rect 14369 27172 14425 27228
rect 14425 27172 14429 27228
rect 14365 27168 14429 27172
rect 14445 27228 14509 27232
rect 14445 27172 14449 27228
rect 14449 27172 14505 27228
rect 14505 27172 14509 27228
rect 14445 27168 14509 27172
rect 14525 27228 14589 27232
rect 14525 27172 14529 27228
rect 14529 27172 14585 27228
rect 14585 27172 14589 27228
rect 14525 27168 14589 27172
rect 6285 26684 6349 26688
rect 6285 26628 6289 26684
rect 6289 26628 6345 26684
rect 6345 26628 6349 26684
rect 6285 26624 6349 26628
rect 6365 26684 6429 26688
rect 6365 26628 6369 26684
rect 6369 26628 6425 26684
rect 6425 26628 6429 26684
rect 6365 26624 6429 26628
rect 6445 26684 6509 26688
rect 6445 26628 6449 26684
rect 6449 26628 6505 26684
rect 6505 26628 6509 26684
rect 6445 26624 6509 26628
rect 6525 26684 6589 26688
rect 6525 26628 6529 26684
rect 6529 26628 6585 26684
rect 6585 26628 6589 26684
rect 6525 26624 6589 26628
rect 11618 26684 11682 26688
rect 11618 26628 11622 26684
rect 11622 26628 11678 26684
rect 11678 26628 11682 26684
rect 11618 26624 11682 26628
rect 11698 26684 11762 26688
rect 11698 26628 11702 26684
rect 11702 26628 11758 26684
rect 11758 26628 11762 26684
rect 11698 26624 11762 26628
rect 11778 26684 11842 26688
rect 11778 26628 11782 26684
rect 11782 26628 11838 26684
rect 11838 26628 11842 26684
rect 11778 26624 11842 26628
rect 11858 26684 11922 26688
rect 11858 26628 11862 26684
rect 11862 26628 11918 26684
rect 11918 26628 11922 26684
rect 11858 26624 11922 26628
rect 3618 26140 3682 26144
rect 3618 26084 3622 26140
rect 3622 26084 3678 26140
rect 3678 26084 3682 26140
rect 3618 26080 3682 26084
rect 3698 26140 3762 26144
rect 3698 26084 3702 26140
rect 3702 26084 3758 26140
rect 3758 26084 3762 26140
rect 3698 26080 3762 26084
rect 3778 26140 3842 26144
rect 3778 26084 3782 26140
rect 3782 26084 3838 26140
rect 3838 26084 3842 26140
rect 3778 26080 3842 26084
rect 3858 26140 3922 26144
rect 3858 26084 3862 26140
rect 3862 26084 3918 26140
rect 3918 26084 3922 26140
rect 3858 26080 3922 26084
rect 8952 26140 9016 26144
rect 8952 26084 8956 26140
rect 8956 26084 9012 26140
rect 9012 26084 9016 26140
rect 8952 26080 9016 26084
rect 9032 26140 9096 26144
rect 9032 26084 9036 26140
rect 9036 26084 9092 26140
rect 9092 26084 9096 26140
rect 9032 26080 9096 26084
rect 9112 26140 9176 26144
rect 9112 26084 9116 26140
rect 9116 26084 9172 26140
rect 9172 26084 9176 26140
rect 9112 26080 9176 26084
rect 9192 26140 9256 26144
rect 9192 26084 9196 26140
rect 9196 26084 9252 26140
rect 9252 26084 9256 26140
rect 9192 26080 9256 26084
rect 14285 26140 14349 26144
rect 14285 26084 14289 26140
rect 14289 26084 14345 26140
rect 14345 26084 14349 26140
rect 14285 26080 14349 26084
rect 14365 26140 14429 26144
rect 14365 26084 14369 26140
rect 14369 26084 14425 26140
rect 14425 26084 14429 26140
rect 14365 26080 14429 26084
rect 14445 26140 14509 26144
rect 14445 26084 14449 26140
rect 14449 26084 14505 26140
rect 14505 26084 14509 26140
rect 14445 26080 14509 26084
rect 14525 26140 14589 26144
rect 14525 26084 14529 26140
rect 14529 26084 14585 26140
rect 14585 26084 14589 26140
rect 14525 26080 14589 26084
rect 6285 25596 6349 25600
rect 6285 25540 6289 25596
rect 6289 25540 6345 25596
rect 6345 25540 6349 25596
rect 6285 25536 6349 25540
rect 6365 25596 6429 25600
rect 6365 25540 6369 25596
rect 6369 25540 6425 25596
rect 6425 25540 6429 25596
rect 6365 25536 6429 25540
rect 6445 25596 6509 25600
rect 6445 25540 6449 25596
rect 6449 25540 6505 25596
rect 6505 25540 6509 25596
rect 6445 25536 6509 25540
rect 6525 25596 6589 25600
rect 6525 25540 6529 25596
rect 6529 25540 6585 25596
rect 6585 25540 6589 25596
rect 6525 25536 6589 25540
rect 11618 25596 11682 25600
rect 11618 25540 11622 25596
rect 11622 25540 11678 25596
rect 11678 25540 11682 25596
rect 11618 25536 11682 25540
rect 11698 25596 11762 25600
rect 11698 25540 11702 25596
rect 11702 25540 11758 25596
rect 11758 25540 11762 25596
rect 11698 25536 11762 25540
rect 11778 25596 11842 25600
rect 11778 25540 11782 25596
rect 11782 25540 11838 25596
rect 11838 25540 11842 25596
rect 11778 25536 11842 25540
rect 11858 25596 11922 25600
rect 11858 25540 11862 25596
rect 11862 25540 11918 25596
rect 11918 25540 11922 25596
rect 11858 25536 11922 25540
rect 3618 25052 3682 25056
rect 3618 24996 3622 25052
rect 3622 24996 3678 25052
rect 3678 24996 3682 25052
rect 3618 24992 3682 24996
rect 3698 25052 3762 25056
rect 3698 24996 3702 25052
rect 3702 24996 3758 25052
rect 3758 24996 3762 25052
rect 3698 24992 3762 24996
rect 3778 25052 3842 25056
rect 3778 24996 3782 25052
rect 3782 24996 3838 25052
rect 3838 24996 3842 25052
rect 3778 24992 3842 24996
rect 3858 25052 3922 25056
rect 3858 24996 3862 25052
rect 3862 24996 3918 25052
rect 3918 24996 3922 25052
rect 3858 24992 3922 24996
rect 8952 25052 9016 25056
rect 8952 24996 8956 25052
rect 8956 24996 9012 25052
rect 9012 24996 9016 25052
rect 8952 24992 9016 24996
rect 9032 25052 9096 25056
rect 9032 24996 9036 25052
rect 9036 24996 9092 25052
rect 9092 24996 9096 25052
rect 9032 24992 9096 24996
rect 9112 25052 9176 25056
rect 9112 24996 9116 25052
rect 9116 24996 9172 25052
rect 9172 24996 9176 25052
rect 9112 24992 9176 24996
rect 9192 25052 9256 25056
rect 9192 24996 9196 25052
rect 9196 24996 9252 25052
rect 9252 24996 9256 25052
rect 9192 24992 9256 24996
rect 14285 25052 14349 25056
rect 14285 24996 14289 25052
rect 14289 24996 14345 25052
rect 14345 24996 14349 25052
rect 14285 24992 14349 24996
rect 14365 25052 14429 25056
rect 14365 24996 14369 25052
rect 14369 24996 14425 25052
rect 14425 24996 14429 25052
rect 14365 24992 14429 24996
rect 14445 25052 14509 25056
rect 14445 24996 14449 25052
rect 14449 24996 14505 25052
rect 14505 24996 14509 25052
rect 14445 24992 14509 24996
rect 14525 25052 14589 25056
rect 14525 24996 14529 25052
rect 14529 24996 14585 25052
rect 14585 24996 14589 25052
rect 14525 24992 14589 24996
rect 5764 24984 5828 24988
rect 5764 24928 5778 24984
rect 5778 24928 5828 24984
rect 5764 24924 5828 24928
rect 6285 24508 6349 24512
rect 6285 24452 6289 24508
rect 6289 24452 6345 24508
rect 6345 24452 6349 24508
rect 6285 24448 6349 24452
rect 6365 24508 6429 24512
rect 6365 24452 6369 24508
rect 6369 24452 6425 24508
rect 6425 24452 6429 24508
rect 6365 24448 6429 24452
rect 6445 24508 6509 24512
rect 6445 24452 6449 24508
rect 6449 24452 6505 24508
rect 6505 24452 6509 24508
rect 6445 24448 6509 24452
rect 6525 24508 6589 24512
rect 6525 24452 6529 24508
rect 6529 24452 6585 24508
rect 6585 24452 6589 24508
rect 6525 24448 6589 24452
rect 11618 24508 11682 24512
rect 11618 24452 11622 24508
rect 11622 24452 11678 24508
rect 11678 24452 11682 24508
rect 11618 24448 11682 24452
rect 11698 24508 11762 24512
rect 11698 24452 11702 24508
rect 11702 24452 11758 24508
rect 11758 24452 11762 24508
rect 11698 24448 11762 24452
rect 11778 24508 11842 24512
rect 11778 24452 11782 24508
rect 11782 24452 11838 24508
rect 11838 24452 11842 24508
rect 11778 24448 11842 24452
rect 11858 24508 11922 24512
rect 11858 24452 11862 24508
rect 11862 24452 11918 24508
rect 11918 24452 11922 24508
rect 11858 24448 11922 24452
rect 3618 23964 3682 23968
rect 3618 23908 3622 23964
rect 3622 23908 3678 23964
rect 3678 23908 3682 23964
rect 3618 23904 3682 23908
rect 3698 23964 3762 23968
rect 3698 23908 3702 23964
rect 3702 23908 3758 23964
rect 3758 23908 3762 23964
rect 3698 23904 3762 23908
rect 3778 23964 3842 23968
rect 3778 23908 3782 23964
rect 3782 23908 3838 23964
rect 3838 23908 3842 23964
rect 3778 23904 3842 23908
rect 3858 23964 3922 23968
rect 3858 23908 3862 23964
rect 3862 23908 3918 23964
rect 3918 23908 3922 23964
rect 3858 23904 3922 23908
rect 8952 23964 9016 23968
rect 8952 23908 8956 23964
rect 8956 23908 9012 23964
rect 9012 23908 9016 23964
rect 8952 23904 9016 23908
rect 9032 23964 9096 23968
rect 9032 23908 9036 23964
rect 9036 23908 9092 23964
rect 9092 23908 9096 23964
rect 9032 23904 9096 23908
rect 9112 23964 9176 23968
rect 9112 23908 9116 23964
rect 9116 23908 9172 23964
rect 9172 23908 9176 23964
rect 9112 23904 9176 23908
rect 9192 23964 9256 23968
rect 9192 23908 9196 23964
rect 9196 23908 9252 23964
rect 9252 23908 9256 23964
rect 9192 23904 9256 23908
rect 14285 23964 14349 23968
rect 14285 23908 14289 23964
rect 14289 23908 14345 23964
rect 14345 23908 14349 23964
rect 14285 23904 14349 23908
rect 14365 23964 14429 23968
rect 14365 23908 14369 23964
rect 14369 23908 14425 23964
rect 14425 23908 14429 23964
rect 14365 23904 14429 23908
rect 14445 23964 14509 23968
rect 14445 23908 14449 23964
rect 14449 23908 14505 23964
rect 14505 23908 14509 23964
rect 14445 23904 14509 23908
rect 14525 23964 14589 23968
rect 14525 23908 14529 23964
rect 14529 23908 14585 23964
rect 14585 23908 14589 23964
rect 14525 23904 14589 23908
rect 6285 23420 6349 23424
rect 6285 23364 6289 23420
rect 6289 23364 6345 23420
rect 6345 23364 6349 23420
rect 6285 23360 6349 23364
rect 6365 23420 6429 23424
rect 6365 23364 6369 23420
rect 6369 23364 6425 23420
rect 6425 23364 6429 23420
rect 6365 23360 6429 23364
rect 6445 23420 6509 23424
rect 6445 23364 6449 23420
rect 6449 23364 6505 23420
rect 6505 23364 6509 23420
rect 6445 23360 6509 23364
rect 6525 23420 6589 23424
rect 6525 23364 6529 23420
rect 6529 23364 6585 23420
rect 6585 23364 6589 23420
rect 6525 23360 6589 23364
rect 11618 23420 11682 23424
rect 11618 23364 11622 23420
rect 11622 23364 11678 23420
rect 11678 23364 11682 23420
rect 11618 23360 11682 23364
rect 11698 23420 11762 23424
rect 11698 23364 11702 23420
rect 11702 23364 11758 23420
rect 11758 23364 11762 23420
rect 11698 23360 11762 23364
rect 11778 23420 11842 23424
rect 11778 23364 11782 23420
rect 11782 23364 11838 23420
rect 11838 23364 11842 23420
rect 11778 23360 11842 23364
rect 11858 23420 11922 23424
rect 11858 23364 11862 23420
rect 11862 23364 11918 23420
rect 11918 23364 11922 23420
rect 11858 23360 11922 23364
rect 3618 22876 3682 22880
rect 3618 22820 3622 22876
rect 3622 22820 3678 22876
rect 3678 22820 3682 22876
rect 3618 22816 3682 22820
rect 3698 22876 3762 22880
rect 3698 22820 3702 22876
rect 3702 22820 3758 22876
rect 3758 22820 3762 22876
rect 3698 22816 3762 22820
rect 3778 22876 3842 22880
rect 3778 22820 3782 22876
rect 3782 22820 3838 22876
rect 3838 22820 3842 22876
rect 3778 22816 3842 22820
rect 3858 22876 3922 22880
rect 3858 22820 3862 22876
rect 3862 22820 3918 22876
rect 3918 22820 3922 22876
rect 3858 22816 3922 22820
rect 8952 22876 9016 22880
rect 8952 22820 8956 22876
rect 8956 22820 9012 22876
rect 9012 22820 9016 22876
rect 8952 22816 9016 22820
rect 9032 22876 9096 22880
rect 9032 22820 9036 22876
rect 9036 22820 9092 22876
rect 9092 22820 9096 22876
rect 9032 22816 9096 22820
rect 9112 22876 9176 22880
rect 9112 22820 9116 22876
rect 9116 22820 9172 22876
rect 9172 22820 9176 22876
rect 9112 22816 9176 22820
rect 9192 22876 9256 22880
rect 9192 22820 9196 22876
rect 9196 22820 9252 22876
rect 9252 22820 9256 22876
rect 9192 22816 9256 22820
rect 14285 22876 14349 22880
rect 14285 22820 14289 22876
rect 14289 22820 14345 22876
rect 14345 22820 14349 22876
rect 14285 22816 14349 22820
rect 14365 22876 14429 22880
rect 14365 22820 14369 22876
rect 14369 22820 14425 22876
rect 14425 22820 14429 22876
rect 14365 22816 14429 22820
rect 14445 22876 14509 22880
rect 14445 22820 14449 22876
rect 14449 22820 14505 22876
rect 14505 22820 14509 22876
rect 14445 22816 14509 22820
rect 14525 22876 14589 22880
rect 14525 22820 14529 22876
rect 14529 22820 14585 22876
rect 14585 22820 14589 22876
rect 14525 22816 14589 22820
rect 6285 22332 6349 22336
rect 6285 22276 6289 22332
rect 6289 22276 6345 22332
rect 6345 22276 6349 22332
rect 6285 22272 6349 22276
rect 6365 22332 6429 22336
rect 6365 22276 6369 22332
rect 6369 22276 6425 22332
rect 6425 22276 6429 22332
rect 6365 22272 6429 22276
rect 6445 22332 6509 22336
rect 6445 22276 6449 22332
rect 6449 22276 6505 22332
rect 6505 22276 6509 22332
rect 6445 22272 6509 22276
rect 6525 22332 6589 22336
rect 6525 22276 6529 22332
rect 6529 22276 6585 22332
rect 6585 22276 6589 22332
rect 6525 22272 6589 22276
rect 11618 22332 11682 22336
rect 11618 22276 11622 22332
rect 11622 22276 11678 22332
rect 11678 22276 11682 22332
rect 11618 22272 11682 22276
rect 11698 22332 11762 22336
rect 11698 22276 11702 22332
rect 11702 22276 11758 22332
rect 11758 22276 11762 22332
rect 11698 22272 11762 22276
rect 11778 22332 11842 22336
rect 11778 22276 11782 22332
rect 11782 22276 11838 22332
rect 11838 22276 11842 22332
rect 11778 22272 11842 22276
rect 11858 22332 11922 22336
rect 11858 22276 11862 22332
rect 11862 22276 11918 22332
rect 11918 22276 11922 22332
rect 11858 22272 11922 22276
rect 3618 21788 3682 21792
rect 3618 21732 3622 21788
rect 3622 21732 3678 21788
rect 3678 21732 3682 21788
rect 3618 21728 3682 21732
rect 3698 21788 3762 21792
rect 3698 21732 3702 21788
rect 3702 21732 3758 21788
rect 3758 21732 3762 21788
rect 3698 21728 3762 21732
rect 3778 21788 3842 21792
rect 3778 21732 3782 21788
rect 3782 21732 3838 21788
rect 3838 21732 3842 21788
rect 3778 21728 3842 21732
rect 3858 21788 3922 21792
rect 3858 21732 3862 21788
rect 3862 21732 3918 21788
rect 3918 21732 3922 21788
rect 3858 21728 3922 21732
rect 8952 21788 9016 21792
rect 8952 21732 8956 21788
rect 8956 21732 9012 21788
rect 9012 21732 9016 21788
rect 8952 21728 9016 21732
rect 9032 21788 9096 21792
rect 9032 21732 9036 21788
rect 9036 21732 9092 21788
rect 9092 21732 9096 21788
rect 9032 21728 9096 21732
rect 9112 21788 9176 21792
rect 9112 21732 9116 21788
rect 9116 21732 9172 21788
rect 9172 21732 9176 21788
rect 9112 21728 9176 21732
rect 9192 21788 9256 21792
rect 9192 21732 9196 21788
rect 9196 21732 9252 21788
rect 9252 21732 9256 21788
rect 9192 21728 9256 21732
rect 14285 21788 14349 21792
rect 14285 21732 14289 21788
rect 14289 21732 14345 21788
rect 14345 21732 14349 21788
rect 14285 21728 14349 21732
rect 14365 21788 14429 21792
rect 14365 21732 14369 21788
rect 14369 21732 14425 21788
rect 14425 21732 14429 21788
rect 14365 21728 14429 21732
rect 14445 21788 14509 21792
rect 14445 21732 14449 21788
rect 14449 21732 14505 21788
rect 14505 21732 14509 21788
rect 14445 21728 14509 21732
rect 14525 21788 14589 21792
rect 14525 21732 14529 21788
rect 14529 21732 14585 21788
rect 14585 21732 14589 21788
rect 14525 21728 14589 21732
rect 5764 21312 5828 21316
rect 5764 21256 5778 21312
rect 5778 21256 5828 21312
rect 5764 21252 5828 21256
rect 6285 21244 6349 21248
rect 6285 21188 6289 21244
rect 6289 21188 6345 21244
rect 6345 21188 6349 21244
rect 6285 21184 6349 21188
rect 6365 21244 6429 21248
rect 6365 21188 6369 21244
rect 6369 21188 6425 21244
rect 6425 21188 6429 21244
rect 6365 21184 6429 21188
rect 6445 21244 6509 21248
rect 6445 21188 6449 21244
rect 6449 21188 6505 21244
rect 6505 21188 6509 21244
rect 6445 21184 6509 21188
rect 6525 21244 6589 21248
rect 6525 21188 6529 21244
rect 6529 21188 6585 21244
rect 6585 21188 6589 21244
rect 6525 21184 6589 21188
rect 11618 21244 11682 21248
rect 11618 21188 11622 21244
rect 11622 21188 11678 21244
rect 11678 21188 11682 21244
rect 11618 21184 11682 21188
rect 11698 21244 11762 21248
rect 11698 21188 11702 21244
rect 11702 21188 11758 21244
rect 11758 21188 11762 21244
rect 11698 21184 11762 21188
rect 11778 21244 11842 21248
rect 11778 21188 11782 21244
rect 11782 21188 11838 21244
rect 11838 21188 11842 21244
rect 11778 21184 11842 21188
rect 11858 21244 11922 21248
rect 11858 21188 11862 21244
rect 11862 21188 11918 21244
rect 11918 21188 11922 21244
rect 11858 21184 11922 21188
rect 3618 20700 3682 20704
rect 3618 20644 3622 20700
rect 3622 20644 3678 20700
rect 3678 20644 3682 20700
rect 3618 20640 3682 20644
rect 3698 20700 3762 20704
rect 3698 20644 3702 20700
rect 3702 20644 3758 20700
rect 3758 20644 3762 20700
rect 3698 20640 3762 20644
rect 3778 20700 3842 20704
rect 3778 20644 3782 20700
rect 3782 20644 3838 20700
rect 3838 20644 3842 20700
rect 3778 20640 3842 20644
rect 3858 20700 3922 20704
rect 3858 20644 3862 20700
rect 3862 20644 3918 20700
rect 3918 20644 3922 20700
rect 3858 20640 3922 20644
rect 8952 20700 9016 20704
rect 8952 20644 8956 20700
rect 8956 20644 9012 20700
rect 9012 20644 9016 20700
rect 8952 20640 9016 20644
rect 9032 20700 9096 20704
rect 9032 20644 9036 20700
rect 9036 20644 9092 20700
rect 9092 20644 9096 20700
rect 9032 20640 9096 20644
rect 9112 20700 9176 20704
rect 9112 20644 9116 20700
rect 9116 20644 9172 20700
rect 9172 20644 9176 20700
rect 9112 20640 9176 20644
rect 9192 20700 9256 20704
rect 9192 20644 9196 20700
rect 9196 20644 9252 20700
rect 9252 20644 9256 20700
rect 9192 20640 9256 20644
rect 14285 20700 14349 20704
rect 14285 20644 14289 20700
rect 14289 20644 14345 20700
rect 14345 20644 14349 20700
rect 14285 20640 14349 20644
rect 14365 20700 14429 20704
rect 14365 20644 14369 20700
rect 14369 20644 14425 20700
rect 14425 20644 14429 20700
rect 14365 20640 14429 20644
rect 14445 20700 14509 20704
rect 14445 20644 14449 20700
rect 14449 20644 14505 20700
rect 14505 20644 14509 20700
rect 14445 20640 14509 20644
rect 14525 20700 14589 20704
rect 14525 20644 14529 20700
rect 14529 20644 14585 20700
rect 14585 20644 14589 20700
rect 14525 20640 14589 20644
rect 9444 20300 9508 20364
rect 6285 20156 6349 20160
rect 6285 20100 6289 20156
rect 6289 20100 6345 20156
rect 6345 20100 6349 20156
rect 6285 20096 6349 20100
rect 6365 20156 6429 20160
rect 6365 20100 6369 20156
rect 6369 20100 6425 20156
rect 6425 20100 6429 20156
rect 6365 20096 6429 20100
rect 6445 20156 6509 20160
rect 6445 20100 6449 20156
rect 6449 20100 6505 20156
rect 6505 20100 6509 20156
rect 6445 20096 6509 20100
rect 6525 20156 6589 20160
rect 6525 20100 6529 20156
rect 6529 20100 6585 20156
rect 6585 20100 6589 20156
rect 6525 20096 6589 20100
rect 11618 20156 11682 20160
rect 11618 20100 11622 20156
rect 11622 20100 11678 20156
rect 11678 20100 11682 20156
rect 11618 20096 11682 20100
rect 11698 20156 11762 20160
rect 11698 20100 11702 20156
rect 11702 20100 11758 20156
rect 11758 20100 11762 20156
rect 11698 20096 11762 20100
rect 11778 20156 11842 20160
rect 11778 20100 11782 20156
rect 11782 20100 11838 20156
rect 11838 20100 11842 20156
rect 11778 20096 11842 20100
rect 11858 20156 11922 20160
rect 11858 20100 11862 20156
rect 11862 20100 11918 20156
rect 11918 20100 11922 20156
rect 11858 20096 11922 20100
rect 12020 19952 12084 19956
rect 12020 19896 12070 19952
rect 12070 19896 12084 19952
rect 12020 19892 12084 19896
rect 3618 19612 3682 19616
rect 3618 19556 3622 19612
rect 3622 19556 3678 19612
rect 3678 19556 3682 19612
rect 3618 19552 3682 19556
rect 3698 19612 3762 19616
rect 3698 19556 3702 19612
rect 3702 19556 3758 19612
rect 3758 19556 3762 19612
rect 3698 19552 3762 19556
rect 3778 19612 3842 19616
rect 3778 19556 3782 19612
rect 3782 19556 3838 19612
rect 3838 19556 3842 19612
rect 3778 19552 3842 19556
rect 3858 19612 3922 19616
rect 3858 19556 3862 19612
rect 3862 19556 3918 19612
rect 3918 19556 3922 19612
rect 3858 19552 3922 19556
rect 8952 19612 9016 19616
rect 8952 19556 8956 19612
rect 8956 19556 9012 19612
rect 9012 19556 9016 19612
rect 8952 19552 9016 19556
rect 9032 19612 9096 19616
rect 9032 19556 9036 19612
rect 9036 19556 9092 19612
rect 9092 19556 9096 19612
rect 9032 19552 9096 19556
rect 9112 19612 9176 19616
rect 9112 19556 9116 19612
rect 9116 19556 9172 19612
rect 9172 19556 9176 19612
rect 9112 19552 9176 19556
rect 9192 19612 9256 19616
rect 9192 19556 9196 19612
rect 9196 19556 9252 19612
rect 9252 19556 9256 19612
rect 9192 19552 9256 19556
rect 14285 19612 14349 19616
rect 14285 19556 14289 19612
rect 14289 19556 14345 19612
rect 14345 19556 14349 19612
rect 14285 19552 14349 19556
rect 14365 19612 14429 19616
rect 14365 19556 14369 19612
rect 14369 19556 14425 19612
rect 14425 19556 14429 19612
rect 14365 19552 14429 19556
rect 14445 19612 14509 19616
rect 14445 19556 14449 19612
rect 14449 19556 14505 19612
rect 14505 19556 14509 19612
rect 14445 19552 14509 19556
rect 14525 19612 14589 19616
rect 14525 19556 14529 19612
rect 14529 19556 14585 19612
rect 14585 19556 14589 19612
rect 14525 19552 14589 19556
rect 6285 19068 6349 19072
rect 6285 19012 6289 19068
rect 6289 19012 6345 19068
rect 6345 19012 6349 19068
rect 6285 19008 6349 19012
rect 6365 19068 6429 19072
rect 6365 19012 6369 19068
rect 6369 19012 6425 19068
rect 6425 19012 6429 19068
rect 6365 19008 6429 19012
rect 6445 19068 6509 19072
rect 6445 19012 6449 19068
rect 6449 19012 6505 19068
rect 6505 19012 6509 19068
rect 6445 19008 6509 19012
rect 6525 19068 6589 19072
rect 6525 19012 6529 19068
rect 6529 19012 6585 19068
rect 6585 19012 6589 19068
rect 6525 19008 6589 19012
rect 11618 19068 11682 19072
rect 11618 19012 11622 19068
rect 11622 19012 11678 19068
rect 11678 19012 11682 19068
rect 11618 19008 11682 19012
rect 11698 19068 11762 19072
rect 11698 19012 11702 19068
rect 11702 19012 11758 19068
rect 11758 19012 11762 19068
rect 11698 19008 11762 19012
rect 11778 19068 11842 19072
rect 11778 19012 11782 19068
rect 11782 19012 11838 19068
rect 11838 19012 11842 19068
rect 11778 19008 11842 19012
rect 11858 19068 11922 19072
rect 11858 19012 11862 19068
rect 11862 19012 11918 19068
rect 11918 19012 11922 19068
rect 11858 19008 11922 19012
rect 3618 18524 3682 18528
rect 3618 18468 3622 18524
rect 3622 18468 3678 18524
rect 3678 18468 3682 18524
rect 3618 18464 3682 18468
rect 3698 18524 3762 18528
rect 3698 18468 3702 18524
rect 3702 18468 3758 18524
rect 3758 18468 3762 18524
rect 3698 18464 3762 18468
rect 3778 18524 3842 18528
rect 3778 18468 3782 18524
rect 3782 18468 3838 18524
rect 3838 18468 3842 18524
rect 3778 18464 3842 18468
rect 3858 18524 3922 18528
rect 3858 18468 3862 18524
rect 3862 18468 3918 18524
rect 3918 18468 3922 18524
rect 3858 18464 3922 18468
rect 8952 18524 9016 18528
rect 8952 18468 8956 18524
rect 8956 18468 9012 18524
rect 9012 18468 9016 18524
rect 8952 18464 9016 18468
rect 9032 18524 9096 18528
rect 9032 18468 9036 18524
rect 9036 18468 9092 18524
rect 9092 18468 9096 18524
rect 9032 18464 9096 18468
rect 9112 18524 9176 18528
rect 9112 18468 9116 18524
rect 9116 18468 9172 18524
rect 9172 18468 9176 18524
rect 9112 18464 9176 18468
rect 9192 18524 9256 18528
rect 9192 18468 9196 18524
rect 9196 18468 9252 18524
rect 9252 18468 9256 18524
rect 9192 18464 9256 18468
rect 14285 18524 14349 18528
rect 14285 18468 14289 18524
rect 14289 18468 14345 18524
rect 14345 18468 14349 18524
rect 14285 18464 14349 18468
rect 14365 18524 14429 18528
rect 14365 18468 14369 18524
rect 14369 18468 14425 18524
rect 14425 18468 14429 18524
rect 14365 18464 14429 18468
rect 14445 18524 14509 18528
rect 14445 18468 14449 18524
rect 14449 18468 14505 18524
rect 14505 18468 14509 18524
rect 14445 18464 14509 18468
rect 14525 18524 14589 18528
rect 14525 18468 14529 18524
rect 14529 18468 14585 18524
rect 14585 18468 14589 18524
rect 14525 18464 14589 18468
rect 6285 17980 6349 17984
rect 6285 17924 6289 17980
rect 6289 17924 6345 17980
rect 6345 17924 6349 17980
rect 6285 17920 6349 17924
rect 6365 17980 6429 17984
rect 6365 17924 6369 17980
rect 6369 17924 6425 17980
rect 6425 17924 6429 17980
rect 6365 17920 6429 17924
rect 6445 17980 6509 17984
rect 6445 17924 6449 17980
rect 6449 17924 6505 17980
rect 6505 17924 6509 17980
rect 6445 17920 6509 17924
rect 6525 17980 6589 17984
rect 6525 17924 6529 17980
rect 6529 17924 6585 17980
rect 6585 17924 6589 17980
rect 6525 17920 6589 17924
rect 11618 17980 11682 17984
rect 11618 17924 11622 17980
rect 11622 17924 11678 17980
rect 11678 17924 11682 17980
rect 11618 17920 11682 17924
rect 11698 17980 11762 17984
rect 11698 17924 11702 17980
rect 11702 17924 11758 17980
rect 11758 17924 11762 17980
rect 11698 17920 11762 17924
rect 11778 17980 11842 17984
rect 11778 17924 11782 17980
rect 11782 17924 11838 17980
rect 11838 17924 11842 17980
rect 11778 17920 11842 17924
rect 11858 17980 11922 17984
rect 11858 17924 11862 17980
rect 11862 17924 11918 17980
rect 11918 17924 11922 17980
rect 11858 17920 11922 17924
rect 3618 17436 3682 17440
rect 3618 17380 3622 17436
rect 3622 17380 3678 17436
rect 3678 17380 3682 17436
rect 3618 17376 3682 17380
rect 3698 17436 3762 17440
rect 3698 17380 3702 17436
rect 3702 17380 3758 17436
rect 3758 17380 3762 17436
rect 3698 17376 3762 17380
rect 3778 17436 3842 17440
rect 3778 17380 3782 17436
rect 3782 17380 3838 17436
rect 3838 17380 3842 17436
rect 3778 17376 3842 17380
rect 3858 17436 3922 17440
rect 3858 17380 3862 17436
rect 3862 17380 3918 17436
rect 3918 17380 3922 17436
rect 3858 17376 3922 17380
rect 8952 17436 9016 17440
rect 8952 17380 8956 17436
rect 8956 17380 9012 17436
rect 9012 17380 9016 17436
rect 8952 17376 9016 17380
rect 9032 17436 9096 17440
rect 9032 17380 9036 17436
rect 9036 17380 9092 17436
rect 9092 17380 9096 17436
rect 9032 17376 9096 17380
rect 9112 17436 9176 17440
rect 9112 17380 9116 17436
rect 9116 17380 9172 17436
rect 9172 17380 9176 17436
rect 9112 17376 9176 17380
rect 9192 17436 9256 17440
rect 9192 17380 9196 17436
rect 9196 17380 9252 17436
rect 9252 17380 9256 17436
rect 9192 17376 9256 17380
rect 14285 17436 14349 17440
rect 14285 17380 14289 17436
rect 14289 17380 14345 17436
rect 14345 17380 14349 17436
rect 14285 17376 14349 17380
rect 14365 17436 14429 17440
rect 14365 17380 14369 17436
rect 14369 17380 14425 17436
rect 14425 17380 14429 17436
rect 14365 17376 14429 17380
rect 14445 17436 14509 17440
rect 14445 17380 14449 17436
rect 14449 17380 14505 17436
rect 14505 17380 14509 17436
rect 14445 17376 14509 17380
rect 14525 17436 14589 17440
rect 14525 17380 14529 17436
rect 14529 17380 14585 17436
rect 14585 17380 14589 17436
rect 14525 17376 14589 17380
rect 5028 17172 5092 17236
rect 6285 16892 6349 16896
rect 6285 16836 6289 16892
rect 6289 16836 6345 16892
rect 6345 16836 6349 16892
rect 6285 16832 6349 16836
rect 6365 16892 6429 16896
rect 6365 16836 6369 16892
rect 6369 16836 6425 16892
rect 6425 16836 6429 16892
rect 6365 16832 6429 16836
rect 6445 16892 6509 16896
rect 6445 16836 6449 16892
rect 6449 16836 6505 16892
rect 6505 16836 6509 16892
rect 6445 16832 6509 16836
rect 6525 16892 6589 16896
rect 6525 16836 6529 16892
rect 6529 16836 6585 16892
rect 6585 16836 6589 16892
rect 6525 16832 6589 16836
rect 11618 16892 11682 16896
rect 11618 16836 11622 16892
rect 11622 16836 11678 16892
rect 11678 16836 11682 16892
rect 11618 16832 11682 16836
rect 11698 16892 11762 16896
rect 11698 16836 11702 16892
rect 11702 16836 11758 16892
rect 11758 16836 11762 16892
rect 11698 16832 11762 16836
rect 11778 16892 11842 16896
rect 11778 16836 11782 16892
rect 11782 16836 11838 16892
rect 11838 16836 11842 16892
rect 11778 16832 11842 16836
rect 11858 16892 11922 16896
rect 11858 16836 11862 16892
rect 11862 16836 11918 16892
rect 11918 16836 11922 16892
rect 11858 16832 11922 16836
rect 3618 16348 3682 16352
rect 3618 16292 3622 16348
rect 3622 16292 3678 16348
rect 3678 16292 3682 16348
rect 3618 16288 3682 16292
rect 3698 16348 3762 16352
rect 3698 16292 3702 16348
rect 3702 16292 3758 16348
rect 3758 16292 3762 16348
rect 3698 16288 3762 16292
rect 3778 16348 3842 16352
rect 3778 16292 3782 16348
rect 3782 16292 3838 16348
rect 3838 16292 3842 16348
rect 3778 16288 3842 16292
rect 3858 16348 3922 16352
rect 3858 16292 3862 16348
rect 3862 16292 3918 16348
rect 3918 16292 3922 16348
rect 3858 16288 3922 16292
rect 8952 16348 9016 16352
rect 8952 16292 8956 16348
rect 8956 16292 9012 16348
rect 9012 16292 9016 16348
rect 8952 16288 9016 16292
rect 9032 16348 9096 16352
rect 9032 16292 9036 16348
rect 9036 16292 9092 16348
rect 9092 16292 9096 16348
rect 9032 16288 9096 16292
rect 9112 16348 9176 16352
rect 9112 16292 9116 16348
rect 9116 16292 9172 16348
rect 9172 16292 9176 16348
rect 9112 16288 9176 16292
rect 9192 16348 9256 16352
rect 9192 16292 9196 16348
rect 9196 16292 9252 16348
rect 9252 16292 9256 16348
rect 9192 16288 9256 16292
rect 14285 16348 14349 16352
rect 14285 16292 14289 16348
rect 14289 16292 14345 16348
rect 14345 16292 14349 16348
rect 14285 16288 14349 16292
rect 14365 16348 14429 16352
rect 14365 16292 14369 16348
rect 14369 16292 14425 16348
rect 14425 16292 14429 16348
rect 14365 16288 14429 16292
rect 14445 16348 14509 16352
rect 14445 16292 14449 16348
rect 14449 16292 14505 16348
rect 14505 16292 14509 16348
rect 14445 16288 14509 16292
rect 14525 16348 14589 16352
rect 14525 16292 14529 16348
rect 14529 16292 14585 16348
rect 14585 16292 14589 16348
rect 14525 16288 14589 16292
rect 6285 15804 6349 15808
rect 6285 15748 6289 15804
rect 6289 15748 6345 15804
rect 6345 15748 6349 15804
rect 6285 15744 6349 15748
rect 6365 15804 6429 15808
rect 6365 15748 6369 15804
rect 6369 15748 6425 15804
rect 6425 15748 6429 15804
rect 6365 15744 6429 15748
rect 6445 15804 6509 15808
rect 6445 15748 6449 15804
rect 6449 15748 6505 15804
rect 6505 15748 6509 15804
rect 6445 15744 6509 15748
rect 6525 15804 6589 15808
rect 6525 15748 6529 15804
rect 6529 15748 6585 15804
rect 6585 15748 6589 15804
rect 6525 15744 6589 15748
rect 11618 15804 11682 15808
rect 11618 15748 11622 15804
rect 11622 15748 11678 15804
rect 11678 15748 11682 15804
rect 11618 15744 11682 15748
rect 11698 15804 11762 15808
rect 11698 15748 11702 15804
rect 11702 15748 11758 15804
rect 11758 15748 11762 15804
rect 11698 15744 11762 15748
rect 11778 15804 11842 15808
rect 11778 15748 11782 15804
rect 11782 15748 11838 15804
rect 11838 15748 11842 15804
rect 11778 15744 11842 15748
rect 11858 15804 11922 15808
rect 11858 15748 11862 15804
rect 11862 15748 11918 15804
rect 11918 15748 11922 15804
rect 11858 15744 11922 15748
rect 3618 15260 3682 15264
rect 3618 15204 3622 15260
rect 3622 15204 3678 15260
rect 3678 15204 3682 15260
rect 3618 15200 3682 15204
rect 3698 15260 3762 15264
rect 3698 15204 3702 15260
rect 3702 15204 3758 15260
rect 3758 15204 3762 15260
rect 3698 15200 3762 15204
rect 3778 15260 3842 15264
rect 3778 15204 3782 15260
rect 3782 15204 3838 15260
rect 3838 15204 3842 15260
rect 3778 15200 3842 15204
rect 3858 15260 3922 15264
rect 3858 15204 3862 15260
rect 3862 15204 3918 15260
rect 3918 15204 3922 15260
rect 3858 15200 3922 15204
rect 8952 15260 9016 15264
rect 8952 15204 8956 15260
rect 8956 15204 9012 15260
rect 9012 15204 9016 15260
rect 8952 15200 9016 15204
rect 9032 15260 9096 15264
rect 9032 15204 9036 15260
rect 9036 15204 9092 15260
rect 9092 15204 9096 15260
rect 9032 15200 9096 15204
rect 9112 15260 9176 15264
rect 9112 15204 9116 15260
rect 9116 15204 9172 15260
rect 9172 15204 9176 15260
rect 9112 15200 9176 15204
rect 9192 15260 9256 15264
rect 9192 15204 9196 15260
rect 9196 15204 9252 15260
rect 9252 15204 9256 15260
rect 9192 15200 9256 15204
rect 14285 15260 14349 15264
rect 14285 15204 14289 15260
rect 14289 15204 14345 15260
rect 14345 15204 14349 15260
rect 14285 15200 14349 15204
rect 14365 15260 14429 15264
rect 14365 15204 14369 15260
rect 14369 15204 14425 15260
rect 14425 15204 14429 15260
rect 14365 15200 14429 15204
rect 14445 15260 14509 15264
rect 14445 15204 14449 15260
rect 14449 15204 14505 15260
rect 14505 15204 14509 15260
rect 14445 15200 14509 15204
rect 14525 15260 14589 15264
rect 14525 15204 14529 15260
rect 14529 15204 14585 15260
rect 14585 15204 14589 15260
rect 14525 15200 14589 15204
rect 6285 14716 6349 14720
rect 6285 14660 6289 14716
rect 6289 14660 6345 14716
rect 6345 14660 6349 14716
rect 6285 14656 6349 14660
rect 6365 14716 6429 14720
rect 6365 14660 6369 14716
rect 6369 14660 6425 14716
rect 6425 14660 6429 14716
rect 6365 14656 6429 14660
rect 6445 14716 6509 14720
rect 6445 14660 6449 14716
rect 6449 14660 6505 14716
rect 6505 14660 6509 14716
rect 6445 14656 6509 14660
rect 6525 14716 6589 14720
rect 6525 14660 6529 14716
rect 6529 14660 6585 14716
rect 6585 14660 6589 14716
rect 6525 14656 6589 14660
rect 11618 14716 11682 14720
rect 11618 14660 11622 14716
rect 11622 14660 11678 14716
rect 11678 14660 11682 14716
rect 11618 14656 11682 14660
rect 11698 14716 11762 14720
rect 11698 14660 11702 14716
rect 11702 14660 11758 14716
rect 11758 14660 11762 14716
rect 11698 14656 11762 14660
rect 11778 14716 11842 14720
rect 11778 14660 11782 14716
rect 11782 14660 11838 14716
rect 11838 14660 11842 14716
rect 11778 14656 11842 14660
rect 11858 14716 11922 14720
rect 11858 14660 11862 14716
rect 11862 14660 11918 14716
rect 11918 14660 11922 14716
rect 11858 14656 11922 14660
rect 3618 14172 3682 14176
rect 3618 14116 3622 14172
rect 3622 14116 3678 14172
rect 3678 14116 3682 14172
rect 3618 14112 3682 14116
rect 3698 14172 3762 14176
rect 3698 14116 3702 14172
rect 3702 14116 3758 14172
rect 3758 14116 3762 14172
rect 3698 14112 3762 14116
rect 3778 14172 3842 14176
rect 3778 14116 3782 14172
rect 3782 14116 3838 14172
rect 3838 14116 3842 14172
rect 3778 14112 3842 14116
rect 3858 14172 3922 14176
rect 3858 14116 3862 14172
rect 3862 14116 3918 14172
rect 3918 14116 3922 14172
rect 3858 14112 3922 14116
rect 8952 14172 9016 14176
rect 8952 14116 8956 14172
rect 8956 14116 9012 14172
rect 9012 14116 9016 14172
rect 8952 14112 9016 14116
rect 9032 14172 9096 14176
rect 9032 14116 9036 14172
rect 9036 14116 9092 14172
rect 9092 14116 9096 14172
rect 9032 14112 9096 14116
rect 9112 14172 9176 14176
rect 9112 14116 9116 14172
rect 9116 14116 9172 14172
rect 9172 14116 9176 14172
rect 9112 14112 9176 14116
rect 9192 14172 9256 14176
rect 9192 14116 9196 14172
rect 9196 14116 9252 14172
rect 9252 14116 9256 14172
rect 9192 14112 9256 14116
rect 14285 14172 14349 14176
rect 14285 14116 14289 14172
rect 14289 14116 14345 14172
rect 14345 14116 14349 14172
rect 14285 14112 14349 14116
rect 14365 14172 14429 14176
rect 14365 14116 14369 14172
rect 14369 14116 14425 14172
rect 14425 14116 14429 14172
rect 14365 14112 14429 14116
rect 14445 14172 14509 14176
rect 14445 14116 14449 14172
rect 14449 14116 14505 14172
rect 14505 14116 14509 14172
rect 14445 14112 14509 14116
rect 14525 14172 14589 14176
rect 14525 14116 14529 14172
rect 14529 14116 14585 14172
rect 14585 14116 14589 14172
rect 14525 14112 14589 14116
rect 6285 13628 6349 13632
rect 6285 13572 6289 13628
rect 6289 13572 6345 13628
rect 6345 13572 6349 13628
rect 6285 13568 6349 13572
rect 6365 13628 6429 13632
rect 6365 13572 6369 13628
rect 6369 13572 6425 13628
rect 6425 13572 6429 13628
rect 6365 13568 6429 13572
rect 6445 13628 6509 13632
rect 6445 13572 6449 13628
rect 6449 13572 6505 13628
rect 6505 13572 6509 13628
rect 6445 13568 6509 13572
rect 6525 13628 6589 13632
rect 6525 13572 6529 13628
rect 6529 13572 6585 13628
rect 6585 13572 6589 13628
rect 6525 13568 6589 13572
rect 11618 13628 11682 13632
rect 11618 13572 11622 13628
rect 11622 13572 11678 13628
rect 11678 13572 11682 13628
rect 11618 13568 11682 13572
rect 11698 13628 11762 13632
rect 11698 13572 11702 13628
rect 11702 13572 11758 13628
rect 11758 13572 11762 13628
rect 11698 13568 11762 13572
rect 11778 13628 11842 13632
rect 11778 13572 11782 13628
rect 11782 13572 11838 13628
rect 11838 13572 11842 13628
rect 11778 13568 11842 13572
rect 11858 13628 11922 13632
rect 11858 13572 11862 13628
rect 11862 13572 11918 13628
rect 11918 13572 11922 13628
rect 11858 13568 11922 13572
rect 3618 13084 3682 13088
rect 3618 13028 3622 13084
rect 3622 13028 3678 13084
rect 3678 13028 3682 13084
rect 3618 13024 3682 13028
rect 3698 13084 3762 13088
rect 3698 13028 3702 13084
rect 3702 13028 3758 13084
rect 3758 13028 3762 13084
rect 3698 13024 3762 13028
rect 3778 13084 3842 13088
rect 3778 13028 3782 13084
rect 3782 13028 3838 13084
rect 3838 13028 3842 13084
rect 3778 13024 3842 13028
rect 3858 13084 3922 13088
rect 3858 13028 3862 13084
rect 3862 13028 3918 13084
rect 3918 13028 3922 13084
rect 3858 13024 3922 13028
rect 8952 13084 9016 13088
rect 8952 13028 8956 13084
rect 8956 13028 9012 13084
rect 9012 13028 9016 13084
rect 8952 13024 9016 13028
rect 9032 13084 9096 13088
rect 9032 13028 9036 13084
rect 9036 13028 9092 13084
rect 9092 13028 9096 13084
rect 9032 13024 9096 13028
rect 9112 13084 9176 13088
rect 9112 13028 9116 13084
rect 9116 13028 9172 13084
rect 9172 13028 9176 13084
rect 9112 13024 9176 13028
rect 9192 13084 9256 13088
rect 9192 13028 9196 13084
rect 9196 13028 9252 13084
rect 9252 13028 9256 13084
rect 9192 13024 9256 13028
rect 14285 13084 14349 13088
rect 14285 13028 14289 13084
rect 14289 13028 14345 13084
rect 14345 13028 14349 13084
rect 14285 13024 14349 13028
rect 14365 13084 14429 13088
rect 14365 13028 14369 13084
rect 14369 13028 14425 13084
rect 14425 13028 14429 13084
rect 14365 13024 14429 13028
rect 14445 13084 14509 13088
rect 14445 13028 14449 13084
rect 14449 13028 14505 13084
rect 14505 13028 14509 13084
rect 14445 13024 14509 13028
rect 14525 13084 14589 13088
rect 14525 13028 14529 13084
rect 14529 13028 14585 13084
rect 14585 13028 14589 13084
rect 14525 13024 14589 13028
rect 6285 12540 6349 12544
rect 6285 12484 6289 12540
rect 6289 12484 6345 12540
rect 6345 12484 6349 12540
rect 6285 12480 6349 12484
rect 6365 12540 6429 12544
rect 6365 12484 6369 12540
rect 6369 12484 6425 12540
rect 6425 12484 6429 12540
rect 6365 12480 6429 12484
rect 6445 12540 6509 12544
rect 6445 12484 6449 12540
rect 6449 12484 6505 12540
rect 6505 12484 6509 12540
rect 6445 12480 6509 12484
rect 6525 12540 6589 12544
rect 6525 12484 6529 12540
rect 6529 12484 6585 12540
rect 6585 12484 6589 12540
rect 6525 12480 6589 12484
rect 11618 12540 11682 12544
rect 11618 12484 11622 12540
rect 11622 12484 11678 12540
rect 11678 12484 11682 12540
rect 11618 12480 11682 12484
rect 11698 12540 11762 12544
rect 11698 12484 11702 12540
rect 11702 12484 11758 12540
rect 11758 12484 11762 12540
rect 11698 12480 11762 12484
rect 11778 12540 11842 12544
rect 11778 12484 11782 12540
rect 11782 12484 11838 12540
rect 11838 12484 11842 12540
rect 11778 12480 11842 12484
rect 11858 12540 11922 12544
rect 11858 12484 11862 12540
rect 11862 12484 11918 12540
rect 11918 12484 11922 12540
rect 11858 12480 11922 12484
rect 3618 11996 3682 12000
rect 3618 11940 3622 11996
rect 3622 11940 3678 11996
rect 3678 11940 3682 11996
rect 3618 11936 3682 11940
rect 3698 11996 3762 12000
rect 3698 11940 3702 11996
rect 3702 11940 3758 11996
rect 3758 11940 3762 11996
rect 3698 11936 3762 11940
rect 3778 11996 3842 12000
rect 3778 11940 3782 11996
rect 3782 11940 3838 11996
rect 3838 11940 3842 11996
rect 3778 11936 3842 11940
rect 3858 11996 3922 12000
rect 3858 11940 3862 11996
rect 3862 11940 3918 11996
rect 3918 11940 3922 11996
rect 3858 11936 3922 11940
rect 8952 11996 9016 12000
rect 8952 11940 8956 11996
rect 8956 11940 9012 11996
rect 9012 11940 9016 11996
rect 8952 11936 9016 11940
rect 9032 11996 9096 12000
rect 9032 11940 9036 11996
rect 9036 11940 9092 11996
rect 9092 11940 9096 11996
rect 9032 11936 9096 11940
rect 9112 11996 9176 12000
rect 9112 11940 9116 11996
rect 9116 11940 9172 11996
rect 9172 11940 9176 11996
rect 9112 11936 9176 11940
rect 9192 11996 9256 12000
rect 9192 11940 9196 11996
rect 9196 11940 9252 11996
rect 9252 11940 9256 11996
rect 9192 11936 9256 11940
rect 14285 11996 14349 12000
rect 14285 11940 14289 11996
rect 14289 11940 14345 11996
rect 14345 11940 14349 11996
rect 14285 11936 14349 11940
rect 14365 11996 14429 12000
rect 14365 11940 14369 11996
rect 14369 11940 14425 11996
rect 14425 11940 14429 11996
rect 14365 11936 14429 11940
rect 14445 11996 14509 12000
rect 14445 11940 14449 11996
rect 14449 11940 14505 11996
rect 14505 11940 14509 11996
rect 14445 11936 14509 11940
rect 14525 11996 14589 12000
rect 14525 11940 14529 11996
rect 14529 11940 14585 11996
rect 14585 11940 14589 11996
rect 14525 11936 14589 11940
rect 5028 11656 5092 11660
rect 5028 11600 5042 11656
rect 5042 11600 5092 11656
rect 5028 11596 5092 11600
rect 6285 11452 6349 11456
rect 6285 11396 6289 11452
rect 6289 11396 6345 11452
rect 6345 11396 6349 11452
rect 6285 11392 6349 11396
rect 6365 11452 6429 11456
rect 6365 11396 6369 11452
rect 6369 11396 6425 11452
rect 6425 11396 6429 11452
rect 6365 11392 6429 11396
rect 6445 11452 6509 11456
rect 6445 11396 6449 11452
rect 6449 11396 6505 11452
rect 6505 11396 6509 11452
rect 6445 11392 6509 11396
rect 6525 11452 6589 11456
rect 6525 11396 6529 11452
rect 6529 11396 6585 11452
rect 6585 11396 6589 11452
rect 6525 11392 6589 11396
rect 11618 11452 11682 11456
rect 11618 11396 11622 11452
rect 11622 11396 11678 11452
rect 11678 11396 11682 11452
rect 11618 11392 11682 11396
rect 11698 11452 11762 11456
rect 11698 11396 11702 11452
rect 11702 11396 11758 11452
rect 11758 11396 11762 11452
rect 11698 11392 11762 11396
rect 11778 11452 11842 11456
rect 11778 11396 11782 11452
rect 11782 11396 11838 11452
rect 11838 11396 11842 11452
rect 11778 11392 11842 11396
rect 11858 11452 11922 11456
rect 11858 11396 11862 11452
rect 11862 11396 11918 11452
rect 11918 11396 11922 11452
rect 11858 11392 11922 11396
rect 3618 10908 3682 10912
rect 3618 10852 3622 10908
rect 3622 10852 3678 10908
rect 3678 10852 3682 10908
rect 3618 10848 3682 10852
rect 3698 10908 3762 10912
rect 3698 10852 3702 10908
rect 3702 10852 3758 10908
rect 3758 10852 3762 10908
rect 3698 10848 3762 10852
rect 3778 10908 3842 10912
rect 3778 10852 3782 10908
rect 3782 10852 3838 10908
rect 3838 10852 3842 10908
rect 3778 10848 3842 10852
rect 3858 10908 3922 10912
rect 3858 10852 3862 10908
rect 3862 10852 3918 10908
rect 3918 10852 3922 10908
rect 3858 10848 3922 10852
rect 8952 10908 9016 10912
rect 8952 10852 8956 10908
rect 8956 10852 9012 10908
rect 9012 10852 9016 10908
rect 8952 10848 9016 10852
rect 9032 10908 9096 10912
rect 9032 10852 9036 10908
rect 9036 10852 9092 10908
rect 9092 10852 9096 10908
rect 9032 10848 9096 10852
rect 9112 10908 9176 10912
rect 9112 10852 9116 10908
rect 9116 10852 9172 10908
rect 9172 10852 9176 10908
rect 9112 10848 9176 10852
rect 9192 10908 9256 10912
rect 9192 10852 9196 10908
rect 9196 10852 9252 10908
rect 9252 10852 9256 10908
rect 9192 10848 9256 10852
rect 14285 10908 14349 10912
rect 14285 10852 14289 10908
rect 14289 10852 14345 10908
rect 14345 10852 14349 10908
rect 14285 10848 14349 10852
rect 14365 10908 14429 10912
rect 14365 10852 14369 10908
rect 14369 10852 14425 10908
rect 14425 10852 14429 10908
rect 14365 10848 14429 10852
rect 14445 10908 14509 10912
rect 14445 10852 14449 10908
rect 14449 10852 14505 10908
rect 14505 10852 14509 10908
rect 14445 10848 14509 10852
rect 14525 10908 14589 10912
rect 14525 10852 14529 10908
rect 14529 10852 14585 10908
rect 14585 10852 14589 10908
rect 14525 10848 14589 10852
rect 6285 10364 6349 10368
rect 6285 10308 6289 10364
rect 6289 10308 6345 10364
rect 6345 10308 6349 10364
rect 6285 10304 6349 10308
rect 6365 10364 6429 10368
rect 6365 10308 6369 10364
rect 6369 10308 6425 10364
rect 6425 10308 6429 10364
rect 6365 10304 6429 10308
rect 6445 10364 6509 10368
rect 6445 10308 6449 10364
rect 6449 10308 6505 10364
rect 6505 10308 6509 10364
rect 6445 10304 6509 10308
rect 6525 10364 6589 10368
rect 6525 10308 6529 10364
rect 6529 10308 6585 10364
rect 6585 10308 6589 10364
rect 6525 10304 6589 10308
rect 11618 10364 11682 10368
rect 11618 10308 11622 10364
rect 11622 10308 11678 10364
rect 11678 10308 11682 10364
rect 11618 10304 11682 10308
rect 11698 10364 11762 10368
rect 11698 10308 11702 10364
rect 11702 10308 11758 10364
rect 11758 10308 11762 10364
rect 11698 10304 11762 10308
rect 11778 10364 11842 10368
rect 11778 10308 11782 10364
rect 11782 10308 11838 10364
rect 11838 10308 11842 10364
rect 11778 10304 11842 10308
rect 11858 10364 11922 10368
rect 11858 10308 11862 10364
rect 11862 10308 11918 10364
rect 11918 10308 11922 10364
rect 11858 10304 11922 10308
rect 3618 9820 3682 9824
rect 3618 9764 3622 9820
rect 3622 9764 3678 9820
rect 3678 9764 3682 9820
rect 3618 9760 3682 9764
rect 3698 9820 3762 9824
rect 3698 9764 3702 9820
rect 3702 9764 3758 9820
rect 3758 9764 3762 9820
rect 3698 9760 3762 9764
rect 3778 9820 3842 9824
rect 3778 9764 3782 9820
rect 3782 9764 3838 9820
rect 3838 9764 3842 9820
rect 3778 9760 3842 9764
rect 3858 9820 3922 9824
rect 3858 9764 3862 9820
rect 3862 9764 3918 9820
rect 3918 9764 3922 9820
rect 3858 9760 3922 9764
rect 8952 9820 9016 9824
rect 8952 9764 8956 9820
rect 8956 9764 9012 9820
rect 9012 9764 9016 9820
rect 8952 9760 9016 9764
rect 9032 9820 9096 9824
rect 9032 9764 9036 9820
rect 9036 9764 9092 9820
rect 9092 9764 9096 9820
rect 9032 9760 9096 9764
rect 9112 9820 9176 9824
rect 9112 9764 9116 9820
rect 9116 9764 9172 9820
rect 9172 9764 9176 9820
rect 9112 9760 9176 9764
rect 9192 9820 9256 9824
rect 9192 9764 9196 9820
rect 9196 9764 9252 9820
rect 9252 9764 9256 9820
rect 9192 9760 9256 9764
rect 14285 9820 14349 9824
rect 14285 9764 14289 9820
rect 14289 9764 14345 9820
rect 14345 9764 14349 9820
rect 14285 9760 14349 9764
rect 14365 9820 14429 9824
rect 14365 9764 14369 9820
rect 14369 9764 14425 9820
rect 14425 9764 14429 9820
rect 14365 9760 14429 9764
rect 14445 9820 14509 9824
rect 14445 9764 14449 9820
rect 14449 9764 14505 9820
rect 14505 9764 14509 9820
rect 14445 9760 14509 9764
rect 14525 9820 14589 9824
rect 14525 9764 14529 9820
rect 14529 9764 14585 9820
rect 14585 9764 14589 9820
rect 14525 9760 14589 9764
rect 6285 9276 6349 9280
rect 6285 9220 6289 9276
rect 6289 9220 6345 9276
rect 6345 9220 6349 9276
rect 6285 9216 6349 9220
rect 6365 9276 6429 9280
rect 6365 9220 6369 9276
rect 6369 9220 6425 9276
rect 6425 9220 6429 9276
rect 6365 9216 6429 9220
rect 6445 9276 6509 9280
rect 6445 9220 6449 9276
rect 6449 9220 6505 9276
rect 6505 9220 6509 9276
rect 6445 9216 6509 9220
rect 6525 9276 6589 9280
rect 6525 9220 6529 9276
rect 6529 9220 6585 9276
rect 6585 9220 6589 9276
rect 6525 9216 6589 9220
rect 11618 9276 11682 9280
rect 11618 9220 11622 9276
rect 11622 9220 11678 9276
rect 11678 9220 11682 9276
rect 11618 9216 11682 9220
rect 11698 9276 11762 9280
rect 11698 9220 11702 9276
rect 11702 9220 11758 9276
rect 11758 9220 11762 9276
rect 11698 9216 11762 9220
rect 11778 9276 11842 9280
rect 11778 9220 11782 9276
rect 11782 9220 11838 9276
rect 11838 9220 11842 9276
rect 11778 9216 11842 9220
rect 11858 9276 11922 9280
rect 11858 9220 11862 9276
rect 11862 9220 11918 9276
rect 11918 9220 11922 9276
rect 11858 9216 11922 9220
rect 7972 9012 8036 9076
rect 3618 8732 3682 8736
rect 3618 8676 3622 8732
rect 3622 8676 3678 8732
rect 3678 8676 3682 8732
rect 3618 8672 3682 8676
rect 3698 8732 3762 8736
rect 3698 8676 3702 8732
rect 3702 8676 3758 8732
rect 3758 8676 3762 8732
rect 3698 8672 3762 8676
rect 3778 8732 3842 8736
rect 3778 8676 3782 8732
rect 3782 8676 3838 8732
rect 3838 8676 3842 8732
rect 3778 8672 3842 8676
rect 3858 8732 3922 8736
rect 3858 8676 3862 8732
rect 3862 8676 3918 8732
rect 3918 8676 3922 8732
rect 3858 8672 3922 8676
rect 8952 8732 9016 8736
rect 8952 8676 8956 8732
rect 8956 8676 9012 8732
rect 9012 8676 9016 8732
rect 8952 8672 9016 8676
rect 9032 8732 9096 8736
rect 9032 8676 9036 8732
rect 9036 8676 9092 8732
rect 9092 8676 9096 8732
rect 9032 8672 9096 8676
rect 9112 8732 9176 8736
rect 9112 8676 9116 8732
rect 9116 8676 9172 8732
rect 9172 8676 9176 8732
rect 9112 8672 9176 8676
rect 9192 8732 9256 8736
rect 9192 8676 9196 8732
rect 9196 8676 9252 8732
rect 9252 8676 9256 8732
rect 9192 8672 9256 8676
rect 14285 8732 14349 8736
rect 14285 8676 14289 8732
rect 14289 8676 14345 8732
rect 14345 8676 14349 8732
rect 14285 8672 14349 8676
rect 14365 8732 14429 8736
rect 14365 8676 14369 8732
rect 14369 8676 14425 8732
rect 14425 8676 14429 8732
rect 14365 8672 14429 8676
rect 14445 8732 14509 8736
rect 14445 8676 14449 8732
rect 14449 8676 14505 8732
rect 14505 8676 14509 8732
rect 14445 8672 14509 8676
rect 14525 8732 14589 8736
rect 14525 8676 14529 8732
rect 14529 8676 14585 8732
rect 14585 8676 14589 8732
rect 14525 8672 14589 8676
rect 6285 8188 6349 8192
rect 6285 8132 6289 8188
rect 6289 8132 6345 8188
rect 6345 8132 6349 8188
rect 6285 8128 6349 8132
rect 6365 8188 6429 8192
rect 6365 8132 6369 8188
rect 6369 8132 6425 8188
rect 6425 8132 6429 8188
rect 6365 8128 6429 8132
rect 6445 8188 6509 8192
rect 6445 8132 6449 8188
rect 6449 8132 6505 8188
rect 6505 8132 6509 8188
rect 6445 8128 6509 8132
rect 6525 8188 6589 8192
rect 6525 8132 6529 8188
rect 6529 8132 6585 8188
rect 6585 8132 6589 8188
rect 6525 8128 6589 8132
rect 11618 8188 11682 8192
rect 11618 8132 11622 8188
rect 11622 8132 11678 8188
rect 11678 8132 11682 8188
rect 11618 8128 11682 8132
rect 11698 8188 11762 8192
rect 11698 8132 11702 8188
rect 11702 8132 11758 8188
rect 11758 8132 11762 8188
rect 11698 8128 11762 8132
rect 11778 8188 11842 8192
rect 11778 8132 11782 8188
rect 11782 8132 11838 8188
rect 11838 8132 11842 8188
rect 11778 8128 11842 8132
rect 11858 8188 11922 8192
rect 11858 8132 11862 8188
rect 11862 8132 11918 8188
rect 11918 8132 11922 8188
rect 11858 8128 11922 8132
rect 7420 7984 7484 7988
rect 7420 7928 7434 7984
rect 7434 7928 7484 7984
rect 7420 7924 7484 7928
rect 3618 7644 3682 7648
rect 3618 7588 3622 7644
rect 3622 7588 3678 7644
rect 3678 7588 3682 7644
rect 3618 7584 3682 7588
rect 3698 7644 3762 7648
rect 3698 7588 3702 7644
rect 3702 7588 3758 7644
rect 3758 7588 3762 7644
rect 3698 7584 3762 7588
rect 3778 7644 3842 7648
rect 3778 7588 3782 7644
rect 3782 7588 3838 7644
rect 3838 7588 3842 7644
rect 3778 7584 3842 7588
rect 3858 7644 3922 7648
rect 3858 7588 3862 7644
rect 3862 7588 3918 7644
rect 3918 7588 3922 7644
rect 3858 7584 3922 7588
rect 8952 7644 9016 7648
rect 8952 7588 8956 7644
rect 8956 7588 9012 7644
rect 9012 7588 9016 7644
rect 8952 7584 9016 7588
rect 9032 7644 9096 7648
rect 9032 7588 9036 7644
rect 9036 7588 9092 7644
rect 9092 7588 9096 7644
rect 9032 7584 9096 7588
rect 9112 7644 9176 7648
rect 9112 7588 9116 7644
rect 9116 7588 9172 7644
rect 9172 7588 9176 7644
rect 9112 7584 9176 7588
rect 9192 7644 9256 7648
rect 9192 7588 9196 7644
rect 9196 7588 9252 7644
rect 9252 7588 9256 7644
rect 9192 7584 9256 7588
rect 14285 7644 14349 7648
rect 14285 7588 14289 7644
rect 14289 7588 14345 7644
rect 14345 7588 14349 7644
rect 14285 7584 14349 7588
rect 14365 7644 14429 7648
rect 14365 7588 14369 7644
rect 14369 7588 14425 7644
rect 14425 7588 14429 7644
rect 14365 7584 14429 7588
rect 14445 7644 14509 7648
rect 14445 7588 14449 7644
rect 14449 7588 14505 7644
rect 14505 7588 14509 7644
rect 14445 7584 14509 7588
rect 14525 7644 14589 7648
rect 14525 7588 14529 7644
rect 14529 7588 14585 7644
rect 14585 7588 14589 7644
rect 14525 7584 14589 7588
rect 6285 7100 6349 7104
rect 6285 7044 6289 7100
rect 6289 7044 6345 7100
rect 6345 7044 6349 7100
rect 6285 7040 6349 7044
rect 6365 7100 6429 7104
rect 6365 7044 6369 7100
rect 6369 7044 6425 7100
rect 6425 7044 6429 7100
rect 6365 7040 6429 7044
rect 6445 7100 6509 7104
rect 6445 7044 6449 7100
rect 6449 7044 6505 7100
rect 6505 7044 6509 7100
rect 6445 7040 6509 7044
rect 6525 7100 6589 7104
rect 6525 7044 6529 7100
rect 6529 7044 6585 7100
rect 6585 7044 6589 7100
rect 6525 7040 6589 7044
rect 11618 7100 11682 7104
rect 11618 7044 11622 7100
rect 11622 7044 11678 7100
rect 11678 7044 11682 7100
rect 11618 7040 11682 7044
rect 11698 7100 11762 7104
rect 11698 7044 11702 7100
rect 11702 7044 11758 7100
rect 11758 7044 11762 7100
rect 11698 7040 11762 7044
rect 11778 7100 11842 7104
rect 11778 7044 11782 7100
rect 11782 7044 11838 7100
rect 11838 7044 11842 7100
rect 11778 7040 11842 7044
rect 11858 7100 11922 7104
rect 11858 7044 11862 7100
rect 11862 7044 11918 7100
rect 11918 7044 11922 7100
rect 11858 7040 11922 7044
rect 3618 6556 3682 6560
rect 3618 6500 3622 6556
rect 3622 6500 3678 6556
rect 3678 6500 3682 6556
rect 3618 6496 3682 6500
rect 3698 6556 3762 6560
rect 3698 6500 3702 6556
rect 3702 6500 3758 6556
rect 3758 6500 3762 6556
rect 3698 6496 3762 6500
rect 3778 6556 3842 6560
rect 3778 6500 3782 6556
rect 3782 6500 3838 6556
rect 3838 6500 3842 6556
rect 3778 6496 3842 6500
rect 3858 6556 3922 6560
rect 3858 6500 3862 6556
rect 3862 6500 3918 6556
rect 3918 6500 3922 6556
rect 3858 6496 3922 6500
rect 8952 6556 9016 6560
rect 8952 6500 8956 6556
rect 8956 6500 9012 6556
rect 9012 6500 9016 6556
rect 8952 6496 9016 6500
rect 9032 6556 9096 6560
rect 9032 6500 9036 6556
rect 9036 6500 9092 6556
rect 9092 6500 9096 6556
rect 9032 6496 9096 6500
rect 9112 6556 9176 6560
rect 9112 6500 9116 6556
rect 9116 6500 9172 6556
rect 9172 6500 9176 6556
rect 9112 6496 9176 6500
rect 9192 6556 9256 6560
rect 9192 6500 9196 6556
rect 9196 6500 9252 6556
rect 9252 6500 9256 6556
rect 9192 6496 9256 6500
rect 14285 6556 14349 6560
rect 14285 6500 14289 6556
rect 14289 6500 14345 6556
rect 14345 6500 14349 6556
rect 14285 6496 14349 6500
rect 14365 6556 14429 6560
rect 14365 6500 14369 6556
rect 14369 6500 14425 6556
rect 14425 6500 14429 6556
rect 14365 6496 14429 6500
rect 14445 6556 14509 6560
rect 14445 6500 14449 6556
rect 14449 6500 14505 6556
rect 14505 6500 14509 6556
rect 14445 6496 14509 6500
rect 14525 6556 14589 6560
rect 14525 6500 14529 6556
rect 14529 6500 14585 6556
rect 14585 6500 14589 6556
rect 14525 6496 14589 6500
rect 6285 6012 6349 6016
rect 6285 5956 6289 6012
rect 6289 5956 6345 6012
rect 6345 5956 6349 6012
rect 6285 5952 6349 5956
rect 6365 6012 6429 6016
rect 6365 5956 6369 6012
rect 6369 5956 6425 6012
rect 6425 5956 6429 6012
rect 6365 5952 6429 5956
rect 6445 6012 6509 6016
rect 6445 5956 6449 6012
rect 6449 5956 6505 6012
rect 6505 5956 6509 6012
rect 6445 5952 6509 5956
rect 6525 6012 6589 6016
rect 6525 5956 6529 6012
rect 6529 5956 6585 6012
rect 6585 5956 6589 6012
rect 6525 5952 6589 5956
rect 11618 6012 11682 6016
rect 11618 5956 11622 6012
rect 11622 5956 11678 6012
rect 11678 5956 11682 6012
rect 11618 5952 11682 5956
rect 11698 6012 11762 6016
rect 11698 5956 11702 6012
rect 11702 5956 11758 6012
rect 11758 5956 11762 6012
rect 11698 5952 11762 5956
rect 11778 6012 11842 6016
rect 11778 5956 11782 6012
rect 11782 5956 11838 6012
rect 11838 5956 11842 6012
rect 11778 5952 11842 5956
rect 11858 6012 11922 6016
rect 11858 5956 11862 6012
rect 11862 5956 11918 6012
rect 11918 5956 11922 6012
rect 11858 5952 11922 5956
rect 3618 5468 3682 5472
rect 3618 5412 3622 5468
rect 3622 5412 3678 5468
rect 3678 5412 3682 5468
rect 3618 5408 3682 5412
rect 3698 5468 3762 5472
rect 3698 5412 3702 5468
rect 3702 5412 3758 5468
rect 3758 5412 3762 5468
rect 3698 5408 3762 5412
rect 3778 5468 3842 5472
rect 3778 5412 3782 5468
rect 3782 5412 3838 5468
rect 3838 5412 3842 5468
rect 3778 5408 3842 5412
rect 3858 5468 3922 5472
rect 3858 5412 3862 5468
rect 3862 5412 3918 5468
rect 3918 5412 3922 5468
rect 3858 5408 3922 5412
rect 8952 5468 9016 5472
rect 8952 5412 8956 5468
rect 8956 5412 9012 5468
rect 9012 5412 9016 5468
rect 8952 5408 9016 5412
rect 9032 5468 9096 5472
rect 9032 5412 9036 5468
rect 9036 5412 9092 5468
rect 9092 5412 9096 5468
rect 9032 5408 9096 5412
rect 9112 5468 9176 5472
rect 9112 5412 9116 5468
rect 9116 5412 9172 5468
rect 9172 5412 9176 5468
rect 9112 5408 9176 5412
rect 9192 5468 9256 5472
rect 9192 5412 9196 5468
rect 9196 5412 9252 5468
rect 9252 5412 9256 5468
rect 9192 5408 9256 5412
rect 14285 5468 14349 5472
rect 14285 5412 14289 5468
rect 14289 5412 14345 5468
rect 14345 5412 14349 5468
rect 14285 5408 14349 5412
rect 14365 5468 14429 5472
rect 14365 5412 14369 5468
rect 14369 5412 14425 5468
rect 14425 5412 14429 5468
rect 14365 5408 14429 5412
rect 14445 5468 14509 5472
rect 14445 5412 14449 5468
rect 14449 5412 14505 5468
rect 14505 5412 14509 5468
rect 14445 5408 14509 5412
rect 14525 5468 14589 5472
rect 14525 5412 14529 5468
rect 14529 5412 14585 5468
rect 14585 5412 14589 5468
rect 14525 5408 14589 5412
rect 6285 4924 6349 4928
rect 6285 4868 6289 4924
rect 6289 4868 6345 4924
rect 6345 4868 6349 4924
rect 6285 4864 6349 4868
rect 6365 4924 6429 4928
rect 6365 4868 6369 4924
rect 6369 4868 6425 4924
rect 6425 4868 6429 4924
rect 6365 4864 6429 4868
rect 6445 4924 6509 4928
rect 6445 4868 6449 4924
rect 6449 4868 6505 4924
rect 6505 4868 6509 4924
rect 6445 4864 6509 4868
rect 6525 4924 6589 4928
rect 6525 4868 6529 4924
rect 6529 4868 6585 4924
rect 6585 4868 6589 4924
rect 6525 4864 6589 4868
rect 11618 4924 11682 4928
rect 11618 4868 11622 4924
rect 11622 4868 11678 4924
rect 11678 4868 11682 4924
rect 11618 4864 11682 4868
rect 11698 4924 11762 4928
rect 11698 4868 11702 4924
rect 11702 4868 11758 4924
rect 11758 4868 11762 4924
rect 11698 4864 11762 4868
rect 11778 4924 11842 4928
rect 11778 4868 11782 4924
rect 11782 4868 11838 4924
rect 11838 4868 11842 4924
rect 11778 4864 11842 4868
rect 11858 4924 11922 4928
rect 11858 4868 11862 4924
rect 11862 4868 11918 4924
rect 11918 4868 11922 4924
rect 11858 4864 11922 4868
rect 3618 4380 3682 4384
rect 3618 4324 3622 4380
rect 3622 4324 3678 4380
rect 3678 4324 3682 4380
rect 3618 4320 3682 4324
rect 3698 4380 3762 4384
rect 3698 4324 3702 4380
rect 3702 4324 3758 4380
rect 3758 4324 3762 4380
rect 3698 4320 3762 4324
rect 3778 4380 3842 4384
rect 3778 4324 3782 4380
rect 3782 4324 3838 4380
rect 3838 4324 3842 4380
rect 3778 4320 3842 4324
rect 3858 4380 3922 4384
rect 3858 4324 3862 4380
rect 3862 4324 3918 4380
rect 3918 4324 3922 4380
rect 3858 4320 3922 4324
rect 8952 4380 9016 4384
rect 8952 4324 8956 4380
rect 8956 4324 9012 4380
rect 9012 4324 9016 4380
rect 8952 4320 9016 4324
rect 9032 4380 9096 4384
rect 9032 4324 9036 4380
rect 9036 4324 9092 4380
rect 9092 4324 9096 4380
rect 9032 4320 9096 4324
rect 9112 4380 9176 4384
rect 9112 4324 9116 4380
rect 9116 4324 9172 4380
rect 9172 4324 9176 4380
rect 9112 4320 9176 4324
rect 9192 4380 9256 4384
rect 9192 4324 9196 4380
rect 9196 4324 9252 4380
rect 9252 4324 9256 4380
rect 9192 4320 9256 4324
rect 14285 4380 14349 4384
rect 14285 4324 14289 4380
rect 14289 4324 14345 4380
rect 14345 4324 14349 4380
rect 14285 4320 14349 4324
rect 14365 4380 14429 4384
rect 14365 4324 14369 4380
rect 14369 4324 14425 4380
rect 14425 4324 14429 4380
rect 14365 4320 14429 4324
rect 14445 4380 14509 4384
rect 14445 4324 14449 4380
rect 14449 4324 14505 4380
rect 14505 4324 14509 4380
rect 14445 4320 14509 4324
rect 14525 4380 14589 4384
rect 14525 4324 14529 4380
rect 14529 4324 14585 4380
rect 14585 4324 14589 4380
rect 14525 4320 14589 4324
rect 6285 3836 6349 3840
rect 6285 3780 6289 3836
rect 6289 3780 6345 3836
rect 6345 3780 6349 3836
rect 6285 3776 6349 3780
rect 6365 3836 6429 3840
rect 6365 3780 6369 3836
rect 6369 3780 6425 3836
rect 6425 3780 6429 3836
rect 6365 3776 6429 3780
rect 6445 3836 6509 3840
rect 6445 3780 6449 3836
rect 6449 3780 6505 3836
rect 6505 3780 6509 3836
rect 6445 3776 6509 3780
rect 6525 3836 6589 3840
rect 6525 3780 6529 3836
rect 6529 3780 6585 3836
rect 6585 3780 6589 3836
rect 6525 3776 6589 3780
rect 11618 3836 11682 3840
rect 11618 3780 11622 3836
rect 11622 3780 11678 3836
rect 11678 3780 11682 3836
rect 11618 3776 11682 3780
rect 11698 3836 11762 3840
rect 11698 3780 11702 3836
rect 11702 3780 11758 3836
rect 11758 3780 11762 3836
rect 11698 3776 11762 3780
rect 11778 3836 11842 3840
rect 11778 3780 11782 3836
rect 11782 3780 11838 3836
rect 11838 3780 11842 3836
rect 11778 3776 11842 3780
rect 11858 3836 11922 3840
rect 11858 3780 11862 3836
rect 11862 3780 11918 3836
rect 11918 3780 11922 3836
rect 11858 3776 11922 3780
rect 3618 3292 3682 3296
rect 3618 3236 3622 3292
rect 3622 3236 3678 3292
rect 3678 3236 3682 3292
rect 3618 3232 3682 3236
rect 3698 3292 3762 3296
rect 3698 3236 3702 3292
rect 3702 3236 3758 3292
rect 3758 3236 3762 3292
rect 3698 3232 3762 3236
rect 3778 3292 3842 3296
rect 3778 3236 3782 3292
rect 3782 3236 3838 3292
rect 3838 3236 3842 3292
rect 3778 3232 3842 3236
rect 3858 3292 3922 3296
rect 3858 3236 3862 3292
rect 3862 3236 3918 3292
rect 3918 3236 3922 3292
rect 3858 3232 3922 3236
rect 8952 3292 9016 3296
rect 8952 3236 8956 3292
rect 8956 3236 9012 3292
rect 9012 3236 9016 3292
rect 8952 3232 9016 3236
rect 9032 3292 9096 3296
rect 9032 3236 9036 3292
rect 9036 3236 9092 3292
rect 9092 3236 9096 3292
rect 9032 3232 9096 3236
rect 9112 3292 9176 3296
rect 9112 3236 9116 3292
rect 9116 3236 9172 3292
rect 9172 3236 9176 3292
rect 9112 3232 9176 3236
rect 9192 3292 9256 3296
rect 9192 3236 9196 3292
rect 9196 3236 9252 3292
rect 9252 3236 9256 3292
rect 9192 3232 9256 3236
rect 14285 3292 14349 3296
rect 14285 3236 14289 3292
rect 14289 3236 14345 3292
rect 14345 3236 14349 3292
rect 14285 3232 14349 3236
rect 14365 3292 14429 3296
rect 14365 3236 14369 3292
rect 14369 3236 14425 3292
rect 14425 3236 14429 3292
rect 14365 3232 14429 3236
rect 14445 3292 14509 3296
rect 14445 3236 14449 3292
rect 14449 3236 14505 3292
rect 14505 3236 14509 3292
rect 14445 3232 14509 3236
rect 14525 3292 14589 3296
rect 14525 3236 14529 3292
rect 14529 3236 14585 3292
rect 14585 3236 14589 3292
rect 14525 3232 14589 3236
rect 7972 3224 8036 3228
rect 7972 3168 7986 3224
rect 7986 3168 8036 3224
rect 7972 3164 8036 3168
rect 6285 2748 6349 2752
rect 6285 2692 6289 2748
rect 6289 2692 6345 2748
rect 6345 2692 6349 2748
rect 6285 2688 6349 2692
rect 6365 2748 6429 2752
rect 6365 2692 6369 2748
rect 6369 2692 6425 2748
rect 6425 2692 6429 2748
rect 6365 2688 6429 2692
rect 6445 2748 6509 2752
rect 6445 2692 6449 2748
rect 6449 2692 6505 2748
rect 6505 2692 6509 2748
rect 6445 2688 6509 2692
rect 6525 2748 6589 2752
rect 6525 2692 6529 2748
rect 6529 2692 6585 2748
rect 6585 2692 6589 2748
rect 6525 2688 6589 2692
rect 11618 2748 11682 2752
rect 11618 2692 11622 2748
rect 11622 2692 11678 2748
rect 11678 2692 11682 2748
rect 11618 2688 11682 2692
rect 11698 2748 11762 2752
rect 11698 2692 11702 2748
rect 11702 2692 11758 2748
rect 11758 2692 11762 2748
rect 11698 2688 11762 2692
rect 11778 2748 11842 2752
rect 11778 2692 11782 2748
rect 11782 2692 11838 2748
rect 11838 2692 11842 2748
rect 11778 2688 11842 2692
rect 11858 2748 11922 2752
rect 11858 2692 11862 2748
rect 11862 2692 11918 2748
rect 11918 2692 11922 2748
rect 11858 2688 11922 2692
rect 7420 2680 7484 2684
rect 7420 2624 7470 2680
rect 7470 2624 7484 2680
rect 7420 2620 7484 2624
rect 3618 2204 3682 2208
rect 3618 2148 3622 2204
rect 3622 2148 3678 2204
rect 3678 2148 3682 2204
rect 3618 2144 3682 2148
rect 3698 2204 3762 2208
rect 3698 2148 3702 2204
rect 3702 2148 3758 2204
rect 3758 2148 3762 2204
rect 3698 2144 3762 2148
rect 3778 2204 3842 2208
rect 3778 2148 3782 2204
rect 3782 2148 3838 2204
rect 3838 2148 3842 2204
rect 3778 2144 3842 2148
rect 3858 2204 3922 2208
rect 3858 2148 3862 2204
rect 3862 2148 3918 2204
rect 3918 2148 3922 2204
rect 3858 2144 3922 2148
rect 8952 2204 9016 2208
rect 8952 2148 8956 2204
rect 8956 2148 9012 2204
rect 9012 2148 9016 2204
rect 8952 2144 9016 2148
rect 9032 2204 9096 2208
rect 9032 2148 9036 2204
rect 9036 2148 9092 2204
rect 9092 2148 9096 2204
rect 9032 2144 9096 2148
rect 9112 2204 9176 2208
rect 9112 2148 9116 2204
rect 9116 2148 9172 2204
rect 9172 2148 9176 2204
rect 9112 2144 9176 2148
rect 9192 2204 9256 2208
rect 9192 2148 9196 2204
rect 9196 2148 9252 2204
rect 9252 2148 9256 2204
rect 9192 2144 9256 2148
rect 14285 2204 14349 2208
rect 14285 2148 14289 2204
rect 14289 2148 14345 2204
rect 14345 2148 14349 2204
rect 14285 2144 14349 2148
rect 14365 2204 14429 2208
rect 14365 2148 14369 2204
rect 14369 2148 14425 2204
rect 14425 2148 14429 2204
rect 14365 2144 14429 2148
rect 14445 2204 14509 2208
rect 14445 2148 14449 2204
rect 14449 2148 14505 2204
rect 14505 2148 14509 2204
rect 14445 2144 14509 2148
rect 14525 2204 14589 2208
rect 14525 2148 14529 2204
rect 14529 2148 14585 2204
rect 14585 2148 14589 2204
rect 14525 2144 14589 2148
<< metal4 >>
rect 3610 37024 3931 37584
rect 3610 36960 3618 37024
rect 3682 36960 3698 37024
rect 3762 36960 3778 37024
rect 3842 36960 3858 37024
rect 3922 36960 3931 37024
rect 3610 35936 3931 36960
rect 3610 35872 3618 35936
rect 3682 35872 3698 35936
rect 3762 35872 3778 35936
rect 3842 35872 3858 35936
rect 3922 35872 3931 35936
rect 3610 34848 3931 35872
rect 3610 34784 3618 34848
rect 3682 34784 3698 34848
rect 3762 34784 3778 34848
rect 3842 34784 3858 34848
rect 3922 34784 3931 34848
rect 3610 33760 3931 34784
rect 3610 33696 3618 33760
rect 3682 33696 3698 33760
rect 3762 33696 3778 33760
rect 3842 33696 3858 33760
rect 3922 33696 3931 33760
rect 3610 32672 3931 33696
rect 3610 32608 3618 32672
rect 3682 32608 3698 32672
rect 3762 32608 3778 32672
rect 3842 32608 3858 32672
rect 3922 32608 3931 32672
rect 3610 31584 3931 32608
rect 3610 31520 3618 31584
rect 3682 31520 3698 31584
rect 3762 31520 3778 31584
rect 3842 31520 3858 31584
rect 3922 31520 3931 31584
rect 3610 30496 3931 31520
rect 3610 30432 3618 30496
rect 3682 30432 3698 30496
rect 3762 30432 3778 30496
rect 3842 30432 3858 30496
rect 3922 30432 3931 30496
rect 3610 29408 3931 30432
rect 3610 29344 3618 29408
rect 3682 29344 3698 29408
rect 3762 29344 3778 29408
rect 3842 29344 3858 29408
rect 3922 29344 3931 29408
rect 3610 28320 3931 29344
rect 3610 28256 3618 28320
rect 3682 28256 3698 28320
rect 3762 28256 3778 28320
rect 3842 28256 3858 28320
rect 3922 28256 3931 28320
rect 3610 27232 3931 28256
rect 3610 27168 3618 27232
rect 3682 27168 3698 27232
rect 3762 27168 3778 27232
rect 3842 27168 3858 27232
rect 3922 27168 3931 27232
rect 3610 26144 3931 27168
rect 3610 26080 3618 26144
rect 3682 26080 3698 26144
rect 3762 26080 3778 26144
rect 3842 26080 3858 26144
rect 3922 26080 3931 26144
rect 3610 25056 3931 26080
rect 3610 24992 3618 25056
rect 3682 24992 3698 25056
rect 3762 24992 3778 25056
rect 3842 24992 3858 25056
rect 3922 24992 3931 25056
rect 3610 23968 3931 24992
rect 6277 37568 6597 37584
rect 6277 37504 6285 37568
rect 6349 37504 6365 37568
rect 6429 37504 6445 37568
rect 6509 37504 6525 37568
rect 6589 37504 6597 37568
rect 6277 36480 6597 37504
rect 6277 36416 6285 36480
rect 6349 36416 6365 36480
rect 6429 36416 6445 36480
rect 6509 36416 6525 36480
rect 6589 36416 6597 36480
rect 6277 35392 6597 36416
rect 6277 35328 6285 35392
rect 6349 35328 6365 35392
rect 6429 35328 6445 35392
rect 6509 35328 6525 35392
rect 6589 35328 6597 35392
rect 6277 34304 6597 35328
rect 6277 34240 6285 34304
rect 6349 34240 6365 34304
rect 6429 34240 6445 34304
rect 6509 34240 6525 34304
rect 6589 34240 6597 34304
rect 6277 33216 6597 34240
rect 6277 33152 6285 33216
rect 6349 33152 6365 33216
rect 6429 33152 6445 33216
rect 6509 33152 6525 33216
rect 6589 33152 6597 33216
rect 6277 32128 6597 33152
rect 6277 32064 6285 32128
rect 6349 32064 6365 32128
rect 6429 32064 6445 32128
rect 6509 32064 6525 32128
rect 6589 32064 6597 32128
rect 6277 31040 6597 32064
rect 6277 30976 6285 31040
rect 6349 30976 6365 31040
rect 6429 30976 6445 31040
rect 6509 30976 6525 31040
rect 6589 30976 6597 31040
rect 6277 29952 6597 30976
rect 6277 29888 6285 29952
rect 6349 29888 6365 29952
rect 6429 29888 6445 29952
rect 6509 29888 6525 29952
rect 6589 29888 6597 29952
rect 6277 28864 6597 29888
rect 6277 28800 6285 28864
rect 6349 28800 6365 28864
rect 6429 28800 6445 28864
rect 6509 28800 6525 28864
rect 6589 28800 6597 28864
rect 6277 27776 6597 28800
rect 6277 27712 6285 27776
rect 6349 27712 6365 27776
rect 6429 27712 6445 27776
rect 6509 27712 6525 27776
rect 6589 27712 6597 27776
rect 6277 26688 6597 27712
rect 6277 26624 6285 26688
rect 6349 26624 6365 26688
rect 6429 26624 6445 26688
rect 6509 26624 6525 26688
rect 6589 26624 6597 26688
rect 6277 25600 6597 26624
rect 6277 25536 6285 25600
rect 6349 25536 6365 25600
rect 6429 25536 6445 25600
rect 6509 25536 6525 25600
rect 6589 25536 6597 25600
rect 5763 24988 5829 24989
rect 5763 24924 5764 24988
rect 5828 24924 5829 24988
rect 5763 24923 5829 24924
rect 3610 23904 3618 23968
rect 3682 23904 3698 23968
rect 3762 23904 3778 23968
rect 3842 23904 3858 23968
rect 3922 23904 3931 23968
rect 3610 22880 3931 23904
rect 3610 22816 3618 22880
rect 3682 22816 3698 22880
rect 3762 22816 3778 22880
rect 3842 22816 3858 22880
rect 3922 22816 3931 22880
rect 3610 21792 3931 22816
rect 3610 21728 3618 21792
rect 3682 21728 3698 21792
rect 3762 21728 3778 21792
rect 3842 21728 3858 21792
rect 3922 21728 3931 21792
rect 3610 20704 3931 21728
rect 5766 21317 5826 24923
rect 6277 24512 6597 25536
rect 6277 24448 6285 24512
rect 6349 24448 6365 24512
rect 6429 24448 6445 24512
rect 6509 24448 6525 24512
rect 6589 24448 6597 24512
rect 6277 23424 6597 24448
rect 6277 23360 6285 23424
rect 6349 23360 6365 23424
rect 6429 23360 6445 23424
rect 6509 23360 6525 23424
rect 6589 23360 6597 23424
rect 6277 22336 6597 23360
rect 6277 22272 6285 22336
rect 6349 22272 6365 22336
rect 6429 22272 6445 22336
rect 6509 22272 6525 22336
rect 6589 22272 6597 22336
rect 5763 21316 5829 21317
rect 5763 21252 5764 21316
rect 5828 21252 5829 21316
rect 5763 21251 5829 21252
rect 3610 20640 3618 20704
rect 3682 20640 3698 20704
rect 3762 20640 3778 20704
rect 3842 20640 3858 20704
rect 3922 20640 3931 20704
rect 3610 19616 3931 20640
rect 3610 19552 3618 19616
rect 3682 19552 3698 19616
rect 3762 19552 3778 19616
rect 3842 19552 3858 19616
rect 3922 19552 3931 19616
rect 3610 18528 3931 19552
rect 3610 18464 3618 18528
rect 3682 18464 3698 18528
rect 3762 18464 3778 18528
rect 3842 18464 3858 18528
rect 3922 18464 3931 18528
rect 3610 17440 3931 18464
rect 3610 17376 3618 17440
rect 3682 17376 3698 17440
rect 3762 17376 3778 17440
rect 3842 17376 3858 17440
rect 3922 17376 3931 17440
rect 3610 16352 3931 17376
rect 6277 21248 6597 22272
rect 6277 21184 6285 21248
rect 6349 21184 6365 21248
rect 6429 21184 6445 21248
rect 6509 21184 6525 21248
rect 6589 21184 6597 21248
rect 6277 20160 6597 21184
rect 6277 20096 6285 20160
rect 6349 20096 6365 20160
rect 6429 20096 6445 20160
rect 6509 20096 6525 20160
rect 6589 20096 6597 20160
rect 6277 19072 6597 20096
rect 6277 19008 6285 19072
rect 6349 19008 6365 19072
rect 6429 19008 6445 19072
rect 6509 19008 6525 19072
rect 6589 19008 6597 19072
rect 6277 17984 6597 19008
rect 6277 17920 6285 17984
rect 6349 17920 6365 17984
rect 6429 17920 6445 17984
rect 6509 17920 6525 17984
rect 6589 17920 6597 17984
rect 5027 17236 5093 17237
rect 5027 17172 5028 17236
rect 5092 17172 5093 17236
rect 5027 17171 5093 17172
rect 3610 16288 3618 16352
rect 3682 16288 3698 16352
rect 3762 16288 3778 16352
rect 3842 16288 3858 16352
rect 3922 16288 3931 16352
rect 3610 15264 3931 16288
rect 3610 15200 3618 15264
rect 3682 15200 3698 15264
rect 3762 15200 3778 15264
rect 3842 15200 3858 15264
rect 3922 15200 3931 15264
rect 3610 14176 3931 15200
rect 3610 14112 3618 14176
rect 3682 14112 3698 14176
rect 3762 14112 3778 14176
rect 3842 14112 3858 14176
rect 3922 14112 3931 14176
rect 3610 13088 3931 14112
rect 3610 13024 3618 13088
rect 3682 13024 3698 13088
rect 3762 13024 3778 13088
rect 3842 13024 3858 13088
rect 3922 13024 3931 13088
rect 3610 12000 3931 13024
rect 3610 11936 3618 12000
rect 3682 11936 3698 12000
rect 3762 11936 3778 12000
rect 3842 11936 3858 12000
rect 3922 11936 3931 12000
rect 3610 10912 3931 11936
rect 5030 11661 5090 17171
rect 6277 16896 6597 17920
rect 6277 16832 6285 16896
rect 6349 16832 6365 16896
rect 6429 16832 6445 16896
rect 6509 16832 6525 16896
rect 6589 16832 6597 16896
rect 6277 15808 6597 16832
rect 6277 15744 6285 15808
rect 6349 15744 6365 15808
rect 6429 15744 6445 15808
rect 6509 15744 6525 15808
rect 6589 15744 6597 15808
rect 6277 14720 6597 15744
rect 6277 14656 6285 14720
rect 6349 14656 6365 14720
rect 6429 14656 6445 14720
rect 6509 14656 6525 14720
rect 6589 14656 6597 14720
rect 6277 13632 6597 14656
rect 6277 13568 6285 13632
rect 6349 13568 6365 13632
rect 6429 13568 6445 13632
rect 6509 13568 6525 13632
rect 6589 13568 6597 13632
rect 6277 12544 6597 13568
rect 6277 12480 6285 12544
rect 6349 12480 6365 12544
rect 6429 12480 6445 12544
rect 6509 12480 6525 12544
rect 6589 12480 6597 12544
rect 5027 11660 5093 11661
rect 5027 11596 5028 11660
rect 5092 11596 5093 11660
rect 5027 11595 5093 11596
rect 3610 10848 3618 10912
rect 3682 10848 3698 10912
rect 3762 10848 3778 10912
rect 3842 10848 3858 10912
rect 3922 10848 3931 10912
rect 3610 9824 3931 10848
rect 3610 9760 3618 9824
rect 3682 9760 3698 9824
rect 3762 9760 3778 9824
rect 3842 9760 3858 9824
rect 3922 9760 3931 9824
rect 3610 8736 3931 9760
rect 3610 8672 3618 8736
rect 3682 8672 3698 8736
rect 3762 8672 3778 8736
rect 3842 8672 3858 8736
rect 3922 8672 3931 8736
rect 3610 7648 3931 8672
rect 3610 7584 3618 7648
rect 3682 7584 3698 7648
rect 3762 7584 3778 7648
rect 3842 7584 3858 7648
rect 3922 7584 3931 7648
rect 3610 6560 3931 7584
rect 3610 6496 3618 6560
rect 3682 6496 3698 6560
rect 3762 6496 3778 6560
rect 3842 6496 3858 6560
rect 3922 6496 3931 6560
rect 3610 5472 3931 6496
rect 3610 5408 3618 5472
rect 3682 5408 3698 5472
rect 3762 5408 3778 5472
rect 3842 5408 3858 5472
rect 3922 5408 3931 5472
rect 3610 4384 3931 5408
rect 3610 4320 3618 4384
rect 3682 4320 3698 4384
rect 3762 4320 3778 4384
rect 3842 4320 3858 4384
rect 3922 4320 3931 4384
rect 3610 3296 3931 4320
rect 3610 3232 3618 3296
rect 3682 3232 3698 3296
rect 3762 3232 3778 3296
rect 3842 3232 3858 3296
rect 3922 3232 3931 3296
rect 3610 2208 3931 3232
rect 3610 2144 3618 2208
rect 3682 2144 3698 2208
rect 3762 2144 3778 2208
rect 3842 2144 3858 2208
rect 3922 2144 3931 2208
rect 3610 2128 3931 2144
rect 6277 11456 6597 12480
rect 6277 11392 6285 11456
rect 6349 11392 6365 11456
rect 6429 11392 6445 11456
rect 6509 11392 6525 11456
rect 6589 11392 6597 11456
rect 6277 10368 6597 11392
rect 6277 10304 6285 10368
rect 6349 10304 6365 10368
rect 6429 10304 6445 10368
rect 6509 10304 6525 10368
rect 6589 10304 6597 10368
rect 6277 9280 6597 10304
rect 6277 9216 6285 9280
rect 6349 9216 6365 9280
rect 6429 9216 6445 9280
rect 6509 9216 6525 9280
rect 6589 9216 6597 9280
rect 6277 8192 6597 9216
rect 8944 37024 9264 37584
rect 8944 36960 8952 37024
rect 9016 36960 9032 37024
rect 9096 36960 9112 37024
rect 9176 36960 9192 37024
rect 9256 36960 9264 37024
rect 8944 35936 9264 36960
rect 8944 35872 8952 35936
rect 9016 35872 9032 35936
rect 9096 35872 9112 35936
rect 9176 35872 9192 35936
rect 9256 35872 9264 35936
rect 8944 34848 9264 35872
rect 8944 34784 8952 34848
rect 9016 34784 9032 34848
rect 9096 34784 9112 34848
rect 9176 34784 9192 34848
rect 9256 34784 9264 34848
rect 8944 33760 9264 34784
rect 8944 33696 8952 33760
rect 9016 33696 9032 33760
rect 9096 33696 9112 33760
rect 9176 33696 9192 33760
rect 9256 33696 9264 33760
rect 8944 32672 9264 33696
rect 8944 32608 8952 32672
rect 9016 32608 9032 32672
rect 9096 32608 9112 32672
rect 9176 32608 9192 32672
rect 9256 32608 9264 32672
rect 8944 31584 9264 32608
rect 8944 31520 8952 31584
rect 9016 31520 9032 31584
rect 9096 31520 9112 31584
rect 9176 31520 9192 31584
rect 9256 31520 9264 31584
rect 8944 30496 9264 31520
rect 8944 30432 8952 30496
rect 9016 30432 9032 30496
rect 9096 30432 9112 30496
rect 9176 30432 9192 30496
rect 9256 30432 9264 30496
rect 8944 29408 9264 30432
rect 8944 29344 8952 29408
rect 9016 29344 9032 29408
rect 9096 29344 9112 29408
rect 9176 29344 9192 29408
rect 9256 29344 9264 29408
rect 8944 28320 9264 29344
rect 11610 37568 11930 37584
rect 11610 37504 11618 37568
rect 11682 37504 11698 37568
rect 11762 37504 11778 37568
rect 11842 37504 11858 37568
rect 11922 37504 11930 37568
rect 11610 36480 11930 37504
rect 11610 36416 11618 36480
rect 11682 36416 11698 36480
rect 11762 36416 11778 36480
rect 11842 36416 11858 36480
rect 11922 36416 11930 36480
rect 11610 35392 11930 36416
rect 11610 35328 11618 35392
rect 11682 35328 11698 35392
rect 11762 35328 11778 35392
rect 11842 35328 11858 35392
rect 11922 35328 11930 35392
rect 11610 34304 11930 35328
rect 11610 34240 11618 34304
rect 11682 34240 11698 34304
rect 11762 34240 11778 34304
rect 11842 34240 11858 34304
rect 11922 34240 11930 34304
rect 11610 33216 11930 34240
rect 11610 33152 11618 33216
rect 11682 33152 11698 33216
rect 11762 33152 11778 33216
rect 11842 33152 11858 33216
rect 11922 33152 11930 33216
rect 11610 32128 11930 33152
rect 11610 32064 11618 32128
rect 11682 32064 11698 32128
rect 11762 32064 11778 32128
rect 11842 32064 11858 32128
rect 11922 32064 11930 32128
rect 11610 31040 11930 32064
rect 11610 30976 11618 31040
rect 11682 30976 11698 31040
rect 11762 30976 11778 31040
rect 11842 30976 11858 31040
rect 11922 30976 11930 31040
rect 11610 29952 11930 30976
rect 11610 29888 11618 29952
rect 11682 29888 11698 29952
rect 11762 29888 11778 29952
rect 11842 29888 11858 29952
rect 11922 29888 11930 29952
rect 11610 28864 11930 29888
rect 11610 28800 11618 28864
rect 11682 28800 11698 28864
rect 11762 28800 11778 28864
rect 11842 28800 11858 28864
rect 11922 28800 11930 28864
rect 9443 28796 9509 28797
rect 9443 28732 9444 28796
rect 9508 28732 9509 28796
rect 9443 28731 9509 28732
rect 8944 28256 8952 28320
rect 9016 28256 9032 28320
rect 9096 28256 9112 28320
rect 9176 28256 9192 28320
rect 9256 28256 9264 28320
rect 8944 27232 9264 28256
rect 8944 27168 8952 27232
rect 9016 27168 9032 27232
rect 9096 27168 9112 27232
rect 9176 27168 9192 27232
rect 9256 27168 9264 27232
rect 8944 26144 9264 27168
rect 8944 26080 8952 26144
rect 9016 26080 9032 26144
rect 9096 26080 9112 26144
rect 9176 26080 9192 26144
rect 9256 26080 9264 26144
rect 8944 25056 9264 26080
rect 8944 24992 8952 25056
rect 9016 24992 9032 25056
rect 9096 24992 9112 25056
rect 9176 24992 9192 25056
rect 9256 24992 9264 25056
rect 8944 23968 9264 24992
rect 8944 23904 8952 23968
rect 9016 23904 9032 23968
rect 9096 23904 9112 23968
rect 9176 23904 9192 23968
rect 9256 23904 9264 23968
rect 8944 22880 9264 23904
rect 8944 22816 8952 22880
rect 9016 22816 9032 22880
rect 9096 22816 9112 22880
rect 9176 22816 9192 22880
rect 9256 22816 9264 22880
rect 8944 21792 9264 22816
rect 8944 21728 8952 21792
rect 9016 21728 9032 21792
rect 9096 21728 9112 21792
rect 9176 21728 9192 21792
rect 9256 21728 9264 21792
rect 8944 20704 9264 21728
rect 8944 20640 8952 20704
rect 9016 20640 9032 20704
rect 9096 20640 9112 20704
rect 9176 20640 9192 20704
rect 9256 20640 9264 20704
rect 8944 19616 9264 20640
rect 9446 20365 9506 28731
rect 11610 27776 11930 28800
rect 11610 27712 11618 27776
rect 11682 27712 11698 27776
rect 11762 27712 11778 27776
rect 11842 27712 11858 27776
rect 11922 27712 11930 27776
rect 11610 26688 11930 27712
rect 14277 37024 14597 37584
rect 14277 36960 14285 37024
rect 14349 36960 14365 37024
rect 14429 36960 14445 37024
rect 14509 36960 14525 37024
rect 14589 36960 14597 37024
rect 14277 35936 14597 36960
rect 14277 35872 14285 35936
rect 14349 35872 14365 35936
rect 14429 35872 14445 35936
rect 14509 35872 14525 35936
rect 14589 35872 14597 35936
rect 14277 34848 14597 35872
rect 14277 34784 14285 34848
rect 14349 34784 14365 34848
rect 14429 34784 14445 34848
rect 14509 34784 14525 34848
rect 14589 34784 14597 34848
rect 14277 33760 14597 34784
rect 14277 33696 14285 33760
rect 14349 33696 14365 33760
rect 14429 33696 14445 33760
rect 14509 33696 14525 33760
rect 14589 33696 14597 33760
rect 14277 32672 14597 33696
rect 14277 32608 14285 32672
rect 14349 32608 14365 32672
rect 14429 32608 14445 32672
rect 14509 32608 14525 32672
rect 14589 32608 14597 32672
rect 14277 31584 14597 32608
rect 14277 31520 14285 31584
rect 14349 31520 14365 31584
rect 14429 31520 14445 31584
rect 14509 31520 14525 31584
rect 14589 31520 14597 31584
rect 14277 30496 14597 31520
rect 14277 30432 14285 30496
rect 14349 30432 14365 30496
rect 14429 30432 14445 30496
rect 14509 30432 14525 30496
rect 14589 30432 14597 30496
rect 14277 29408 14597 30432
rect 14277 29344 14285 29408
rect 14349 29344 14365 29408
rect 14429 29344 14445 29408
rect 14509 29344 14525 29408
rect 14589 29344 14597 29408
rect 14277 28320 14597 29344
rect 14277 28256 14285 28320
rect 14349 28256 14365 28320
rect 14429 28256 14445 28320
rect 14509 28256 14525 28320
rect 14589 28256 14597 28320
rect 12019 27708 12085 27709
rect 12019 27644 12020 27708
rect 12084 27644 12085 27708
rect 12019 27643 12085 27644
rect 11610 26624 11618 26688
rect 11682 26624 11698 26688
rect 11762 26624 11778 26688
rect 11842 26624 11858 26688
rect 11922 26624 11930 26688
rect 11610 25600 11930 26624
rect 11610 25536 11618 25600
rect 11682 25536 11698 25600
rect 11762 25536 11778 25600
rect 11842 25536 11858 25600
rect 11922 25536 11930 25600
rect 11610 24512 11930 25536
rect 11610 24448 11618 24512
rect 11682 24448 11698 24512
rect 11762 24448 11778 24512
rect 11842 24448 11858 24512
rect 11922 24448 11930 24512
rect 11610 23424 11930 24448
rect 11610 23360 11618 23424
rect 11682 23360 11698 23424
rect 11762 23360 11778 23424
rect 11842 23360 11858 23424
rect 11922 23360 11930 23424
rect 11610 22336 11930 23360
rect 11610 22272 11618 22336
rect 11682 22272 11698 22336
rect 11762 22272 11778 22336
rect 11842 22272 11858 22336
rect 11922 22272 11930 22336
rect 11610 21248 11930 22272
rect 11610 21184 11618 21248
rect 11682 21184 11698 21248
rect 11762 21184 11778 21248
rect 11842 21184 11858 21248
rect 11922 21184 11930 21248
rect 9443 20364 9509 20365
rect 9443 20300 9444 20364
rect 9508 20300 9509 20364
rect 9443 20299 9509 20300
rect 8944 19552 8952 19616
rect 9016 19552 9032 19616
rect 9096 19552 9112 19616
rect 9176 19552 9192 19616
rect 9256 19552 9264 19616
rect 8944 18528 9264 19552
rect 8944 18464 8952 18528
rect 9016 18464 9032 18528
rect 9096 18464 9112 18528
rect 9176 18464 9192 18528
rect 9256 18464 9264 18528
rect 8944 17440 9264 18464
rect 8944 17376 8952 17440
rect 9016 17376 9032 17440
rect 9096 17376 9112 17440
rect 9176 17376 9192 17440
rect 9256 17376 9264 17440
rect 8944 16352 9264 17376
rect 8944 16288 8952 16352
rect 9016 16288 9032 16352
rect 9096 16288 9112 16352
rect 9176 16288 9192 16352
rect 9256 16288 9264 16352
rect 8944 15264 9264 16288
rect 8944 15200 8952 15264
rect 9016 15200 9032 15264
rect 9096 15200 9112 15264
rect 9176 15200 9192 15264
rect 9256 15200 9264 15264
rect 8944 14176 9264 15200
rect 8944 14112 8952 14176
rect 9016 14112 9032 14176
rect 9096 14112 9112 14176
rect 9176 14112 9192 14176
rect 9256 14112 9264 14176
rect 8944 13088 9264 14112
rect 8944 13024 8952 13088
rect 9016 13024 9032 13088
rect 9096 13024 9112 13088
rect 9176 13024 9192 13088
rect 9256 13024 9264 13088
rect 8944 12000 9264 13024
rect 8944 11936 8952 12000
rect 9016 11936 9032 12000
rect 9096 11936 9112 12000
rect 9176 11936 9192 12000
rect 9256 11936 9264 12000
rect 8944 10912 9264 11936
rect 8944 10848 8952 10912
rect 9016 10848 9032 10912
rect 9096 10848 9112 10912
rect 9176 10848 9192 10912
rect 9256 10848 9264 10912
rect 8944 9824 9264 10848
rect 8944 9760 8952 9824
rect 9016 9760 9032 9824
rect 9096 9760 9112 9824
rect 9176 9760 9192 9824
rect 9256 9760 9264 9824
rect 7971 9076 8037 9077
rect 7971 9012 7972 9076
rect 8036 9012 8037 9076
rect 7971 9011 8037 9012
rect 6277 8128 6285 8192
rect 6349 8128 6365 8192
rect 6429 8128 6445 8192
rect 6509 8128 6525 8192
rect 6589 8128 6597 8192
rect 6277 7104 6597 8128
rect 7419 7988 7485 7989
rect 7419 7924 7420 7988
rect 7484 7924 7485 7988
rect 7419 7923 7485 7924
rect 6277 7040 6285 7104
rect 6349 7040 6365 7104
rect 6429 7040 6445 7104
rect 6509 7040 6525 7104
rect 6589 7040 6597 7104
rect 6277 6016 6597 7040
rect 6277 5952 6285 6016
rect 6349 5952 6365 6016
rect 6429 5952 6445 6016
rect 6509 5952 6525 6016
rect 6589 5952 6597 6016
rect 6277 4928 6597 5952
rect 6277 4864 6285 4928
rect 6349 4864 6365 4928
rect 6429 4864 6445 4928
rect 6509 4864 6525 4928
rect 6589 4864 6597 4928
rect 6277 3840 6597 4864
rect 6277 3776 6285 3840
rect 6349 3776 6365 3840
rect 6429 3776 6445 3840
rect 6509 3776 6525 3840
rect 6589 3776 6597 3840
rect 6277 2752 6597 3776
rect 6277 2688 6285 2752
rect 6349 2688 6365 2752
rect 6429 2688 6445 2752
rect 6509 2688 6525 2752
rect 6589 2688 6597 2752
rect 6277 2128 6597 2688
rect 7422 2685 7482 7923
rect 7974 3229 8034 9011
rect 8944 8736 9264 9760
rect 8944 8672 8952 8736
rect 9016 8672 9032 8736
rect 9096 8672 9112 8736
rect 9176 8672 9192 8736
rect 9256 8672 9264 8736
rect 8944 7648 9264 8672
rect 8944 7584 8952 7648
rect 9016 7584 9032 7648
rect 9096 7584 9112 7648
rect 9176 7584 9192 7648
rect 9256 7584 9264 7648
rect 8944 6560 9264 7584
rect 8944 6496 8952 6560
rect 9016 6496 9032 6560
rect 9096 6496 9112 6560
rect 9176 6496 9192 6560
rect 9256 6496 9264 6560
rect 8944 5472 9264 6496
rect 8944 5408 8952 5472
rect 9016 5408 9032 5472
rect 9096 5408 9112 5472
rect 9176 5408 9192 5472
rect 9256 5408 9264 5472
rect 8944 4384 9264 5408
rect 8944 4320 8952 4384
rect 9016 4320 9032 4384
rect 9096 4320 9112 4384
rect 9176 4320 9192 4384
rect 9256 4320 9264 4384
rect 8944 3296 9264 4320
rect 8944 3232 8952 3296
rect 9016 3232 9032 3296
rect 9096 3232 9112 3296
rect 9176 3232 9192 3296
rect 9256 3232 9264 3296
rect 7971 3228 8037 3229
rect 7971 3164 7972 3228
rect 8036 3164 8037 3228
rect 7971 3163 8037 3164
rect 7419 2684 7485 2685
rect 7419 2620 7420 2684
rect 7484 2620 7485 2684
rect 7419 2619 7485 2620
rect 8944 2208 9264 3232
rect 8944 2144 8952 2208
rect 9016 2144 9032 2208
rect 9096 2144 9112 2208
rect 9176 2144 9192 2208
rect 9256 2144 9264 2208
rect 8944 2128 9264 2144
rect 11610 20160 11930 21184
rect 11610 20096 11618 20160
rect 11682 20096 11698 20160
rect 11762 20096 11778 20160
rect 11842 20096 11858 20160
rect 11922 20096 11930 20160
rect 11610 19072 11930 20096
rect 12022 19957 12082 27643
rect 14277 27232 14597 28256
rect 14277 27168 14285 27232
rect 14349 27168 14365 27232
rect 14429 27168 14445 27232
rect 14509 27168 14525 27232
rect 14589 27168 14597 27232
rect 14277 26144 14597 27168
rect 14277 26080 14285 26144
rect 14349 26080 14365 26144
rect 14429 26080 14445 26144
rect 14509 26080 14525 26144
rect 14589 26080 14597 26144
rect 14277 25056 14597 26080
rect 14277 24992 14285 25056
rect 14349 24992 14365 25056
rect 14429 24992 14445 25056
rect 14509 24992 14525 25056
rect 14589 24992 14597 25056
rect 14277 23968 14597 24992
rect 14277 23904 14285 23968
rect 14349 23904 14365 23968
rect 14429 23904 14445 23968
rect 14509 23904 14525 23968
rect 14589 23904 14597 23968
rect 14277 22880 14597 23904
rect 14277 22816 14285 22880
rect 14349 22816 14365 22880
rect 14429 22816 14445 22880
rect 14509 22816 14525 22880
rect 14589 22816 14597 22880
rect 14277 21792 14597 22816
rect 14277 21728 14285 21792
rect 14349 21728 14365 21792
rect 14429 21728 14445 21792
rect 14509 21728 14525 21792
rect 14589 21728 14597 21792
rect 14277 20704 14597 21728
rect 14277 20640 14285 20704
rect 14349 20640 14365 20704
rect 14429 20640 14445 20704
rect 14509 20640 14525 20704
rect 14589 20640 14597 20704
rect 12019 19956 12085 19957
rect 12019 19892 12020 19956
rect 12084 19892 12085 19956
rect 12019 19891 12085 19892
rect 11610 19008 11618 19072
rect 11682 19008 11698 19072
rect 11762 19008 11778 19072
rect 11842 19008 11858 19072
rect 11922 19008 11930 19072
rect 11610 17984 11930 19008
rect 11610 17920 11618 17984
rect 11682 17920 11698 17984
rect 11762 17920 11778 17984
rect 11842 17920 11858 17984
rect 11922 17920 11930 17984
rect 11610 16896 11930 17920
rect 11610 16832 11618 16896
rect 11682 16832 11698 16896
rect 11762 16832 11778 16896
rect 11842 16832 11858 16896
rect 11922 16832 11930 16896
rect 11610 15808 11930 16832
rect 11610 15744 11618 15808
rect 11682 15744 11698 15808
rect 11762 15744 11778 15808
rect 11842 15744 11858 15808
rect 11922 15744 11930 15808
rect 11610 14720 11930 15744
rect 11610 14656 11618 14720
rect 11682 14656 11698 14720
rect 11762 14656 11778 14720
rect 11842 14656 11858 14720
rect 11922 14656 11930 14720
rect 11610 13632 11930 14656
rect 11610 13568 11618 13632
rect 11682 13568 11698 13632
rect 11762 13568 11778 13632
rect 11842 13568 11858 13632
rect 11922 13568 11930 13632
rect 11610 12544 11930 13568
rect 11610 12480 11618 12544
rect 11682 12480 11698 12544
rect 11762 12480 11778 12544
rect 11842 12480 11858 12544
rect 11922 12480 11930 12544
rect 11610 11456 11930 12480
rect 11610 11392 11618 11456
rect 11682 11392 11698 11456
rect 11762 11392 11778 11456
rect 11842 11392 11858 11456
rect 11922 11392 11930 11456
rect 11610 10368 11930 11392
rect 11610 10304 11618 10368
rect 11682 10304 11698 10368
rect 11762 10304 11778 10368
rect 11842 10304 11858 10368
rect 11922 10304 11930 10368
rect 11610 9280 11930 10304
rect 11610 9216 11618 9280
rect 11682 9216 11698 9280
rect 11762 9216 11778 9280
rect 11842 9216 11858 9280
rect 11922 9216 11930 9280
rect 11610 8192 11930 9216
rect 11610 8128 11618 8192
rect 11682 8128 11698 8192
rect 11762 8128 11778 8192
rect 11842 8128 11858 8192
rect 11922 8128 11930 8192
rect 11610 7104 11930 8128
rect 11610 7040 11618 7104
rect 11682 7040 11698 7104
rect 11762 7040 11778 7104
rect 11842 7040 11858 7104
rect 11922 7040 11930 7104
rect 11610 6016 11930 7040
rect 11610 5952 11618 6016
rect 11682 5952 11698 6016
rect 11762 5952 11778 6016
rect 11842 5952 11858 6016
rect 11922 5952 11930 6016
rect 11610 4928 11930 5952
rect 11610 4864 11618 4928
rect 11682 4864 11698 4928
rect 11762 4864 11778 4928
rect 11842 4864 11858 4928
rect 11922 4864 11930 4928
rect 11610 3840 11930 4864
rect 11610 3776 11618 3840
rect 11682 3776 11698 3840
rect 11762 3776 11778 3840
rect 11842 3776 11858 3840
rect 11922 3776 11930 3840
rect 11610 2752 11930 3776
rect 11610 2688 11618 2752
rect 11682 2688 11698 2752
rect 11762 2688 11778 2752
rect 11842 2688 11858 2752
rect 11922 2688 11930 2752
rect 11610 2128 11930 2688
rect 14277 19616 14597 20640
rect 14277 19552 14285 19616
rect 14349 19552 14365 19616
rect 14429 19552 14445 19616
rect 14509 19552 14525 19616
rect 14589 19552 14597 19616
rect 14277 18528 14597 19552
rect 14277 18464 14285 18528
rect 14349 18464 14365 18528
rect 14429 18464 14445 18528
rect 14509 18464 14525 18528
rect 14589 18464 14597 18528
rect 14277 17440 14597 18464
rect 14277 17376 14285 17440
rect 14349 17376 14365 17440
rect 14429 17376 14445 17440
rect 14509 17376 14525 17440
rect 14589 17376 14597 17440
rect 14277 16352 14597 17376
rect 14277 16288 14285 16352
rect 14349 16288 14365 16352
rect 14429 16288 14445 16352
rect 14509 16288 14525 16352
rect 14589 16288 14597 16352
rect 14277 15264 14597 16288
rect 14277 15200 14285 15264
rect 14349 15200 14365 15264
rect 14429 15200 14445 15264
rect 14509 15200 14525 15264
rect 14589 15200 14597 15264
rect 14277 14176 14597 15200
rect 14277 14112 14285 14176
rect 14349 14112 14365 14176
rect 14429 14112 14445 14176
rect 14509 14112 14525 14176
rect 14589 14112 14597 14176
rect 14277 13088 14597 14112
rect 14277 13024 14285 13088
rect 14349 13024 14365 13088
rect 14429 13024 14445 13088
rect 14509 13024 14525 13088
rect 14589 13024 14597 13088
rect 14277 12000 14597 13024
rect 14277 11936 14285 12000
rect 14349 11936 14365 12000
rect 14429 11936 14445 12000
rect 14509 11936 14525 12000
rect 14589 11936 14597 12000
rect 14277 10912 14597 11936
rect 14277 10848 14285 10912
rect 14349 10848 14365 10912
rect 14429 10848 14445 10912
rect 14509 10848 14525 10912
rect 14589 10848 14597 10912
rect 14277 9824 14597 10848
rect 14277 9760 14285 9824
rect 14349 9760 14365 9824
rect 14429 9760 14445 9824
rect 14509 9760 14525 9824
rect 14589 9760 14597 9824
rect 14277 8736 14597 9760
rect 14277 8672 14285 8736
rect 14349 8672 14365 8736
rect 14429 8672 14445 8736
rect 14509 8672 14525 8736
rect 14589 8672 14597 8736
rect 14277 7648 14597 8672
rect 14277 7584 14285 7648
rect 14349 7584 14365 7648
rect 14429 7584 14445 7648
rect 14509 7584 14525 7648
rect 14589 7584 14597 7648
rect 14277 6560 14597 7584
rect 14277 6496 14285 6560
rect 14349 6496 14365 6560
rect 14429 6496 14445 6560
rect 14509 6496 14525 6560
rect 14589 6496 14597 6560
rect 14277 5472 14597 6496
rect 14277 5408 14285 5472
rect 14349 5408 14365 5472
rect 14429 5408 14445 5472
rect 14509 5408 14525 5472
rect 14589 5408 14597 5472
rect 14277 4384 14597 5408
rect 14277 4320 14285 4384
rect 14349 4320 14365 4384
rect 14429 4320 14445 4384
rect 14509 4320 14525 4384
rect 14589 4320 14597 4384
rect 14277 3296 14597 4320
rect 14277 3232 14285 3296
rect 14349 3232 14365 3296
rect 14429 3232 14445 3296
rect 14509 3232 14525 3296
rect 14589 3232 14597 3296
rect 14277 2208 14597 3232
rect 14277 2144 14285 2208
rect 14349 2144 14365 2208
rect 14429 2144 14445 2208
rect 14509 2144 14525 2208
rect 14589 2144 14597 2208
rect 14277 2128 14597 2144
use sky130_fd_sc_hd__decap_4  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_9 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1932 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_14 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2392 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11
timestamp 1604666999
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604666999
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604666999
transform 1 0 2024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1604666999
transform 1 0 2760 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604666999
transform 1 0 2576 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604666999
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1604666999
transform 1 0 3496 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23
timestamp 1604666999
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604666999
transform 1 0 2944 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604666999
transform 1 0 3680 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604666999
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604666999
transform 1 0 3128 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_30
timestamp 1604666999
transform 1 0 3864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1604666999
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4232 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4600 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 4232 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 4784 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604666999
transform 1 0 6256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1604666999
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53
timestamp 1604666999
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1604666999
transform 1 0 6348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1604666999
transform 1 0 5980 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1604666999
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67
timestamp 1604666999
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604666999
transform 1 0 7452 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7176 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_79
timestamp 1604666999
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_75
timestamp 1604666999
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_71
timestamp 1604666999
transform 1 0 7636 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 8096 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8740 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9108 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1604666999
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1604666999
transform 1 0 9292 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1604666999
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604666999
transform 1 0 10672 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_106
timestamp 1604666999
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604666999
transform 1 0 11040 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1604666999
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1604666999
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_114
timestamp 1604666999
transform 1 0 11592 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_117
timestamp 1604666999
transform 1 0 11868 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11684 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 11776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_121
timestamp 1604666999
transform 1 0 12236 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_1_136 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 13616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_132
timestamp 1604666999
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1604666999
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_134
timestamp 1604666999
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13432 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 14812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 14812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_142
timestamp 1604666999
transform 1 0 14168 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1604666999
transform 1 0 14352 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604666999
transform 1 0 2852 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604666999
transform 1 0 1748 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2392 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_11
timestamp 1604666999
transform 1 0 2116 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_16
timestamp 1604666999
transform 1 0 2576 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4692 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4508 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3404 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_23
timestamp 1604666999
transform 1 0 3220 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_36
timestamp 1604666999
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5704 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_48
timestamp 1604666999
transform 1 0 5520 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_52
timestamp 1604666999
transform 1 0 5888 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7636 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7176 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1604666999
transform 1 0 6624 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1604666999
transform 1 0 6992 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1604666999
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8648 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_88
timestamp 1604666999
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9016 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1604666999
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11132 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1604666999
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 13064 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_128
timestamp 1604666999
transform 1 0 12880 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_132 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 13248 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 14812 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1604666999
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604666999
transform 1 0 1472 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2576 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604666999
transform 1 0 2024 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2392 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_8
timestamp 1604666999
transform 1 0 1840 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_12
timestamp 1604666999
transform 1 0 2208 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1604666999
transform 1 0 4324 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 5060 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 6072 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_41
timestamp 1604666999
transform 1 0 4876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_52
timestamp 1604666999
transform 1 0 5888 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_56
timestamp 1604666999
transform 1 0 6256 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1604666999
transform 1 0 7636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_77
timestamp 1604666999
transform 1 0 8188 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10028 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8464 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 9844 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1604666999
transform 1 0 9292 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_93
timestamp 1604666999
transform 1 0 9660 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_106
timestamp 1604666999
transform 1 0 10856 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_114
timestamp 1604666999
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_118
timestamp 1604666999
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_132
timestamp 1604666999
transform 1 0 13248 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_136
timestamp 1604666999
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 14812 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_140 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 13984 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _30_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2208 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 1840 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1604666999
transform 1 0 1656 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1604666999
transform 1 0 2024 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 3404 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1604666999
transform 1 0 3220 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 6072 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 5888 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 5428 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_41
timestamp 1604666999
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1604666999
transform 1 0 5244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_49
timestamp 1604666999
transform 1 0 5612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1604666999
transform 1 0 6900 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1604666999
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1604666999
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1604666999
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1604666999
transform 1 0 9200 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_99
timestamp 1604666999
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10580 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 10396 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_112
timestamp 1604666999
transform 1 0 11408 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12144 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_133
timestamp 1604666999
transform 1 0 13340 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 14812 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_145
timestamp 1604666999
transform 1 0 14444 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604666999
transform 1 0 1748 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604666999
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604666999
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604666999
transform 1 0 2300 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1604666999
transform 1 0 2116 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 1604666999
transform 1 0 2484 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 2944 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1604666999
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604666999
transform 1 0 5612 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4876 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 5244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_43
timestamp 1604666999
transform 1 0 5060 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1604666999
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_53
timestamp 1604666999
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1604666999
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8096 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604666999
transform 1 0 7360 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_66
timestamp 1604666999
transform 1 0 7176 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_70
timestamp 1604666999
transform 1 0 7544 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10212 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_95
timestamp 1604666999
transform 1 0 9844 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10580 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1604666999
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_114
timestamp 1604666999
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1604666999
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_126
timestamp 1604666999
transform 1 0 12696 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_138
timestamp 1604666999
transform 1 0 13800 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 14812 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604666999
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604666999
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_13
timestamp 1604666999
transform 1 0 2300 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_7
timestamp 1604666999
transform 1 0 1748 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604666999
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1604666999
transform 1 0 2760 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_16
timestamp 1604666999
transform 1 0 2576 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2392 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604666999
transform 1 0 2852 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_29
timestamp 1604666999
transform 1 0 3772 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1604666999
transform 1 0 3496 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp 1604666999
transform 1 0 3128 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_27
timestamp 1604666999
transform 1 0 3588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 1604666999
transform 1 0 3220 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2944 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 3404 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_33
timestamp 1604666999
transform 1 0 4140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4232 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3956 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4324 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4416 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4508 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1604666999
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1604666999
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1604666999
transform 1 0 5244 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 5520 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_54
timestamp 1604666999
transform 1 0 6072 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_50
timestamp 1604666999
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5888 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 5980 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604666999
transform 1 0 6992 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604666999
transform 1 0 7176 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1604666999
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1604666999
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_72
timestamp 1604666999
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7728 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8280 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1604666999
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_84
timestamp 1604666999
transform 1 0 8832 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1604666999
transform 1 0 9292 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_91
timestamp 1604666999
transform 1 0 9476 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_97
timestamp 1604666999
transform 1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10212 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11776 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 12052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 11224 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_108
timestamp 1604666999
transform 1 0 11040 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_112
timestamp 1604666999
transform 1 0 11408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1604666999
transform 1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_108
timestamp 1604666999
transform 1 0 11040 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_116
timestamp 1604666999
transform 1 0 11776 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 12604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_135
timestamp 1604666999
transform 1 0 13524 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1604666999
transform 1 0 12236 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_127
timestamp 1604666999
transform 1 0 12788 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 14812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_143
timestamp 1604666999
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_139
timestamp 1604666999
transform 1 0 13892 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_145
timestamp 1604666999
transform 1 0 14444 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2392 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_6
timestamp 1604666999
transform 1 0 1656 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_17
timestamp 1604666999
transform 1 0 2668 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4508 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_21
timestamp 1604666999
transform 1 0 3036 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1604666999
transform 1 0 3772 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_36
timestamp 1604666999
transform 1 0 4416 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_39
timestamp 1604666999
transform 1 0 4692 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5428 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_45
timestamp 1604666999
transform 1 0 5244 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7912 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_66
timestamp 1604666999
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_70
timestamp 1604666999
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8924 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_83
timestamp 1604666999
transform 1 0 8740 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1604666999
transform 1 0 9108 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1604666999
transform 1 0 9476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_97
timestamp 1604666999
transform 1 0 10028 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 12052 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 10304 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_102
timestamp 1604666999
transform 1 0 10488 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp 1604666999
transform 1 0 10856 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_110
timestamp 1604666999
transform 1 0 11224 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_118
timestamp 1604666999
transform 1 0 11960 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_138
timestamp 1604666999
transform 1 0 13800 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 14812 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1748 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 1564 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_26
timestamp 1604666999
transform 1 0 3496 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_32
timestamp 1604666999
transform 1 0 4048 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_35
timestamp 1604666999
transform 1 0 4324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1604666999
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5060 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_52
timestamp 1604666999
transform 1 0 5888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604666999
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 6992 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1604666999
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_77
timestamp 1604666999
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8556 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10120 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_90
timestamp 1604666999
transform 1 0 9384 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_94
timestamp 1604666999
transform 1 0 9752 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10304 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11316 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11684 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_109
timestamp 1604666999
transform 1 0 11132 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 1604666999
transform 1 0 11500 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_117
timestamp 1604666999
transform 1 0 11868 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1604666999
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 14812 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_143
timestamp 1604666999
transform 1 0 14260 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_9
timestamp 1604666999
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4508 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 3312 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp 1604666999
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1604666999
transform 1 0 3496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1604666999
transform 1 0 3864 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp 1604666999
transform 1 0 4416 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6440 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1604666999
transform 1 0 6256 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6992 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1604666999
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_83
timestamp 1604666999
transform 1 0 8740 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1604666999
transform 1 0 9108 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1604666999
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_96
timestamp 1604666999
transform 1 0 9936 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10672 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10488 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_100
timestamp 1604666999
transform 1 0 10304 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_113
timestamp 1604666999
transform 1 0 11500 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 12788 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1604666999
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_125
timestamp 1604666999
transform 1 0 12604 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 14812 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_145
timestamp 1604666999
transform 1 0 14444 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_15
timestamp 1604666999
transform 1 0 2484 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 3312 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4692 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_21
timestamp 1604666999
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_33
timestamp 1604666999
transform 1 0 4140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_37
timestamp 1604666999
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_41
timestamp 1604666999
transform 1 0 4876 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7268 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1604666999
transform 1 0 8096 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8832 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1604666999
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11316 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1604666999
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1604666999
transform 1 0 10948 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1604666999
transform 1 0 11500 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_117
timestamp 1604666999
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_132
timestamp 1604666999
transform 1 0 13248 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 14812 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_144
timestamp 1604666999
transform 1 0 14352 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 2392 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_7
timestamp 1604666999
transform 1 0 1748 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_13
timestamp 1604666999
transform 1 0 2300 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_16
timestamp 1604666999
transform 1 0 2576 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_21
timestamp 1604666999
transform 1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_26
timestamp 1604666999
transform 1 0 3496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1604666999
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_51
timestamp 1604666999
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 7268 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_63
timestamp 1604666999
transform 1 0 6900 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1604666999
transform 1 0 7452 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9016 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1604666999
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1604666999
transform 1 0 9200 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11684 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 11500 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_102
timestamp 1604666999
transform 1 0 10488 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_107
timestamp 1604666999
transform 1 0 10948 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_111
timestamp 1604666999
transform 1 0 11316 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_134
timestamp 1604666999
transform 1 0 13432 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 14812 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_6
timestamp 1604666999
transform 1 0 1656 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1604666999
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_15
timestamp 1604666999
transform 1 0 2484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_11
timestamp 1604666999
transform 1 0 2116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2208 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2300 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 1604666999
transform 1 0 3680 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3404 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_38
timestamp 1604666999
transform 1 0 4600 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_32
timestamp 1604666999
transform 1 0 4048 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 4416 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4416 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_46
timestamp 1604666999
transform 1 0 5336 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1604666999
transform 1 0 4968 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 5520 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 5152 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 4784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1604666999
transform 1 0 6440 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1604666999
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1604666999
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604666999
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 5888 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_45
timestamp 1604666999
transform 1 0 5244 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 6992 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7360 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1604666999
transform 1 0 7176 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_70
timestamp 1604666999
transform 1 0 7544 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_72
timestamp 1604666999
transform 1 0 7728 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_84
timestamp 1604666999
transform 1 0 8832 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_84
timestamp 1604666999
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9200 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1604666999
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1604666999
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_97
timestamp 1604666999
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10488 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 10764 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10488 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_101
timestamp 1604666999
transform 1 0 10396 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_104
timestamp 1604666999
transform 1 0 10672 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1604666999
transform 1 0 11960 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_125
timestamp 1604666999
transform 1 0 12604 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1604666999
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 12788 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_14_138
timestamp 1604666999
transform 1 0 13800 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1604666999
transform 1 0 13616 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_132
timestamp 1604666999
transform 1 0 13248 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12972 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 14812 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_140
timestamp 1604666999
transform 1 0 13984 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 2760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 2024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 1656 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_8
timestamp 1604666999
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_12
timestamp 1604666999
transform 1 0 2208 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_16
timestamp 1604666999
transform 1 0 2576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4508 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 2944 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 3956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_29
timestamp 1604666999
transform 1 0 3772 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1604666999
transform 1 0 4140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 5796 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_46
timestamp 1604666999
transform 1 0 5336 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_50
timestamp 1604666999
transform 1 0 5704 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604666999
transform 1 0 8372 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7820 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1604666999
transform 1 0 7636 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_75
timestamp 1604666999
transform 1 0 8004 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_82
timestamp 1604666999
transform 1 0 8648 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_94
timestamp 1604666999
transform 1 0 9752 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_106
timestamp 1604666999
transform 1 0 10856 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_126
timestamp 1604666999
transform 1 0 12696 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_138
timestamp 1604666999
transform 1 0 13800 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 14812 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_11
timestamp 1604666999
transform 1 0 2116 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604666999
transform 1 0 4140 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1604666999
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 5152 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4968 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_40
timestamp 1604666999
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_53
timestamp 1604666999
transform 1 0 5980 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6716 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1604666999
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1604666999
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1604666999
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1604666999
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 14812 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1604666999
transform 1 0 14076 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_145
timestamp 1604666999
transform 1 0 14444 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2484 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2300 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1604666999
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 1604666999
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1604666999
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1604666999
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_55
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7360 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_87
timestamp 1604666999
transform 1 0 9108 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1604666999
transform 1 0 10212 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10672 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_102
timestamp 1604666999
transform 1 0 10488 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_106
timestamp 1604666999
transform 1 0 10856 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1604666999
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 14812 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_143
timestamp 1604666999
transform 1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2484 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_17
timestamp 1604666999
transform 1 0 2668 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 5980 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 6348 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_51
timestamp 1604666999
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1604666999
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 8004 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_72
timestamp 1604666999
transform 1 0 7728 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1604666999
transform 1 0 8188 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10028 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1604666999
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1604666999
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_99
timestamp 1604666999
transform 1 0 10212 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10304 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_119
timestamp 1604666999
transform 1 0 12052 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_131
timestamp 1604666999
transform 1 0 13156 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 14812 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_143
timestamp 1604666999
transform 1 0 14260 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_6
timestamp 1604666999
transform 1 0 1656 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_7
timestamp 1604666999
transform 1 0 1748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_14
timestamp 1604666999
transform 1 0 2392 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_13
timestamp 1604666999
transform 1 0 2300 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2392 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_18
timestamp 1604666999
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2576 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_35
timestamp 1604666999
transform 1 0 4324 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1604666999
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5888 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5520 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_47
timestamp 1604666999
transform 1 0 5428 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_50
timestamp 1604666999
transform 1 0 5704 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_54
timestamp 1604666999
transform 1 0 6072 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_58
timestamp 1604666999
transform 1 0 6440 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_44
timestamp 1604666999
transform 1 0 5152 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1604666999
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_61
timestamp 1604666999
transform 1 0 6716 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7360 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_70
timestamp 1604666999
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1604666999
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 7820 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8372 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_88
timestamp 1604666999
transform 1 0 9200 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604666999
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_81
timestamp 1604666999
transform 1 0 8556 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 8740 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9844 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10028 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8924 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1604666999
transform 1 0 10856 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_108
timestamp 1604666999
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1604666999
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 11040 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_110
timestamp 1604666999
transform 1 0 11224 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1604666999
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 11592 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_127
timestamp 1604666999
transform 1 0 12788 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1604666999
transform 1 0 12420 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_127
timestamp 1604666999
transform 1 0 12788 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 14812 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 14812 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_139
timestamp 1604666999
transform 1 0 13892 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1604666999
transform 1 0 14444 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_139
timestamp 1604666999
transform 1 0 13892 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1604666999
transform 1 0 14444 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1604666999
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1604666999
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 5060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_41
timestamp 1604666999
transform 1 0 4876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_45
timestamp 1604666999
transform 1 0 5244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_49
timestamp 1604666999
transform 1 0 5612 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1604666999
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10212 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9844 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9476 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_88
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_93
timestamp 1604666999
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_97
timestamp 1604666999
transform 1 0 10028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10396 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1604666999
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13432 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1604666999
transform 1 0 13248 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_136
timestamp 1604666999
transform 1 0 13616 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 14812 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1604666999
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1604666999
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 4692 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 4232 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_32
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_36
timestamp 1604666999
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_48
timestamp 1604666999
transform 1 0 5520 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_56
timestamp 1604666999
transform 1 0 6256 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6992 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 8004 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6808 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8372 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 1604666999
transform 1 0 6624 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1604666999
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_77
timestamp 1604666999
transform 1 0 8188 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10212 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10028 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8740 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_81
timestamp 1604666999
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_85
timestamp 1604666999
transform 1 0 8924 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_89
timestamp 1604666999
transform 1 0 9292 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11776 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11408 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_108
timestamp 1604666999
transform 1 0 11040 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1604666999
transform 1 0 11592 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_135
timestamp 1604666999
transform 1 0 13524 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 14812 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_143
timestamp 1604666999
transform 1 0 14260 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_6
timestamp 1604666999
transform 1 0 1656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_10
timestamp 1604666999
transform 1 0 2024 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 4048 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3864 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_22
timestamp 1604666999
transform 1 0 3128 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_28
timestamp 1604666999
transform 1 0 3680 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 5060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_41
timestamp 1604666999
transform 1 0 4876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_45
timestamp 1604666999
transform 1 0 5244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_49
timestamp 1604666999
transform 1 0 5612 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7820 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6992 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1604666999
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_70
timestamp 1604666999
transform 1 0 7544 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 9844 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_92
timestamp 1604666999
transform 1 0 9568 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1604666999
transform 1 0 10028 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604666999
transform 1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 11132 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1604666999
transform 1 0 10396 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_107
timestamp 1604666999
transform 1 0 10948 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_114
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1604666999
transform 1 0 11960 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_132
timestamp 1604666999
transform 1 0 13248 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 14812 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_144
timestamp 1604666999
transform 1 0 14352 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2392 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_7
timestamp 1604666999
transform 1 0 1748 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_13
timestamp 1604666999
transform 1 0 2300 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_16
timestamp 1604666999
transform 1 0 2576 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4232 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_21
timestamp 1604666999
transform 1 0 3036 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4876 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_24_40
timestamp 1604666999
transform 1 0 4784 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7360 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_60
timestamp 1604666999
transform 1 0 6624 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_64
timestamp 1604666999
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_77
timestamp 1604666999
transform 1 0 8188 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9844 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9292 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1604666999
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1604666999
transform 1 0 11408 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 10856 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1604666999
transform 1 0 10672 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_108
timestamp 1604666999
transform 1 0 11040 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12420 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1604666999
transform 1 0 12236 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_125
timestamp 1604666999
transform 1 0 12604 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_137
timestamp 1604666999
transform 1 0 13708 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 14812 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1604666999
transform 1 0 14444 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 2852 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 2668 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2300 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 1932 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_6
timestamp 1604666999
transform 1 0 1656 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1604666999
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_15
timestamp 1604666999
transform 1 0 2484 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1604666999
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_42
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_50
timestamp 1604666999
transform 1 0 5704 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_53
timestamp 1604666999
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1604666999
transform 1 0 6348 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 7820 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1604666999
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_75
timestamp 1604666999
transform 1 0 8004 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9292 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11224 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1604666999
transform 1 0 11040 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_112
timestamp 1604666999
transform 1 0 11408 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_120
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp 1604666999
transform 1 0 13524 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 14812 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_143
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_16
timestamp 1604666999
transform 1 0 2576 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_11
timestamp 1604666999
transform 1 0 2116 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1604666999
transform 1 0 2116 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2760 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_29
timestamp 1604666999
transform 1 0 3772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2944 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1604666999
transform 1 0 4508 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1604666999
transform 1 0 4140 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 3956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4324 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4692 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_26_49
timestamp 1604666999
transform 1 0 5612 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_45
timestamp 1604666999
transform 1 0 5244 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_41
timestamp 1604666999
transform 1 0 4876 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 5060 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4876 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_27_58
timestamp 1604666999
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_54
timestamp 1604666999
transform 1 0 6072 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1604666999
transform 1 0 5704 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_55
timestamp 1604666999
transform 1 0 6164 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 5888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6256 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 8372 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1604666999
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1604666999
transform 1 0 7636 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_75
timestamp 1604666999
transform 1 0 8004 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_89
timestamp 1604666999
transform 1 0 9292 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_83
timestamp 1604666999
transform 1 0 8740 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8556 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8556 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9568 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_90
timestamp 1604666999
transform 1 0 9384 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_94
timestamp 1604666999
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9844 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1604666999
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10120 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 10212 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_118
timestamp 1604666999
transform 1 0 11960 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_107
timestamp 1604666999
transform 1 0 10948 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_111
timestamp 1604666999
transform 1 0 11316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1604666999
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_130
timestamp 1604666999
transform 1 0 13064 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_135
timestamp 1604666999
transform 1 0 13524 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 14812 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_142
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_143
timestamp 1604666999
transform 1 0 14260 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp 1604666999
transform 1 0 2852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 2944 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_22
timestamp 1604666999
transform 1 0 3128 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604666999
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4876 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_28_40
timestamp 1604666999
transform 1 0 4784 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_50
timestamp 1604666999
transform 1 0 5704 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7728 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6808 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 7176 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 7544 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_64
timestamp 1604666999
transform 1 0 6992 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1604666999
transform 1 0 7360 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8740 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_81
timestamp 1604666999
transform 1 0 8556 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_85
timestamp 1604666999
transform 1 0 8924 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1604666999
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11592 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1604666999
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_106
timestamp 1604666999
transform 1 0 10856 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_133
timestamp 1604666999
transform 1 0 13340 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 14812 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_145
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_6
timestamp 1604666999
transform 1 0 1656 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_10
timestamp 1604666999
transform 1 0 2024 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3864 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_22
timestamp 1604666999
transform 1 0 3128 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_32
timestamp 1604666999
transform 1 0 4048 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1604666999
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4784 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1604666999
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_53
timestamp 1604666999
transform 1 0 5980 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1604666999
transform 1 0 6348 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8004 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1604666999
transform 1 0 7268 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604666999
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1604666999
transform 1 0 9752 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_106
timestamp 1604666999
transform 1 0 10856 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_135
timestamp 1604666999
transform 1 0 13524 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 14812 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_143
timestamp 1604666999
transform 1 0 14260 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2852 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_15
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 4508 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_21
timestamp 1604666999
transform 1 0 3036 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1604666999
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_36
timestamp 1604666999
transform 1 0 4416 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_39
timestamp 1604666999
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4876 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7176 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7544 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_60
timestamp 1604666999
transform 1 0 6624 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_68
timestamp 1604666999
transform 1 0 7360 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_72
timestamp 1604666999
transform 1 0 7728 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_84
timestamp 1604666999
transform 1 0 8832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_89
timestamp 1604666999
transform 1 0 9292 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_93
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_98
timestamp 1604666999
transform 1 0 10120 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10304 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_102
timestamp 1604666999
transform 1 0 10488 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_114
timestamp 1604666999
transform 1 0 11592 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_126
timestamp 1604666999
transform 1 0 12696 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_138
timestamp 1604666999
transform 1 0 13800 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 14812 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2852 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2668 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_15
timestamp 1604666999
transform 1 0 2484 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604666999
transform 1 0 5336 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_42
timestamp 1604666999
transform 1 0 4968 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_49
timestamp 1604666999
transform 1 0 5612 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7176 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6992 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8188 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_75
timestamp 1604666999
transform 1 0 8004 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_79
timestamp 1604666999
transform 1 0 8372 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9108 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8924 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11500 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11040 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 11868 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1604666999
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_110
timestamp 1604666999
transform 1 0 11224 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1604666999
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1604666999
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1604666999
transform 1 0 13524 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 14812 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1604666999
transform 1 0 14260 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4508 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 3680 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1604666999
transform 1 0 3864 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_36
timestamp 1604666999
transform 1 0 4416 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 6348 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_32_46
timestamp 1604666999
transform 1 0 5336 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_54
timestamp 1604666999
transform 1 0 6072 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_32_76
timestamp 1604666999
transform 1 0 8096 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9936 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1604666999
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_88
timestamp 1604666999
transform 1 0 9200 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11500 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 11040 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_105
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_110
timestamp 1604666999
transform 1 0 11224 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_132
timestamp 1604666999
transform 1 0 13248 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 14812 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1604666999
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_15
timestamp 1604666999
transform 1 0 2484 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1604666999
transform 1 0 3312 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_21
timestamp 1604666999
transform 1 0 3036 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_23
timestamp 1604666999
transform 1 0 3220 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3680 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 3128 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 3680 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_38
timestamp 1604666999
transform 1 0 4600 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_30
timestamp 1604666999
transform 1 0 3864 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4692 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_37
timestamp 1604666999
transform 1 0 4508 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_41
timestamp 1604666999
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_49
timestamp 1604666999
transform 1 0 5612 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5060 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_57
timestamp 1604666999
transform 1 0 6348 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1604666999
transform 1 0 6348 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_53
timestamp 1604666999
transform 1 0 5980 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1604666999
transform 1 0 5704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_45
timestamp 1604666999
transform 1 0 5244 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_64
timestamp 1604666999
transform 1 0 6992 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_60
timestamp 1604666999
transform 1 0 6624 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 6808 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 7084 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_34_79
timestamp 1604666999
transform 1 0 8372 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_34_74
timestamp 1604666999
transform 1 0 7912 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_79
timestamp 1604666999
transform 1 0 8372 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1604666999
transform 1 0 8004 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_71
timestamp 1604666999
transform 1 0 7636 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8188 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 7820 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_88
timestamp 1604666999
transform 1 0 9200 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_85
timestamp 1604666999
transform 1 0 8924 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1604666999
transform 1 0 8740 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9016 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_34_99
timestamp 1604666999
transform 1 0 10212 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1604666999
transform 1 0 10212 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_95
timestamp 1604666999
transform 1 0 9844 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10028 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 10580 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 10396 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 11040 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 10580 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_116
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1604666999
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 11960 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 12052 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_135
timestamp 1604666999
transform 1 0 13524 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_121
timestamp 1604666999
transform 1 0 12236 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_125
timestamp 1604666999
transform 1 0 12604 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_137
timestamp 1604666999
transform 1 0 13708 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 14812 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 14812 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_143
timestamp 1604666999
transform 1 0 14260 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_145
timestamp 1604666999
transform 1 0 14444 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_6
timestamp 1604666999
transform 1 0 1656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_10
timestamp 1604666999
transform 1 0 2024 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1604666999
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4692 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1604666999
transform 1 0 3128 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 2944 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_31
timestamp 1604666999
transform 1 0 3956 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 5704 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_48
timestamp 1604666999
transform 1 0 5520 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_52
timestamp 1604666999
transform 1 0 5888 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_58
timestamp 1604666999
transform 1 0 6440 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8188 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7268 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_62
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_66
timestamp 1604666999
transform 1 0 7176 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_69
timestamp 1604666999
transform 1 0 7452 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_73
timestamp 1604666999
transform 1 0 7820 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 10028 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 9660 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 9292 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_86
timestamp 1604666999
transform 1 0 9016 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_91
timestamp 1604666999
transform 1 0 9476 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_95
timestamp 1604666999
transform 1 0 9844 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_112
timestamp 1604666999
transform 1 0 11408 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_132
timestamp 1604666999
transform 1 0 13248 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 14812 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_144
timestamp 1604666999
transform 1 0 14352 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1604666999
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 2668 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1604666999
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_7
timestamp 1604666999
transform 1 0 1748 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_36_15
timestamp 1604666999
transform 1 0 2484 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_19
timestamp 1604666999
transform 1 0 2852 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4692 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3128 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 4324 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_24
timestamp 1604666999
transform 1 0 3312 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_30
timestamp 1604666999
transform 1 0 3864 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_36_32
timestamp 1604666999
transform 1 0 4048 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_37
timestamp 1604666999
transform 1 0 4508 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4968 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_36_41
timestamp 1604666999
transform 1 0 4876 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7544 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6992 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 7360 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_61
timestamp 1604666999
transform 1 0 6716 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_66
timestamp 1604666999
transform 1 0 7176 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_79
timestamp 1604666999
transform 1 0 8372 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9384 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_85
timestamp 1604666999
transform 1 0 8924 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_88
timestamp 1604666999
transform 1 0 9200 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 11224 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 10672 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 11040 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_102
timestamp 1604666999
transform 1 0 10488 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_106
timestamp 1604666999
transform 1 0 10856 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_119
timestamp 1604666999
transform 1 0 12052 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604666999
transform 1 0 12788 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12420 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_125
timestamp 1604666999
transform 1 0 12604 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_130
timestamp 1604666999
transform 1 0 13064 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1604666999
transform -1 0 14812 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_142
timestamp 1604666999
transform 1 0 14168 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2668 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1604666999
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2484 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2116 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 1748 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1604666999
transform 1 0 1380 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_9
timestamp 1604666999
transform 1 0 1932 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_13
timestamp 1604666999
transform 1 0 2300 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4600 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1604666999
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 4968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6164 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_40
timestamp 1604666999
transform 1 0 4784 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1604666999
transform 1 0 5980 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1604666999
transform 1 0 6348 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 6808 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9476 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9292 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 8924 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_81
timestamp 1604666999
transform 1 0 8556 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_87
timestamp 1604666999
transform 1 0 9108 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11408 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_110
timestamp 1604666999
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_114
timestamp 1604666999
transform 1 0 11592 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1604666999
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12420 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13432 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 13800 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_132
timestamp 1604666999
transform 1 0 13248 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_136
timestamp 1604666999
transform 1 0 13616 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1604666999
transform -1 0 14812 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_37_140
timestamp 1604666999
transform 1 0 13984 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1604666999
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 2208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 1840 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_6
timestamp 1604666999
transform 1 0 1656 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_10
timestamp 1604666999
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4508 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4324 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3772 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_23
timestamp 1604666999
transform 1 0 3220 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_32
timestamp 1604666999
transform 1 0 4048 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6440 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_56
timestamp 1604666999
transform 1 0 6256 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6992 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8004 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 6808 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8372 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_60
timestamp 1604666999
transform 1 0 6624 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_73
timestamp 1604666999
transform 1 0 7820 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_77
timestamp 1604666999
transform 1 0 8188 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_81
timestamp 1604666999
transform 1 0 8556 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_89
timestamp 1604666999
transform 1 0 9292 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_112
timestamp 1604666999
transform 1 0 11408 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12144 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13156 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_129
timestamp 1604666999
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_133
timestamp 1604666999
transform 1 0 13340 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1604666999
transform -1 0 14812 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_145
timestamp 1604666999
transform 1 0 14444 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_7
timestamp 1604666999
transform 1 0 1748 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_3
timestamp 1604666999
transform 1 0 1380 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1604666999
transform 1 0 1748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1604666999
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 1932 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1604666999
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1604666999
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_11
timestamp 1604666999
transform 1 0 2116 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_14
timestamp 1604666999
transform 1 0 2392 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_10
timestamp 1604666999
transform 1 0 2024 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2208 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2576 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2300 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2760 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_40_26
timestamp 1604666999
transform 1 0 3496 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_22
timestamp 1604666999
transform 1 0 3128 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_27
timestamp 1604666999
transform 1 0 3588 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3312 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 3772 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_30
timestamp 1604666999
transform 1 0 3864 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_31
timestamp 1604666999
transform 1 0 3956 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4140 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4048 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4324 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_40_41
timestamp 1604666999
transform 1 0 4876 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_48
timestamp 1604666999
transform 1 0 5520 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_44
timestamp 1604666999
transform 1 0 5152 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 5152 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 5336 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_58
timestamp 1604666999
transform 1 0 6440 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_58
timestamp 1604666999
transform 1 0 6440 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_52
timestamp 1604666999
transform 1 0 5888 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 5704 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6532 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_46
timestamp 1604666999
transform 1 0 5336 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 7728 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7176 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6992 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1604666999
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_68
timestamp 1604666999
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_75
timestamp 1604666999
transform 1 0 8004 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9660 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10028 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_91
timestamp 1604666999
transform 1 0 9476 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_95
timestamp 1604666999
transform 1 0 9844 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_99
timestamp 1604666999
transform 1 0 10212 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_87
timestamp 1604666999
transform 1 0 9108 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_91
timestamp 1604666999
transform 1 0 9476 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1604666999
transform 1 0 10856 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_102
timestamp 1604666999
transform 1 0 10488 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_109
timestamp 1604666999
transform 1 0 11132 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_103
timestamp 1604666999
transform 1 0 10580 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10396 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 10672 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_116
timestamp 1604666999
transform 1 0 11776 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_112
timestamp 1604666999
transform 1 0 11408 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11592 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11224 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11224 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1604666999
transform 1 0 12420 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_135
timestamp 1604666999
transform 1 0 13524 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_129
timestamp 1604666999
transform 1 0 12972 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1604666999
transform -1 0 14812 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1604666999
transform -1 0 14812 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_143
timestamp 1604666999
transform 1 0 14260 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_141
timestamp 1604666999
transform 1 0 14076 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_145
timestamp 1604666999
transform 1 0 14444 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1932 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1604666999
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1748 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_3
timestamp 1604666999
transform 1 0 1380 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4416 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3864 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_28
timestamp 1604666999
transform 1 0 3680 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_32
timestamp 1604666999
transform 1 0 4048 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_45
timestamp 1604666999
transform 1 0 5244 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_49
timestamp 1604666999
transform 1 0 5612 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 7912 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 7728 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_62
timestamp 1604666999
transform 1 0 6808 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_70
timestamp 1604666999
transform 1 0 7544 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1604666999
transform 1 0 10028 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 9660 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9292 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_83
timestamp 1604666999
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_87
timestamp 1604666999
transform 1 0 9108 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_91
timestamp 1604666999
transform 1 0 9476 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_95
timestamp 1604666999
transform 1 0 9844 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_106
timestamp 1604666999
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1604666999
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_114
timestamp 1604666999
transform 1 0 11592 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1604666999
transform 1 0 12420 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_135
timestamp 1604666999
transform 1 0 13524 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1604666999
transform -1 0 14812 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_143
timestamp 1604666999
transform 1 0 14260 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1604666999
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_6
timestamp 1604666999
transform 1 0 1656 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_18
timestamp 1604666999
transform 1 0 2760 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604666999
transform 1 0 4508 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1604666999
transform 1 0 3864 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_32
timestamp 1604666999
transform 1 0 4048 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_36
timestamp 1604666999
transform 1 0 4416 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_40
timestamp 1604666999
transform 1 0 4784 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_52
timestamp 1604666999
transform 1 0 5888 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 7912 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_60
timestamp 1604666999
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_64
timestamp 1604666999
transform 1 0 6992 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_72
timestamp 1604666999
transform 1 0 7728 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_76
timestamp 1604666999
transform 1 0 8096 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_88
timestamp 1604666999
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 10672 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_102
timestamp 1604666999
transform 1 0 10488 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_106
timestamp 1604666999
transform 1 0 10856 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_118
timestamp 1604666999
transform 1 0 11960 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_130
timestamp 1604666999
transform 1 0 13064 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1604666999
transform -1 0 14812 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_142
timestamp 1604666999
transform 1 0 14168 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1604666999
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1604666999
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1604666999
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1604666999
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_39
timestamp 1604666999
transform 1 0 4692 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 6532 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 5152 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5520 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_43
timestamp 1604666999
transform 1 0 5060 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_46
timestamp 1604666999
transform 1 0 5336 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_50
timestamp 1604666999
transform 1 0 5704 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_54
timestamp 1604666999
transform 1 0 6072 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_57
timestamp 1604666999
transform 1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp 1604666999
transform 1 0 7636 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_75
timestamp 1604666999
transform 1 0 8004 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_79
timestamp 1604666999
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9476 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 9292 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8924 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_83
timestamp 1604666999
transform 1 0 8740 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_87
timestamp 1604666999
transform 1 0 9108 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604666999
transform 1 0 11040 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10488 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11868 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10856 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_100
timestamp 1604666999
transform 1 0 10304 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_104
timestamp 1604666999
transform 1 0 10672 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_111
timestamp 1604666999
transform 1 0 11316 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_43_119
timestamp 1604666999
transform 1 0 12052 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 12604 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_123
timestamp 1604666999
transform 1 0 12420 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_127
timestamp 1604666999
transform 1 0 12788 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1604666999
transform -1 0 14812 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_43_139
timestamp 1604666999
transform 1 0 13892 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_145
timestamp 1604666999
transform 1 0 14444 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1604666999
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 2576 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1604666999
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_15
timestamp 1604666999
transform 1 0 2484 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_18
timestamp 1604666999
transform 1 0 2760 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2944 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_22
timestamp 1604666999
transform 1 0 3128 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_30
timestamp 1604666999
transform 1 0 3864 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1604666999
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5152 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 7728 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 7084 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_63
timestamp 1604666999
transform 1 0 6900 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_67
timestamp 1604666999
transform 1 0 7268 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 1604666999
transform 1 0 7636 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 8740 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 9108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_81
timestamp 1604666999
transform 1 0 8556 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1604666999
transform 1 0 8924 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_89
timestamp 1604666999
transform 1 0 9292 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_44_93
timestamp 1604666999
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_98
timestamp 1604666999
transform 1 0 10120 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11868 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1604666999
transform 1 0 10304 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_44_109
timestamp 1604666999
transform 1 0 11132 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_136
timestamp 1604666999
transform 1 0 13616 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1604666999
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_144
timestamp 1604666999
transform 1 0 14352 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 2576 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1604666999
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 2392 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 2024 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 1656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_3
timestamp 1604666999
transform 1 0 1380 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_8
timestamp 1604666999
transform 1 0 1840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_12
timestamp 1604666999
transform 1 0 2208 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_35
timestamp 1604666999
transform 1 0 4324 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 5244 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 6532 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 5612 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 6164 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_43
timestamp 1604666999
transform 1 0 5060 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_47
timestamp 1604666999
transform 1 0 5428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1604666999
transform 1 0 5796 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1604666999
transform 1 0 6348 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1604666999
transform 1 0 8372 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 8004 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_71
timestamp 1604666999
transform 1 0 7636 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_77
timestamp 1604666999
transform 1 0 8188 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1604666999
transform 1 0 9936 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 9384 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_88
timestamp 1604666999
transform 1 0 9200 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_92
timestamp 1604666999
transform 1 0 9568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 10948 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11316 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_105
timestamp 1604666999
transform 1 0 10764 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_109
timestamp 1604666999
transform 1 0 11132 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_113
timestamp 1604666999
transform 1 0 11500 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_118
timestamp 1604666999
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_132
timestamp 1604666999
transform 1 0 13248 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1604666999
transform -1 0 14812 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_144
timestamp 1604666999
transform 1 0 14352 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1604666999
transform 1 0 1380 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp 1604666999
transform 1 0 1380 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1604666999
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1604666999
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_16
timestamp 1604666999
transform 1 0 2576 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_11
timestamp 1604666999
transform 1 0 2116 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_11
timestamp 1604666999
transform 1 0 2116 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 2760 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 2392 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_24
timestamp 1604666999
transform 1 0 3312 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_20
timestamp 1604666999
transform 1 0 2944 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1604666999
transform 1 0 3588 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_23
timestamp 1604666999
transform 1 0 3220 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3128 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3680 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 3496 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_32
timestamp 1604666999
transform 1 0 4048 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_30
timestamp 1604666999
transform 1 0 3864 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 3680 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_47_47
timestamp 1604666999
transform 1 0 5428 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_43
timestamp 1604666999
transform 1 0 5060 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_40
timestamp 1604666999
transform 1 0 4784 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 4876 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 5612 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_55
timestamp 1604666999
transform 1 0 6164 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_51
timestamp 1604666999
transform 1 0 5796 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 5980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 5244 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_47_69
timestamp 1604666999
transform 1 0 7452 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_65
timestamp 1604666999
transform 1 0 7084 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_64
timestamp 1604666999
transform 1 0 6992 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 7268 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604666999
transform 1 0 6808 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_47_73
timestamp 1604666999
transform 1 0 7820 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_72
timestamp 1604666999
transform 1 0 7728 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7820 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 8004 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 8096 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9936 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_84
timestamp 1604666999
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_88
timestamp 1604666999
transform 1 0 9200 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_93
timestamp 1604666999
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_98
timestamp 1604666999
transform 1 0 10120 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_95
timestamp 1604666999
transform 1 0 9844 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_46_105
timestamp 1604666999
transform 1 0 10764 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_102
timestamp 1604666999
transform 1 0 10488 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10580 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10396 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10580 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_116
timestamp 1604666999
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_112
timestamp 1604666999
transform 1 0 11408 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 10948 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 12880 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_126
timestamp 1604666999
transform 1 0 12696 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_130
timestamp 1604666999
transform 1 0 13064 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1604666999
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1604666999
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_135
timestamp 1604666999
transform 1 0 13524 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1604666999
transform -1 0 14812 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1604666999
transform -1 0 14812 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_142
timestamp 1604666999
transform 1 0 14168 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_143
timestamp 1604666999
transform 1 0 14260 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1604666999
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_3
timestamp 1604666999
transform 1 0 1380 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_11
timestamp 1604666999
transform 1 0 2116 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4600 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_23
timestamp 1604666999
transform 1 0 3220 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_48_32
timestamp 1604666999
transform 1 0 4048 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 6532 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1604666999
transform 1 0 4876 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_48_40
timestamp 1604666999
transform 1 0 4784 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_50
timestamp 1604666999
transform 1 0 5704 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_58
timestamp 1604666999
transform 1 0 6440 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_78
timestamp 1604666999
transform 1 0 8280 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8464 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9844 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10212 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_82
timestamp 1604666999
transform 1 0 8648 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_86
timestamp 1604666999
transform 1 0 9016 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1604666999
transform 1 0 9660 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_97
timestamp 1604666999
transform 1 0 10028 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11132 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 10580 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1604666999
transform 1 0 10396 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_105
timestamp 1604666999
transform 1 0 10764 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_128
timestamp 1604666999
transform 1 0 12880 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1604666999
transform -1 0 14812 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_140
timestamp 1604666999
transform 1 0 13984 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1604666999
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2208 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_6
timestamp 1604666999
transform 1 0 1656 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_10
timestamp 1604666999
transform 1 0 2024 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_14
timestamp 1604666999
transform 1 0 2392 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4600 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4416 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 4048 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_26
timestamp 1604666999
transform 1 0 3496 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_34
timestamp 1604666999
transform 1 0 4232 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5612 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 5980 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6348 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_47
timestamp 1604666999
transform 1 0 5428 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_51
timestamp 1604666999
transform 1 0 5796 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_55
timestamp 1604666999
transform 1 0 6164 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_59
timestamp 1604666999
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_1_
timestamp 1604666999
transform 1 0 8004 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7636 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7268 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_62
timestamp 1604666999
transform 1 0 6808 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1604666999
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_69
timestamp 1604666999
transform 1 0 7452 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_73
timestamp 1604666999
transform 1 0 7820 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9568 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 9384 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 9016 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_84
timestamp 1604666999
transform 1 0 8832 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_88
timestamp 1604666999
transform 1 0 9200 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 10580 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10948 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_101
timestamp 1604666999
transform 1 0 10396 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_105
timestamp 1604666999
transform 1 0 10764 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_109
timestamp 1604666999
transform 1 0 11132 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1604666999
transform 1 0 12236 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1604666999
transform 1 0 12420 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_135
timestamp 1604666999
transform 1 0 13524 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1604666999
transform -1 0 14812 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_49_143
timestamp 1604666999
transform 1 0 14260 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1604666999
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_6
timestamp 1604666999
transform 1 0 1656 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_18
timestamp 1604666999
transform 1 0 2760 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 4600 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4232 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1604666999
transform 1 0 3864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_32
timestamp 1604666999
transform 1 0 4048 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_36
timestamp 1604666999
transform 1 0 4416 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5244 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6440 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_40
timestamp 1604666999
transform 1 0 4784 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_44
timestamp 1604666999
transform 1 0 5152 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_54
timestamp 1604666999
transform 1 0 6072 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7636 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6808 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7452 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_60
timestamp 1604666999
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_64
timestamp 1604666999
transform 1 0 6992 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_68
timestamp 1604666999
transform 1 0 7360 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9844 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 8648 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_80
timestamp 1604666999
transform 1 0 8464 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_84
timestamp 1604666999
transform 1 0 8832 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1604666999
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_97
timestamp 1604666999
transform 1 0 10028 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10304 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_119
timestamp 1604666999
transform 1 0 12052 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_131
timestamp 1604666999
transform 1 0 13156 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1604666999
transform -1 0 14812 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_143
timestamp 1604666999
transform 1 0 14260 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1604666999
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1604666999
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_15
timestamp 1604666999
transform 1 0 2484 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1604666999
transform 1 0 4600 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 4416 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 4048 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3680 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3312 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_23
timestamp 1604666999
transform 1 0 3220 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_26
timestamp 1604666999
transform 1 0 3496 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_30
timestamp 1604666999
transform 1 0 3864 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_34
timestamp 1604666999
transform 1 0 4232 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5796 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_47
timestamp 1604666999
transform 1 0 5428 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_53
timestamp 1604666999
transform 1 0 5980 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1604666999
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7820 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_71
timestamp 1604666999
transform 1 0 7636 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_75
timestamp 1604666999
transform 1 0 8004 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 9660 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_89
timestamp 1604666999
transform 1 0 9292 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_102
timestamp 1604666999
transform 1 0 10488 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_116
timestamp 1604666999
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_120
timestamp 1604666999
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_123
timestamp 1604666999
transform 1 0 12420 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_135
timestamp 1604666999
transform 1 0 13524 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1604666999
transform -1 0 14812 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_51_143
timestamp 1604666999
transform 1 0 14260 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_53_9
timestamp 1604666999
transform 1 0 1932 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_3
timestamp 1604666999
transform 1 0 1380 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1604666999
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1604666999
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_16
timestamp 1604666999
transform 1 0 2576 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_12
timestamp 1604666999
transform 1 0 2208 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_19
timestamp 1604666999
transform 1 0 2852 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1604666999
transform 1 0 2484 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2024 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 2392 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2760 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1604666999
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_29
timestamp 1604666999
transform 1 0 3772 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_23
timestamp 1604666999
transform 1 0 3220 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1604666999
transform 1 0 2944 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604666999
transform 1 0 2944 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_34
timestamp 1604666999
transform 1 0 4232 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4048 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4508 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_46
timestamp 1604666999
transform 1 0 5336 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_45
timestamp 1604666999
transform 1 0 5244 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_41
timestamp 1604666999
transform 1 0 4876 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5060 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5520 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1604666999
transform 1 0 6348 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_54
timestamp 1604666999
transform 1 0 6072 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_50
timestamp 1604666999
transform 1 0 5704 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_53
timestamp 1604666999
transform 1 0 5980 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 6256 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6440 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_53_62
timestamp 1604666999
transform 1 0 6808 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_67
timestamp 1604666999
transform 1 0 7268 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7452 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1604666999
transform 1 0 6900 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_76
timestamp 1604666999
transform 1 0 8096 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_72
timestamp 1604666999
transform 1 0 7728 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_79
timestamp 1604666999
transform 1 0 8372 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_71
timestamp 1604666999
transform 1 0 7636 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8280 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 7912 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_89
timestamp 1604666999
transform 1 0 9292 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_82
timestamp 1604666999
transform 1 0 8648 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 8464 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8464 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1604666999
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_99
timestamp 1604666999
transform 1 0 10212 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_93
timestamp 1604666999
transform 1 0 9660 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_90
timestamp 1604666999
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 9476 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 10028 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1604666999
transform 1 0 10028 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 11592 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10396 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 11040 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_103
timestamp 1604666999
transform 1 0 10580 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_107
timestamp 1604666999
transform 1 0 10948 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_113
timestamp 1604666999
transform 1 0 11500 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_106
timestamp 1604666999
transform 1 0 10856 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_110
timestamp 1604666999
transform 1 0 11224 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 13340 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 13800 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_133
timestamp 1604666999
transform 1 0 13340 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_123
timestamp 1604666999
transform 1 0 12420 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_131
timestamp 1604666999
transform 1 0 13156 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_136
timestamp 1604666999
transform 1 0 13616 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1604666999
transform -1 0 14812 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1604666999
transform -1 0 14812 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1604666999
transform 1 0 14444 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_140
timestamp 1604666999
transform 1 0 13984 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1604666999
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1604666999
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_15
timestamp 1604666999
transform 1 0 2484 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4048 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 3220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_25
timestamp 1604666999
transform 1 0 3404 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 6348 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_51
timestamp 1604666999
transform 1 0 5796 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7728 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8096 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_68
timestamp 1604666999
transform 1 0 7360 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_74
timestamp 1604666999
transform 1 0 7912 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_78
timestamp 1604666999
transform 1 0 8280 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1604666999
transform 1 0 9660 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 8464 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_82
timestamp 1604666999
transform 1 0 8648 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_90
timestamp 1604666999
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 10764 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 11132 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 11500 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_102
timestamp 1604666999
transform 1 0 10488 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_107
timestamp 1604666999
transform 1 0 10948 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_111
timestamp 1604666999
transform 1 0 11316 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_115
timestamp 1604666999
transform 1 0 11684 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 12420 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 12788 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_125
timestamp 1604666999
transform 1 0 12604 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_129
timestamp 1604666999
transform 1 0 12972 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1604666999
transform -1 0 14812 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1604666999
transform 1 0 14076 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_145
timestamp 1604666999
transform 1 0 14444 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1604666999
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1564 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1604666999
transform 1 0 1380 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_7
timestamp 1604666999
transform 1 0 1748 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_19
timestamp 1604666999
transform 1 0 2852 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1604666999
transform 1 0 3220 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3036 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_32
timestamp 1604666999
transform 1 0 4048 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_36
timestamp 1604666999
transform 1 0 4416 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_39
timestamp 1604666999
transform 1 0 4692 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5704 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 6072 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5336 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_45
timestamp 1604666999
transform 1 0 5244 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_48
timestamp 1604666999
transform 1 0 5520 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_52
timestamp 1604666999
transform 1 0 5888 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_56
timestamp 1604666999
transform 1 0 6256 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 7728 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7268 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_62
timestamp 1604666999
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_66
timestamp 1604666999
transform 1 0 7176 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_69
timestamp 1604666999
transform 1 0 7452 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 9844 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_91
timestamp 1604666999
transform 1 0 9476 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_97
timestamp 1604666999
transform 1 0 10028 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10580 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_101
timestamp 1604666999
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_114
timestamp 1604666999
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_118
timestamp 1604666999
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1604666999
transform 1 0 12420 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1604666999
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13432 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_132
timestamp 1604666999
transform 1 0 13248 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_136
timestamp 1604666999
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1604666999
transform -1 0 14812 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_140
timestamp 1604666999
transform 1 0 13984 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1604666999
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_6
timestamp 1604666999
transform 1 0 1656 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_18
timestamp 1604666999
transform 1 0 2760 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1604666999
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 4692 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_22
timestamp 1604666999
transform 1 0 3128 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_25
timestamp 1604666999
transform 1 0 3404 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_32
timestamp 1604666999
transform 1 0 4048 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_38
timestamp 1604666999
transform 1 0 4600 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5704 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1604666999
transform 1 0 4876 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_49
timestamp 1604666999
transform 1 0 5612 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_56_59
timestamp 1604666999
transform 1 0 6532 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7268 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6808 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 8280 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_64
timestamp 1604666999
transform 1 0 6992 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_76
timestamp 1604666999
transform 1 0 8096 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604666999
transform 1 0 9660 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1604666999
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10120 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1604666999
transform 1 0 8464 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_96
timestamp 1604666999
transform 1 0 9936 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1604666999
transform 1 0 10672 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 11776 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 10488 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_100
timestamp 1604666999
transform 1 0 10304 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_113
timestamp 1604666999
transform 1 0 11500 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_56_118
timestamp 1604666999
transform 1 0 11960 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1604666999
transform 1 0 12236 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 13248 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_130
timestamp 1604666999
transform 1 0 13064 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_134
timestamp 1604666999
transform 1 0 13432 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1604666999
transform -1 0 14812 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604666999
transform 1 0 2852 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1604666999
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604666999
transform 1 0 2208 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_6
timestamp 1604666999
transform 1 0 1656 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_10
timestamp 1604666999
transform 1 0 2024 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_14
timestamp 1604666999
transform 1 0 2392 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_18
timestamp 1604666999
transform 1 0 2760 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604666999
transform 1 0 3956 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604666999
transform 1 0 3404 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604666999
transform 1 0 4508 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_23
timestamp 1604666999
transform 1 0 3220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_27
timestamp 1604666999
transform 1 0 3588 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_35
timestamp 1604666999
transform 1 0 4324 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_39
timestamp 1604666999
transform 1 0 4692 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604666999
transform 1 0 5060 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604666999
transform 1 0 5612 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 4876 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_47
timestamp 1604666999
transform 1 0 5428 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1604666999
transform 1 0 5796 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1604666999
transform 1 0 6348 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6808 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1604666999
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604666999
transform 1 0 9476 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604666999
transform 1 0 10028 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 9292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_81
timestamp 1604666999
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_85
timestamp 1604666999
transform 1 0 8924 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_95
timestamp 1604666999
transform 1 0 9844 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_99
timestamp 1604666999
transform 1 0 10212 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 10580 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10396 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_112
timestamp 1604666999
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_116
timestamp 1604666999
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1604666999
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 13432 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 13800 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_120
timestamp 1604666999
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_132
timestamp 1604666999
transform 1 0 13248 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_136
timestamp 1604666999
transform 1 0 13616 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1604666999
transform -1 0 14812 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_57_140
timestamp 1604666999
transform 1 0 13984 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604666999
transform 1 0 2208 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1604666999
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604666999
transform 1 0 1564 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1604666999
transform 1 0 1380 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_7
timestamp 1604666999
transform 1 0 1748 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_11
timestamp 1604666999
transform 1 0 2116 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_16
timestamp 1604666999
transform 1 0 2576 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4692 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1604666999
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3496 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_24
timestamp 1604666999
transform 1 0 3312 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_28
timestamp 1604666999
transform 1 0 3680 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_32
timestamp 1604666999
transform 1 0 4048 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_38
timestamp 1604666999
transform 1 0 4600 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_58
timestamp 1604666999
transform 1 0 6440 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7544 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7360 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 6992 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_66
timestamp 1604666999
transform 1 0 7176 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_79
timestamp 1604666999
transform 1 0 8372 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10120 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1604666999
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_87
timestamp 1604666999
transform 1 0 9108 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1604666999
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_97
timestamp 1604666999
transform 1 0 10028 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11776 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11132 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_107
timestamp 1604666999
transform 1 0 10948 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_111
timestamp 1604666999
transform 1 0 11316 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_115
timestamp 1604666999
transform 1 0 11684 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_135
timestamp 1604666999
transform 1 0 13524 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1604666999
transform -1 0 14812 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_143
timestamp 1604666999
transform 1 0 14260 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_7
timestamp 1604666999
transform 1 0 1748 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_7
timestamp 1604666999
transform 1 0 1748 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604666999
transform 1 0 1932 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1604666999
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1604666999
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604666999
transform 1 0 1380 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604666999
transform 1 0 1380 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_18
timestamp 1604666999
transform 1 0 2760 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_11
timestamp 1604666999
transform 1 0 2116 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2300 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604666999
transform 1 0 2484 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_19
timestamp 1604666999
transform 1 0 2852 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 3496 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1604666999
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604666999
transform 1 0 2944 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3312 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_22
timestamp 1604666999
transform 1 0 3128 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_32
timestamp 1604666999
transform 1 0 4048 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_45
timestamp 1604666999
transform 1 0 5244 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_40
timestamp 1604666999
transform 1 0 4784 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_45
timestamp 1604666999
transform 1 0 5244 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604666999
transform 1 0 5428 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604666999
transform 1 0 4876 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_53
timestamp 1604666999
transform 1 0 5980 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1604666999
transform 1 0 6164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_49
timestamp 1604666999
transform 1 0 5612 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604666999
transform 1 0 6256 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604666999
transform 1 0 6256 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_58
timestamp 1604666999
transform 1 0 6440 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604666999
transform 1 0 7360 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7360 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1604666999
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604666999
transform 1 0 7176 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7912 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_62
timestamp 1604666999
transform 1 0 6808 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_60
timestamp 1604666999
transform 1 0 6624 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_72
timestamp 1604666999
transform 1 0 7728 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_76
timestamp 1604666999
transform 1 0 8096 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_84
timestamp 1604666999
transform 1 0 8832 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_87
timestamp 1604666999
transform 1 0 9108 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604666999
transform 1 0 9292 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604666999
transform 1 0 8464 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_91
timestamp 1604666999
transform 1 0 9476 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9660 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1604666999
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 9844 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9660 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_114
timestamp 1604666999
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_118
timestamp 1604666999
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_112
timestamp 1604666999
transform 1 0 11408 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604666999
transform 1 0 12328 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12420 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1604666999
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 12788 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_132
timestamp 1604666999
transform 1 0 13248 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_120
timestamp 1604666999
transform 1 0 12144 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_125
timestamp 1604666999
transform 1 0 12604 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1604666999
transform 1 0 12972 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1604666999
transform -1 0 14812 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1604666999
transform -1 0 14812 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_144
timestamp 1604666999
transform 1 0 14352 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_141
timestamp 1604666999
transform 1 0 14076 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_145
timestamp 1604666999
transform 1 0 14444 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604666999
transform 1 0 2760 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1604666999
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1604666999
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_15
timestamp 1604666999
transform 1 0 2484 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604666999
transform 1 0 3864 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604666999
transform 1 0 4692 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604666999
transform 1 0 3680 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604666999
transform 1 0 3312 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_22
timestamp 1604666999
transform 1 0 3128 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_26
timestamp 1604666999
transform 1 0 3496 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_34
timestamp 1604666999
transform 1 0 4232 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_38
timestamp 1604666999
transform 1 0 4600 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604666999
transform 1 0 4968 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604666999
transform 1 0 5520 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604666999
transform 1 0 5888 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_41
timestamp 1604666999
transform 1 0 4876 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_46
timestamp 1604666999
transform 1 0 5336 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_50
timestamp 1604666999
transform 1 0 5704 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_54
timestamp 1604666999
transform 1 0 6072 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604666999
transform 1 0 7268 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1604666999
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604666999
transform 1 0 7820 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_60
timestamp 1604666999
transform 1 0 6624 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_62
timestamp 1604666999
transform 1 0 6808 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_66
timestamp 1604666999
transform 1 0 7176 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_71
timestamp 1604666999
transform 1 0 7636 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_75
timestamp 1604666999
transform 1 0 8004 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604666999
transform 1 0 9660 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604666999
transform 1 0 10212 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_61_87
timestamp 1604666999
transform 1 0 9108 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_61_97
timestamp 1604666999
transform 1 0 10028 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_101
timestamp 1604666999
transform 1 0 10396 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_113
timestamp 1604666999
transform 1 0 11500 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1604666999
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1604666999
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1604666999
transform 1 0 12420 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_135
timestamp 1604666999
transform 1 0 13524 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1604666999
transform -1 0 14812 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_143
timestamp 1604666999
transform 1 0 14260 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1604666999
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1604666999
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1604666999
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604666999
transform 1 0 4692 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1604666999
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1604666999
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1604666999
transform 1 0 4048 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_38
timestamp 1604666999
transform 1 0 4600 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604666999
transform 1 0 5796 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_43
timestamp 1604666999
transform 1 0 5060 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_55
timestamp 1604666999
transform 1 0 6164 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_67
timestamp 1604666999
transform 1 0 7268 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_79
timestamp 1604666999
transform 1 0 8372 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1604666999
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_91
timestamp 1604666999
transform 1 0 9476 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1604666999
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1604666999
transform 1 0 10764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1604666999
transform 1 0 11868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1604666999
transform 1 0 12972 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1604666999
transform -1 0 14812 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1604666999
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_145
timestamp 1604666999
transform 1 0 14444 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1604666999
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1604666999
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1604666999
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1604666999
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_39
timestamp 1604666999
transform 1 0 4692 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604666999
transform 1 0 5428 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604666999
transform 1 0 5980 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_51
timestamp 1604666999
transform 1 0 5796 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_55
timestamp 1604666999
transform 1 0 6164 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1604666999
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1604666999
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1604666999
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1604666999
transform 1 0 9016 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1604666999
transform 1 0 10120 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1604666999
transform 1 0 11224 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1604666999
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1604666999
transform 1 0 12420 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_135
timestamp 1604666999
transform 1 0 13524 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1604666999
transform -1 0 14812 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_63_143
timestamp 1604666999
transform 1 0 14260 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1604666999
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1604666999
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1604666999
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1604666999
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1604666999
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1604666999
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1604666999
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_56
timestamp 1604666999
transform 1 0 6256 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1604666999
transform 1 0 6808 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_63
timestamp 1604666999
transform 1 0 6900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_75
timestamp 1604666999
transform 1 0 8004 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1604666999
transform 1 0 9660 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_87
timestamp 1604666999
transform 1 0 9108 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_94
timestamp 1604666999
transform 1 0 9752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_106
timestamp 1604666999
transform 1 0 10856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1604666999
transform 1 0 11960 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1604666999
transform 1 0 12512 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_125
timestamp 1604666999
transform 1 0 12604 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_137
timestamp 1604666999
transform 1 0 13708 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1604666999
transform -1 0 14812 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_64_145
timestamp 1604666999
transform 1 0 14444 0 -1 37536
box -38 -48 130 592
<< labels >>
rlabel metal3 s 0 1096 480 1216 6 ccff_head
port 0 nsew default input
rlabel metal3 s 15520 20000 16000 20120 6 ccff_tail
port 1 nsew default tristate
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[0]
port 2 nsew default input
rlabel metal2 s 12162 0 12218 480 6 chany_bottom_in[10]
port 3 nsew default input
rlabel metal2 s 12530 0 12586 480 6 chany_bottom_in[11]
port 4 nsew default input
rlabel metal2 s 12990 0 13046 480 6 chany_bottom_in[12]
port 5 nsew default input
rlabel metal2 s 13358 0 13414 480 6 chany_bottom_in[13]
port 6 nsew default input
rlabel metal2 s 13726 0 13782 480 6 chany_bottom_in[14]
port 7 nsew default input
rlabel metal2 s 14186 0 14242 480 6 chany_bottom_in[15]
port 8 nsew default input
rlabel metal2 s 14554 0 14610 480 6 chany_bottom_in[16]
port 9 nsew default input
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_in[17]
port 10 nsew default input
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_in[18]
port 11 nsew default input
rlabel metal2 s 15750 0 15806 480 6 chany_bottom_in[19]
port 12 nsew default input
rlabel metal2 s 8574 0 8630 480 6 chany_bottom_in[1]
port 13 nsew default input
rlabel metal2 s 8942 0 8998 480 6 chany_bottom_in[2]
port 14 nsew default input
rlabel metal2 s 9402 0 9458 480 6 chany_bottom_in[3]
port 15 nsew default input
rlabel metal2 s 9770 0 9826 480 6 chany_bottom_in[4]
port 16 nsew default input
rlabel metal2 s 10138 0 10194 480 6 chany_bottom_in[5]
port 17 nsew default input
rlabel metal2 s 10598 0 10654 480 6 chany_bottom_in[6]
port 18 nsew default input
rlabel metal2 s 10966 0 11022 480 6 chany_bottom_in[7]
port 19 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[8]
port 20 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[9]
port 21 nsew default input
rlabel metal2 s 202 0 258 480 6 chany_bottom_out[0]
port 22 nsew default tristate
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_out[10]
port 23 nsew default tristate
rlabel metal2 s 4526 0 4582 480 6 chany_bottom_out[11]
port 24 nsew default tristate
rlabel metal2 s 4986 0 5042 480 6 chany_bottom_out[12]
port 25 nsew default tristate
rlabel metal2 s 5354 0 5410 480 6 chany_bottom_out[13]
port 26 nsew default tristate
rlabel metal2 s 5722 0 5778 480 6 chany_bottom_out[14]
port 27 nsew default tristate
rlabel metal2 s 6182 0 6238 480 6 chany_bottom_out[15]
port 28 nsew default tristate
rlabel metal2 s 6550 0 6606 480 6 chany_bottom_out[16]
port 29 nsew default tristate
rlabel metal2 s 6918 0 6974 480 6 chany_bottom_out[17]
port 30 nsew default tristate
rlabel metal2 s 7378 0 7434 480 6 chany_bottom_out[18]
port 31 nsew default tristate
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_out[19]
port 32 nsew default tristate
rlabel metal2 s 570 0 626 480 6 chany_bottom_out[1]
port 33 nsew default tristate
rlabel metal2 s 938 0 994 480 6 chany_bottom_out[2]
port 34 nsew default tristate
rlabel metal2 s 1398 0 1454 480 6 chany_bottom_out[3]
port 35 nsew default tristate
rlabel metal2 s 1766 0 1822 480 6 chany_bottom_out[4]
port 36 nsew default tristate
rlabel metal2 s 2134 0 2190 480 6 chany_bottom_out[5]
port 37 nsew default tristate
rlabel metal2 s 2594 0 2650 480 6 chany_bottom_out[6]
port 38 nsew default tristate
rlabel metal2 s 2962 0 3018 480 6 chany_bottom_out[7]
port 39 nsew default tristate
rlabel metal2 s 3330 0 3386 480 6 chany_bottom_out[8]
port 40 nsew default tristate
rlabel metal2 s 3790 0 3846 480 6 chany_bottom_out[9]
port 41 nsew default tristate
rlabel metal2 s 8206 39520 8262 40000 6 chany_top_in[0]
port 42 nsew default input
rlabel metal2 s 12162 39520 12218 40000 6 chany_top_in[10]
port 43 nsew default input
rlabel metal2 s 12530 39520 12586 40000 6 chany_top_in[11]
port 44 nsew default input
rlabel metal2 s 12990 39520 13046 40000 6 chany_top_in[12]
port 45 nsew default input
rlabel metal2 s 13358 39520 13414 40000 6 chany_top_in[13]
port 46 nsew default input
rlabel metal2 s 13726 39520 13782 40000 6 chany_top_in[14]
port 47 nsew default input
rlabel metal2 s 14186 39520 14242 40000 6 chany_top_in[15]
port 48 nsew default input
rlabel metal2 s 14554 39520 14610 40000 6 chany_top_in[16]
port 49 nsew default input
rlabel metal2 s 14922 39520 14978 40000 6 chany_top_in[17]
port 50 nsew default input
rlabel metal2 s 15382 39520 15438 40000 6 chany_top_in[18]
port 51 nsew default input
rlabel metal2 s 15750 39520 15806 40000 6 chany_top_in[19]
port 52 nsew default input
rlabel metal2 s 8574 39520 8630 40000 6 chany_top_in[1]
port 53 nsew default input
rlabel metal2 s 8942 39520 8998 40000 6 chany_top_in[2]
port 54 nsew default input
rlabel metal2 s 9402 39520 9458 40000 6 chany_top_in[3]
port 55 nsew default input
rlabel metal2 s 9770 39520 9826 40000 6 chany_top_in[4]
port 56 nsew default input
rlabel metal2 s 10138 39520 10194 40000 6 chany_top_in[5]
port 57 nsew default input
rlabel metal2 s 10598 39520 10654 40000 6 chany_top_in[6]
port 58 nsew default input
rlabel metal2 s 10966 39520 11022 40000 6 chany_top_in[7]
port 59 nsew default input
rlabel metal2 s 11334 39520 11390 40000 6 chany_top_in[8]
port 60 nsew default input
rlabel metal2 s 11794 39520 11850 40000 6 chany_top_in[9]
port 61 nsew default input
rlabel metal2 s 202 39520 258 40000 6 chany_top_out[0]
port 62 nsew default tristate
rlabel metal2 s 4158 39520 4214 40000 6 chany_top_out[10]
port 63 nsew default tristate
rlabel metal2 s 4526 39520 4582 40000 6 chany_top_out[11]
port 64 nsew default tristate
rlabel metal2 s 4986 39520 5042 40000 6 chany_top_out[12]
port 65 nsew default tristate
rlabel metal2 s 5354 39520 5410 40000 6 chany_top_out[13]
port 66 nsew default tristate
rlabel metal2 s 5722 39520 5778 40000 6 chany_top_out[14]
port 67 nsew default tristate
rlabel metal2 s 6182 39520 6238 40000 6 chany_top_out[15]
port 68 nsew default tristate
rlabel metal2 s 6550 39520 6606 40000 6 chany_top_out[16]
port 69 nsew default tristate
rlabel metal2 s 6918 39520 6974 40000 6 chany_top_out[17]
port 70 nsew default tristate
rlabel metal2 s 7378 39520 7434 40000 6 chany_top_out[18]
port 71 nsew default tristate
rlabel metal2 s 7746 39520 7802 40000 6 chany_top_out[19]
port 72 nsew default tristate
rlabel metal2 s 570 39520 626 40000 6 chany_top_out[1]
port 73 nsew default tristate
rlabel metal2 s 938 39520 994 40000 6 chany_top_out[2]
port 74 nsew default tristate
rlabel metal2 s 1398 39520 1454 40000 6 chany_top_out[3]
port 75 nsew default tristate
rlabel metal2 s 1766 39520 1822 40000 6 chany_top_out[4]
port 76 nsew default tristate
rlabel metal2 s 2134 39520 2190 40000 6 chany_top_out[5]
port 77 nsew default tristate
rlabel metal2 s 2594 39520 2650 40000 6 chany_top_out[6]
port 78 nsew default tristate
rlabel metal2 s 2962 39520 3018 40000 6 chany_top_out[7]
port 79 nsew default tristate
rlabel metal2 s 3330 39520 3386 40000 6 chany_top_out[8]
port 80 nsew default tristate
rlabel metal2 s 3790 39520 3846 40000 6 chany_top_out[9]
port 81 nsew default tristate
rlabel metal3 s 0 3408 480 3528 6 left_grid_pin_0_
port 82 nsew default tristate
rlabel metal3 s 0 26936 480 27056 6 left_grid_pin_10_
port 83 nsew default tristate
rlabel metal3 s 0 29248 480 29368 6 left_grid_pin_11_
port 84 nsew default tristate
rlabel metal3 s 0 31560 480 31680 6 left_grid_pin_12_
port 85 nsew default tristate
rlabel metal3 s 0 34008 480 34128 6 left_grid_pin_13_
port 86 nsew default tristate
rlabel metal3 s 0 36320 480 36440 6 left_grid_pin_14_
port 87 nsew default tristate
rlabel metal3 s 0 38632 480 38752 6 left_grid_pin_15_
port 88 nsew default tristate
rlabel metal3 s 0 5720 480 5840 6 left_grid_pin_1_
port 89 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 left_grid_pin_2_
port 90 nsew default tristate
rlabel metal3 s 0 10480 480 10600 6 left_grid_pin_3_
port 91 nsew default tristate
rlabel metal3 s 0 12792 480 12912 6 left_grid_pin_4_
port 92 nsew default tristate
rlabel metal3 s 0 15104 480 15224 6 left_grid_pin_5_
port 93 nsew default tristate
rlabel metal3 s 0 17552 480 17672 6 left_grid_pin_6_
port 94 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_grid_pin_7_
port 95 nsew default tristate
rlabel metal3 s 0 22176 480 22296 6 left_grid_pin_8_
port 96 nsew default tristate
rlabel metal3 s 0 24488 480 24608 6 left_grid_pin_9_
port 97 nsew default tristate
rlabel metal3 s 15520 6672 16000 6792 6 prog_clk
port 98 nsew default input
rlabel metal3 s 15520 33328 16000 33448 6 right_grid_pin_52_
port 99 nsew default tristate
rlabel metal4 s 3611 2128 3931 37584 6 VPWR
port 100 nsew default input
rlabel metal4 s 6277 2128 6597 37584 6 VGND
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 16000 40000
<< end >>
