magic
tech sky130A
magscale 1 2
timestamp 1609022864
<< locali >>
rect 3065 10523 3099 10761
rect 7205 9911 7239 10081
rect 2237 9367 2271 9537
rect 13645 9435 13679 9605
rect 8401 8823 8435 9061
rect 7849 7939 7883 8041
rect 15761 7259 15795 7361
rect 18981 7055 19015 7701
rect 14565 5627 14599 5865
<< viali >>
rect 1409 14569 1443 14603
rect 1593 14433 1627 14467
rect 2145 14433 2179 14467
rect 2789 14433 2823 14467
rect 1777 14365 1811 14399
rect 2329 14365 2363 14399
rect 17969 14229 18003 14263
rect 1501 14025 1535 14059
rect 6377 14025 6411 14059
rect 9413 14025 9447 14059
rect 16681 13957 16715 13991
rect 1777 13889 1811 13923
rect 2421 13889 2455 13923
rect 9873 13889 9907 13923
rect 17141 13889 17175 13923
rect 1593 13821 1627 13855
rect 2145 13821 2179 13855
rect 2697 13821 2731 13855
rect 6193 13821 6227 13855
rect 6561 13821 6595 13855
rect 9597 13821 9631 13855
rect 16865 13821 16899 13855
rect 17417 13821 17451 13855
rect 17785 13821 17819 13855
rect 18061 13821 18095 13855
rect 18337 13821 18371 13855
rect 17601 13685 17635 13719
rect 1501 13481 1535 13515
rect 17417 13481 17451 13515
rect 1685 13345 1719 13379
rect 2053 13345 2087 13379
rect 2605 13345 2639 13379
rect 17601 13345 17635 13379
rect 2329 13277 2363 13311
rect 17877 13277 17911 13311
rect 1869 13209 1903 13243
rect 17785 12937 17819 12971
rect 18061 12733 18095 12767
rect 18337 12665 18371 12699
rect 10241 12257 10275 12291
rect 10333 12189 10367 12223
rect 10517 12189 10551 12223
rect 7941 12053 7975 12087
rect 9873 12053 9907 12087
rect 8217 11849 8251 11883
rect 10333 11849 10367 11883
rect 12081 11849 12115 11883
rect 14289 11849 14323 11883
rect 18153 11849 18187 11883
rect 18429 11849 18463 11883
rect 11161 11781 11195 11815
rect 2605 11713 2639 11747
rect 6561 11713 6595 11747
rect 7665 11713 7699 11747
rect 10793 11713 10827 11747
rect 10977 11713 11011 11747
rect 11713 11713 11747 11747
rect 14841 11713 14875 11747
rect 17693 11713 17727 11747
rect 6285 11645 6319 11679
rect 8401 11645 8435 11679
rect 8668 11645 8702 11679
rect 14473 11645 14507 11679
rect 7481 11577 7515 11611
rect 7941 11577 7975 11611
rect 10149 11577 10183 11611
rect 10701 11577 10735 11611
rect 1961 11509 1995 11543
rect 2329 11509 2363 11543
rect 2421 11509 2455 11543
rect 5917 11509 5951 11543
rect 6377 11509 6411 11543
rect 6837 11509 6871 11543
rect 7113 11509 7147 11543
rect 7573 11509 7607 11543
rect 9781 11509 9815 11543
rect 11529 11509 11563 11543
rect 11621 11509 11655 11543
rect 12265 11509 12299 11543
rect 17785 11509 17819 11543
rect 6745 11305 6779 11339
rect 7573 11305 7607 11339
rect 8861 11305 8895 11339
rect 9965 11305 9999 11339
rect 11713 11305 11747 11339
rect 12081 11305 12115 11339
rect 17969 11305 18003 11339
rect 2504 11237 2538 11271
rect 3709 11237 3743 11271
rect 5540 11237 5574 11271
rect 8769 11237 8803 11271
rect 10508 11237 10542 11271
rect 13737 11237 13771 11271
rect 16957 11237 16991 11271
rect 17233 11237 17267 11271
rect 18337 11237 18371 11271
rect 2237 11169 2271 11203
rect 7113 11169 7147 11203
rect 7941 11169 7975 11203
rect 8033 11169 8067 11203
rect 9229 11169 9263 11203
rect 12909 11169 12943 11203
rect 14841 11169 14875 11203
rect 15557 11169 15591 11203
rect 17877 11169 17911 11203
rect 5273 11101 5307 11135
rect 7205 11101 7239 11135
rect 7297 11101 7331 11135
rect 8125 11101 8159 11135
rect 8953 11101 8987 11135
rect 10241 11101 10275 11135
rect 12173 11101 12207 11135
rect 12265 11101 12299 11135
rect 13001 11101 13035 11135
rect 13093 11101 13127 11135
rect 15301 11101 15335 11135
rect 18061 11101 18095 11135
rect 6653 11033 6687 11067
rect 12541 11033 12575 11067
rect 14565 11033 14599 11067
rect 15025 11033 15059 11067
rect 17325 11033 17359 11067
rect 17509 11033 17543 11067
rect 1685 10965 1719 10999
rect 1869 10965 1903 10999
rect 2145 10965 2179 10999
rect 3617 10965 3651 10999
rect 4261 10965 4295 10999
rect 8401 10965 8435 10999
rect 11621 10965 11655 10999
rect 16681 10965 16715 10999
rect 16773 10965 16807 10999
rect 1409 10761 1443 10795
rect 2237 10761 2271 10795
rect 3065 10761 3099 10795
rect 5917 10761 5951 10795
rect 8217 10761 8251 10795
rect 11161 10761 11195 10795
rect 1869 10625 1903 10659
rect 2053 10625 2087 10659
rect 2789 10625 2823 10659
rect 2605 10557 2639 10591
rect 10149 10693 10183 10727
rect 13829 10693 13863 10727
rect 3709 10625 3743 10659
rect 3985 10625 4019 10659
rect 6377 10625 6411 10659
rect 6561 10625 6595 10659
rect 10977 10625 11011 10659
rect 11713 10625 11747 10659
rect 16037 10625 16071 10659
rect 17693 10625 17727 10659
rect 5457 10557 5491 10591
rect 6285 10557 6319 10591
rect 6837 10557 6871 10591
rect 7104 10557 7138 10591
rect 8769 10557 8803 10591
rect 11529 10557 11563 10591
rect 12449 10557 12483 10591
rect 13921 10557 13955 10591
rect 16221 10557 16255 10591
rect 18061 10557 18095 10591
rect 3065 10489 3099 10523
rect 3617 10489 3651 10523
rect 4252 10489 4286 10523
rect 8401 10489 8435 10523
rect 9036 10489 9070 10523
rect 11621 10489 11655 10523
rect 12265 10489 12299 10523
rect 12716 10489 12750 10523
rect 14188 10489 14222 10523
rect 15761 10489 15795 10523
rect 16488 10489 16522 10523
rect 1777 10421 1811 10455
rect 2697 10421 2731 10455
rect 3157 10421 3191 10455
rect 3525 10421 3559 10455
rect 5365 10421 5399 10455
rect 10333 10421 10367 10455
rect 10701 10421 10735 10455
rect 10793 10421 10827 10455
rect 11989 10421 12023 10455
rect 15301 10421 15335 10455
rect 15393 10421 15427 10455
rect 15853 10421 15887 10455
rect 17601 10421 17635 10455
rect 18245 10421 18279 10455
rect 18429 10421 18463 10455
rect 2881 10217 2915 10251
rect 3157 10217 3191 10251
rect 3525 10217 3559 10251
rect 4353 10217 4387 10251
rect 4721 10217 4755 10251
rect 5181 10217 5215 10251
rect 9873 10217 9907 10251
rect 10701 10217 10735 10251
rect 11069 10217 11103 10251
rect 13369 10217 13403 10251
rect 14565 10217 14599 10251
rect 16773 10217 16807 10251
rect 17141 10217 17175 10251
rect 18061 10217 18095 10251
rect 4813 10149 4847 10183
rect 6101 10149 6135 10183
rect 6653 10149 6687 10183
rect 7818 10149 7852 10183
rect 9229 10149 9263 10183
rect 14657 10149 14691 10183
rect 1676 10081 1710 10115
rect 3617 10081 3651 10115
rect 5549 10081 5583 10115
rect 6561 10081 6595 10115
rect 7021 10081 7055 10115
rect 7205 10081 7239 10115
rect 7481 10081 7515 10115
rect 9505 10081 9539 10115
rect 9689 10081 9723 10115
rect 10241 10081 10275 10115
rect 11713 10081 11747 10115
rect 12164 10081 12198 10115
rect 13737 10081 13771 10115
rect 15568 10081 15602 10115
rect 17969 10081 18003 10115
rect 1409 10013 1443 10047
rect 3801 10013 3835 10047
rect 4997 10013 5031 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 6745 10013 6779 10047
rect 7573 10013 7607 10047
rect 10333 10013 10367 10047
rect 10517 10013 10551 10047
rect 11161 10013 11195 10047
rect 11253 10013 11287 10047
rect 11897 10013 11931 10047
rect 13829 10013 13863 10047
rect 13921 10013 13955 10047
rect 14749 10013 14783 10047
rect 15301 10013 15335 10047
rect 17233 10013 17267 10047
rect 17325 10013 17359 10047
rect 18153 10013 18187 10047
rect 7297 9945 7331 9979
rect 8953 9945 8987 9979
rect 2789 9877 2823 9911
rect 4169 9877 4203 9911
rect 6193 9877 6227 9911
rect 7205 9877 7239 9911
rect 9045 9877 9079 9911
rect 11529 9877 11563 9911
rect 13277 9877 13311 9911
rect 14197 9877 14231 9911
rect 15025 9877 15059 9911
rect 16681 9877 16715 9911
rect 17601 9877 17635 9911
rect 18429 9877 18463 9911
rect 3157 9673 3191 9707
rect 6285 9673 6319 9707
rect 9873 9673 9907 9707
rect 10701 9673 10735 9707
rect 13737 9673 13771 9707
rect 2329 9605 2363 9639
rect 3525 9605 3559 9639
rect 4353 9605 4387 9639
rect 6009 9605 6043 9639
rect 8217 9605 8251 9639
rect 9689 9605 9723 9639
rect 11529 9605 11563 9639
rect 13645 9605 13679 9639
rect 14565 9605 14599 9639
rect 15393 9605 15427 9639
rect 15577 9605 15611 9639
rect 16773 9605 16807 9639
rect 18245 9605 18279 9639
rect 2237 9537 2271 9571
rect 2789 9537 2823 9571
rect 2973 9537 3007 9571
rect 4169 9537 4203 9571
rect 4997 9537 5031 9571
rect 5733 9537 5767 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 11253 9537 11287 9571
rect 12173 9537 12207 9571
rect 13369 9537 13403 9571
rect 1685 9469 1719 9503
rect 2697 9469 2731 9503
rect 3341 9469 3375 9503
rect 6193 9469 6227 9503
rect 6837 9469 6871 9503
rect 8309 9469 8343 9503
rect 11989 9469 12023 9503
rect 12541 9469 12575 9503
rect 14289 9537 14323 9571
rect 15117 9537 15151 9571
rect 16129 9537 16163 9571
rect 17325 9537 17359 9571
rect 14933 9469 14967 9503
rect 16589 9469 16623 9503
rect 17601 9469 17635 9503
rect 18061 9469 18095 9503
rect 3893 9401 3927 9435
rect 5641 9401 5675 9435
rect 7082 9401 7116 9435
rect 8576 9401 8610 9435
rect 10241 9401 10275 9435
rect 11161 9401 11195 9435
rect 13185 9401 13219 9435
rect 13645 9401 13679 9435
rect 17141 9401 17175 9435
rect 17233 9401 17267 9435
rect 1501 9333 1535 9367
rect 1869 9333 1903 9367
rect 2145 9333 2179 9367
rect 2237 9333 2271 9367
rect 3985 9333 4019 9367
rect 4721 9333 4755 9367
rect 4813 9333 4847 9367
rect 5181 9333 5215 9367
rect 5549 9333 5583 9367
rect 6561 9333 6595 9367
rect 11069 9333 11103 9367
rect 11897 9333 11931 9367
rect 12817 9333 12851 9367
rect 13277 9333 13311 9367
rect 14105 9333 14139 9367
rect 14197 9333 14231 9367
rect 15025 9333 15059 9367
rect 15945 9333 15979 9367
rect 16037 9333 16071 9367
rect 16405 9333 16439 9367
rect 17785 9333 17819 9367
rect 18429 9333 18463 9367
rect 6193 9129 6227 9163
rect 6285 9129 6319 9163
rect 6745 9129 6779 9163
rect 9413 9129 9447 9163
rect 11161 9129 11195 9163
rect 11989 9129 12023 9163
rect 12357 9129 12391 9163
rect 12449 9129 12483 9163
rect 12817 9129 12851 9163
rect 15025 9129 15059 9163
rect 17417 9129 17451 9163
rect 1952 9061 1986 9095
rect 3433 9061 3467 9095
rect 8033 9061 8067 9095
rect 8401 9061 8435 9095
rect 9934 9061 9968 9095
rect 11529 9061 11563 9095
rect 13890 9061 13924 9095
rect 15660 9061 15694 9095
rect 17325 9061 17359 9095
rect 1685 8993 1719 9027
rect 3525 8993 3559 9027
rect 4813 8993 4847 9027
rect 5080 8993 5114 9027
rect 6653 8993 6687 9027
rect 7941 8993 7975 9027
rect 4169 8925 4203 8959
rect 6929 8925 6963 8959
rect 7481 8925 7515 8959
rect 8217 8925 8251 8959
rect 3065 8857 3099 8891
rect 7573 8857 7607 8891
rect 8861 8993 8895 9027
rect 8953 8993 8987 9027
rect 9689 8993 9723 9027
rect 13185 8993 13219 9027
rect 17877 8993 17911 9027
rect 18245 8993 18279 9027
rect 9137 8925 9171 8959
rect 11621 8925 11655 8959
rect 11713 8925 11747 8959
rect 12541 8925 12575 8959
rect 13277 8925 13311 8959
rect 13461 8925 13495 8959
rect 13645 8925 13679 8959
rect 15393 8925 15427 8959
rect 17509 8925 17543 8959
rect 11069 8857 11103 8891
rect 18429 8857 18463 8891
rect 1501 8789 1535 8823
rect 3157 8789 3191 8823
rect 3709 8789 3743 8823
rect 4353 8789 4387 8823
rect 4629 8789 4663 8823
rect 8401 8789 8435 8823
rect 8493 8789 8527 8823
rect 16773 8789 16807 8823
rect 16957 8789 16991 8823
rect 18061 8789 18095 8823
rect 5917 8585 5951 8619
rect 6193 8585 6227 8619
rect 8217 8585 8251 8619
rect 11897 8585 11931 8619
rect 13185 8585 13219 8619
rect 14105 8585 14139 8619
rect 16129 8585 16163 8619
rect 11989 8517 12023 8551
rect 12725 8517 12759 8551
rect 18245 8517 18279 8551
rect 1593 8449 1627 8483
rect 10241 8449 10275 8483
rect 13829 8449 13863 8483
rect 16313 8449 16347 8483
rect 3065 8381 3099 8415
rect 4537 8381 4571 8415
rect 6837 8381 6871 8415
rect 8309 8381 8343 8415
rect 8576 8381 8610 8415
rect 10333 8381 10367 8415
rect 10517 8381 10551 8415
rect 12173 8381 12207 8415
rect 12909 8381 12943 8415
rect 14197 8381 14231 8415
rect 14381 8381 14415 8415
rect 15945 8381 15979 8415
rect 16580 8381 16614 8415
rect 18061 8381 18095 8415
rect 1860 8313 1894 8347
rect 3310 8313 3344 8347
rect 4782 8313 4816 8347
rect 6377 8313 6411 8347
rect 7104 8313 7138 8347
rect 10057 8313 10091 8347
rect 10784 8313 10818 8347
rect 13645 8313 13679 8347
rect 14648 8313 14682 8347
rect 1409 8245 1443 8279
rect 2973 8245 3007 8279
rect 4445 8245 4479 8279
rect 6469 8245 6503 8279
rect 9689 8245 9723 8279
rect 9873 8245 9907 8279
rect 12449 8245 12483 8279
rect 13001 8245 13035 8279
rect 13553 8245 13587 8279
rect 15761 8245 15795 8279
rect 17693 8245 17727 8279
rect 17785 8245 17819 8279
rect 18429 8245 18463 8279
rect 3065 8041 3099 8075
rect 3893 8041 3927 8075
rect 4445 8041 4479 8075
rect 7389 8041 7423 8075
rect 7849 8041 7883 8075
rect 8125 8041 8159 8075
rect 8493 8041 8527 8075
rect 11529 8041 11563 8075
rect 13921 8041 13955 8075
rect 14289 8041 14323 8075
rect 15761 8041 15795 8075
rect 17693 8041 17727 8075
rect 3157 7973 3191 8007
rect 5273 7973 5307 8007
rect 5733 7973 5767 8007
rect 11989 7973 12023 8007
rect 12716 7973 12750 8007
rect 15853 7973 15887 8007
rect 1593 7905 1627 7939
rect 2237 7905 2271 7939
rect 5917 7905 5951 7939
rect 6184 7905 6218 7939
rect 7849 7905 7883 7939
rect 9413 7905 9447 7939
rect 9689 7905 9723 7939
rect 11897 7905 11931 7939
rect 16313 7905 16347 7939
rect 16865 7905 16899 7939
rect 18153 7905 18187 7939
rect 2329 7837 2363 7871
rect 2513 7837 2547 7871
rect 3249 7837 3283 7871
rect 4537 7837 4571 7871
rect 4629 7837 4663 7871
rect 5365 7837 5399 7871
rect 5457 7837 5491 7871
rect 7665 7837 7699 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 12081 7837 12115 7871
rect 12449 7837 12483 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 15945 7837 15979 7871
rect 16957 7837 16991 7871
rect 17049 7837 17083 7871
rect 17785 7837 17819 7871
rect 17877 7837 17911 7871
rect 7297 7769 7331 7803
rect 13829 7769 13863 7803
rect 1685 7701 1719 7735
rect 1869 7701 1903 7735
rect 2697 7701 2731 7735
rect 3617 7701 3651 7735
rect 4077 7701 4111 7735
rect 4905 7701 4939 7735
rect 8033 7701 8067 7735
rect 8953 7701 8987 7735
rect 10977 7701 11011 7735
rect 14841 7701 14875 7735
rect 15025 7701 15059 7735
rect 15393 7701 15427 7735
rect 16497 7701 16531 7735
rect 17325 7701 17359 7735
rect 18337 7701 18371 7735
rect 18981 7701 19015 7735
rect 2605 7497 2639 7531
rect 2789 7497 2823 7531
rect 6561 7497 6595 7531
rect 8125 7497 8159 7531
rect 8953 7497 8987 7531
rect 13829 7497 13863 7531
rect 14197 7497 14231 7531
rect 6837 7429 6871 7463
rect 9781 7429 9815 7463
rect 11529 7429 11563 7463
rect 2237 7361 2271 7395
rect 2421 7361 2455 7395
rect 3341 7361 3375 7395
rect 4169 7361 4203 7395
rect 4537 7361 4571 7395
rect 5181 7361 5215 7395
rect 5917 7361 5951 7395
rect 6009 7361 6043 7395
rect 7389 7361 7423 7395
rect 8677 7361 8711 7395
rect 9505 7361 9539 7395
rect 10241 7361 10275 7395
rect 10333 7361 10367 7395
rect 11161 7361 11195 7395
rect 12173 7361 12207 7395
rect 14289 7361 14323 7395
rect 15761 7361 15795 7395
rect 16589 7361 16623 7395
rect 16681 7361 16715 7395
rect 17509 7361 17543 7395
rect 1409 7293 1443 7327
rect 2145 7293 2179 7327
rect 3249 7293 3283 7327
rect 3985 7293 4019 7327
rect 4997 7293 5031 7327
rect 6285 7293 6319 7327
rect 7297 7293 7331 7327
rect 7665 7293 7699 7327
rect 9321 7293 9355 7327
rect 9413 7293 9447 7327
rect 10977 7293 11011 7327
rect 12449 7293 12483 7327
rect 12705 7293 12739 7327
rect 14013 7293 14047 7327
rect 17325 7293 17359 7327
rect 17785 7293 17819 7327
rect 18061 7293 18095 7327
rect 18429 7293 18463 7327
rect 4077 7225 4111 7259
rect 5825 7225 5859 7259
rect 7205 7225 7239 7259
rect 7941 7225 7975 7259
rect 8493 7225 8527 7259
rect 10149 7225 10183 7259
rect 11069 7225 11103 7259
rect 14556 7225 14590 7259
rect 15761 7225 15795 7259
rect 16497 7225 16531 7259
rect 17417 7225 17451 7259
rect 1593 7157 1627 7191
rect 1777 7157 1811 7191
rect 3157 7157 3191 7191
rect 3617 7157 3651 7191
rect 4629 7157 4663 7191
rect 5089 7157 5123 7191
rect 5457 7157 5491 7191
rect 8585 7157 8619 7191
rect 10609 7157 10643 7191
rect 11897 7157 11931 7191
rect 11989 7157 12023 7191
rect 15669 7157 15703 7191
rect 15853 7157 15887 7191
rect 16129 7157 16163 7191
rect 16957 7157 16991 7191
rect 18245 7157 18279 7191
rect 18981 7021 19015 7055
rect 9413 6953 9447 6987
rect 12909 6953 12943 6987
rect 13369 6953 13403 6987
rect 13737 6953 13771 6987
rect 14105 6953 14139 6987
rect 14749 6953 14783 6987
rect 17325 6953 17359 6987
rect 3525 6885 3559 6919
rect 6653 6885 6687 6919
rect 12449 6885 12483 6919
rect 14933 6885 14967 6919
rect 15730 6885 15764 6919
rect 17417 6885 17451 6919
rect 18153 6885 18187 6919
rect 1860 6817 1894 6851
rect 3617 6817 3651 6851
rect 4445 6817 4479 6851
rect 4537 6817 4571 6851
rect 5172 6817 5206 6851
rect 6561 6817 6595 6851
rect 7205 6817 7239 6851
rect 8024 6817 8058 6851
rect 10425 6817 10459 6851
rect 10517 6817 10551 6851
rect 11152 6817 11186 6851
rect 13277 6817 13311 6851
rect 18245 6817 18279 6851
rect 1593 6749 1627 6783
rect 3801 6749 3835 6783
rect 4629 6749 4663 6783
rect 4905 6749 4939 6783
rect 7297 6749 7331 6783
rect 7389 6749 7423 6783
rect 7757 6749 7791 6783
rect 9781 6749 9815 6783
rect 10701 6749 10735 6783
rect 10885 6749 10919 6783
rect 12633 6749 12667 6783
rect 13553 6749 13587 6783
rect 14197 6749 14231 6783
rect 14289 6749 14323 6783
rect 15485 6749 15519 6783
rect 17509 6749 17543 6783
rect 18337 6749 18371 6783
rect 3157 6681 3191 6715
rect 6837 6681 6871 6715
rect 9321 6681 9355 6715
rect 15393 6681 15427 6715
rect 17785 6681 17819 6715
rect 1409 6613 1443 6647
rect 2973 6613 3007 6647
rect 4077 6613 4111 6647
rect 6285 6613 6319 6647
rect 6377 6613 6411 6647
rect 9137 6613 9171 6647
rect 10057 6613 10091 6647
rect 12265 6613 12299 6647
rect 12725 6613 12759 6647
rect 15117 6613 15151 6647
rect 16865 6613 16899 6647
rect 16957 6613 16991 6647
rect 4629 6409 4663 6443
rect 6469 6409 6503 6443
rect 9873 6409 9907 6443
rect 11529 6409 11563 6443
rect 15669 6409 15703 6443
rect 15209 6341 15243 6375
rect 15393 6341 15427 6375
rect 2697 6273 2731 6307
rect 2973 6273 3007 6307
rect 4813 6273 4847 6307
rect 5089 6273 5123 6307
rect 8401 6273 8435 6307
rect 10517 6273 10551 6307
rect 11345 6273 11379 6307
rect 12173 6273 12207 6307
rect 13645 6273 13679 6307
rect 16221 6273 16255 6307
rect 16313 6273 16347 6307
rect 17049 6273 17083 6307
rect 17141 6273 17175 6307
rect 1685 6205 1719 6239
rect 2513 6205 2547 6239
rect 3229 6205 3263 6239
rect 4445 6205 4479 6239
rect 6561 6205 6595 6239
rect 6837 6205 6871 6239
rect 11069 6205 11103 6239
rect 12449 6205 12483 6239
rect 12817 6205 12851 6239
rect 13461 6205 13495 6239
rect 13829 6205 13863 6239
rect 16957 6205 16991 6239
rect 17601 6205 17635 6239
rect 18061 6205 18095 6239
rect 18429 6205 18463 6239
rect 1593 6137 1627 6171
rect 5356 6137 5390 6171
rect 7104 6137 7138 6171
rect 8668 6137 8702 6171
rect 10241 6137 10275 6171
rect 11161 6137 11195 6171
rect 11989 6137 12023 6171
rect 14096 6137 14130 6171
rect 16129 6137 16163 6171
rect 17417 6137 17451 6171
rect 1869 6069 1903 6103
rect 2145 6069 2179 6103
rect 2605 6069 2639 6103
rect 4353 6069 4387 6103
rect 8217 6069 8251 6103
rect 9781 6069 9815 6103
rect 10333 6069 10367 6103
rect 10701 6069 10735 6103
rect 11897 6069 11931 6103
rect 13001 6069 13035 6103
rect 13369 6069 13403 6103
rect 15761 6069 15795 6103
rect 16589 6069 16623 6103
rect 17785 6069 17819 6103
rect 18245 6069 18279 6103
rect 1961 5865 1995 5899
rect 2329 5865 2363 5899
rect 3157 5865 3191 5899
rect 5917 5865 5951 5899
rect 6009 5865 6043 5899
rect 6377 5865 6411 5899
rect 7389 5865 7423 5899
rect 8217 5865 8251 5899
rect 11253 5865 11287 5899
rect 12081 5865 12115 5899
rect 13737 5865 13771 5899
rect 14105 5865 14139 5899
rect 14565 5865 14599 5899
rect 14933 5865 14967 5899
rect 15761 5865 15795 5899
rect 3525 5797 3559 5831
rect 6837 5797 6871 5831
rect 8677 5797 8711 5831
rect 9045 5797 9079 5831
rect 13553 5797 13587 5831
rect 1869 5729 1903 5763
rect 2697 5729 2731 5763
rect 4344 5729 4378 5763
rect 6745 5729 6779 5763
rect 7757 5729 7791 5763
rect 8585 5729 8619 5763
rect 10048 5729 10082 5763
rect 11621 5729 11655 5763
rect 12449 5729 12483 5763
rect 12909 5729 12943 5763
rect 13001 5729 13035 5763
rect 14197 5729 14231 5763
rect 2145 5661 2179 5695
rect 2789 5661 2823 5695
rect 2973 5661 3007 5695
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 6193 5661 6227 5695
rect 6929 5661 6963 5695
rect 7297 5661 7331 5695
rect 7849 5661 7883 5695
rect 8033 5661 8067 5695
rect 8769 5661 8803 5695
rect 9229 5661 9263 5695
rect 9781 5661 9815 5695
rect 11713 5661 11747 5695
rect 11897 5661 11931 5695
rect 13185 5661 13219 5695
rect 14289 5661 14323 5695
rect 14657 5797 14691 5831
rect 15669 5797 15703 5831
rect 16672 5797 16706 5831
rect 15025 5729 15059 5763
rect 16405 5729 16439 5763
rect 17877 5729 17911 5763
rect 18245 5729 18279 5763
rect 15853 5661 15887 5695
rect 16129 5661 16163 5695
rect 5549 5593 5583 5627
rect 9413 5593 9447 5627
rect 13369 5593 13403 5627
rect 14565 5593 14599 5627
rect 1501 5525 1535 5559
rect 5457 5525 5491 5559
rect 11161 5525 11195 5559
rect 12265 5525 12299 5559
rect 12541 5525 12575 5559
rect 15301 5525 15335 5559
rect 17785 5525 17819 5559
rect 18061 5525 18095 5559
rect 18429 5525 18463 5559
rect 2605 5321 2639 5355
rect 3433 5321 3467 5355
rect 6929 5321 6963 5355
rect 7757 5321 7791 5355
rect 10333 5321 10367 5355
rect 13921 5321 13955 5355
rect 15025 5321 15059 5355
rect 18429 5321 18463 5355
rect 4445 5253 4479 5287
rect 13829 5253 13863 5287
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 3249 5185 3283 5219
rect 3985 5185 4019 5219
rect 7389 5185 7423 5219
rect 7573 5185 7607 5219
rect 8309 5185 8343 5219
rect 8585 5185 8619 5219
rect 10885 5185 10919 5219
rect 12449 5185 12483 5219
rect 14473 5185 14507 5219
rect 16129 5185 16163 5219
rect 16773 5185 16807 5219
rect 16865 5185 16899 5219
rect 17693 5185 17727 5219
rect 1409 5117 1443 5151
rect 2145 5117 2179 5151
rect 3801 5117 3835 5151
rect 4261 5117 4295 5151
rect 4721 5117 4755 5151
rect 4988 5117 5022 5151
rect 6377 5117 6411 5151
rect 6653 5117 6687 5151
rect 8217 5117 8251 5151
rect 8953 5117 8987 5151
rect 9220 5117 9254 5151
rect 10609 5117 10643 5151
rect 11152 5117 11186 5151
rect 12705 5117 12739 5151
rect 14933 5117 14967 5151
rect 15945 5117 15979 5151
rect 18061 5117 18095 5151
rect 8125 5049 8159 5083
rect 15393 5049 15427 5083
rect 16681 5049 16715 5083
rect 1593 4981 1627 5015
rect 1777 4981 1811 5015
rect 2973 4981 3007 5015
rect 3065 4981 3099 5015
rect 3893 4981 3927 5015
rect 6101 4981 6135 5015
rect 6193 4981 6227 5015
rect 6469 4981 6503 5015
rect 7297 4981 7331 5015
rect 10425 4981 10459 5015
rect 10793 4981 10827 5015
rect 12265 4981 12299 5015
rect 14289 4981 14323 5015
rect 14381 4981 14415 5015
rect 14749 4981 14783 5015
rect 15485 4981 15519 5015
rect 15853 4981 15887 5015
rect 16313 4981 16347 5015
rect 17141 4981 17175 5015
rect 17509 4981 17543 5015
rect 17601 4981 17635 5015
rect 18245 4981 18279 5015
rect 1593 4777 1627 4811
rect 3893 4777 3927 4811
rect 7113 4777 7147 4811
rect 8585 4777 8619 4811
rect 9137 4777 9171 4811
rect 10333 4777 10367 4811
rect 10885 4777 10919 4811
rect 11713 4777 11747 4811
rect 12081 4777 12115 4811
rect 12909 4777 12943 4811
rect 13369 4777 13403 4811
rect 2780 4709 2814 4743
rect 4537 4709 4571 4743
rect 6561 4709 6595 4743
rect 11621 4709 11655 4743
rect 13277 4709 13311 4743
rect 15568 4709 15602 4743
rect 16957 4709 16991 4743
rect 17509 4709 17543 4743
rect 1685 4641 1719 4675
rect 2053 4641 2087 4675
rect 4261 4641 4295 4675
rect 4813 4641 4847 4675
rect 5365 4641 5399 4675
rect 5825 4641 5859 4675
rect 6377 4641 6411 4675
rect 7472 4641 7506 4675
rect 9229 4641 9263 4675
rect 9689 4641 9723 4675
rect 10793 4641 10827 4675
rect 12449 4641 12483 4675
rect 13993 4641 14027 4675
rect 16773 4641 16807 4675
rect 17969 4641 18003 4675
rect 18337 4641 18371 4675
rect 2513 4573 2547 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 7205 4573 7239 4607
rect 9413 4573 9447 4607
rect 11069 4573 11103 4607
rect 11897 4573 11931 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 15301 4573 15335 4607
rect 17601 4573 17635 4607
rect 17693 4573 17727 4607
rect 6193 4505 6227 4539
rect 1869 4437 1903 4471
rect 2237 4437 2271 4471
rect 4077 4437 4111 4471
rect 4445 4437 4479 4471
rect 4997 4437 5031 4471
rect 6009 4437 6043 4471
rect 6745 4437 6779 4471
rect 8769 4437 8803 4471
rect 9873 4437 9907 4471
rect 10149 4437 10183 4471
rect 10425 4437 10459 4471
rect 11253 4437 11287 4471
rect 15117 4437 15151 4471
rect 16681 4437 16715 4471
rect 17141 4437 17175 4471
rect 18153 4437 18187 4471
rect 8217 4233 8251 4267
rect 12173 4233 12207 4267
rect 13737 4233 13771 4267
rect 3433 4165 3467 4199
rect 10149 4165 10183 4199
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 4537 4097 4571 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 6101 4097 6135 4131
rect 9873 4097 9907 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 11529 4097 11563 4131
rect 12449 4097 12483 4131
rect 12817 4097 12851 4131
rect 13461 4097 13495 4131
rect 14289 4097 14323 4131
rect 14565 4097 14599 4131
rect 15301 4097 15335 4131
rect 17233 4097 17267 4131
rect 17417 4097 17451 4131
rect 1501 4029 1535 4063
rect 1869 4029 1903 4063
rect 2237 4029 2271 4063
rect 2973 4029 3007 4063
rect 6837 4029 6871 4063
rect 8309 4029 8343 4063
rect 13369 4029 13403 4063
rect 14105 4029 14139 4063
rect 14841 4029 14875 4063
rect 15568 4029 15602 4063
rect 17141 4029 17175 4063
rect 17601 4029 17635 4063
rect 18061 4029 18095 4063
rect 18429 4029 18463 4063
rect 4261 3961 4295 3995
rect 5917 3961 5951 3995
rect 7082 3961 7116 3995
rect 8576 3961 8610 3995
rect 11437 3961 11471 3995
rect 11989 3961 12023 3995
rect 15025 3961 15059 3995
rect 1685 3893 1719 3927
rect 2053 3893 2087 3927
rect 2421 3893 2455 3927
rect 2605 3893 2639 3927
rect 3709 3893 3743 3927
rect 3893 3893 3927 3927
rect 4353 3893 4387 3927
rect 4721 3893 4755 3927
rect 5089 3893 5123 3927
rect 5549 3893 5583 3927
rect 6009 3893 6043 3927
rect 6377 3893 6411 3927
rect 9689 3893 9723 3927
rect 10057 3893 10091 3927
rect 10517 3893 10551 3927
rect 10977 3893 11011 3927
rect 11345 3893 11379 3927
rect 11805 3893 11839 3927
rect 12909 3893 12943 3927
rect 13277 3893 13311 3927
rect 14197 3893 14231 3927
rect 16681 3893 16715 3927
rect 16773 3893 16807 3927
rect 17785 3893 17819 3927
rect 18245 3893 18279 3927
rect 2789 3689 2823 3723
rect 3617 3689 3651 3723
rect 7297 3689 7331 3723
rect 9137 3689 9171 3723
rect 9229 3689 9263 3723
rect 15945 3689 15979 3723
rect 16865 3689 16899 3723
rect 17325 3689 17359 3723
rect 17509 3689 17543 3723
rect 5794 3621 5828 3655
rect 7757 3621 7791 3655
rect 8493 3621 8527 3655
rect 13176 3621 13210 3655
rect 14381 3621 14415 3655
rect 15393 3621 15427 3655
rect 16773 3621 16807 3655
rect 1665 3553 1699 3587
rect 2881 3553 2915 3587
rect 3525 3553 3559 3587
rect 4077 3553 4111 3587
rect 4344 3553 4378 3587
rect 7205 3553 7239 3587
rect 7665 3553 7699 3587
rect 8217 3553 8251 3587
rect 9689 3553 9723 3587
rect 9956 3553 9990 3587
rect 11693 3553 11727 3587
rect 12909 3553 12943 3587
rect 14657 3553 14691 3587
rect 16037 3553 16071 3587
rect 17877 3553 17911 3587
rect 18245 3553 18279 3587
rect 1409 3485 1443 3519
rect 3801 3485 3835 3519
rect 5549 3485 5583 3519
rect 7941 3485 7975 3519
rect 9413 3485 9447 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 14933 3485 14967 3519
rect 16129 3485 16163 3519
rect 16957 3485 16991 3519
rect 17785 3485 17819 3519
rect 5457 3417 5491 3451
rect 12817 3417 12851 3451
rect 3157 3349 3191 3383
rect 6929 3349 6963 3383
rect 8769 3349 8803 3383
rect 11069 3349 11103 3383
rect 14289 3349 14323 3383
rect 15577 3349 15611 3383
rect 16405 3349 16439 3383
rect 18061 3349 18095 3383
rect 18429 3349 18463 3383
rect 4261 3145 4295 3179
rect 8217 3145 8251 3179
rect 9045 3145 9079 3179
rect 12725 3145 12759 3179
rect 17417 3145 17451 3179
rect 17601 3145 17635 3179
rect 7297 3077 7331 3111
rect 10609 3077 10643 3111
rect 14749 3077 14783 3111
rect 17785 3077 17819 3111
rect 4905 3009 4939 3043
rect 5641 3009 5675 3043
rect 6469 3009 6503 3043
rect 8861 3009 8895 3043
rect 9505 3009 9539 3043
rect 9597 3009 9631 3043
rect 11161 3009 11195 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 13369 3009 13403 3043
rect 13737 3009 13771 3043
rect 14289 3009 14323 3043
rect 15117 3009 15151 3043
rect 16037 3009 16071 3043
rect 16681 3009 16715 3043
rect 16865 3009 16899 3043
rect 17049 3009 17083 3043
rect 1409 2941 1443 2975
rect 1777 2941 1811 2975
rect 2145 2941 2179 2975
rect 2513 2941 2547 2975
rect 2973 2941 3007 2975
rect 3525 2941 3559 2975
rect 3893 2941 3927 2975
rect 5457 2941 5491 2975
rect 6285 2941 6319 2975
rect 6377 2941 6411 2975
rect 6837 2941 6871 2975
rect 7665 2941 7699 2975
rect 7941 2941 7975 2975
rect 9413 2941 9447 2975
rect 10057 2941 10091 2975
rect 11069 2941 11103 2975
rect 11805 2941 11839 2975
rect 13093 2941 13127 2975
rect 13553 2941 13587 2975
rect 14105 2941 14139 2975
rect 15209 2941 15243 2975
rect 15761 2941 15795 2975
rect 17233 2941 17267 2975
rect 18061 2941 18095 2975
rect 3249 2873 3283 2907
rect 4629 2873 4663 2907
rect 7573 2873 7607 2907
rect 8677 2873 8711 2907
rect 9965 2873 9999 2907
rect 10517 2873 10551 2907
rect 14841 2873 14875 2907
rect 16589 2873 16623 2907
rect 18337 2873 18371 2907
rect 1593 2805 1627 2839
rect 1961 2805 1995 2839
rect 2329 2805 2363 2839
rect 2697 2805 2731 2839
rect 3709 2805 3743 2839
rect 4077 2805 4111 2839
rect 4721 2805 4755 2839
rect 5089 2805 5123 2839
rect 5549 2805 5583 2839
rect 5917 2805 5951 2839
rect 7113 2805 7147 2839
rect 8585 2805 8619 2839
rect 10241 2805 10275 2839
rect 10977 2805 11011 2839
rect 11437 2805 11471 2839
rect 11897 2805 11931 2839
rect 12541 2805 12575 2839
rect 15393 2805 15427 2839
rect 15853 2805 15887 2839
rect 16221 2805 16255 2839
rect 1501 2601 1535 2635
rect 6009 2601 6043 2635
rect 6193 2601 6227 2635
rect 8033 2601 8067 2635
rect 8401 2601 8435 2635
rect 8861 2601 8895 2635
rect 9321 2601 9355 2635
rect 11069 2601 11103 2635
rect 11161 2601 11195 2635
rect 11989 2601 12023 2635
rect 13001 2601 13035 2635
rect 15209 2601 15243 2635
rect 17049 2601 17083 2635
rect 18429 2601 18463 2635
rect 5825 2533 5859 2567
rect 8493 2533 8527 2567
rect 9229 2533 9263 2567
rect 10241 2533 10275 2567
rect 10333 2533 10367 2567
rect 14289 2533 14323 2567
rect 17141 2533 17175 2567
rect 1593 2465 1627 2499
rect 1961 2465 1995 2499
rect 2513 2465 2547 2499
rect 2881 2465 2915 2499
rect 3433 2465 3467 2499
rect 4169 2465 4203 2499
rect 4721 2465 4755 2499
rect 5273 2465 5307 2499
rect 6929 2465 6963 2499
rect 7481 2465 7515 2499
rect 11897 2465 11931 2499
rect 13461 2465 13495 2499
rect 14013 2465 14047 2499
rect 14565 2465 14599 2499
rect 15485 2465 15519 2499
rect 17325 2465 17359 2499
rect 17693 2465 17727 2499
rect 2145 2397 2179 2431
rect 3617 2397 3651 2431
rect 4353 2397 4387 2431
rect 4905 2397 4939 2431
rect 5549 2397 5583 2431
rect 7113 2397 7147 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9413 2397 9447 2431
rect 10425 2397 10459 2431
rect 11253 2397 11287 2431
rect 12081 2397 12115 2431
rect 12449 2397 12483 2431
rect 13093 2397 13127 2431
rect 13185 2397 13219 2431
rect 13645 2397 13679 2431
rect 14749 2397 14783 2431
rect 15669 2397 15703 2431
rect 17969 2397 18003 2431
rect 2697 2329 2731 2363
rect 6377 2329 6411 2363
rect 9873 2329 9907 2363
rect 10701 2329 10735 2363
rect 1777 2261 1811 2295
rect 3065 2261 3099 2295
rect 3341 2261 3375 2295
rect 6561 2261 6595 2295
rect 11529 2261 11563 2295
rect 12633 2261 12667 2295
rect 17509 2261 17543 2295
<< metal1 >>
rect 4062 15172 4068 15224
rect 4120 15212 4126 15224
rect 9398 15212 9404 15224
rect 4120 15184 9404 15212
rect 4120 15172 4126 15184
rect 9398 15172 9404 15184
rect 9456 15172 9462 15224
rect 1104 14714 18860 14736
rect 1104 14662 6912 14714
rect 6964 14662 6976 14714
rect 7028 14662 7040 14714
rect 7092 14662 7104 14714
rect 7156 14662 12843 14714
rect 12895 14662 12907 14714
rect 12959 14662 12971 14714
rect 13023 14662 13035 14714
rect 13087 14662 18860 14714
rect 1104 14640 18860 14662
rect 1394 14600 1400 14612
rect 1355 14572 1400 14600
rect 1394 14560 1400 14572
rect 1452 14560 1458 14612
rect 1412 14464 1440 14560
rect 1581 14467 1639 14473
rect 1581 14464 1593 14467
rect 1412 14436 1593 14464
rect 1581 14433 1593 14436
rect 1627 14464 1639 14467
rect 2038 14464 2044 14476
rect 1627 14436 2044 14464
rect 1627 14433 1639 14436
rect 1581 14427 1639 14433
rect 2038 14424 2044 14436
rect 2096 14424 2102 14476
rect 2133 14467 2191 14473
rect 2133 14433 2145 14467
rect 2179 14464 2191 14467
rect 2777 14467 2835 14473
rect 2777 14464 2789 14467
rect 2179 14436 2789 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 2777 14433 2789 14436
rect 2823 14464 2835 14467
rect 2866 14464 2872 14476
rect 2823 14436 2872 14464
rect 2823 14433 2835 14436
rect 2777 14427 2835 14433
rect 2866 14424 2872 14436
rect 2924 14464 2930 14476
rect 3694 14464 3700 14476
rect 2924 14436 3700 14464
rect 2924 14424 2930 14436
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 1762 14396 1768 14408
rect 1723 14368 1768 14396
rect 1762 14356 1768 14368
rect 1820 14356 1826 14408
rect 2314 14396 2320 14408
rect 2275 14368 2320 14396
rect 2314 14356 2320 14368
rect 2372 14356 2378 14408
rect 1946 14288 1952 14340
rect 2004 14328 2010 14340
rect 17310 14328 17316 14340
rect 2004 14300 17316 14328
rect 2004 14288 2010 14300
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 3786 14220 3792 14272
rect 3844 14260 3850 14272
rect 17957 14263 18015 14269
rect 17957 14260 17969 14263
rect 3844 14232 17969 14260
rect 3844 14220 3850 14232
rect 17957 14229 17969 14232
rect 18003 14260 18015 14263
rect 18046 14260 18052 14272
rect 18003 14232 18052 14260
rect 18003 14229 18015 14232
rect 17957 14223 18015 14229
rect 18046 14220 18052 14232
rect 18104 14220 18110 14272
rect 1104 14170 18860 14192
rect 1104 14118 3947 14170
rect 3999 14118 4011 14170
rect 4063 14118 4075 14170
rect 4127 14118 4139 14170
rect 4191 14118 9878 14170
rect 9930 14118 9942 14170
rect 9994 14118 10006 14170
rect 10058 14118 10070 14170
rect 10122 14118 15808 14170
rect 15860 14118 15872 14170
rect 15924 14118 15936 14170
rect 15988 14118 16000 14170
rect 16052 14118 18860 14170
rect 1104 14096 18860 14118
rect 1489 14059 1547 14065
rect 1489 14025 1501 14059
rect 1535 14056 1547 14059
rect 2958 14056 2964 14068
rect 1535 14028 2964 14056
rect 1535 14025 1547 14028
rect 1489 14019 1547 14025
rect 1596 13861 1624 14028
rect 2958 14016 2964 14028
rect 3016 14056 3022 14068
rect 3786 14056 3792 14068
rect 3016 14028 3792 14056
rect 3016 14016 3022 14028
rect 3786 14016 3792 14028
rect 3844 14016 3850 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 5960 14028 6377 14056
rect 5960 14016 5966 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 9398 14056 9404 14068
rect 9359 14028 9404 14056
rect 6365 14019 6423 14025
rect 9398 14016 9404 14028
rect 9456 14056 9462 14068
rect 17402 14056 17408 14068
rect 9456 14028 17408 14056
rect 9456 14016 9462 14028
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 13906 13948 13912 14000
rect 13964 13988 13970 14000
rect 16669 13991 16727 13997
rect 16669 13988 16681 13991
rect 13964 13960 16681 13988
rect 13964 13948 13970 13960
rect 16669 13957 16681 13960
rect 16715 13957 16727 13991
rect 16669 13951 16727 13957
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1765 13923 1823 13929
rect 1765 13920 1777 13923
rect 1728 13892 1777 13920
rect 1728 13880 1734 13892
rect 1765 13889 1777 13892
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13920 2467 13923
rect 2774 13920 2780 13932
rect 2455 13892 2780 13920
rect 2455 13889 2467 13892
rect 2409 13883 2467 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 9674 13920 9680 13932
rect 3068 13892 9680 13920
rect 1581 13855 1639 13861
rect 1581 13821 1593 13855
rect 1627 13821 1639 13855
rect 2130 13852 2136 13864
rect 2043 13824 2136 13852
rect 1581 13815 1639 13821
rect 2130 13812 2136 13824
rect 2188 13852 2194 13864
rect 2685 13855 2743 13861
rect 2685 13852 2697 13855
rect 2188 13824 2697 13852
rect 2188 13812 2194 13824
rect 2685 13821 2697 13824
rect 2731 13852 2743 13855
rect 3068 13852 3096 13892
rect 9674 13880 9680 13892
rect 9732 13880 9738 13932
rect 9858 13920 9864 13932
rect 9819 13892 9864 13920
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 2731 13824 3096 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6181 13855 6239 13861
rect 6181 13852 6193 13855
rect 6144 13824 6193 13852
rect 6144 13812 6150 13824
rect 6181 13821 6193 13824
rect 6227 13852 6239 13855
rect 6549 13855 6607 13861
rect 6549 13852 6561 13855
rect 6227 13824 6561 13852
rect 6227 13821 6239 13824
rect 6181 13815 6239 13821
rect 6549 13821 6561 13824
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 9398 13812 9404 13864
rect 9456 13852 9462 13864
rect 9585 13855 9643 13861
rect 9585 13852 9597 13855
rect 9456 13824 9597 13852
rect 9456 13812 9462 13824
rect 9585 13821 9597 13824
rect 9631 13821 9643 13855
rect 16684 13852 16712 13951
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17862 13920 17868 13932
rect 17175 13892 17868 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16684 13824 16865 13852
rect 9585 13815 9643 13821
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 17310 13812 17316 13864
rect 17368 13852 17374 13864
rect 17405 13855 17463 13861
rect 17405 13852 17417 13855
rect 17368 13824 17417 13852
rect 17368 13812 17374 13824
rect 17405 13821 17417 13824
rect 17451 13852 17463 13855
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17451 13824 17785 13852
rect 17451 13821 17463 13824
rect 17405 13815 17463 13821
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 17773 13815 17831 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18322 13852 18328 13864
rect 18283 13824 18328 13852
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 17494 13676 17500 13728
rect 17552 13716 17558 13728
rect 17589 13719 17647 13725
rect 17589 13716 17601 13719
rect 17552 13688 17601 13716
rect 17552 13676 17558 13688
rect 17589 13685 17601 13688
rect 17635 13685 17647 13719
rect 17589 13679 17647 13685
rect 1104 13626 18860 13648
rect 1104 13574 6912 13626
rect 6964 13574 6976 13626
rect 7028 13574 7040 13626
rect 7092 13574 7104 13626
rect 7156 13574 12843 13626
rect 12895 13574 12907 13626
rect 12959 13574 12971 13626
rect 13023 13574 13035 13626
rect 13087 13574 18860 13626
rect 1104 13552 18860 13574
rect 1486 13512 1492 13524
rect 1447 13484 1492 13512
rect 1486 13472 1492 13484
rect 1544 13472 1550 13524
rect 17402 13512 17408 13524
rect 17363 13484 17408 13512
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 1504 13376 1532 13472
rect 1673 13379 1731 13385
rect 1673 13376 1685 13379
rect 1504 13348 1685 13376
rect 1673 13345 1685 13348
rect 1719 13345 1731 13379
rect 2038 13376 2044 13388
rect 1999 13348 2044 13376
rect 1673 13339 1731 13345
rect 2038 13336 2044 13348
rect 2096 13376 2102 13388
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2096 13348 2605 13376
rect 2096 13336 2102 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 17420 13376 17448 13472
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 17420 13348 17601 13376
rect 2593 13339 2651 13345
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 2314 13308 2320 13320
rect 2275 13280 2320 13308
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 17865 13311 17923 13317
rect 17865 13277 17877 13311
rect 17911 13308 17923 13311
rect 18046 13308 18052 13320
rect 17911 13280 18052 13308
rect 17911 13277 17923 13280
rect 17865 13271 17923 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 1854 13240 1860 13252
rect 1815 13212 1860 13240
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 1104 13082 18860 13104
rect 1104 13030 3947 13082
rect 3999 13030 4011 13082
rect 4063 13030 4075 13082
rect 4127 13030 4139 13082
rect 4191 13030 9878 13082
rect 9930 13030 9942 13082
rect 9994 13030 10006 13082
rect 10058 13030 10070 13082
rect 10122 13030 15808 13082
rect 15860 13030 15872 13082
rect 15924 13030 15936 13082
rect 15988 13030 16000 13082
rect 16052 13030 18860 13082
rect 1104 13008 18860 13030
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 17773 12971 17831 12977
rect 17773 12968 17785 12971
rect 9732 12940 17785 12968
rect 9732 12928 9738 12940
rect 17773 12937 17785 12940
rect 17819 12937 17831 12971
rect 17773 12931 17831 12937
rect 17788 12764 17816 12931
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17788 12736 18061 12764
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 5902 12696 5908 12708
rect 4028 12668 5908 12696
rect 4028 12656 4034 12668
rect 5902 12656 5908 12668
rect 5960 12656 5966 12708
rect 18325 12699 18383 12705
rect 18325 12665 18337 12699
rect 18371 12696 18383 12699
rect 18598 12696 18604 12708
rect 18371 12668 18604 12696
rect 18371 12665 18383 12668
rect 18325 12659 18383 12665
rect 18598 12656 18604 12668
rect 18656 12656 18662 12708
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 15746 12628 15752 12640
rect 9640 12600 15752 12628
rect 9640 12588 9646 12600
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 1104 12538 18860 12560
rect 1104 12486 6912 12538
rect 6964 12486 6976 12538
rect 7028 12486 7040 12538
rect 7092 12486 7104 12538
rect 7156 12486 12843 12538
rect 12895 12486 12907 12538
rect 12959 12486 12971 12538
rect 13023 12486 13035 12538
rect 13087 12486 18860 12538
rect 1104 12464 18860 12486
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 16942 12424 16948 12436
rect 6788 12396 16948 12424
rect 6788 12384 6794 12396
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 9214 12316 9220 12368
rect 9272 12356 9278 12368
rect 11054 12356 11060 12368
rect 9272 12328 11060 12356
rect 9272 12316 9278 12328
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3694 12288 3700 12300
rect 3108 12260 3700 12288
rect 3108 12248 3114 12260
rect 3694 12248 3700 12260
rect 3752 12248 3758 12300
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12288 10287 12291
rect 10962 12288 10968 12300
rect 10275 12260 10968 12288
rect 10275 12257 10287 12260
rect 10229 12251 10287 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 10134 12220 10140 12232
rect 3476 12192 10140 12220
rect 3476 12180 3482 12192
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10318 12220 10324 12232
rect 10279 12192 10324 12220
rect 10318 12180 10324 12192
rect 10376 12180 10382 12232
rect 10502 12220 10508 12232
rect 10463 12192 10508 12220
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 15746 12220 15752 12232
rect 10652 12192 15752 12220
rect 10652 12180 10658 12192
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 15194 12152 15200 12164
rect 3752 12124 15200 12152
rect 3752 12112 3758 12124
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 7929 12087 7987 12093
rect 7929 12084 7941 12087
rect 7800 12056 7941 12084
rect 7800 12044 7806 12056
rect 7929 12053 7941 12056
rect 7975 12053 7987 12087
rect 7929 12047 7987 12053
rect 9861 12087 9919 12093
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 12066 12084 12072 12096
rect 9907 12056 12072 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 1104 11994 18860 12016
rect 1104 11942 3947 11994
rect 3999 11942 4011 11994
rect 4063 11942 4075 11994
rect 4127 11942 4139 11994
rect 4191 11942 9878 11994
rect 9930 11942 9942 11994
rect 9994 11942 10006 11994
rect 10058 11942 10070 11994
rect 10122 11942 15808 11994
rect 15860 11942 15872 11994
rect 15924 11942 15936 11994
rect 15988 11942 16000 11994
rect 16052 11942 18860 11994
rect 1104 11920 18860 11942
rect 3786 11840 3792 11892
rect 3844 11880 3850 11892
rect 7926 11880 7932 11892
rect 3844 11852 7932 11880
rect 3844 11840 3850 11852
rect 7926 11840 7932 11852
rect 7984 11880 7990 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7984 11852 8217 11880
rect 7984 11840 7990 11852
rect 8205 11849 8217 11852
rect 8251 11880 8263 11883
rect 10318 11880 10324 11892
rect 8251 11852 10088 11880
rect 10279 11852 10324 11880
rect 8251 11849 8263 11852
rect 8205 11843 8263 11849
rect 10060 11824 10088 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 10962 11840 10968 11892
rect 11020 11880 11026 11892
rect 12069 11883 12127 11889
rect 11020 11852 11100 11880
rect 11020 11840 11026 11852
rect 10042 11772 10048 11824
rect 10100 11772 10106 11824
rect 11072 11812 11100 11852
rect 11256 11852 11744 11880
rect 11149 11815 11207 11821
rect 11149 11812 11161 11815
rect 11072 11784 11161 11812
rect 11149 11781 11161 11784
rect 11195 11781 11207 11815
rect 11149 11775 11207 11781
rect 2593 11747 2651 11753
rect 2593 11713 2605 11747
rect 2639 11744 2651 11747
rect 3602 11744 3608 11756
rect 2639 11716 3608 11744
rect 2639 11713 2651 11716
rect 2593 11707 2651 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 7558 11744 7564 11756
rect 6595 11716 7564 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 10778 11744 10784 11756
rect 7708 11716 7753 11744
rect 10739 11716 10784 11744
rect 7708 11704 7714 11716
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 10962 11744 10968 11756
rect 10875 11716 10968 11744
rect 10962 11704 10968 11716
rect 11020 11744 11026 11756
rect 11256 11744 11284 11852
rect 11716 11753 11744 11852
rect 12069 11849 12081 11883
rect 12115 11880 12127 11883
rect 12158 11880 12164 11892
rect 12115 11852 12164 11880
rect 12115 11849 12127 11852
rect 12069 11843 12127 11849
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 13964 11852 14289 11880
rect 13964 11840 13970 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 11020 11716 11284 11744
rect 11701 11747 11759 11753
rect 11020 11704 11026 11716
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11676 6331 11679
rect 8110 11676 8116 11688
rect 6319 11648 8116 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 8386 11636 8392 11688
rect 8444 11676 8450 11688
rect 8656 11679 8714 11685
rect 8444 11648 8489 11676
rect 8444 11636 8450 11648
rect 8656 11645 8668 11679
rect 8702 11676 8714 11679
rect 10502 11676 10508 11688
rect 8702 11648 10508 11676
rect 8702 11645 8714 11648
rect 8656 11639 8714 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 11606 11676 11612 11688
rect 10560 11648 11612 11676
rect 10560 11636 10566 11648
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 14292 11676 14320 11843
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18138 11880 18144 11892
rect 18012 11852 18144 11880
rect 18012 11840 18018 11852
rect 18138 11840 18144 11852
rect 18196 11840 18202 11892
rect 18414 11880 18420 11892
rect 18375 11852 18420 11880
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 16298 11812 16304 11824
rect 14516 11784 16304 11812
rect 14516 11772 14522 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 14366 11704 14372 11756
rect 14424 11744 14430 11756
rect 14829 11747 14887 11753
rect 14829 11744 14841 11747
rect 14424 11716 14841 11744
rect 14424 11704 14430 11716
rect 14829 11713 14841 11716
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 18230 11744 18236 11756
rect 17727 11716 18236 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 18230 11704 18236 11716
rect 18288 11704 18294 11756
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 14292 11648 14473 11676
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 14918 11636 14924 11688
rect 14976 11676 14982 11688
rect 14976 11648 17724 11676
rect 14976 11636 14982 11648
rect 7282 11608 7288 11620
rect 5920 11580 7288 11608
rect 1946 11540 1952 11552
rect 1907 11512 1952 11540
rect 1946 11500 1952 11512
rect 2004 11500 2010 11552
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 2096 11512 2329 11540
rect 2096 11500 2102 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2317 11503 2375 11509
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 5920 11549 5948 11580
rect 7282 11568 7288 11580
rect 7340 11568 7346 11620
rect 7469 11611 7527 11617
rect 7469 11577 7481 11611
rect 7515 11608 7527 11611
rect 7929 11611 7987 11617
rect 7929 11608 7941 11611
rect 7515 11580 7941 11608
rect 7515 11577 7527 11580
rect 7469 11571 7527 11577
rect 7929 11577 7941 11580
rect 7975 11577 7987 11611
rect 10042 11608 10048 11620
rect 7929 11571 7987 11577
rect 9048 11580 10048 11608
rect 5905 11543 5963 11549
rect 2464 11512 2509 11540
rect 2464 11500 2470 11512
rect 5905 11509 5917 11543
rect 5951 11509 5963 11543
rect 5905 11503 5963 11509
rect 6362 11500 6368 11552
rect 6420 11540 6426 11552
rect 6420 11512 6465 11540
rect 6420 11500 6426 11512
rect 6730 11500 6736 11552
rect 6788 11540 6794 11552
rect 6825 11543 6883 11549
rect 6825 11540 6837 11543
rect 6788 11512 6837 11540
rect 6788 11500 6794 11512
rect 6825 11509 6837 11512
rect 6871 11509 6883 11543
rect 6825 11503 6883 11509
rect 7101 11543 7159 11549
rect 7101 11509 7113 11543
rect 7147 11540 7159 11543
rect 7374 11540 7380 11552
rect 7147 11512 7380 11540
rect 7147 11509 7159 11512
rect 7101 11503 7159 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 7561 11543 7619 11549
rect 7561 11509 7573 11543
rect 7607 11540 7619 11543
rect 7742 11540 7748 11552
rect 7607 11512 7748 11540
rect 7607 11509 7619 11512
rect 7561 11503 7619 11509
rect 7742 11500 7748 11512
rect 7800 11540 7806 11552
rect 9048 11540 9076 11580
rect 10042 11568 10048 11580
rect 10100 11568 10106 11620
rect 10134 11568 10140 11620
rect 10192 11608 10198 11620
rect 10689 11611 10747 11617
rect 10689 11608 10701 11611
rect 10192 11580 10701 11608
rect 10192 11568 10198 11580
rect 10689 11577 10701 11580
rect 10735 11608 10747 11611
rect 15194 11608 15200 11620
rect 10735 11580 15200 11608
rect 10735 11577 10747 11580
rect 10689 11571 10747 11577
rect 15194 11568 15200 11580
rect 15252 11568 15258 11620
rect 17696 11552 17724 11648
rect 9766 11540 9772 11552
rect 7800 11512 9076 11540
rect 9727 11512 9772 11540
rect 7800 11500 7806 11512
rect 9766 11500 9772 11512
rect 9824 11500 9830 11552
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 11238 11540 11244 11552
rect 10284 11512 11244 11540
rect 10284 11500 10290 11512
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11330 11500 11336 11552
rect 11388 11540 11394 11552
rect 11517 11543 11575 11549
rect 11517 11540 11529 11543
rect 11388 11512 11529 11540
rect 11388 11500 11394 11512
rect 11517 11509 11529 11512
rect 11563 11509 11575 11543
rect 11517 11503 11575 11509
rect 11609 11543 11667 11549
rect 11609 11509 11621 11543
rect 11655 11540 11667 11543
rect 11698 11540 11704 11552
rect 11655 11512 11704 11540
rect 11655 11509 11667 11512
rect 11609 11503 11667 11509
rect 11698 11500 11704 11512
rect 11756 11540 11762 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 11756 11512 12265 11540
rect 11756 11500 11762 11512
rect 12253 11509 12265 11512
rect 12299 11540 12311 11543
rect 15746 11540 15752 11552
rect 12299 11512 15752 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 17678 11500 17684 11552
rect 17736 11540 17742 11552
rect 17773 11543 17831 11549
rect 17773 11540 17785 11543
rect 17736 11512 17785 11540
rect 17736 11500 17742 11512
rect 17773 11509 17785 11512
rect 17819 11509 17831 11543
rect 17773 11503 17831 11509
rect 1104 11450 18860 11472
rect 1104 11398 6912 11450
rect 6964 11398 6976 11450
rect 7028 11398 7040 11450
rect 7092 11398 7104 11450
rect 7156 11398 12843 11450
rect 12895 11398 12907 11450
rect 12959 11398 12971 11450
rect 13023 11398 13035 11450
rect 13087 11398 18860 11450
rect 1104 11376 18860 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 2280 11308 4200 11336
rect 2280 11296 2286 11308
rect 2498 11277 2504 11280
rect 2492 11268 2504 11277
rect 2459 11240 2504 11268
rect 2492 11231 2504 11240
rect 2498 11228 2504 11231
rect 2556 11228 2562 11280
rect 3694 11268 3700 11280
rect 3655 11240 3700 11268
rect 3694 11228 3700 11240
rect 3752 11228 3758 11280
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 4172 11200 4200 11308
rect 6270 11296 6276 11348
rect 6328 11336 6334 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6328 11308 6745 11336
rect 6328 11296 6334 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7561 11339 7619 11345
rect 7561 11305 7573 11339
rect 7607 11336 7619 11339
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 7607 11308 8861 11336
rect 7607 11305 7619 11308
rect 7561 11299 7619 11305
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9953 11339 10011 11345
rect 9953 11305 9965 11339
rect 9999 11336 10011 11339
rect 11330 11336 11336 11348
rect 9999 11308 11336 11336
rect 9999 11305 10011 11308
rect 9953 11299 10011 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11698 11336 11704 11348
rect 11659 11308 11704 11336
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12066 11336 12072 11348
rect 12027 11308 12072 11336
rect 12066 11296 12072 11308
rect 12124 11296 12130 11348
rect 12158 11296 12164 11348
rect 12216 11336 12222 11348
rect 15562 11336 15568 11348
rect 12216 11308 15568 11336
rect 12216 11296 12222 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 17957 11339 18015 11345
rect 17957 11336 17969 11339
rect 15804 11308 17969 11336
rect 15804 11296 15810 11308
rect 17957 11305 17969 11308
rect 18003 11336 18015 11339
rect 18414 11336 18420 11348
rect 18003 11308 18420 11336
rect 18003 11305 18015 11308
rect 17957 11299 18015 11305
rect 18414 11296 18420 11308
rect 18472 11296 18478 11348
rect 5528 11271 5586 11277
rect 5528 11237 5540 11271
rect 5574 11268 5586 11271
rect 5574 11240 7328 11268
rect 5574 11237 5586 11240
rect 5528 11231 5586 11237
rect 6730 11200 6736 11212
rect 2271 11172 3832 11200
rect 4172 11172 6736 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 3804 11144 3832 11172
rect 6730 11160 6736 11172
rect 6788 11200 6794 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 6788 11172 7113 11200
rect 6788 11160 6794 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 7101 11163 7159 11169
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 3844 11104 5273 11132
rect 3844 11092 3850 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7300 11141 7328 11240
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 8757 11271 8815 11277
rect 8757 11268 8769 11271
rect 7432 11240 8769 11268
rect 7432 11228 7438 11240
rect 8757 11237 8769 11240
rect 8803 11237 8815 11271
rect 8757 11231 8815 11237
rect 10496 11271 10554 11277
rect 10496 11237 10508 11271
rect 10542 11268 10554 11271
rect 10962 11268 10968 11280
rect 10542 11240 10968 11268
rect 10542 11237 10554 11240
rect 10496 11231 10554 11237
rect 10962 11228 10968 11240
rect 11020 11228 11026 11280
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 11848 11240 13124 11268
rect 11848 11228 11854 11240
rect 7926 11200 7932 11212
rect 7887 11172 7932 11200
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 9214 11200 9220 11212
rect 8076 11172 9220 11200
rect 8076 11160 8082 11172
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 12897 11203 12955 11209
rect 12897 11200 12909 11203
rect 11480 11172 12909 11200
rect 11480 11160 11486 11172
rect 12897 11169 12909 11172
rect 12943 11169 12955 11203
rect 12897 11163 12955 11169
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 6880 11104 7205 11132
rect 6880 11092 6886 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7193 11095 7251 11101
rect 7285 11135 7343 11141
rect 7285 11101 7297 11135
rect 7331 11132 7343 11135
rect 7650 11132 7656 11144
rect 7331 11104 7656 11132
rect 7331 11101 7343 11104
rect 7285 11095 7343 11101
rect 7650 11092 7656 11104
rect 7708 11132 7714 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7708 11104 8125 11132
rect 7708 11092 7714 11104
rect 8113 11101 8125 11104
rect 8159 11132 8171 11135
rect 8202 11132 8208 11144
rect 8159 11104 8208 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8938 11132 8944 11144
rect 8899 11104 8944 11132
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 10226 11132 10232 11144
rect 10187 11104 10232 11132
rect 10226 11092 10232 11104
rect 10284 11092 10290 11144
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 12158 11132 12164 11144
rect 12119 11104 12164 11132
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 3510 11024 3516 11076
rect 3568 11064 3574 11076
rect 4798 11064 4804 11076
rect 3568 11036 4804 11064
rect 3568 11024 3574 11036
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 6641 11067 6699 11073
rect 6641 11033 6653 11067
rect 6687 11064 6699 11067
rect 7098 11064 7104 11076
rect 6687 11036 7104 11064
rect 6687 11033 6699 11036
rect 6641 11027 6699 11033
rect 7098 11024 7104 11036
rect 7156 11064 7162 11076
rect 8294 11064 8300 11076
rect 7156 11036 8300 11064
rect 7156 11024 7162 11036
rect 8294 11024 8300 11036
rect 8352 11024 8358 11076
rect 1670 10996 1676 11008
rect 1631 10968 1676 10996
rect 1670 10956 1676 10968
rect 1728 10956 1734 11008
rect 1854 10996 1860 11008
rect 1815 10968 1860 10996
rect 1854 10956 1860 10968
rect 1912 10956 1918 11008
rect 2130 10996 2136 11008
rect 2091 10968 2136 10996
rect 2130 10956 2136 10968
rect 2188 10956 2194 11008
rect 3602 10996 3608 11008
rect 3563 10968 3608 10996
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 4246 10996 4252 11008
rect 4207 10968 4252 10996
rect 4246 10956 4252 10968
rect 4304 10956 4310 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8389 10999 8447 11005
rect 8389 10996 8401 10999
rect 8168 10968 8401 10996
rect 8168 10956 8174 10968
rect 8389 10965 8401 10968
rect 8435 10965 8447 10999
rect 8389 10959 8447 10965
rect 8570 10956 8576 11008
rect 8628 10996 8634 11008
rect 11514 10996 11520 11008
rect 8628 10968 11520 10996
rect 8628 10956 8634 10968
rect 11514 10956 11520 10968
rect 11572 10956 11578 11008
rect 11624 11005 11652 11092
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12268 11064 12296 11095
rect 12342 11092 12348 11144
rect 12400 11132 12406 11144
rect 13096 11141 13124 11240
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13725 11271 13783 11277
rect 13725 11268 13737 11271
rect 13228 11240 13737 11268
rect 13228 11228 13234 11240
rect 13725 11237 13737 11240
rect 13771 11268 13783 11271
rect 14458 11268 14464 11280
rect 13771 11240 14464 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 14458 11228 14464 11240
rect 14516 11228 14522 11280
rect 16206 11268 16212 11280
rect 14568 11240 16212 11268
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12400 11104 13001 11132
rect 12400 11092 12406 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 13081 11095 13139 11101
rect 12124 11036 12296 11064
rect 12529 11067 12587 11073
rect 12124 11024 12130 11036
rect 12529 11033 12541 11067
rect 12575 11064 12587 11067
rect 12710 11064 12716 11076
rect 12575 11036 12716 11064
rect 12575 11033 12587 11036
rect 12529 11027 12587 11033
rect 12710 11024 12716 11036
rect 12768 11024 12774 11076
rect 14182 11024 14188 11076
rect 14240 11064 14246 11076
rect 14568 11073 14596 11240
rect 16206 11228 16212 11240
rect 16264 11228 16270 11280
rect 16942 11268 16948 11280
rect 16903 11240 16948 11268
rect 16942 11228 16948 11240
rect 17000 11228 17006 11280
rect 17218 11268 17224 11280
rect 17179 11240 17224 11268
rect 17218 11228 17224 11240
rect 17276 11228 17282 11280
rect 18138 11268 18144 11280
rect 17328 11240 18144 11268
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 14918 11200 14924 11212
rect 14875 11172 14924 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 14844 11132 14872 11163
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15545 11203 15603 11209
rect 15545 11200 15557 11203
rect 15436 11172 15557 11200
rect 15436 11160 15442 11172
rect 15545 11169 15557 11172
rect 15591 11169 15603 11203
rect 17328 11200 17356 11240
rect 18138 11228 18144 11240
rect 18196 11268 18202 11280
rect 18325 11271 18383 11277
rect 18325 11268 18337 11271
rect 18196 11240 18337 11268
rect 18196 11228 18202 11240
rect 18325 11237 18337 11240
rect 18371 11237 18383 11271
rect 18325 11231 18383 11237
rect 17862 11200 17868 11212
rect 15545 11163 15603 11169
rect 16500 11172 17356 11200
rect 17823 11172 17868 11200
rect 14660 11104 14872 11132
rect 14553 11067 14611 11073
rect 14553 11064 14565 11067
rect 14240 11036 14565 11064
rect 14240 11024 14246 11036
rect 14553 11033 14565 11036
rect 14599 11033 14611 11067
rect 14553 11027 14611 11033
rect 11609 10999 11667 11005
rect 11609 10965 11621 10999
rect 11655 10965 11667 10999
rect 11609 10959 11667 10965
rect 14458 10956 14464 11008
rect 14516 10996 14522 11008
rect 14660 10996 14688 11104
rect 15102 11092 15108 11144
rect 15160 11132 15166 11144
rect 15289 11135 15347 11141
rect 15289 11132 15301 11135
rect 15160 11104 15301 11132
rect 15160 11092 15166 11104
rect 15289 11101 15301 11104
rect 15335 11101 15347 11135
rect 15289 11095 15347 11101
rect 14826 11024 14832 11076
rect 14884 11064 14890 11076
rect 15010 11064 15016 11076
rect 14884 11036 15016 11064
rect 14884 11024 14890 11036
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 14516 10968 14688 10996
rect 14516 10956 14522 10968
rect 14918 10956 14924 11008
rect 14976 10996 14982 11008
rect 16500 10996 16528 11172
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 18049 11135 18107 11141
rect 16684 11104 17908 11132
rect 14976 10968 16528 10996
rect 14976 10956 14982 10968
rect 16574 10956 16580 11008
rect 16632 10996 16638 11008
rect 16684 11005 16712 11104
rect 16850 11024 16856 11076
rect 16908 11064 16914 11076
rect 17313 11067 17371 11073
rect 17313 11064 17325 11067
rect 16908 11036 17325 11064
rect 16908 11024 16914 11036
rect 17313 11033 17325 11036
rect 17359 11033 17371 11067
rect 17494 11064 17500 11076
rect 17455 11036 17500 11064
rect 17313 11027 17371 11033
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 17880 11064 17908 11104
rect 18049 11101 18061 11135
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18064 11064 18092 11095
rect 17880 11036 18092 11064
rect 16669 10999 16727 11005
rect 16669 10996 16681 10999
rect 16632 10968 16681 10996
rect 16632 10956 16638 10968
rect 16669 10965 16681 10968
rect 16715 10965 16727 10999
rect 16669 10959 16727 10965
rect 16761 10999 16819 11005
rect 16761 10965 16773 10999
rect 16807 10996 16819 10999
rect 17126 10996 17132 11008
rect 16807 10968 17132 10996
rect 16807 10965 16819 10968
rect 16761 10959 16819 10965
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 1104 10906 18860 10928
rect 1104 10854 3947 10906
rect 3999 10854 4011 10906
rect 4063 10854 4075 10906
rect 4127 10854 4139 10906
rect 4191 10854 9878 10906
rect 9930 10854 9942 10906
rect 9994 10854 10006 10906
rect 10058 10854 10070 10906
rect 10122 10854 15808 10906
rect 15860 10854 15872 10906
rect 15924 10854 15936 10906
rect 15988 10854 16000 10906
rect 16052 10854 18860 10906
rect 1104 10832 18860 10854
rect 1397 10795 1455 10801
rect 1397 10761 1409 10795
rect 1443 10792 1455 10795
rect 2038 10792 2044 10804
rect 1443 10764 2044 10792
rect 1443 10761 1455 10764
rect 1397 10755 1455 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2225 10795 2283 10801
rect 2225 10761 2237 10795
rect 2271 10792 2283 10795
rect 2406 10792 2412 10804
rect 2271 10764 2412 10792
rect 2271 10761 2283 10764
rect 2225 10755 2283 10761
rect 2406 10752 2412 10764
rect 2464 10752 2470 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 4890 10792 4896 10804
rect 3099 10764 4896 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6362 10792 6368 10804
rect 5951 10764 6368 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7616 10764 8217 10792
rect 7616 10752 7622 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 11149 10795 11207 10801
rect 8536 10764 10272 10792
rect 8536 10752 8542 10764
rect 6822 10724 6828 10736
rect 5460 10696 6828 10724
rect 1854 10656 1860 10668
rect 1815 10628 1860 10656
rect 1854 10616 1860 10628
rect 1912 10616 1918 10668
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2498 10656 2504 10668
rect 2087 10628 2504 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2498 10616 2504 10628
rect 2556 10656 2562 10668
rect 2777 10659 2835 10665
rect 2777 10656 2789 10659
rect 2556 10628 2789 10656
rect 2556 10616 2562 10628
rect 2777 10625 2789 10628
rect 2823 10656 2835 10659
rect 2958 10656 2964 10668
rect 2823 10628 2964 10656
rect 2823 10625 2835 10628
rect 2777 10619 2835 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3697 10659 3755 10665
rect 3697 10656 3709 10659
rect 3660 10628 3709 10656
rect 3660 10616 3666 10628
rect 3697 10625 3709 10628
rect 3743 10625 3755 10659
rect 3697 10619 3755 10625
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3844 10628 3985 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 1872 10520 1900 10616
rect 2130 10548 2136 10600
rect 2188 10588 2194 10600
rect 2593 10591 2651 10597
rect 2593 10588 2605 10591
rect 2188 10560 2605 10588
rect 2188 10548 2194 10560
rect 2593 10557 2605 10560
rect 2639 10588 2651 10591
rect 4522 10588 4528 10600
rect 2639 10560 4528 10588
rect 2639 10557 2651 10560
rect 2593 10551 2651 10557
rect 4522 10548 4528 10560
rect 4580 10548 4586 10600
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 5460 10597 5488 10696
rect 6822 10684 6828 10696
rect 6880 10684 6886 10736
rect 10137 10727 10195 10733
rect 10137 10693 10149 10727
rect 10183 10693 10195 10727
rect 10244 10724 10272 10764
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 12158 10792 12164 10804
rect 11195 10764 12164 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 14918 10792 14924 10804
rect 12492 10764 14924 10792
rect 12492 10752 12498 10764
rect 14918 10752 14924 10764
rect 14976 10752 14982 10804
rect 17218 10792 17224 10804
rect 16040 10764 17224 10792
rect 12250 10724 12256 10736
rect 10244 10696 12256 10724
rect 10137 10687 10195 10693
rect 6362 10656 6368 10668
rect 6323 10628 6368 10656
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 10152 10656 10180 10687
rect 12250 10684 12256 10696
rect 12308 10684 12314 10736
rect 13817 10727 13875 10733
rect 13817 10693 13829 10727
rect 13863 10693 13875 10727
rect 13817 10687 13875 10693
rect 10502 10656 10508 10668
rect 6595 10628 6960 10656
rect 10152 10628 10508 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 5445 10591 5503 10597
rect 5445 10588 5457 10591
rect 4764 10560 5457 10588
rect 4764 10548 4770 10560
rect 5445 10557 5457 10560
rect 5491 10557 5503 10591
rect 6270 10588 6276 10600
rect 6231 10560 6276 10588
rect 5445 10551 5503 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6932 10588 6960 10628
rect 10502 10616 10508 10628
rect 10560 10656 10566 10668
rect 10962 10656 10968 10668
rect 10560 10628 10968 10656
rect 10560 10616 10566 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 11606 10616 11612 10668
rect 11664 10656 11670 10668
rect 11701 10659 11759 10665
rect 11701 10656 11713 10659
rect 11664 10628 11713 10656
rect 11664 10616 11670 10628
rect 11701 10625 11713 10628
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 7098 10597 7104 10600
rect 7092 10588 7104 10597
rect 6932 10560 7104 10588
rect 6825 10551 6883 10557
rect 7092 10551 7104 10560
rect 3053 10523 3111 10529
rect 3053 10520 3065 10523
rect 1872 10492 3065 10520
rect 3053 10489 3065 10492
rect 3099 10489 3111 10523
rect 3053 10483 3111 10489
rect 3234 10480 3240 10532
rect 3292 10520 3298 10532
rect 3605 10523 3663 10529
rect 3605 10520 3617 10523
rect 3292 10492 3617 10520
rect 3292 10480 3298 10492
rect 3605 10489 3617 10492
rect 3651 10489 3663 10523
rect 3605 10483 3663 10489
rect 4240 10523 4298 10529
rect 4240 10489 4252 10523
rect 4286 10520 4298 10523
rect 5074 10520 5080 10532
rect 4286 10492 5080 10520
rect 4286 10489 4298 10492
rect 4240 10483 4298 10489
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 6546 10480 6552 10532
rect 6604 10520 6610 10532
rect 6840 10520 6868 10551
rect 7098 10548 7104 10551
rect 7156 10548 7162 10600
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8757 10591 8815 10597
rect 8757 10588 8769 10591
rect 8352 10560 8769 10588
rect 8352 10548 8358 10560
rect 8757 10557 8769 10560
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 9916 10560 11529 10588
rect 9916 10548 9922 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 11517 10551 11575 10557
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 11940 10560 12449 10588
rect 11940 10548 11946 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 6604 10492 6868 10520
rect 6604 10480 6610 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 6972 10492 8401 10520
rect 6972 10480 6978 10492
rect 8389 10489 8401 10492
rect 8435 10520 8447 10523
rect 8846 10520 8852 10532
rect 8435 10492 8852 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 8846 10480 8852 10492
rect 8904 10480 8910 10532
rect 9024 10523 9082 10529
rect 9024 10489 9036 10523
rect 9070 10520 9082 10523
rect 9674 10520 9680 10532
rect 9070 10492 9680 10520
rect 9070 10489 9082 10492
rect 9024 10483 9082 10489
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 11609 10523 11667 10529
rect 11609 10520 11621 10523
rect 10336 10492 11621 10520
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 2590 10412 2596 10464
rect 2648 10452 2654 10464
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 2648 10424 2697 10452
rect 2648 10412 2654 10424
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 2685 10415 2743 10421
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 2832 10424 3157 10452
rect 2832 10412 2838 10424
rect 3145 10421 3157 10424
rect 3191 10421 3203 10455
rect 3145 10415 3203 10421
rect 3513 10455 3571 10461
rect 3513 10421 3525 10455
rect 3559 10452 3571 10455
rect 4614 10452 4620 10464
rect 3559 10424 4620 10452
rect 3559 10421 3571 10424
rect 3513 10415 3571 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 5350 10452 5356 10464
rect 5311 10424 5356 10452
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 10336 10461 10364 10492
rect 11609 10489 11621 10492
rect 11655 10489 11667 10523
rect 12250 10520 12256 10532
rect 12211 10492 12256 10520
rect 11609 10483 11667 10489
rect 12250 10480 12256 10492
rect 12308 10480 12314 10532
rect 12704 10523 12762 10529
rect 12704 10489 12716 10523
rect 12750 10520 12762 10523
rect 13262 10520 13268 10532
rect 12750 10492 13268 10520
rect 12750 10489 12762 10492
rect 12704 10483 12762 10489
rect 13262 10480 13268 10492
rect 13320 10480 13326 10532
rect 13832 10520 13860 10687
rect 16040 10668 16068 10764
rect 17218 10752 17224 10764
rect 17276 10752 17282 10804
rect 16022 10656 16028 10668
rect 15935 10628 16028 10656
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 17681 10659 17739 10665
rect 17681 10625 17693 10659
rect 17727 10656 17739 10659
rect 17862 10656 17868 10668
rect 17727 10628 17868 10656
rect 17727 10625 17739 10628
rect 17681 10619 17739 10625
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10588 13967 10591
rect 15102 10588 15108 10600
rect 13955 10560 15108 10588
rect 13955 10557 13967 10560
rect 13909 10551 13967 10557
rect 15102 10548 15108 10560
rect 15160 10588 15166 10600
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15160 10560 16221 10588
rect 15160 10548 15166 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 18049 10591 18107 10597
rect 16209 10551 16267 10557
rect 16408 10560 16712 10588
rect 14176 10523 14234 10529
rect 14176 10520 14188 10523
rect 13832 10492 14188 10520
rect 14176 10489 14188 10492
rect 14222 10520 14234 10523
rect 14734 10520 14740 10532
rect 14222 10492 14740 10520
rect 14222 10489 14234 10492
rect 14176 10483 14234 10489
rect 14734 10480 14740 10492
rect 14792 10480 14798 10532
rect 15749 10523 15807 10529
rect 15749 10489 15761 10523
rect 15795 10520 15807 10523
rect 16408 10520 16436 10560
rect 16684 10532 16712 10560
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 15795 10492 16436 10520
rect 16476 10523 16534 10529
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 16476 10489 16488 10523
rect 16522 10520 16534 10523
rect 16574 10520 16580 10532
rect 16522 10492 16580 10520
rect 16522 10489 16534 10492
rect 16476 10483 16534 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 16666 10480 16672 10532
rect 16724 10480 16730 10532
rect 10321 10455 10379 10461
rect 10321 10421 10333 10455
rect 10367 10421 10379 10455
rect 10686 10452 10692 10464
rect 10647 10424 10692 10452
rect 10321 10415 10379 10421
rect 10686 10412 10692 10424
rect 10744 10412 10750 10464
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 10836 10424 10881 10452
rect 10836 10412 10842 10424
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11977 10455 12035 10461
rect 11977 10452 11989 10455
rect 11572 10424 11989 10452
rect 11572 10412 11578 10424
rect 11977 10421 11989 10424
rect 12023 10452 12035 10455
rect 12066 10452 12072 10464
rect 12023 10424 12072 10452
rect 12023 10421 12035 10424
rect 11977 10415 12035 10421
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 15286 10452 15292 10464
rect 15247 10424 15292 10452
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15378 10412 15384 10464
rect 15436 10452 15442 10464
rect 15841 10455 15899 10461
rect 15436 10424 15481 10452
rect 15436 10412 15442 10424
rect 15841 10421 15853 10455
rect 15887 10452 15899 10455
rect 16758 10452 16764 10464
rect 15887 10424 16764 10452
rect 15887 10421 15899 10424
rect 15841 10415 15899 10421
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 17218 10412 17224 10464
rect 17276 10452 17282 10464
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 17276 10424 17601 10452
rect 17276 10412 17282 10424
rect 17589 10421 17601 10424
rect 17635 10421 17647 10455
rect 17589 10415 17647 10421
rect 17862 10412 17868 10464
rect 17920 10452 17926 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 17920 10424 18245 10452
rect 17920 10412 17926 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18414 10452 18420 10464
rect 18375 10424 18420 10452
rect 18233 10415 18291 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 1104 10362 18860 10384
rect 1104 10310 6912 10362
rect 6964 10310 6976 10362
rect 7028 10310 7040 10362
rect 7092 10310 7104 10362
rect 7156 10310 12843 10362
rect 12895 10310 12907 10362
rect 12959 10310 12971 10362
rect 13023 10310 13035 10362
rect 13087 10310 18860 10362
rect 1104 10288 18860 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 2869 10251 2927 10257
rect 2869 10248 2881 10251
rect 1820 10220 2881 10248
rect 1820 10208 1826 10220
rect 2869 10217 2881 10220
rect 2915 10217 2927 10251
rect 2869 10211 2927 10217
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3234 10248 3240 10260
rect 3191 10220 3240 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3234 10208 3240 10220
rect 3292 10208 3298 10260
rect 3513 10251 3571 10257
rect 3513 10217 3525 10251
rect 3559 10248 3571 10251
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 3559 10220 4353 10248
rect 3559 10217 3571 10220
rect 3513 10211 3571 10217
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 4706 10248 4712 10260
rect 4667 10220 4712 10248
rect 4341 10211 4399 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 5169 10251 5227 10257
rect 5169 10217 5181 10251
rect 5215 10217 5227 10251
rect 5169 10211 5227 10217
rect 2038 10140 2044 10192
rect 2096 10180 2102 10192
rect 2590 10180 2596 10192
rect 2096 10152 2596 10180
rect 2096 10140 2102 10152
rect 2590 10140 2596 10152
rect 2648 10180 2654 10192
rect 3694 10180 3700 10192
rect 2648 10152 3700 10180
rect 2648 10140 2654 10152
rect 3694 10140 3700 10152
rect 3752 10140 3758 10192
rect 4246 10140 4252 10192
rect 4304 10180 4310 10192
rect 4801 10183 4859 10189
rect 4801 10180 4813 10183
rect 4304 10152 4813 10180
rect 4304 10140 4310 10152
rect 1664 10115 1722 10121
rect 1664 10081 1676 10115
rect 1710 10112 1722 10115
rect 3510 10112 3516 10124
rect 1710 10084 3516 10112
rect 1710 10081 1722 10084
rect 1664 10075 1722 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 3605 10115 3663 10121
rect 3605 10081 3617 10115
rect 3651 10112 3663 10115
rect 4338 10112 4344 10124
rect 3651 10084 4344 10112
rect 3651 10081 3663 10084
rect 3605 10075 3663 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10004 1458 10056
rect 2958 10004 2964 10056
rect 3016 10044 3022 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3016 10016 3801 10044
rect 3016 10004 3022 10016
rect 3789 10013 3801 10016
rect 3835 10044 3847 10047
rect 4430 10044 4436 10056
rect 3835 10016 4436 10044
rect 3835 10013 3847 10016
rect 3789 10007 3847 10013
rect 4430 10004 4436 10016
rect 4488 10004 4494 10056
rect 4540 10044 4568 10152
rect 4801 10149 4813 10152
rect 4847 10149 4859 10183
rect 4801 10143 4859 10149
rect 4614 10072 4620 10124
rect 4672 10112 4678 10124
rect 5184 10112 5212 10211
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 9858 10248 9864 10260
rect 5592 10220 9720 10248
rect 9819 10220 9864 10248
rect 5592 10208 5598 10220
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 6089 10183 6147 10189
rect 6089 10180 6101 10183
rect 5500 10152 6101 10180
rect 5500 10140 5506 10152
rect 6089 10149 6101 10152
rect 6135 10180 6147 10183
rect 6641 10183 6699 10189
rect 6641 10180 6653 10183
rect 6135 10152 6653 10180
rect 6135 10149 6147 10152
rect 6089 10143 6147 10149
rect 6641 10149 6653 10152
rect 6687 10180 6699 10183
rect 6822 10180 6828 10192
rect 6687 10152 6828 10180
rect 6687 10149 6699 10152
rect 6641 10143 6699 10149
rect 6822 10140 6828 10152
rect 6880 10140 6886 10192
rect 7558 10140 7564 10192
rect 7616 10180 7622 10192
rect 7806 10183 7864 10189
rect 7806 10180 7818 10183
rect 7616 10152 7818 10180
rect 7616 10140 7622 10152
rect 7806 10149 7818 10152
rect 7852 10149 7864 10183
rect 7806 10143 7864 10149
rect 8846 10140 8852 10192
rect 8904 10180 8910 10192
rect 9217 10183 9275 10189
rect 9217 10180 9229 10183
rect 8904 10152 9229 10180
rect 8904 10140 8910 10152
rect 9217 10149 9229 10152
rect 9263 10180 9275 10183
rect 9263 10152 9628 10180
rect 9263 10149 9275 10152
rect 9217 10143 9275 10149
rect 5534 10112 5540 10124
rect 4672 10084 5212 10112
rect 5495 10084 5540 10112
rect 4672 10072 4678 10084
rect 5534 10072 5540 10084
rect 5592 10072 5598 10124
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6328 10084 6561 10112
rect 6328 10072 6334 10084
rect 6549 10081 6561 10084
rect 6595 10112 6607 10115
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6595 10084 7021 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 7009 10081 7021 10084
rect 7055 10112 7067 10115
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 7055 10084 7205 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7193 10081 7205 10084
rect 7239 10081 7251 10115
rect 7466 10112 7472 10124
rect 7427 10084 7472 10112
rect 7193 10075 7251 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7650 10072 7656 10124
rect 7708 10112 7714 10124
rect 9490 10112 9496 10124
rect 7708 10084 9496 10112
rect 7708 10072 7714 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 4706 10044 4712 10056
rect 4540 10016 4712 10044
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4985 10047 5043 10053
rect 4985 10013 4997 10047
rect 5031 10044 5043 10047
rect 5074 10044 5080 10056
rect 5031 10016 5080 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 5074 10004 5080 10016
rect 5132 10004 5138 10056
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5316 10016 5641 10044
rect 5316 10004 5322 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3234 9976 3240 9988
rect 2740 9948 3240 9976
rect 2740 9936 2746 9948
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5736 9976 5764 10007
rect 6638 10004 6644 10056
rect 6696 10044 6702 10056
rect 6733 10047 6791 10053
rect 6733 10044 6745 10047
rect 6696 10016 6745 10044
rect 6696 10004 6702 10016
rect 6733 10013 6745 10016
rect 6779 10013 6791 10047
rect 6733 10007 6791 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10013 7619 10047
rect 9306 10044 9312 10056
rect 7561 10007 7619 10013
rect 8864 10016 9312 10044
rect 5408 9948 5764 9976
rect 5408 9936 5414 9948
rect 6546 9936 6552 9988
rect 6604 9976 6610 9988
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 6604 9948 7297 9976
rect 6604 9936 6610 9948
rect 7285 9945 7297 9948
rect 7331 9976 7343 9979
rect 7576 9976 7604 10007
rect 7331 9948 7604 9976
rect 7331 9945 7343 9948
rect 7285 9939 7343 9945
rect 2777 9911 2835 9917
rect 2777 9877 2789 9911
rect 2823 9908 2835 9911
rect 2958 9908 2964 9920
rect 2823 9880 2964 9908
rect 2823 9877 2835 9880
rect 2777 9871 2835 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 3418 9868 3424 9920
rect 3476 9908 3482 9920
rect 4157 9911 4215 9917
rect 4157 9908 4169 9911
rect 3476 9880 4169 9908
rect 3476 9868 3482 9880
rect 4157 9877 4169 9880
rect 4203 9908 4215 9911
rect 5534 9908 5540 9920
rect 4203 9880 5540 9908
rect 4203 9877 4215 9880
rect 4157 9871 4215 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 6181 9911 6239 9917
rect 6181 9877 6193 9911
rect 6227 9908 6239 9911
rect 6730 9908 6736 9920
rect 6227 9880 6736 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 7193 9911 7251 9917
rect 7193 9877 7205 9911
rect 7239 9908 7251 9911
rect 8864 9908 8892 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9600 10044 9628 10152
rect 9692 10121 9720 10220
rect 9858 10208 9864 10220
rect 9916 10208 9922 10260
rect 10686 10248 10692 10260
rect 10647 10220 10692 10248
rect 10686 10208 10692 10220
rect 10744 10208 10750 10260
rect 11054 10248 11060 10260
rect 11015 10220 11060 10248
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 13357 10251 13415 10257
rect 13357 10217 13369 10251
rect 13403 10248 13415 10251
rect 14553 10251 14611 10257
rect 14553 10248 14565 10251
rect 13403 10220 14565 10248
rect 13403 10217 13415 10220
rect 13357 10211 13415 10217
rect 14553 10217 14565 10220
rect 14599 10217 14611 10251
rect 14553 10211 14611 10217
rect 16206 10208 16212 10260
rect 16264 10248 16270 10260
rect 16482 10248 16488 10260
rect 16264 10220 16488 10248
rect 16264 10208 16270 10220
rect 16482 10208 16488 10220
rect 16540 10208 16546 10260
rect 16758 10248 16764 10260
rect 16719 10220 16764 10248
rect 16758 10208 16764 10220
rect 16816 10208 16822 10260
rect 17126 10248 17132 10260
rect 17087 10220 17132 10248
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 18012 10220 18061 10248
rect 18012 10208 18018 10220
rect 18049 10217 18061 10220
rect 18095 10248 18107 10251
rect 18690 10248 18696 10260
rect 18095 10220 18696 10248
rect 18095 10217 18107 10220
rect 18049 10211 18107 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 11072 10180 11100 10208
rect 10100 10152 11100 10180
rect 11532 10152 11836 10180
rect 10100 10140 10106 10152
rect 9677 10115 9735 10121
rect 9677 10081 9689 10115
rect 9723 10112 9735 10115
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 9723 10084 10241 10112
rect 9723 10081 9735 10084
rect 9677 10075 9735 10081
rect 10229 10081 10241 10084
rect 10275 10112 10287 10115
rect 11330 10112 11336 10124
rect 10275 10084 11336 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 11330 10072 11336 10084
rect 11388 10072 11394 10124
rect 10042 10044 10048 10056
rect 9600 10016 10048 10044
rect 10042 10004 10048 10016
rect 10100 10004 10106 10056
rect 10318 10044 10324 10056
rect 10279 10016 10324 10044
rect 10318 10004 10324 10016
rect 10376 10004 10382 10056
rect 10502 10044 10508 10056
rect 10463 10016 10508 10044
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 11241 10047 11299 10053
rect 11241 10013 11253 10047
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 8941 9979 8999 9985
rect 8941 9945 8953 9979
rect 8987 9976 8999 9979
rect 9122 9976 9128 9988
rect 8987 9948 9128 9976
rect 8987 9945 8999 9948
rect 8941 9939 8999 9945
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9950 9976 9956 9988
rect 9548 9948 9956 9976
rect 9548 9936 9554 9948
rect 9950 9936 9956 9948
rect 10008 9936 10014 9988
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 11256 9976 11284 10007
rect 11020 9948 11284 9976
rect 11020 9936 11026 9948
rect 9030 9908 9036 9920
rect 7239 9880 8892 9908
rect 8991 9880 9036 9908
rect 7239 9877 7251 9880
rect 7193 9871 7251 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 10502 9908 10508 9920
rect 10284 9880 10508 9908
rect 10284 9868 10290 9880
rect 10502 9868 10508 9880
rect 10560 9908 10566 9920
rect 11532 9917 11560 10152
rect 11701 10115 11759 10121
rect 11701 10081 11713 10115
rect 11747 10081 11759 10115
rect 11701 10075 11759 10081
rect 11517 9911 11575 9917
rect 11517 9908 11529 9911
rect 10560 9880 11529 9908
rect 10560 9868 10566 9880
rect 11517 9877 11529 9880
rect 11563 9877 11575 9911
rect 11716 9908 11744 10075
rect 11808 10044 11836 10152
rect 13078 10140 13084 10192
rect 13136 10180 13142 10192
rect 14645 10183 14703 10189
rect 14645 10180 14657 10183
rect 13136 10152 14657 10180
rect 13136 10140 13142 10152
rect 14645 10149 14657 10152
rect 14691 10149 14703 10183
rect 14645 10143 14703 10149
rect 16574 10140 16580 10192
rect 16632 10180 16638 10192
rect 16632 10152 17264 10180
rect 16632 10140 16638 10152
rect 12158 10121 12164 10124
rect 12152 10075 12164 10121
rect 12216 10112 12222 10124
rect 13725 10115 13783 10121
rect 12216 10084 12252 10112
rect 12158 10072 12164 10075
rect 12216 10072 12222 10084
rect 13725 10081 13737 10115
rect 13771 10112 13783 10115
rect 14550 10112 14556 10124
rect 13771 10084 14556 10112
rect 13771 10081 13783 10084
rect 13725 10075 13783 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 15556 10115 15614 10121
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 16022 10112 16028 10124
rect 15602 10084 16028 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 17236 10112 17264 10152
rect 17236 10084 17356 10112
rect 17328 10056 17356 10084
rect 17770 10072 17776 10124
rect 17828 10112 17834 10124
rect 17957 10115 18015 10121
rect 17957 10112 17969 10115
rect 17828 10084 17969 10112
rect 17828 10072 17834 10084
rect 17957 10081 17969 10084
rect 18003 10112 18015 10115
rect 18414 10112 18420 10124
rect 18003 10084 18420 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 18414 10072 18420 10084
rect 18472 10072 18478 10124
rect 11882 10044 11888 10056
rect 11795 10016 11888 10044
rect 11882 10004 11888 10016
rect 11940 10004 11946 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13740 10016 13829 10044
rect 13740 9988 13768 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10013 13967 10047
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 13909 10007 13967 10013
rect 13354 9976 13360 9988
rect 13096 9948 13360 9976
rect 13096 9908 13124 9948
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 13722 9936 13728 9988
rect 13780 9936 13786 9988
rect 13262 9908 13268 9920
rect 11716 9880 13124 9908
rect 13223 9880 13268 9908
rect 11517 9871 11575 9877
rect 13262 9868 13268 9880
rect 13320 9908 13326 9920
rect 13924 9908 13952 10007
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15289 10047 15347 10053
rect 15289 10044 15301 10047
rect 15160 10016 15301 10044
rect 15160 10004 15166 10016
rect 15289 10013 15301 10016
rect 15335 10013 15347 10047
rect 15289 10007 15347 10013
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 16632 9948 16804 9976
rect 16632 9936 16638 9948
rect 13320 9880 13952 9908
rect 13320 9868 13326 9880
rect 13998 9868 14004 9920
rect 14056 9908 14062 9920
rect 14185 9911 14243 9917
rect 14185 9908 14197 9911
rect 14056 9880 14197 9908
rect 14056 9868 14062 9880
rect 14185 9877 14197 9880
rect 14231 9877 14243 9911
rect 15010 9908 15016 9920
rect 14971 9880 15016 9908
rect 14185 9871 14243 9877
rect 15010 9868 15016 9880
rect 15068 9868 15074 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16669 9911 16727 9917
rect 16669 9908 16681 9911
rect 15712 9880 16681 9908
rect 15712 9868 15718 9880
rect 16669 9877 16681 9880
rect 16715 9877 16727 9911
rect 16776 9908 16804 9948
rect 17236 9908 17264 10007
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 18141 10047 18199 10053
rect 17368 10016 17461 10044
rect 17368 10004 17374 10016
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 17328 9976 17356 10004
rect 18156 9976 18184 10007
rect 17328 9948 18184 9976
rect 17586 9908 17592 9920
rect 16776 9880 17264 9908
rect 17547 9880 17592 9908
rect 16669 9871 16727 9877
rect 17586 9868 17592 9880
rect 17644 9868 17650 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 18230 9908 18236 9920
rect 18012 9880 18236 9908
rect 18012 9868 18018 9880
rect 18230 9868 18236 9880
rect 18288 9868 18294 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 1104 9818 18860 9840
rect 1104 9766 3947 9818
rect 3999 9766 4011 9818
rect 4063 9766 4075 9818
rect 4127 9766 4139 9818
rect 4191 9766 9878 9818
rect 9930 9766 9942 9818
rect 9994 9766 10006 9818
rect 10058 9766 10070 9818
rect 10122 9766 15808 9818
rect 15860 9766 15872 9818
rect 15924 9766 15936 9818
rect 15988 9766 16000 9818
rect 16052 9766 18860 9818
rect 1104 9744 18860 9766
rect 3145 9707 3203 9713
rect 3145 9673 3157 9707
rect 3191 9704 3203 9707
rect 3786 9704 3792 9716
rect 3191 9676 3792 9704
rect 3191 9673 3203 9676
rect 3145 9667 3203 9673
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 5166 9704 5172 9716
rect 4172 9676 5172 9704
rect 2317 9639 2375 9645
rect 2317 9605 2329 9639
rect 2363 9636 2375 9639
rect 3513 9639 3571 9645
rect 2363 9608 3464 9636
rect 2363 9605 2375 9608
rect 2317 9599 2375 9605
rect 2225 9571 2283 9577
rect 2225 9568 2237 9571
rect 1688 9540 2237 9568
rect 1688 9509 1716 9540
rect 2225 9537 2237 9540
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 2958 9568 2964 9580
rect 2832 9540 2877 9568
rect 2919 9540 2964 9568
rect 2832 9528 2838 9540
rect 2958 9528 2964 9540
rect 3016 9528 3022 9580
rect 3436 9568 3464 9608
rect 3513 9605 3525 9639
rect 3559 9636 3571 9639
rect 4172 9636 4200 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 6270 9704 6276 9716
rect 5316 9676 6276 9704
rect 5316 9664 5322 9676
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 7466 9704 7472 9716
rect 6840 9676 7472 9704
rect 4338 9636 4344 9648
rect 3559 9608 4200 9636
rect 4299 9608 4344 9636
rect 3559 9605 3571 9608
rect 3513 9599 3571 9605
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 5810 9636 5816 9648
rect 4488 9608 5816 9636
rect 4488 9596 4494 9608
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 5997 9639 6055 9645
rect 5997 9605 6009 9639
rect 6043 9636 6055 9639
rect 6840 9636 6868 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 9861 9707 9919 9713
rect 9861 9673 9873 9707
rect 9907 9704 9919 9707
rect 10318 9704 10324 9716
rect 9907 9676 10324 9704
rect 9907 9673 9919 9676
rect 9861 9667 9919 9673
rect 10318 9664 10324 9676
rect 10376 9664 10382 9716
rect 10689 9707 10747 9713
rect 10689 9673 10701 9707
rect 10735 9704 10747 9707
rect 10778 9704 10784 9716
rect 10735 9676 10784 9704
rect 10735 9673 10747 9676
rect 10689 9667 10747 9673
rect 10778 9664 10784 9676
rect 10836 9664 10842 9716
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 13722 9704 13728 9716
rect 12216 9676 13400 9704
rect 13683 9676 13728 9704
rect 12216 9664 12222 9676
rect 8202 9636 8208 9648
rect 6043 9608 6868 9636
rect 7852 9608 8208 9636
rect 6043 9605 6055 9608
rect 5997 9599 6055 9605
rect 4062 9568 4068 9580
rect 3436 9540 4068 9568
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4985 9571 5043 9577
rect 4985 9568 4997 9571
rect 4203 9540 4997 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4985 9537 4997 9540
rect 5031 9568 5043 9571
rect 5074 9568 5080 9580
rect 5031 9540 5080 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5718 9568 5724 9580
rect 5679 9540 5724 9568
rect 5718 9528 5724 9540
rect 5776 9528 5782 9580
rect 6012 9568 6040 9599
rect 5828 9540 6040 9568
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9469 1731 9503
rect 1673 9463 1731 9469
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2004 9472 2697 9500
rect 2004 9460 2010 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 3329 9503 3387 9509
rect 3329 9469 3341 9503
rect 3375 9500 3387 9503
rect 5828 9500 5856 9540
rect 3375 9472 5856 9500
rect 6181 9503 6239 9509
rect 3375 9469 3387 9472
rect 3329 9463 3387 9469
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6270 9500 6276 9512
rect 6227 9472 6276 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6825 9503 6883 9509
rect 6825 9500 6837 9503
rect 6604 9472 6837 9500
rect 6604 9460 6610 9472
rect 6825 9469 6837 9472
rect 6871 9469 6883 9503
rect 6825 9463 6883 9469
rect 6914 9460 6920 9512
rect 6972 9500 6978 9512
rect 6972 9472 7236 9500
rect 6972 9460 6978 9472
rect 3234 9432 3240 9444
rect 1872 9404 3240 9432
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 1872 9373 1900 9404
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 3881 9435 3939 9441
rect 3881 9401 3893 9435
rect 3927 9432 3939 9435
rect 3927 9404 4292 9432
rect 3927 9401 3939 9404
rect 3881 9395 3939 9401
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9333 1915 9367
rect 1857 9327 1915 9333
rect 2133 9367 2191 9373
rect 2133 9333 2145 9367
rect 2179 9364 2191 9367
rect 2222 9364 2228 9376
rect 2179 9336 2228 9364
rect 2179 9333 2191 9336
rect 2133 9327 2191 9333
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 2406 9324 2412 9376
rect 2464 9364 2470 9376
rect 3896 9364 3924 9395
rect 2464 9336 3924 9364
rect 2464 9324 2470 9336
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4264 9364 4292 9404
rect 4338 9392 4344 9444
rect 4396 9432 4402 9444
rect 5629 9435 5687 9441
rect 5629 9432 5641 9435
rect 4396 9404 5641 9432
rect 4396 9392 4402 9404
rect 5629 9401 5641 9404
rect 5675 9401 5687 9435
rect 5629 9395 5687 9401
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 6638 9432 6644 9444
rect 6052 9404 6644 9432
rect 6052 9392 6058 9404
rect 6638 9392 6644 9404
rect 6696 9432 6702 9444
rect 7070 9435 7128 9441
rect 7070 9432 7082 9435
rect 6696 9404 7082 9432
rect 6696 9392 6702 9404
rect 7070 9401 7082 9404
rect 7116 9401 7128 9435
rect 7208 9432 7236 9472
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 7852 9500 7880 9608
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 9674 9636 9680 9648
rect 9635 9608 9680 9636
rect 9674 9596 9680 9608
rect 9732 9636 9738 9648
rect 11517 9639 11575 9645
rect 9732 9608 10456 9636
rect 9732 9596 9738 9608
rect 10134 9568 10140 9580
rect 9324 9540 10140 9568
rect 8294 9500 8300 9512
rect 7432 9472 7880 9500
rect 8255 9472 8300 9500
rect 7432 9460 7438 9472
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 9324 9500 9352 9540
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10318 9568 10324 9580
rect 10279 9540 10324 9568
rect 10318 9528 10324 9540
rect 10376 9528 10382 9580
rect 10428 9577 10456 9608
rect 11517 9605 11529 9639
rect 11563 9636 11575 9639
rect 13078 9636 13084 9648
rect 11563 9608 13084 9636
rect 11563 9605 11575 9608
rect 11517 9599 11575 9605
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9568 10471 9571
rect 10962 9568 10968 9580
rect 10459 9540 10968 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10962 9528 10968 9540
rect 11020 9568 11026 9580
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11020 9540 11253 9568
rect 11020 9528 11026 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 13262 9568 13268 9580
rect 12207 9540 13268 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13372 9577 13400 9676
rect 13722 9664 13728 9676
rect 13780 9664 13786 9716
rect 13814 9664 13820 9716
rect 13872 9704 13878 9716
rect 14458 9704 14464 9716
rect 13872 9676 14464 9704
rect 13872 9664 13878 9676
rect 14458 9664 14464 9676
rect 14516 9704 14522 9716
rect 14734 9704 14740 9716
rect 14516 9676 14740 9704
rect 14516 9664 14522 9676
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 15010 9664 15016 9716
rect 15068 9704 15074 9716
rect 16114 9704 16120 9716
rect 15068 9676 16120 9704
rect 15068 9664 15074 9676
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 17402 9664 17408 9716
rect 17460 9664 17466 9716
rect 13633 9639 13691 9645
rect 13633 9605 13645 9639
rect 13679 9636 13691 9639
rect 13906 9636 13912 9648
rect 13679 9608 13912 9636
rect 13679 9605 13691 9608
rect 13633 9599 13691 9605
rect 13906 9596 13912 9608
rect 13964 9596 13970 9648
rect 14550 9636 14556 9648
rect 14511 9608 14556 9636
rect 14550 9596 14556 9608
rect 14608 9596 14614 9648
rect 15194 9596 15200 9648
rect 15252 9636 15258 9648
rect 15381 9639 15439 9645
rect 15381 9636 15393 9639
rect 15252 9608 15393 9636
rect 15252 9596 15258 9608
rect 15381 9605 15393 9608
rect 15427 9605 15439 9639
rect 15381 9599 15439 9605
rect 15565 9639 15623 9645
rect 15565 9605 15577 9639
rect 15611 9636 15623 9639
rect 16574 9636 16580 9648
rect 15611 9608 16580 9636
rect 15611 9605 15623 9608
rect 15565 9599 15623 9605
rect 16574 9596 16580 9608
rect 16632 9596 16638 9648
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16761 9639 16819 9645
rect 16761 9636 16773 9639
rect 16724 9608 16773 9636
rect 16724 9596 16730 9608
rect 16761 9605 16773 9608
rect 16807 9605 16819 9639
rect 16761 9599 16819 9605
rect 13357 9571 13415 9577
rect 13357 9537 13369 9571
rect 13403 9568 13415 9571
rect 14277 9571 14335 9577
rect 14277 9568 14289 9571
rect 13403 9540 14289 9568
rect 13403 9537 13415 9540
rect 13357 9531 13415 9537
rect 14277 9537 14289 9540
rect 14323 9568 14335 9571
rect 15010 9568 15016 9580
rect 14323 9540 15016 9568
rect 14323 9537 14335 9540
rect 14277 9531 14335 9537
rect 15010 9528 15016 9540
rect 15068 9568 15074 9580
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 15068 9540 15117 9568
rect 15068 9528 15074 9540
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 8404 9472 9352 9500
rect 8404 9432 8432 9472
rect 9398 9460 9404 9512
rect 9456 9500 9462 9512
rect 10336 9500 10364 9528
rect 9456 9472 10364 9500
rect 11977 9503 12035 9509
rect 9456 9460 9462 9472
rect 11977 9469 11989 9503
rect 12023 9500 12035 9503
rect 12529 9503 12587 9509
rect 12023 9472 12388 9500
rect 12023 9469 12035 9472
rect 11977 9463 12035 9469
rect 7208 9404 8432 9432
rect 8564 9435 8622 9441
rect 7070 9395 7128 9401
rect 8564 9401 8576 9435
rect 8610 9432 8622 9435
rect 9674 9432 9680 9444
rect 8610 9404 9680 9432
rect 8610 9401 8622 9404
rect 8564 9395 8622 9401
rect 9674 9392 9680 9404
rect 9732 9392 9738 9444
rect 10229 9435 10287 9441
rect 10229 9401 10241 9435
rect 10275 9432 10287 9435
rect 10594 9432 10600 9444
rect 10275 9404 10600 9432
rect 10275 9401 10287 9404
rect 10229 9395 10287 9401
rect 4430 9364 4436 9376
rect 4028 9336 4073 9364
rect 4264 9336 4436 9364
rect 4028 9324 4034 9336
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 4709 9367 4767 9373
rect 4709 9364 4721 9367
rect 4672 9336 4721 9364
rect 4672 9324 4678 9336
rect 4709 9333 4721 9336
rect 4755 9333 4767 9367
rect 4709 9327 4767 9333
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 4982 9364 4988 9376
rect 4847 9336 4988 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5442 9324 5448 9376
rect 5500 9364 5506 9376
rect 5537 9367 5595 9373
rect 5537 9364 5549 9367
rect 5500 9336 5549 9364
rect 5500 9324 5506 9336
rect 5537 9333 5549 9336
rect 5583 9333 5595 9367
rect 5537 9327 5595 9333
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 5868 9336 6561 9364
rect 5868 9324 5874 9336
rect 6549 9333 6561 9336
rect 6595 9364 6607 9367
rect 9030 9364 9036 9376
rect 6595 9336 9036 9364
rect 6595 9333 6607 9336
rect 6549 9327 6607 9333
rect 9030 9324 9036 9336
rect 9088 9364 9094 9376
rect 10244 9364 10272 9395
rect 10594 9392 10600 9404
rect 10652 9392 10658 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 10888 9404 11161 9432
rect 9088 9336 10272 9364
rect 9088 9324 9094 9336
rect 10318 9324 10324 9376
rect 10376 9364 10382 9376
rect 10888 9364 10916 9404
rect 11149 9401 11161 9404
rect 11195 9432 11207 9435
rect 12360 9432 12388 9472
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 12575 9472 14933 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 15212 9500 15240 9596
rect 17420 9580 17448 9664
rect 17678 9596 17684 9648
rect 17736 9636 17742 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17736 9608 18245 9636
rect 17736 9596 17742 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 16117 9571 16175 9577
rect 16117 9568 16129 9571
rect 15344 9540 16129 9568
rect 15344 9528 15350 9540
rect 16117 9537 16129 9540
rect 16163 9537 16175 9571
rect 17310 9568 17316 9580
rect 16117 9531 16175 9537
rect 16500 9540 16712 9568
rect 17271 9540 17316 9568
rect 16500 9500 16528 9540
rect 15212 9472 16528 9500
rect 16577 9503 16635 9509
rect 14921 9463 14979 9469
rect 16577 9469 16589 9503
rect 16623 9469 16635 9503
rect 16684 9500 16712 9540
rect 17310 9528 17316 9540
rect 17368 9528 17374 9580
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 17589 9503 17647 9509
rect 17589 9500 17601 9503
rect 16684 9472 17601 9500
rect 16577 9463 16635 9469
rect 17589 9469 17601 9472
rect 17635 9500 17647 9503
rect 17770 9500 17776 9512
rect 17635 9472 17776 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 13173 9435 13231 9441
rect 11195 9404 12296 9432
rect 12360 9404 12848 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 11054 9364 11060 9376
rect 10376 9336 10916 9364
rect 11015 9336 11060 9364
rect 10376 9324 10382 9336
rect 11054 9324 11060 9336
rect 11112 9364 11118 9376
rect 11606 9364 11612 9376
rect 11112 9336 11612 9364
rect 11112 9324 11118 9336
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 11882 9364 11888 9376
rect 11843 9336 11888 9364
rect 11882 9324 11888 9336
rect 11940 9324 11946 9376
rect 12268 9364 12296 9404
rect 12526 9364 12532 9376
rect 12268 9336 12532 9364
rect 12526 9324 12532 9336
rect 12584 9324 12590 9376
rect 12820 9373 12848 9404
rect 13173 9401 13185 9435
rect 13219 9432 13231 9435
rect 13633 9435 13691 9441
rect 13633 9432 13645 9435
rect 13219 9404 13645 9432
rect 13219 9401 13231 9404
rect 13173 9395 13231 9401
rect 13633 9401 13645 9404
rect 13679 9401 13691 9435
rect 16592 9432 16620 9463
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18049 9503 18107 9509
rect 18049 9469 18061 9503
rect 18095 9500 18107 9503
rect 18414 9500 18420 9512
rect 18095 9472 18420 9500
rect 18095 9469 18107 9472
rect 18049 9463 18107 9469
rect 18414 9460 18420 9472
rect 18472 9460 18478 9512
rect 13633 9395 13691 9401
rect 13924 9404 16620 9432
rect 12805 9367 12863 9373
rect 12805 9333 12817 9367
rect 12851 9333 12863 9367
rect 13262 9364 13268 9376
rect 13223 9336 13268 9364
rect 12805 9327 12863 9333
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13924 9364 13952 9404
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 16942 9432 16948 9444
rect 16816 9404 16948 9432
rect 16816 9392 16822 9404
rect 16942 9392 16948 9404
rect 17000 9432 17006 9444
rect 17129 9435 17187 9441
rect 17129 9432 17141 9435
rect 17000 9404 17141 9432
rect 17000 9392 17006 9404
rect 17129 9401 17141 9404
rect 17175 9401 17187 9435
rect 17129 9395 17187 9401
rect 17221 9435 17279 9441
rect 17221 9401 17233 9435
rect 17267 9432 17279 9435
rect 17310 9432 17316 9444
rect 17267 9404 17316 9432
rect 17267 9401 17279 9404
rect 17221 9395 17279 9401
rect 17310 9392 17316 9404
rect 17368 9432 17374 9444
rect 17954 9432 17960 9444
rect 17368 9404 17960 9432
rect 17368 9392 17374 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 14090 9364 14096 9376
rect 13412 9336 13952 9364
rect 14051 9336 14096 9364
rect 13412 9324 13418 9336
rect 14090 9324 14096 9336
rect 14148 9324 14154 9376
rect 14182 9324 14188 9376
rect 14240 9364 14246 9376
rect 14240 9336 14285 9364
rect 14240 9324 14246 9336
rect 14826 9324 14832 9376
rect 14884 9364 14890 9376
rect 15013 9367 15071 9373
rect 15013 9364 15025 9367
rect 14884 9336 15025 9364
rect 14884 9324 14890 9336
rect 15013 9333 15025 9336
rect 15059 9333 15071 9367
rect 15930 9364 15936 9376
rect 15891 9336 15936 9364
rect 15013 9327 15071 9333
rect 15930 9324 15936 9336
rect 15988 9324 15994 9376
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16114 9364 16120 9376
rect 16071 9336 16120 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 16356 9336 16405 9364
rect 16356 9324 16362 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 17770 9364 17776 9376
rect 17731 9336 17776 9364
rect 16393 9327 16451 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 18230 9324 18236 9376
rect 18288 9364 18294 9376
rect 18417 9367 18475 9373
rect 18417 9364 18429 9367
rect 18288 9336 18429 9364
rect 18288 9324 18294 9336
rect 18417 9333 18429 9336
rect 18463 9333 18475 9367
rect 18417 9327 18475 9333
rect 1104 9274 18860 9296
rect 1104 9222 6912 9274
rect 6964 9222 6976 9274
rect 7028 9222 7040 9274
rect 7092 9222 7104 9274
rect 7156 9222 12843 9274
rect 12895 9222 12907 9274
rect 12959 9222 12971 9274
rect 13023 9222 13035 9274
rect 13087 9222 18860 9274
rect 1104 9200 18860 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 2406 9160 2412 9172
rect 1544 9132 2412 9160
rect 1544 9120 1550 9132
rect 2406 9120 2412 9132
rect 2464 9120 2470 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4982 9160 4988 9172
rect 4212 9132 4988 9160
rect 4212 9120 4218 9132
rect 4982 9120 4988 9132
rect 5040 9160 5046 9172
rect 5350 9160 5356 9172
rect 5040 9132 5356 9160
rect 5040 9120 5046 9132
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6181 9163 6239 9169
rect 6181 9160 6193 9163
rect 6052 9132 6193 9160
rect 6052 9120 6058 9132
rect 6181 9129 6193 9132
rect 6227 9129 6239 9163
rect 6181 9123 6239 9129
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 6362 9160 6368 9172
rect 6319 9132 6368 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6730 9160 6736 9172
rect 6691 9132 6736 9160
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 9398 9160 9404 9172
rect 6840 9132 9404 9160
rect 1940 9095 1998 9101
rect 1940 9061 1952 9095
rect 1986 9092 1998 9095
rect 2958 9092 2964 9104
rect 1986 9064 2964 9092
rect 1986 9061 1998 9064
rect 1940 9055 1998 9061
rect 2958 9052 2964 9064
rect 3016 9052 3022 9104
rect 3418 9092 3424 9104
rect 3379 9064 3424 9092
rect 3418 9052 3424 9064
rect 3476 9092 3482 9104
rect 3970 9092 3976 9104
rect 3476 9064 3976 9092
rect 3476 9052 3482 9064
rect 3970 9052 3976 9064
rect 4028 9092 4034 9104
rect 6840 9092 6868 9132
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 10962 9160 10968 9172
rect 9600 9132 10968 9160
rect 4028 9064 6868 9092
rect 4028 9052 4034 9064
rect 8018 9052 8024 9104
rect 8076 9092 8082 9104
rect 8389 9095 8447 9101
rect 8076 9064 8121 9092
rect 8076 9052 8082 9064
rect 8389 9061 8401 9095
rect 8435 9092 8447 9095
rect 9600 9092 9628 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11149 9163 11207 9169
rect 11149 9129 11161 9163
rect 11195 9160 11207 9163
rect 11422 9160 11428 9172
rect 11195 9132 11428 9160
rect 11195 9129 11207 9132
rect 11149 9123 11207 9129
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 11977 9163 12035 9169
rect 11977 9160 11989 9163
rect 11940 9132 11989 9160
rect 11940 9120 11946 9132
rect 11977 9129 11989 9132
rect 12023 9129 12035 9163
rect 11977 9123 12035 9129
rect 12066 9120 12072 9172
rect 12124 9160 12130 9172
rect 12345 9163 12403 9169
rect 12345 9160 12357 9163
rect 12124 9132 12357 9160
rect 12124 9120 12130 9132
rect 12345 9129 12357 9132
rect 12391 9129 12403 9163
rect 12345 9123 12403 9129
rect 12437 9163 12495 9169
rect 12437 9129 12449 9163
rect 12483 9160 12495 9163
rect 12805 9163 12863 9169
rect 12805 9160 12817 9163
rect 12483 9132 12817 9160
rect 12483 9129 12495 9132
rect 12437 9123 12495 9129
rect 12805 9129 12817 9132
rect 12851 9129 12863 9163
rect 14826 9160 14832 9172
rect 12805 9123 12863 9129
rect 13372 9132 14832 9160
rect 8435 9064 9628 9092
rect 8435 9061 8447 9064
rect 8389 9055 8447 9061
rect 9766 9052 9772 9104
rect 9824 9092 9830 9104
rect 9922 9095 9980 9101
rect 9922 9092 9934 9095
rect 9824 9064 9934 9092
rect 9824 9052 9830 9064
rect 9922 9061 9934 9064
rect 9968 9061 9980 9095
rect 9922 9055 9980 9061
rect 10226 9052 10232 9104
rect 10284 9092 10290 9104
rect 11517 9095 11575 9101
rect 11517 9092 11529 9095
rect 10284 9064 11529 9092
rect 10284 9052 10290 9064
rect 11517 9061 11529 9064
rect 11563 9092 11575 9095
rect 12526 9092 12532 9104
rect 11563 9064 12532 9092
rect 11563 9061 11575 9064
rect 11517 9055 11575 9061
rect 12526 9052 12532 9064
rect 12584 9052 12590 9104
rect 1394 8984 1400 9036
rect 1452 9024 1458 9036
rect 1673 9027 1731 9033
rect 1673 9024 1685 9027
rect 1452 8996 1685 9024
rect 1452 8984 1458 8996
rect 1673 8993 1685 8996
rect 1719 8993 1731 9027
rect 1673 8987 1731 8993
rect 2774 8984 2780 9036
rect 2832 9024 2838 9036
rect 3513 9027 3571 9033
rect 3513 9024 3525 9027
rect 2832 8996 3525 9024
rect 2832 8984 2838 8996
rect 3513 8993 3525 8996
rect 3559 8993 3571 9027
rect 3513 8987 3571 8993
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 4801 9027 4859 9033
rect 4801 9024 4813 9027
rect 3844 8996 4813 9024
rect 3844 8984 3850 8996
rect 4801 8993 4813 8996
rect 4847 8993 4859 9027
rect 4801 8987 4859 8993
rect 5068 9027 5126 9033
rect 5068 8993 5080 9027
rect 5114 9024 5126 9027
rect 5810 9024 5816 9036
rect 5114 8996 5816 9024
rect 5114 8993 5126 8996
rect 5068 8987 5126 8993
rect 5810 8984 5816 8996
rect 5868 8984 5874 9036
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6641 9027 6699 9033
rect 6641 9024 6653 9027
rect 6236 8996 6653 9024
rect 6236 8984 6242 8996
rect 6641 8993 6653 8996
rect 6687 9024 6699 9027
rect 7650 9024 7656 9036
rect 6687 8996 7656 9024
rect 6687 8993 6699 8996
rect 6641 8987 6699 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 7926 9024 7932 9036
rect 7887 8996 7932 9024
rect 7926 8984 7932 8996
rect 7984 8984 7990 9036
rect 8846 9024 8852 9036
rect 8036 8996 8340 9024
rect 8807 8996 8852 9024
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3418 8956 3424 8968
rect 3200 8928 3424 8956
rect 3200 8916 3206 8928
rect 3418 8916 3424 8928
rect 3476 8916 3482 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 4154 8956 4160 8968
rect 3752 8928 4160 8956
rect 3752 8916 3758 8928
rect 4154 8916 4160 8928
rect 4212 8916 4218 8968
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4614 8956 4620 8968
rect 4488 8928 4620 8956
rect 4488 8916 4494 8928
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 6917 8959 6975 8965
rect 6917 8925 6929 8959
rect 6963 8956 6975 8959
rect 7374 8956 7380 8968
rect 6963 8928 7380 8956
rect 6963 8925 6975 8928
rect 6917 8919 6975 8925
rect 7374 8916 7380 8928
rect 7432 8916 7438 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 8036 8956 8064 8996
rect 8202 8956 8208 8968
rect 7515 8928 8064 8956
rect 8163 8928 8208 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 8312 8956 8340 8996
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 9024 8999 9027
rect 9582 9024 9588 9036
rect 8987 8996 9588 9024
rect 8987 8993 8999 8996
rect 8941 8987 8999 8993
rect 8386 8956 8392 8968
rect 8299 8928 8392 8956
rect 8386 8916 8392 8928
rect 8444 8956 8450 8968
rect 8956 8956 8984 8987
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 10502 9024 10508 9036
rect 9723 8996 10508 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11204 8996 11836 9024
rect 11204 8984 11210 8996
rect 9122 8956 9128 8968
rect 8444 8928 8984 8956
rect 9083 8928 9128 8956
rect 8444 8916 8450 8928
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 11514 8916 11520 8968
rect 11572 8956 11578 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11572 8928 11621 8956
rect 11572 8916 11578 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8925 11759 8959
rect 11701 8919 11759 8925
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 3053 8891 3111 8897
rect 3053 8888 3065 8891
rect 2740 8860 3065 8888
rect 2740 8848 2746 8860
rect 3053 8857 3065 8860
rect 3099 8857 3111 8891
rect 3053 8851 3111 8857
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 4706 8888 4712 8900
rect 4120 8860 4712 8888
rect 4120 8848 4126 8860
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 7561 8891 7619 8897
rect 7561 8857 7573 8891
rect 7607 8888 7619 8891
rect 11057 8891 11115 8897
rect 7607 8860 9720 8888
rect 7607 8857 7619 8860
rect 7561 8851 7619 8857
rect 1118 8780 1124 8832
rect 1176 8820 1182 8832
rect 1489 8823 1547 8829
rect 1489 8820 1501 8823
rect 1176 8792 1501 8820
rect 1176 8780 1182 8792
rect 1489 8789 1501 8792
rect 1535 8789 1547 8823
rect 3142 8820 3148 8832
rect 3103 8792 3148 8820
rect 1489 8783 1547 8789
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3602 8780 3608 8832
rect 3660 8820 3666 8832
rect 3697 8823 3755 8829
rect 3697 8820 3709 8823
rect 3660 8792 3709 8820
rect 3660 8780 3666 8792
rect 3697 8789 3709 8792
rect 3743 8789 3755 8823
rect 3697 8783 3755 8789
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 4304 8792 4353 8820
rect 4304 8780 4310 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4614 8820 4620 8832
rect 4527 8792 4620 8820
rect 4341 8783 4399 8789
rect 4614 8780 4620 8792
rect 4672 8820 4678 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 4672 8792 8401 8820
rect 4672 8780 4678 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8820 8539 8823
rect 8570 8820 8576 8832
rect 8527 8792 8576 8820
rect 8527 8789 8539 8792
rect 8481 8783 8539 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 8846 8780 8852 8832
rect 8904 8820 8910 8832
rect 9490 8820 9496 8832
rect 8904 8792 9496 8820
rect 8904 8780 8910 8792
rect 9490 8780 9496 8792
rect 9548 8780 9554 8832
rect 9692 8820 9720 8860
rect 11057 8857 11069 8891
rect 11103 8888 11115 8891
rect 11330 8888 11336 8900
rect 11103 8860 11336 8888
rect 11103 8857 11115 8860
rect 11057 8851 11115 8857
rect 11330 8848 11336 8860
rect 11388 8888 11394 8900
rect 11716 8888 11744 8919
rect 11388 8860 11744 8888
rect 11808 8888 11836 8996
rect 13078 8984 13084 9036
rect 13136 9024 13142 9036
rect 13173 9027 13231 9033
rect 13173 9024 13185 9027
rect 13136 8996 13185 9024
rect 13136 8984 13142 8996
rect 13173 8993 13185 8996
rect 13219 8993 13231 9027
rect 13173 8987 13231 8993
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 12216 8928 12541 8956
rect 12216 8916 12222 8928
rect 12529 8925 12541 8928
rect 12575 8925 12587 8959
rect 12529 8919 12587 8925
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8925 13323 8959
rect 13265 8919 13323 8925
rect 13170 8888 13176 8900
rect 11808 8860 13176 8888
rect 11388 8848 11394 8860
rect 13170 8848 13176 8860
rect 13228 8888 13234 8900
rect 13280 8888 13308 8919
rect 13228 8860 13308 8888
rect 13228 8848 13234 8860
rect 10870 8820 10876 8832
rect 9692 8792 10876 8820
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 13372 8820 13400 9132
rect 14826 9120 14832 9132
rect 14884 9120 14890 9172
rect 15010 9160 15016 9172
rect 14971 9132 15016 9160
rect 15010 9120 15016 9132
rect 15068 9120 15074 9172
rect 15930 9160 15936 9172
rect 15120 9132 15936 9160
rect 13814 9052 13820 9104
rect 13872 9101 13878 9104
rect 13872 9095 13936 9101
rect 13872 9061 13890 9095
rect 13924 9061 13936 9095
rect 13872 9055 13936 9061
rect 13872 9052 13878 9055
rect 14090 9052 14096 9104
rect 14148 9092 14154 9104
rect 14148 9064 14228 9092
rect 14148 9052 14154 9064
rect 13832 9024 13860 9052
rect 13464 8996 13860 9024
rect 14200 9024 14228 9064
rect 14274 9052 14280 9104
rect 14332 9092 14338 9104
rect 14550 9092 14556 9104
rect 14332 9064 14556 9092
rect 14332 9052 14338 9064
rect 14550 9052 14556 9064
rect 14608 9092 14614 9104
rect 15120 9092 15148 9132
rect 15930 9120 15936 9132
rect 15988 9160 15994 9172
rect 16482 9160 16488 9172
rect 15988 9132 16488 9160
rect 15988 9120 15994 9132
rect 16482 9120 16488 9132
rect 16540 9120 16546 9172
rect 17405 9163 17463 9169
rect 17405 9129 17417 9163
rect 17451 9160 17463 9163
rect 17586 9160 17592 9172
rect 17451 9132 17592 9160
rect 17451 9129 17463 9132
rect 17405 9123 17463 9129
rect 17586 9120 17592 9132
rect 17644 9120 17650 9172
rect 15654 9101 15660 9104
rect 15648 9092 15660 9101
rect 14608 9064 15148 9092
rect 15615 9064 15660 9092
rect 14608 9052 14614 9064
rect 15648 9055 15660 9064
rect 15654 9052 15660 9055
rect 15712 9052 15718 9104
rect 17313 9095 17371 9101
rect 17313 9061 17325 9095
rect 17359 9092 17371 9095
rect 17494 9092 17500 9104
rect 17359 9064 17500 9092
rect 17359 9061 17371 9064
rect 17313 9055 17371 9061
rect 17494 9052 17500 9064
rect 17552 9052 17558 9104
rect 18414 9092 18420 9104
rect 17604 9064 18420 9092
rect 17604 9024 17632 9064
rect 18414 9052 18420 9064
rect 18472 9052 18478 9104
rect 14200 8996 17632 9024
rect 17865 9027 17923 9033
rect 13464 8965 13492 8996
rect 17865 8993 17877 9027
rect 17911 9024 17923 9027
rect 17954 9024 17960 9036
rect 17911 8996 17960 9024
rect 17911 8993 17923 8996
rect 17865 8987 17923 8993
rect 17954 8984 17960 8996
rect 18012 8984 18018 9036
rect 18230 9024 18236 9036
rect 18191 8996 18236 9024
rect 18230 8984 18236 8996
rect 18288 8984 18294 9036
rect 13449 8959 13507 8965
rect 13449 8925 13461 8959
rect 13495 8925 13507 8959
rect 13449 8919 13507 8925
rect 13633 8959 13691 8965
rect 13633 8925 13645 8959
rect 13679 8925 13691 8959
rect 13633 8919 13691 8925
rect 15381 8959 15439 8965
rect 15381 8925 15393 8959
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 11020 8792 13400 8820
rect 13648 8820 13676 8919
rect 14274 8820 14280 8832
rect 13648 8792 14280 8820
rect 11020 8780 11026 8792
rect 14274 8780 14280 8792
rect 14332 8820 14338 8832
rect 15102 8820 15108 8832
rect 14332 8792 15108 8820
rect 14332 8780 14338 8792
rect 15102 8780 15108 8792
rect 15160 8820 15166 8832
rect 15396 8820 15424 8919
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17276 8928 17509 8956
rect 17276 8916 17282 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17862 8848 17868 8900
rect 17920 8888 17926 8900
rect 18417 8891 18475 8897
rect 18417 8888 18429 8891
rect 17920 8860 18429 8888
rect 17920 8848 17926 8860
rect 18417 8857 18429 8860
rect 18463 8857 18475 8891
rect 18417 8851 18475 8857
rect 16298 8820 16304 8832
rect 15160 8792 16304 8820
rect 15160 8780 15166 8792
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 16761 8823 16819 8829
rect 16761 8820 16773 8823
rect 16632 8792 16773 8820
rect 16632 8780 16638 8792
rect 16761 8789 16773 8792
rect 16807 8789 16819 8823
rect 16942 8820 16948 8832
rect 16903 8792 16948 8820
rect 16761 8783 16819 8789
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 18049 8823 18107 8829
rect 18049 8820 18061 8823
rect 17644 8792 18061 8820
rect 17644 8780 17650 8792
rect 18049 8789 18061 8792
rect 18095 8789 18107 8823
rect 18049 8783 18107 8789
rect 1104 8730 18860 8752
rect 1104 8678 3947 8730
rect 3999 8678 4011 8730
rect 4063 8678 4075 8730
rect 4127 8678 4139 8730
rect 4191 8678 9878 8730
rect 9930 8678 9942 8730
rect 9994 8678 10006 8730
rect 10058 8678 10070 8730
rect 10122 8678 15808 8730
rect 15860 8678 15872 8730
rect 15924 8678 15936 8730
rect 15988 8678 16000 8730
rect 16052 8678 18860 8730
rect 1104 8656 18860 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2280 8588 5764 8616
rect 2280 8576 2286 8588
rect 5736 8548 5764 8588
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5868 8588 5917 8616
rect 5868 8576 5874 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 6178 8616 6184 8628
rect 6139 8588 6184 8616
rect 5905 8579 5963 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 7742 8616 7748 8628
rect 6840 8588 7748 8616
rect 6840 8548 6868 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 8205 8619 8263 8625
rect 8205 8585 8217 8619
rect 8251 8616 8263 8619
rect 9674 8616 9680 8628
rect 8251 8588 9680 8616
rect 8251 8585 8263 8588
rect 8205 8579 8263 8585
rect 9674 8576 9680 8588
rect 9732 8616 9738 8628
rect 10410 8616 10416 8628
rect 9732 8588 10416 8616
rect 9732 8576 9738 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 11146 8616 11152 8628
rect 10520 8588 11152 8616
rect 5736 8520 6868 8548
rect 9398 8508 9404 8560
rect 9456 8548 9462 8560
rect 10520 8548 10548 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11790 8616 11796 8628
rect 11664 8588 11796 8616
rect 11664 8576 11670 8588
rect 11790 8576 11796 8588
rect 11848 8616 11854 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11848 8588 11897 8616
rect 11848 8576 11854 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13262 8616 13268 8628
rect 13219 8588 13268 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13262 8576 13268 8588
rect 13320 8576 13326 8628
rect 14090 8616 14096 8628
rect 14051 8588 14096 8616
rect 14090 8576 14096 8588
rect 14148 8576 14154 8628
rect 16114 8616 16120 8628
rect 16075 8588 16120 8616
rect 16114 8576 16120 8588
rect 16172 8576 16178 8628
rect 17494 8616 17500 8628
rect 16316 8588 17500 8616
rect 9456 8520 10548 8548
rect 11977 8551 12035 8557
rect 9456 8508 9462 8520
rect 11977 8517 11989 8551
rect 12023 8548 12035 8551
rect 12526 8548 12532 8560
rect 12023 8520 12532 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 12713 8551 12771 8557
rect 12713 8517 12725 8551
rect 12759 8548 12771 8551
rect 13354 8548 13360 8560
rect 12759 8520 13360 8548
rect 12759 8517 12771 8520
rect 12713 8511 12771 8517
rect 13354 8508 13360 8520
rect 13412 8508 13418 8560
rect 16316 8548 16344 8588
rect 17494 8576 17500 8588
rect 17552 8576 17558 8628
rect 15948 8520 16344 8548
rect 18233 8551 18291 8557
rect 1394 8440 1400 8492
rect 1452 8480 1458 8492
rect 1581 8483 1639 8489
rect 1581 8480 1593 8483
rect 1452 8452 1593 8480
rect 1452 8440 1458 8452
rect 1581 8449 1593 8452
rect 1627 8449 1639 8483
rect 1581 8443 1639 8449
rect 1596 8412 1624 8443
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9858 8480 9864 8492
rect 9548 8452 9864 8480
rect 9548 8440 9554 8452
rect 9858 8440 9864 8452
rect 9916 8440 9922 8492
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8480 10287 8483
rect 10275 8452 10640 8480
rect 10275 8449 10287 8452
rect 10229 8443 10287 8449
rect 10612 8424 10640 8452
rect 3053 8415 3111 8421
rect 3053 8412 3065 8415
rect 1596 8384 3065 8412
rect 3053 8381 3065 8384
rect 3099 8412 3111 8415
rect 3786 8412 3792 8424
rect 3099 8384 3792 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3786 8372 3792 8384
rect 3844 8412 3850 8424
rect 4525 8415 4583 8421
rect 4525 8412 4537 8415
rect 3844 8384 4537 8412
rect 3844 8372 3850 8384
rect 4525 8381 4537 8384
rect 4571 8381 4583 8415
rect 4525 8375 4583 8381
rect 5902 8372 5908 8424
rect 5960 8412 5966 8424
rect 6546 8412 6552 8424
rect 5960 8384 6552 8412
rect 5960 8372 5966 8384
rect 6546 8372 6552 8384
rect 6604 8412 6610 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6604 8384 6837 8412
rect 6604 8372 6610 8384
rect 6825 8381 6837 8384
rect 6871 8412 6883 8415
rect 8294 8412 8300 8424
rect 6871 8384 8300 8412
rect 6871 8381 6883 8384
rect 6825 8375 6883 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 8564 8415 8622 8421
rect 8564 8381 8576 8415
rect 8610 8412 8622 8415
rect 9122 8412 9128 8424
rect 8610 8384 9128 8412
rect 8610 8381 8622 8384
rect 8564 8375 8622 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 10318 8412 10324 8424
rect 10279 8384 10324 8412
rect 10318 8372 10324 8384
rect 10376 8372 10382 8424
rect 10502 8412 10508 8424
rect 10415 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 11054 8372 11060 8424
rect 11112 8412 11118 8424
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11112 8384 12173 8412
rect 11112 8372 11118 8384
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12544 8412 12572 8508
rect 13170 8440 13176 8492
rect 13228 8440 13234 8492
rect 13814 8480 13820 8492
rect 13775 8452 13820 8480
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12544 8384 12909 8412
rect 12161 8375 12219 8381
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 13188 8412 13216 8440
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13188 8384 14197 8412
rect 12897 8375 12955 8381
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 1848 8347 1906 8353
rect 1848 8313 1860 8347
rect 1894 8344 1906 8347
rect 2682 8344 2688 8356
rect 1894 8316 2688 8344
rect 1894 8313 1906 8316
rect 1848 8307 1906 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 3298 8347 3356 8353
rect 3298 8344 3310 8347
rect 2976 8316 3310 8344
rect 2976 8288 3004 8316
rect 3298 8313 3310 8316
rect 3344 8313 3356 8347
rect 4770 8347 4828 8353
rect 4770 8344 4782 8347
rect 3298 8307 3356 8313
rect 4448 8316 4782 8344
rect 4448 8288 4476 8316
rect 4770 8313 4782 8316
rect 4816 8313 4828 8347
rect 4770 8307 4828 8313
rect 4982 8304 4988 8356
rect 5040 8344 5046 8356
rect 6362 8344 6368 8356
rect 5040 8316 6368 8344
rect 5040 8304 5046 8316
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 7092 8347 7150 8353
rect 7092 8313 7104 8347
rect 7138 8344 7150 8347
rect 7282 8344 7288 8356
rect 7138 8316 7288 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 9508 8316 10057 8344
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 2958 8276 2964 8288
rect 2919 8248 2964 8276
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3786 8276 3792 8288
rect 3660 8248 3792 8276
rect 3660 8236 3666 8248
rect 3786 8236 3792 8248
rect 3844 8236 3850 8288
rect 4430 8276 4436 8288
rect 4391 8248 4436 8276
rect 4430 8236 4436 8248
rect 4488 8236 4494 8288
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 5776 8248 6469 8276
rect 5776 8236 5782 8248
rect 6457 8245 6469 8248
rect 6503 8276 6515 8279
rect 7374 8276 7380 8288
rect 6503 8248 7380 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 7374 8236 7380 8248
rect 7432 8236 7438 8288
rect 8846 8236 8852 8288
rect 8904 8276 8910 8288
rect 9508 8276 9536 8316
rect 10045 8313 10057 8316
rect 10091 8344 10103 8347
rect 10226 8344 10232 8356
rect 10091 8316 10232 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 9674 8276 9680 8288
rect 8904 8248 9536 8276
rect 9635 8248 9680 8276
rect 8904 8236 8910 8248
rect 9674 8236 9680 8248
rect 9732 8236 9738 8288
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 10520 8276 10548 8372
rect 10772 8347 10830 8353
rect 10772 8313 10784 8347
rect 10818 8344 10830 8347
rect 11330 8344 11336 8356
rect 10818 8316 11336 8344
rect 10818 8313 10830 8316
rect 10772 8307 10830 8313
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 13170 8344 13176 8356
rect 13004 8316 13176 8344
rect 12158 8276 12164 8288
rect 10520 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12437 8279 12495 8285
rect 12437 8276 12449 8279
rect 12308 8248 12449 8276
rect 12308 8236 12314 8248
rect 12437 8245 12449 8248
rect 12483 8276 12495 8279
rect 12618 8276 12624 8288
rect 12483 8248 12624 8276
rect 12483 8245 12495 8248
rect 12437 8239 12495 8245
rect 12618 8236 12624 8248
rect 12676 8276 12682 8288
rect 13004 8285 13032 8316
rect 13170 8304 13176 8316
rect 13228 8344 13234 8356
rect 13633 8347 13691 8353
rect 13633 8344 13645 8347
rect 13228 8316 13645 8344
rect 13228 8304 13234 8316
rect 13633 8313 13645 8316
rect 13679 8344 13691 8347
rect 13722 8344 13728 8356
rect 13679 8316 13728 8344
rect 13679 8313 13691 8316
rect 13633 8307 13691 8313
rect 13722 8304 13728 8316
rect 13780 8304 13786 8356
rect 14200 8344 14228 8375
rect 14274 8372 14280 8424
rect 14332 8412 14338 8424
rect 14369 8415 14427 8421
rect 14369 8412 14381 8415
rect 14332 8384 14381 8412
rect 14332 8372 14338 8384
rect 14369 8381 14381 8384
rect 14415 8381 14427 8415
rect 14369 8375 14427 8381
rect 15010 8372 15016 8424
rect 15068 8412 15074 8424
rect 15948 8421 15976 8520
rect 18233 8517 18245 8551
rect 18279 8548 18291 8551
rect 18782 8548 18788 8560
rect 18279 8520 18788 8548
rect 18279 8517 18291 8520
rect 18233 8511 18291 8517
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 16298 8480 16304 8492
rect 16259 8452 16304 8480
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 16574 8421 16580 8424
rect 15933 8415 15991 8421
rect 15933 8412 15945 8415
rect 15068 8384 15945 8412
rect 15068 8372 15074 8384
rect 15933 8381 15945 8384
rect 15979 8381 15991 8415
rect 16568 8412 16580 8421
rect 16535 8384 16580 8412
rect 15933 8375 15991 8381
rect 16568 8375 16580 8384
rect 16574 8372 16580 8375
rect 16632 8372 16638 8424
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 18049 8415 18107 8421
rect 18049 8412 18061 8415
rect 16908 8384 18061 8412
rect 16908 8372 16914 8384
rect 18049 8381 18061 8384
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 14458 8344 14464 8356
rect 14200 8316 14464 8344
rect 14458 8304 14464 8316
rect 14516 8304 14522 8356
rect 14636 8347 14694 8353
rect 14636 8313 14648 8347
rect 14682 8344 14694 8347
rect 16666 8344 16672 8356
rect 14682 8316 16672 8344
rect 14682 8313 14694 8316
rect 14636 8307 14694 8313
rect 16666 8304 16672 8316
rect 16724 8344 16730 8356
rect 16724 8316 17724 8344
rect 16724 8304 16730 8316
rect 12989 8279 13047 8285
rect 12989 8276 13001 8279
rect 12676 8248 13001 8276
rect 12676 8236 12682 8248
rect 12989 8245 13001 8248
rect 13035 8245 13047 8279
rect 13538 8276 13544 8288
rect 13499 8248 13544 8276
rect 12989 8239 13047 8245
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 15749 8279 15807 8285
rect 15749 8245 15761 8279
rect 15795 8276 15807 8279
rect 16390 8276 16396 8288
rect 15795 8248 16396 8276
rect 15795 8245 15807 8248
rect 15749 8239 15807 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 17696 8285 17724 8316
rect 17681 8279 17739 8285
rect 17681 8245 17693 8279
rect 17727 8245 17739 8279
rect 17681 8239 17739 8245
rect 17770 8236 17776 8288
rect 17828 8276 17834 8288
rect 17954 8276 17960 8288
rect 17828 8248 17960 8276
rect 17828 8236 17834 8248
rect 17954 8236 17960 8248
rect 18012 8236 18018 8288
rect 18138 8236 18144 8288
rect 18196 8276 18202 8288
rect 18417 8279 18475 8285
rect 18417 8276 18429 8279
rect 18196 8248 18429 8276
rect 18196 8236 18202 8248
rect 18417 8245 18429 8248
rect 18463 8245 18475 8279
rect 18417 8239 18475 8245
rect 1104 8186 18860 8208
rect 1104 8134 6912 8186
rect 6964 8134 6976 8186
rect 7028 8134 7040 8186
rect 7092 8134 7104 8186
rect 7156 8134 12843 8186
rect 12895 8134 12907 8186
rect 12959 8134 12971 8186
rect 13023 8134 13035 8186
rect 13087 8134 18860 8186
rect 1104 8112 18860 8134
rect 2774 8032 2780 8084
rect 2832 8072 2838 8084
rect 3050 8072 3056 8084
rect 2832 8044 3056 8072
rect 2832 8032 2838 8044
rect 3050 8032 3056 8044
rect 3108 8032 3114 8084
rect 3878 8072 3884 8084
rect 3839 8044 3884 8072
rect 3878 8032 3884 8044
rect 3936 8032 3942 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4304 8044 4445 8072
rect 4304 8032 4310 8044
rect 4433 8041 4445 8044
rect 4479 8072 4491 8075
rect 4890 8072 4896 8084
rect 4479 8044 4896 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4890 8032 4896 8044
rect 4948 8032 4954 8084
rect 7374 8072 7380 8084
rect 5276 8044 7236 8072
rect 7335 8044 7380 8072
rect 2406 7964 2412 8016
rect 2464 8004 2470 8016
rect 3145 8007 3203 8013
rect 3145 8004 3157 8007
rect 2464 7976 3157 8004
rect 2464 7964 2470 7976
rect 3145 7973 3157 7976
rect 3191 7973 3203 8007
rect 3896 8004 3924 8032
rect 5276 8013 5304 8044
rect 7208 8016 7236 8044
rect 7374 8032 7380 8044
rect 7432 8072 7438 8084
rect 7837 8075 7895 8081
rect 7837 8072 7849 8075
rect 7432 8044 7849 8072
rect 7432 8032 7438 8044
rect 7837 8041 7849 8044
rect 7883 8041 7895 8075
rect 7837 8035 7895 8041
rect 8018 8032 8024 8084
rect 8076 8072 8082 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 8076 8044 8125 8072
rect 8076 8032 8082 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8478 8072 8484 8084
rect 8439 8044 8484 8072
rect 8113 8035 8171 8041
rect 8478 8032 8484 8044
rect 8536 8072 8542 8084
rect 10594 8072 10600 8084
rect 8536 8044 10600 8072
rect 8536 8032 8542 8044
rect 10594 8032 10600 8044
rect 10652 8032 10658 8084
rect 11517 8075 11575 8081
rect 11517 8041 11529 8075
rect 11563 8072 11575 8075
rect 11790 8072 11796 8084
rect 11563 8044 11796 8072
rect 11563 8041 11575 8044
rect 11517 8035 11575 8041
rect 11790 8032 11796 8044
rect 11848 8032 11854 8084
rect 12618 8072 12624 8084
rect 12360 8044 12624 8072
rect 5261 8007 5319 8013
rect 5261 8004 5273 8007
rect 3896 7976 5273 8004
rect 3145 7967 3203 7973
rect 5261 7973 5273 7976
rect 5307 7973 5319 8007
rect 5261 7967 5319 7973
rect 5350 7964 5356 8016
rect 5408 8004 5414 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 5408 7976 5733 8004
rect 5408 7964 5414 7976
rect 5721 7973 5733 7976
rect 5767 7973 5779 8007
rect 5721 7967 5779 7973
rect 7190 7964 7196 8016
rect 7248 7964 7254 8016
rect 10502 8004 10508 8016
rect 7668 7976 10508 8004
rect 1581 7939 1639 7945
rect 1581 7905 1593 7939
rect 1627 7936 1639 7939
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 1627 7908 2237 7936
rect 1627 7905 1639 7908
rect 1581 7899 1639 7905
rect 2225 7905 2237 7908
rect 2271 7936 2283 7939
rect 2590 7936 2596 7948
rect 2271 7908 2596 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 5902 7936 5908 7948
rect 5368 7908 5764 7936
rect 5863 7908 5908 7936
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 1688 7840 2329 7868
rect 1688 7744 1716 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2682 7868 2688 7880
rect 2547 7840 2688 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 2682 7828 2688 7840
rect 2740 7868 2746 7880
rect 2866 7868 2872 7880
rect 2740 7840 2872 7868
rect 2740 7828 2746 7840
rect 2866 7828 2872 7840
rect 2924 7868 2930 7880
rect 3237 7871 3295 7877
rect 3237 7868 3249 7871
rect 2924 7840 3249 7868
rect 2924 7828 2930 7840
rect 3237 7837 3249 7840
rect 3283 7837 3295 7871
rect 4522 7868 4528 7880
rect 4483 7840 4528 7868
rect 3237 7831 3295 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 5368 7877 5396 7908
rect 5736 7880 5764 7908
rect 5902 7896 5908 7908
rect 5960 7896 5966 7948
rect 6172 7939 6230 7945
rect 6172 7905 6184 7939
rect 6218 7936 6230 7939
rect 7374 7936 7380 7948
rect 6218 7908 7380 7936
rect 6218 7905 6230 7908
rect 6172 7899 6230 7905
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 5353 7871 5411 7877
rect 5353 7837 5365 7871
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5445 7871 5503 7877
rect 5445 7837 5457 7871
rect 5491 7837 5503 7871
rect 5445 7831 5503 7837
rect 2958 7760 2964 7812
rect 3016 7800 3022 7812
rect 4632 7800 4660 7831
rect 5166 7800 5172 7812
rect 3016 7772 5172 7800
rect 3016 7760 3022 7772
rect 5166 7760 5172 7772
rect 5224 7800 5230 7812
rect 5460 7800 5488 7831
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7668 7877 7696 7976
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 11977 8007 12035 8013
rect 11977 7973 11989 8007
rect 12023 8004 12035 8007
rect 12023 7976 12112 8004
rect 12023 7973 12035 7976
rect 11977 7967 12035 7973
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 9306 7936 9312 7948
rect 7883 7908 9312 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 9306 7896 9312 7908
rect 9364 7936 9370 7948
rect 9401 7939 9459 7945
rect 9401 7936 9413 7939
rect 9364 7908 9413 7936
rect 9364 7896 9370 7908
rect 9401 7905 9413 7908
rect 9447 7936 9459 7939
rect 9490 7936 9496 7948
rect 9447 7908 9496 7936
rect 9447 7905 9459 7908
rect 9401 7899 9459 7905
rect 9490 7896 9496 7908
rect 9548 7896 9554 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 7653 7871 7711 7877
rect 7653 7868 7665 7871
rect 7156 7840 7665 7868
rect 7156 7828 7162 7840
rect 7653 7837 7665 7840
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 8754 7868 8760 7880
rect 8628 7840 8673 7868
rect 8715 7840 8760 7868
rect 8628 7828 8634 7840
rect 8754 7828 8760 7840
rect 8812 7828 8818 7880
rect 9692 7868 9720 7899
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12084 7936 12112 7976
rect 12360 7936 12388 8044
rect 12618 8032 12624 8044
rect 12676 8032 12682 8084
rect 13906 8072 13912 8084
rect 13867 8044 13912 8072
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 14182 8032 14188 8084
rect 14240 8072 14246 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 14240 8044 14289 8072
rect 14240 8032 14246 8044
rect 14277 8041 14289 8044
rect 14323 8072 14335 8075
rect 14734 8072 14740 8084
rect 14323 8044 14740 8072
rect 14323 8041 14335 8044
rect 14277 8035 14335 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 15749 8075 15807 8081
rect 15749 8041 15761 8075
rect 15795 8072 15807 8075
rect 16942 8072 16948 8084
rect 15795 8044 16948 8072
rect 15795 8041 15807 8044
rect 15749 8035 15807 8041
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17681 8075 17739 8081
rect 17681 8072 17693 8075
rect 17552 8044 17693 8072
rect 17552 8032 17558 8044
rect 17681 8041 17693 8044
rect 17727 8041 17739 8075
rect 17681 8035 17739 8041
rect 12704 8007 12762 8013
rect 12704 7973 12716 8007
rect 12750 8004 12762 8007
rect 12802 8004 12808 8016
rect 12750 7976 12808 8004
rect 12750 7973 12762 7976
rect 12704 7967 12762 7973
rect 12802 7964 12808 7976
rect 12860 7964 12866 8016
rect 15378 7964 15384 8016
rect 15436 8004 15442 8016
rect 15841 8007 15899 8013
rect 15841 8004 15853 8007
rect 15436 7976 15853 8004
rect 15436 7964 15442 7976
rect 15841 7973 15853 7976
rect 15887 7973 15899 8007
rect 15841 7967 15899 7973
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16632 7976 16988 8004
rect 16632 7964 16638 7976
rect 11940 7908 11985 7936
rect 12084 7908 12388 7936
rect 11940 7896 11946 7908
rect 13722 7896 13728 7948
rect 13780 7936 13786 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 13780 7908 16313 7936
rect 13780 7896 13786 7908
rect 16301 7905 16313 7908
rect 16347 7936 16359 7939
rect 16850 7936 16856 7948
rect 16347 7908 16611 7936
rect 16811 7908 16856 7936
rect 16347 7905 16359 7908
rect 16301 7899 16359 7905
rect 9692 7840 9812 7868
rect 7282 7800 7288 7812
rect 5224 7772 5488 7800
rect 7195 7772 7288 7800
rect 5224 7760 5230 7772
rect 7282 7760 7288 7772
rect 7340 7800 7346 7812
rect 8202 7800 8208 7812
rect 7340 7772 8208 7800
rect 7340 7760 7346 7772
rect 8202 7760 8208 7772
rect 8260 7800 8266 7812
rect 9784 7800 9812 7840
rect 11330 7828 11336 7880
rect 11388 7868 11394 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11388 7840 12081 7868
rect 11388 7828 11394 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12437 7871 12495 7877
rect 12437 7868 12449 7871
rect 12216 7840 12449 7868
rect 12216 7828 12222 7840
rect 12437 7837 12449 7840
rect 12483 7837 12495 7871
rect 12437 7831 12495 7837
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 13906 7868 13912 7880
rect 13688 7840 13912 7868
rect 13688 7828 13694 7840
rect 13906 7828 13912 7840
rect 13964 7868 13970 7880
rect 14369 7871 14427 7877
rect 14369 7868 14381 7871
rect 13964 7840 14381 7868
rect 13964 7828 13970 7840
rect 14369 7837 14381 7840
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 14461 7871 14519 7877
rect 14461 7837 14473 7871
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 13814 7800 13820 7812
rect 8260 7772 9076 7800
rect 9784 7772 12388 7800
rect 13727 7772 13820 7800
rect 8260 7760 8266 7772
rect 1670 7732 1676 7744
rect 1631 7704 1676 7732
rect 1670 7692 1676 7704
rect 1728 7692 1734 7744
rect 1857 7735 1915 7741
rect 1857 7701 1869 7735
rect 1903 7732 1915 7735
rect 2222 7732 2228 7744
rect 1903 7704 2228 7732
rect 1903 7701 1915 7704
rect 1857 7695 1915 7701
rect 2222 7692 2228 7704
rect 2280 7692 2286 7744
rect 2682 7732 2688 7744
rect 2643 7704 2688 7732
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 3602 7732 3608 7744
rect 3563 7704 3608 7732
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 4065 7735 4123 7741
rect 4065 7701 4077 7735
rect 4111 7732 4123 7735
rect 4246 7732 4252 7744
rect 4111 7704 4252 7732
rect 4111 7701 4123 7704
rect 4065 7695 4123 7701
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7732 4951 7735
rect 5626 7732 5632 7744
rect 4939 7704 5632 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 5626 7692 5632 7704
rect 5684 7692 5690 7744
rect 8018 7732 8024 7744
rect 7979 7704 8024 7732
rect 8018 7692 8024 7704
rect 8076 7732 8082 7744
rect 8478 7732 8484 7744
rect 8076 7704 8484 7732
rect 8076 7692 8082 7704
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 8846 7692 8852 7744
rect 8904 7732 8910 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8904 7704 8953 7732
rect 8904 7692 8910 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 9048 7732 9076 7772
rect 10318 7732 10324 7744
rect 9048 7704 10324 7732
rect 8941 7695 8999 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 12360 7732 12388 7772
rect 13814 7760 13820 7772
rect 13872 7800 13878 7812
rect 14476 7800 14504 7831
rect 15654 7828 15660 7880
rect 15712 7868 15718 7880
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 15712 7840 15945 7868
rect 15712 7828 15718 7840
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 16583 7868 16611 7908
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 16960 7936 16988 7976
rect 18138 7936 18144 7948
rect 16960 7908 17080 7936
rect 18099 7908 18144 7936
rect 17052 7877 17080 7908
rect 18138 7896 18144 7908
rect 18196 7896 18202 7948
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16583 7840 16957 7868
rect 15933 7831 15991 7837
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 17037 7831 17095 7837
rect 17678 7828 17684 7880
rect 17736 7868 17742 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 17736 7840 17785 7868
rect 17736 7828 17742 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7837 17923 7871
rect 17865 7831 17923 7837
rect 13872 7772 14504 7800
rect 13872 7760 13878 7772
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 16206 7800 16212 7812
rect 14792 7772 16212 7800
rect 14792 7760 14798 7772
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 17494 7760 17500 7812
rect 17552 7800 17558 7812
rect 17880 7800 17908 7831
rect 17552 7772 17908 7800
rect 17552 7760 17558 7772
rect 14366 7732 14372 7744
rect 12360 7704 14372 7732
rect 14366 7692 14372 7704
rect 14424 7692 14430 7744
rect 14826 7732 14832 7744
rect 14787 7704 14832 7732
rect 14826 7692 14832 7704
rect 14884 7732 14890 7744
rect 15010 7732 15016 7744
rect 14884 7704 15016 7732
rect 14884 7692 14890 7704
rect 15010 7692 15016 7704
rect 15068 7692 15074 7744
rect 15102 7692 15108 7744
rect 15160 7732 15166 7744
rect 15381 7735 15439 7741
rect 15381 7732 15393 7735
rect 15160 7704 15393 7732
rect 15160 7692 15166 7704
rect 15381 7701 15393 7704
rect 15427 7701 15439 7735
rect 15381 7695 15439 7701
rect 16485 7735 16543 7741
rect 16485 7701 16497 7735
rect 16531 7732 16543 7735
rect 16574 7732 16580 7744
rect 16531 7704 16580 7732
rect 16531 7701 16543 7704
rect 16485 7695 16543 7701
rect 16574 7692 16580 7704
rect 16632 7692 16638 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17092 7704 17325 7732
rect 17092 7692 17098 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18969 7735 19027 7741
rect 18969 7732 18981 7735
rect 18371 7704 18981 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18969 7701 18981 7704
rect 19015 7701 19027 7735
rect 18969 7695 19027 7701
rect 1104 7642 18860 7664
rect 1104 7590 3947 7642
rect 3999 7590 4011 7642
rect 4063 7590 4075 7642
rect 4127 7590 4139 7642
rect 4191 7590 9878 7642
rect 9930 7590 9942 7642
rect 9994 7590 10006 7642
rect 10058 7590 10070 7642
rect 10122 7590 15808 7642
rect 15860 7590 15872 7642
rect 15924 7590 15936 7642
rect 15988 7590 16000 7642
rect 16052 7590 18860 7642
rect 1104 7568 18860 7590
rect 2406 7488 2412 7540
rect 2464 7528 2470 7540
rect 2593 7531 2651 7537
rect 2593 7528 2605 7531
rect 2464 7500 2605 7528
rect 2464 7488 2470 7500
rect 2593 7497 2605 7500
rect 2639 7497 2651 7531
rect 2593 7491 2651 7497
rect 2777 7531 2835 7537
rect 2777 7497 2789 7531
rect 2823 7528 2835 7531
rect 4522 7528 4528 7540
rect 2823 7500 4528 7528
rect 2823 7497 2835 7500
rect 2777 7491 2835 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6052 7500 6561 7528
rect 6052 7488 6058 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 2958 7460 2964 7472
rect 2424 7432 2964 7460
rect 2222 7392 2228 7404
rect 2183 7364 2228 7392
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2424 7401 2452 7432
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 4430 7460 4436 7472
rect 4172 7432 4436 7460
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2866 7352 2872 7404
rect 2924 7392 2930 7404
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 2924 7364 3341 7392
rect 2924 7352 2930 7364
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3786 7392 3792 7404
rect 3476 7364 3792 7392
rect 3476 7352 3482 7364
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4172 7401 4200 7432
rect 4430 7420 4436 7432
rect 4488 7460 4494 7472
rect 4488 7432 6040 7460
rect 4488 7420 4494 7432
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4525 7395 4583 7401
rect 4525 7392 4537 7395
rect 4157 7355 4215 7361
rect 4448 7364 4537 7392
rect 4448 7336 4476 7364
rect 4525 7361 4537 7364
rect 4571 7392 4583 7395
rect 4798 7392 4804 7404
rect 4571 7364 4804 7392
rect 4571 7361 4583 7364
rect 4525 7355 4583 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 5166 7392 5172 7404
rect 5127 7364 5172 7392
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 6012 7401 6040 7432
rect 5905 7395 5963 7401
rect 5905 7392 5917 7395
rect 5684 7364 5917 7392
rect 5684 7352 5690 7364
rect 5905 7361 5917 7364
rect 5951 7361 5963 7395
rect 5905 7355 5963 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 1394 7324 1400 7336
rect 1355 7296 1400 7324
rect 1394 7284 1400 7296
rect 1452 7284 1458 7336
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2682 7324 2688 7336
rect 2179 7296 2688 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 3237 7327 3295 7333
rect 3237 7293 3249 7327
rect 3283 7324 3295 7327
rect 3602 7324 3608 7336
rect 3283 7296 3608 7324
rect 3283 7293 3295 7296
rect 3237 7287 3295 7293
rect 3602 7284 3608 7296
rect 3660 7284 3666 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7324 4031 7327
rect 4246 7324 4252 7336
rect 4019 7296 4252 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 4985 7327 5043 7333
rect 4985 7293 4997 7327
rect 5031 7324 5043 7327
rect 6273 7327 6331 7333
rect 6273 7324 6285 7327
rect 5031 7296 6285 7324
rect 5031 7293 5043 7296
rect 4985 7287 5043 7293
rect 6273 7293 6285 7296
rect 6319 7293 6331 7327
rect 6273 7287 6331 7293
rect 4065 7259 4123 7265
rect 4065 7256 4077 7259
rect 1780 7228 4077 7256
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 1780 7197 1808 7228
rect 4065 7225 4077 7228
rect 4111 7225 4123 7259
rect 5813 7259 5871 7265
rect 5813 7256 5825 7259
rect 4065 7219 4123 7225
rect 4632 7228 5825 7256
rect 1765 7191 1823 7197
rect 1765 7157 1777 7191
rect 1811 7157 1823 7191
rect 1765 7151 1823 7157
rect 2866 7148 2872 7200
rect 2924 7188 2930 7200
rect 3145 7191 3203 7197
rect 3145 7188 3157 7191
rect 2924 7160 3157 7188
rect 2924 7148 2930 7160
rect 3145 7157 3157 7160
rect 3191 7188 3203 7191
rect 3418 7188 3424 7200
rect 3191 7160 3424 7188
rect 3191 7157 3203 7160
rect 3145 7151 3203 7157
rect 3418 7148 3424 7160
rect 3476 7148 3482 7200
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 4338 7188 4344 7200
rect 3651 7160 4344 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4632 7197 4660 7228
rect 5813 7225 5825 7228
rect 5859 7225 5871 7259
rect 6564 7256 6592 7491
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 7984 7500 8125 7528
rect 7984 7488 7990 7500
rect 8113 7497 8125 7500
rect 8159 7497 8171 7531
rect 8113 7491 8171 7497
rect 8941 7531 8999 7537
rect 8941 7497 8953 7531
rect 8987 7528 8999 7531
rect 9582 7528 9588 7540
rect 8987 7500 9588 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9692 7500 9904 7528
rect 6825 7463 6883 7469
rect 6825 7429 6837 7463
rect 6871 7460 6883 7463
rect 9692 7460 9720 7500
rect 6871 7432 9720 7460
rect 9769 7463 9827 7469
rect 6871 7429 6883 7432
rect 6825 7423 6883 7429
rect 9769 7429 9781 7463
rect 9815 7429 9827 7463
rect 9769 7423 9827 7429
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 7374 7352 7380 7364
rect 7432 7392 7438 7404
rect 8665 7395 8723 7401
rect 8665 7392 8677 7395
rect 7432 7364 8677 7392
rect 7432 7352 7438 7364
rect 8665 7361 8677 7364
rect 8711 7392 8723 7395
rect 8754 7392 8760 7404
rect 8711 7364 8760 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8754 7352 8760 7364
rect 8812 7392 8818 7404
rect 9493 7395 9551 7401
rect 9493 7392 9505 7395
rect 8812 7364 9505 7392
rect 8812 7352 8818 7364
rect 9493 7361 9505 7364
rect 9539 7392 9551 7395
rect 9674 7392 9680 7404
rect 9539 7364 9680 7392
rect 9539 7361 9551 7364
rect 9493 7355 9551 7361
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 7098 7324 7104 7336
rect 6788 7296 7104 7324
rect 6788 7284 6794 7296
rect 7098 7284 7104 7296
rect 7156 7324 7162 7336
rect 7285 7327 7343 7333
rect 7285 7324 7297 7327
rect 7156 7296 7297 7324
rect 7156 7284 7162 7296
rect 7285 7293 7297 7296
rect 7331 7293 7343 7327
rect 7285 7287 7343 7293
rect 7653 7327 7711 7333
rect 7653 7293 7665 7327
rect 7699 7324 7711 7327
rect 9309 7327 9367 7333
rect 9309 7324 9321 7327
rect 7699 7296 9321 7324
rect 7699 7293 7711 7296
rect 7653 7287 7711 7293
rect 9309 7293 9321 7296
rect 9355 7293 9367 7327
rect 9309 7287 9367 7293
rect 9398 7284 9404 7336
rect 9456 7324 9462 7336
rect 9784 7324 9812 7423
rect 9876 7392 9904 7500
rect 10318 7488 10324 7540
rect 10376 7488 10382 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 12802 7528 12808 7540
rect 11112 7500 12808 7528
rect 11112 7488 11118 7500
rect 12802 7488 12808 7500
rect 12860 7528 12866 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 12860 7500 13829 7528
rect 12860 7488 12866 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 15010 7528 15016 7540
rect 14231 7500 15016 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 10336 7401 10364 7488
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10560 7432 11529 7460
rect 10560 7420 10566 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 11517 7423 11575 7429
rect 13538 7420 13544 7472
rect 13596 7460 13602 7472
rect 14200 7460 14228 7491
rect 15010 7488 15016 7500
rect 15068 7528 15074 7540
rect 16850 7528 16856 7540
rect 15068 7500 16856 7528
rect 15068 7488 15074 7500
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18506 7528 18512 7540
rect 18104 7500 18512 7528
rect 18104 7488 18110 7500
rect 18506 7488 18512 7500
rect 18564 7488 18570 7540
rect 13596 7432 14228 7460
rect 13596 7420 13602 7432
rect 10229 7395 10287 7401
rect 10229 7392 10241 7395
rect 9876 7364 10241 7392
rect 10229 7361 10241 7364
rect 10275 7361 10287 7395
rect 10229 7355 10287 7361
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10468 7364 11161 7392
rect 10468 7352 10474 7364
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 14274 7392 14280 7404
rect 12207 7364 12572 7392
rect 14235 7364 14280 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 10965 7327 11023 7333
rect 10965 7324 10977 7327
rect 9456 7296 9501 7324
rect 9784 7296 10977 7324
rect 9456 7284 9462 7296
rect 10965 7293 10977 7296
rect 11011 7293 11023 7327
rect 12176 7324 12204 7355
rect 12250 7324 12256 7336
rect 12176 7296 12256 7324
rect 10965 7287 11023 7293
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 12437 7327 12495 7333
rect 12437 7293 12449 7327
rect 12483 7293 12495 7327
rect 12544 7324 12572 7364
rect 14274 7352 14280 7364
rect 14332 7352 14338 7404
rect 15749 7395 15807 7401
rect 15749 7361 15761 7395
rect 15795 7392 15807 7395
rect 16390 7392 16396 7404
rect 15795 7364 16396 7392
rect 15795 7361 15807 7364
rect 15749 7355 15807 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 16574 7392 16580 7404
rect 16535 7364 16580 7392
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16666 7352 16672 7404
rect 16724 7392 16730 7404
rect 17494 7392 17500 7404
rect 16724 7364 17500 7392
rect 16724 7352 16730 7364
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18230 7392 18236 7404
rect 18012 7364 18236 7392
rect 18012 7352 18018 7364
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 12693 7327 12751 7333
rect 12693 7324 12705 7327
rect 12544 7296 12705 7324
rect 12437 7287 12495 7293
rect 12693 7293 12705 7296
rect 12739 7293 12751 7327
rect 12693 7287 12751 7293
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 6564 7228 7205 7256
rect 5813 7219 5871 7225
rect 7193 7225 7205 7228
rect 7239 7225 7251 7259
rect 7193 7219 7251 7225
rect 4617 7191 4675 7197
rect 4617 7157 4629 7191
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 4890 7148 4896 7200
rect 4948 7188 4954 7200
rect 5077 7191 5135 7197
rect 5077 7188 5089 7191
rect 4948 7160 5089 7188
rect 4948 7148 4954 7160
rect 5077 7157 5089 7160
rect 5123 7188 5135 7191
rect 5350 7188 5356 7200
rect 5123 7160 5356 7188
rect 5123 7157 5135 7160
rect 5077 7151 5135 7157
rect 5350 7148 5356 7160
rect 5408 7148 5414 7200
rect 5445 7191 5503 7197
rect 5445 7157 5457 7191
rect 5491 7188 5503 7191
rect 5626 7188 5632 7200
rect 5491 7160 5632 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 5626 7148 5632 7160
rect 5684 7148 5690 7200
rect 7208 7188 7236 7219
rect 7834 7216 7840 7268
rect 7892 7256 7898 7268
rect 7929 7259 7987 7265
rect 7929 7256 7941 7259
rect 7892 7228 7941 7256
rect 7892 7216 7898 7228
rect 7929 7225 7941 7228
rect 7975 7256 7987 7259
rect 8481 7259 8539 7265
rect 8481 7256 8493 7259
rect 7975 7228 8493 7256
rect 7975 7225 7987 7228
rect 7929 7219 7987 7225
rect 8481 7225 8493 7228
rect 8527 7256 8539 7259
rect 8527 7228 8984 7256
rect 8527 7225 8539 7228
rect 8481 7219 8539 7225
rect 8386 7188 8392 7200
rect 7208 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 8846 7188 8852 7200
rect 8619 7160 8852 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 8846 7148 8852 7160
rect 8904 7148 8910 7200
rect 8956 7188 8984 7228
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 10137 7259 10195 7265
rect 10137 7256 10149 7259
rect 9640 7228 10149 7256
rect 9640 7216 9646 7228
rect 10137 7225 10149 7228
rect 10183 7225 10195 7259
rect 10137 7219 10195 7225
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 11057 7259 11115 7265
rect 11057 7256 11069 7259
rect 10928 7228 11069 7256
rect 10928 7216 10934 7228
rect 11057 7225 11069 7228
rect 11103 7225 11115 7259
rect 11057 7219 11115 7225
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 12452 7256 12480 7287
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13964 7296 14013 7324
rect 13964 7284 13970 7296
rect 14001 7293 14013 7296
rect 14047 7324 14059 7327
rect 15378 7324 15384 7336
rect 14047 7296 15384 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 15378 7284 15384 7296
rect 15436 7324 15442 7336
rect 15436 7296 16436 7324
rect 15436 7284 15442 7296
rect 12216 7228 12480 7256
rect 14544 7259 14602 7265
rect 12216 7216 12222 7228
rect 14544 7225 14556 7259
rect 14590 7256 14602 7259
rect 15749 7259 15807 7265
rect 15749 7256 15761 7259
rect 14590 7228 15761 7256
rect 14590 7225 14602 7228
rect 14544 7219 14602 7225
rect 15749 7225 15761 7228
rect 15795 7225 15807 7259
rect 16408 7256 16436 7296
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 17000 7296 17325 7324
rect 17000 7284 17006 7296
rect 17313 7293 17325 7296
rect 17359 7324 17371 7327
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 17359 7296 17785 7324
rect 17359 7293 17371 7296
rect 17313 7287 17371 7293
rect 17773 7293 17785 7296
rect 17819 7324 17831 7327
rect 17862 7324 17868 7336
rect 17819 7296 17868 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 17862 7284 17868 7296
rect 17920 7284 17926 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7324 18110 7336
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18104 7296 18429 7324
rect 18104 7284 18110 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 16485 7259 16543 7265
rect 16485 7256 16497 7259
rect 16408 7228 16497 7256
rect 15749 7219 15807 7225
rect 16485 7225 16497 7228
rect 16531 7225 16543 7259
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 16485 7219 16543 7225
rect 16583 7228 17417 7256
rect 10318 7188 10324 7200
rect 8956 7160 10324 7188
rect 10318 7148 10324 7160
rect 10376 7148 10382 7200
rect 10410 7148 10416 7200
rect 10468 7188 10474 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10468 7160 10609 7188
rect 10468 7148 10474 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 11882 7188 11888 7200
rect 11843 7160 11888 7188
rect 10597 7151 10655 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 11977 7191 12035 7197
rect 11977 7157 11989 7191
rect 12023 7188 12035 7191
rect 12618 7188 12624 7200
rect 12023 7160 12624 7188
rect 12023 7157 12035 7160
rect 11977 7151 12035 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 15930 7188 15936 7200
rect 15887 7160 15936 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16114 7188 16120 7200
rect 16075 7160 16120 7188
rect 16114 7148 16120 7160
rect 16172 7148 16178 7200
rect 16206 7148 16212 7200
rect 16264 7188 16270 7200
rect 16583 7188 16611 7228
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 17405 7219 17463 7225
rect 16264 7160 16611 7188
rect 16264 7148 16270 7160
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 16724 7160 16957 7188
rect 16724 7148 16730 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 18230 7188 18236 7200
rect 18191 7160 18236 7188
rect 16945 7151 17003 7157
rect 18230 7148 18236 7160
rect 18288 7148 18294 7200
rect 1104 7098 18860 7120
rect 1104 7046 6912 7098
rect 6964 7046 6976 7098
rect 7028 7046 7040 7098
rect 7092 7046 7104 7098
rect 7156 7046 12843 7098
rect 12895 7046 12907 7098
rect 12959 7046 12971 7098
rect 13023 7046 13035 7098
rect 13087 7046 18860 7098
rect 18966 7052 18972 7064
rect 1104 7024 18860 7046
rect 18927 7024 18972 7052
rect 18966 7012 18972 7024
rect 19024 7012 19030 7064
rect 2682 6944 2688 6996
rect 2740 6984 2746 6996
rect 3050 6984 3056 6996
rect 2740 6956 3056 6984
rect 2740 6944 2746 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 9398 6984 9404 6996
rect 3436 6956 9404 6984
rect 1394 6876 1400 6928
rect 1452 6916 1458 6928
rect 3436 6916 3464 6956
rect 9398 6944 9404 6956
rect 9456 6984 9462 6996
rect 12342 6984 12348 6996
rect 9456 6956 12348 6984
rect 9456 6944 9462 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12676 6956 12909 6984
rect 12676 6944 12682 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 13357 6987 13415 6993
rect 13357 6953 13369 6987
rect 13403 6984 13415 6987
rect 13725 6987 13783 6993
rect 13725 6984 13737 6987
rect 13403 6956 13737 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 13725 6953 13737 6956
rect 13771 6953 13783 6987
rect 13725 6947 13783 6953
rect 14093 6987 14151 6993
rect 14093 6953 14105 6987
rect 14139 6984 14151 6987
rect 14366 6984 14372 6996
rect 14139 6956 14372 6984
rect 14139 6953 14151 6956
rect 14093 6947 14151 6953
rect 14366 6944 14372 6956
rect 14424 6984 14430 6996
rect 14550 6984 14556 6996
rect 14424 6956 14556 6984
rect 14424 6944 14430 6956
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14734 6984 14740 6996
rect 14695 6956 14740 6984
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 17313 6987 17371 6993
rect 17313 6984 17325 6987
rect 15988 6956 17325 6984
rect 15988 6944 15994 6956
rect 17313 6953 17325 6956
rect 17359 6953 17371 6987
rect 17313 6947 17371 6953
rect 1452 6888 3464 6916
rect 3513 6919 3571 6925
rect 1452 6876 1458 6888
rect 3513 6885 3525 6919
rect 3559 6916 3571 6919
rect 4798 6916 4804 6928
rect 3559 6888 4804 6916
rect 3559 6885 3571 6888
rect 3513 6879 3571 6885
rect 4798 6876 4804 6888
rect 4856 6876 4862 6928
rect 5442 6916 5448 6928
rect 5092 6888 5448 6916
rect 1848 6851 1906 6857
rect 1848 6817 1860 6851
rect 1894 6848 1906 6851
rect 3605 6851 3663 6857
rect 1894 6820 3556 6848
rect 1894 6817 1906 6820
rect 1848 6811 1906 6817
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 1581 6783 1639 6789
rect 1581 6780 1593 6783
rect 1268 6752 1593 6780
rect 1268 6740 1274 6752
rect 1581 6749 1593 6752
rect 1627 6749 1639 6783
rect 1581 6743 1639 6749
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3528 6780 3556 6820
rect 3605 6817 3617 6851
rect 3651 6848 3663 6851
rect 3651 6820 4016 6848
rect 3651 6817 3663 6820
rect 3605 6811 3663 6817
rect 3786 6780 3792 6792
rect 3528 6752 3792 6780
rect 3786 6740 3792 6752
rect 3844 6740 3850 6792
rect 3988 6780 4016 6820
rect 4246 6808 4252 6860
rect 4304 6848 4310 6860
rect 4433 6851 4491 6857
rect 4433 6848 4445 6851
rect 4304 6820 4445 6848
rect 4304 6808 4310 6820
rect 4433 6817 4445 6820
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6848 4583 6851
rect 5092 6848 5120 6888
rect 5442 6876 5448 6888
rect 5500 6916 5506 6928
rect 6641 6919 6699 6925
rect 6641 6916 6653 6919
rect 5500 6888 6653 6916
rect 5500 6876 5506 6888
rect 6641 6885 6653 6888
rect 6687 6916 6699 6919
rect 6730 6916 6736 6928
rect 6687 6888 6736 6916
rect 6687 6885 6699 6888
rect 6641 6879 6699 6885
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 10962 6916 10968 6928
rect 7085 6888 8248 6916
rect 4571 6820 5120 6848
rect 5160 6851 5218 6857
rect 4571 6817 4583 6820
rect 4525 6811 4583 6817
rect 5160 6817 5172 6851
rect 5206 6848 5218 6851
rect 6454 6848 6460 6860
rect 5206 6820 6460 6848
rect 5206 6817 5218 6820
rect 5160 6811 5218 6817
rect 6454 6808 6460 6820
rect 6512 6808 6518 6860
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7085 6848 7113 6888
rect 8018 6857 8024 6860
rect 6595 6820 7113 6848
rect 7193 6851 7251 6857
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7239 6820 7604 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 4338 6780 4344 6792
rect 3988 6752 4344 6780
rect 4338 6740 4344 6752
rect 4396 6740 4402 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6749 4675 6783
rect 4890 6780 4896 6792
rect 4851 6752 4896 6780
rect 4617 6743 4675 6749
rect 2590 6672 2596 6724
rect 2648 6712 2654 6724
rect 3145 6715 3203 6721
rect 3145 6712 3157 6715
rect 2648 6684 3157 6712
rect 2648 6672 2654 6684
rect 3145 6681 3157 6684
rect 3191 6681 3203 6715
rect 3436 6712 3464 6740
rect 3145 6675 3203 6681
rect 3252 6684 3464 6712
rect 3804 6712 3832 6740
rect 4632 6712 4660 6743
rect 4890 6740 4896 6752
rect 4948 6740 4954 6792
rect 6638 6740 6644 6792
rect 6696 6780 6702 6792
rect 7282 6780 7288 6792
rect 6696 6752 7144 6780
rect 7243 6752 7288 6780
rect 6696 6740 6702 6752
rect 3804 6684 4660 6712
rect 1394 6644 1400 6656
rect 1355 6616 1400 6644
rect 1394 6604 1400 6616
rect 1452 6604 1458 6656
rect 2682 6604 2688 6656
rect 2740 6644 2746 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2740 6616 2973 6644
rect 2740 6604 2746 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3252 6644 3280 6684
rect 5902 6672 5908 6724
rect 5960 6712 5966 6724
rect 6825 6715 6883 6721
rect 6825 6712 6837 6715
rect 5960 6684 6837 6712
rect 5960 6672 5966 6684
rect 6825 6681 6837 6684
rect 6871 6681 6883 6715
rect 7116 6712 7144 6752
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 7392 6712 7420 6743
rect 7116 6684 7420 6712
rect 6825 6675 6883 6681
rect 3108 6616 3280 6644
rect 3108 6604 3114 6616
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 4065 6647 4123 6653
rect 4065 6644 4077 6647
rect 3476 6616 4077 6644
rect 3476 6604 3482 6616
rect 4065 6613 4077 6616
rect 4111 6613 4123 6647
rect 4065 6607 4123 6613
rect 4338 6604 4344 6656
rect 4396 6644 4402 6656
rect 4614 6644 4620 6656
rect 4396 6616 4620 6644
rect 4396 6604 4402 6616
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5074 6604 5080 6656
rect 5132 6644 5138 6656
rect 6273 6647 6331 6653
rect 6273 6644 6285 6647
rect 5132 6616 6285 6644
rect 5132 6604 5138 6616
rect 6273 6613 6285 6616
rect 6319 6613 6331 6647
rect 6273 6607 6331 6613
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 7576 6644 7604 6820
rect 8012 6811 8024 6857
rect 8076 6848 8082 6860
rect 8220 6848 8248 6888
rect 10244 6888 10968 6916
rect 10244 6848 10272 6888
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11054 6876 11060 6928
rect 11112 6876 11118 6928
rect 11790 6876 11796 6928
rect 11848 6876 11854 6928
rect 12437 6919 12495 6925
rect 12437 6885 12449 6919
rect 12483 6916 12495 6919
rect 13538 6916 13544 6928
rect 12483 6888 13544 6916
rect 12483 6885 12495 6888
rect 12437 6879 12495 6885
rect 13538 6876 13544 6888
rect 13596 6916 13602 6928
rect 13814 6916 13820 6928
rect 13596 6888 13820 6916
rect 13596 6876 13602 6888
rect 13814 6876 13820 6888
rect 13872 6876 13878 6928
rect 14921 6919 14979 6925
rect 14921 6885 14933 6919
rect 14967 6916 14979 6919
rect 15010 6916 15016 6928
rect 14967 6888 15016 6916
rect 14967 6885 14979 6888
rect 14921 6879 14979 6885
rect 15010 6876 15016 6888
rect 15068 6876 15074 6928
rect 15470 6876 15476 6928
rect 15528 6876 15534 6928
rect 15654 6876 15660 6928
rect 15712 6925 15718 6928
rect 15712 6919 15776 6925
rect 15712 6885 15730 6919
rect 15764 6885 15776 6919
rect 17405 6919 17463 6925
rect 17405 6916 17417 6919
rect 15712 6879 15776 6885
rect 15856 6888 17417 6916
rect 15712 6876 15718 6879
rect 10410 6848 10416 6860
rect 8076 6820 8112 6848
rect 8220 6820 10272 6848
rect 10371 6820 10416 6848
rect 8018 6808 8024 6811
rect 8076 6808 8082 6820
rect 10410 6808 10416 6820
rect 10468 6808 10474 6860
rect 10502 6808 10508 6860
rect 10560 6848 10566 6860
rect 11072 6848 11100 6876
rect 11146 6857 11152 6860
rect 10560 6820 10605 6848
rect 10704 6820 11100 6848
rect 10560 6808 10566 6820
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9766 6780 9772 6792
rect 9727 6752 9772 6780
rect 9766 6740 9772 6752
rect 9824 6740 9830 6792
rect 10226 6740 10232 6792
rect 10284 6780 10290 6792
rect 10594 6780 10600 6792
rect 10284 6752 10600 6780
rect 10284 6740 10290 6752
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10704 6789 10732 6820
rect 11140 6811 11152 6857
rect 11204 6848 11210 6860
rect 11808 6848 11836 6876
rect 13262 6848 13268 6860
rect 11204 6820 11240 6848
rect 11808 6820 12664 6848
rect 13223 6820 13268 6848
rect 11146 6808 11152 6811
rect 11204 6808 11210 6820
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6749 10747 6783
rect 10870 6780 10876 6792
rect 10831 6752 10876 6780
rect 10689 6743 10747 6749
rect 10870 6740 10876 6752
rect 10928 6740 10934 6792
rect 12636 6789 12664 6820
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 15488 6848 15516 6876
rect 13372 6820 15516 6848
rect 12621 6783 12679 6789
rect 12621 6749 12633 6783
rect 12667 6780 12679 6783
rect 13372 6780 13400 6820
rect 15562 6808 15568 6860
rect 15620 6848 15626 6860
rect 15856 6848 15884 6888
rect 17405 6885 17417 6888
rect 17451 6885 17463 6919
rect 17405 6879 17463 6885
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6916 18199 6919
rect 18690 6916 18696 6928
rect 18187 6888 18696 6916
rect 18187 6885 18199 6888
rect 18141 6879 18199 6885
rect 18690 6876 18696 6888
rect 18748 6876 18754 6928
rect 15620 6820 15884 6848
rect 15620 6808 15626 6820
rect 16850 6808 16856 6860
rect 16908 6848 16914 6860
rect 18233 6851 18291 6857
rect 16908 6820 17908 6848
rect 16908 6808 16914 6820
rect 13538 6780 13544 6792
rect 12667 6752 13400 6780
rect 13451 6752 13544 6780
rect 12667 6749 12679 6752
rect 12621 6743 12679 6749
rect 13538 6740 13544 6752
rect 13596 6780 13602 6792
rect 13596 6752 13676 6780
rect 13596 6740 13602 6752
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 10502 6712 10508 6724
rect 9355 6684 10508 6712
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 13648 6712 13676 6752
rect 13906 6740 13912 6792
rect 13964 6780 13970 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 13964 6752 14197 6780
rect 13964 6740 13970 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 14185 6743 14243 6749
rect 14274 6740 14280 6792
rect 14332 6780 14338 6792
rect 14332 6752 14377 6780
rect 14332 6740 14338 6752
rect 14918 6740 14924 6792
rect 14976 6780 14982 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 14976 6752 15485 6780
rect 14976 6740 14982 6752
rect 15473 6749 15485 6752
rect 15519 6749 15531 6783
rect 15473 6743 15531 6749
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17310 6780 17316 6792
rect 16632 6752 17316 6780
rect 16632 6740 16638 6752
rect 17310 6740 17316 6752
rect 17368 6740 17374 6792
rect 17494 6780 17500 6792
rect 17455 6752 17500 6780
rect 17494 6740 17500 6752
rect 17552 6740 17558 6792
rect 15194 6712 15200 6724
rect 11808 6684 13400 6712
rect 13648 6684 15200 6712
rect 8110 6644 8116 6656
rect 6420 6616 6465 6644
rect 7576 6616 8116 6644
rect 6420 6604 6426 6616
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9398 6644 9404 6656
rect 9171 6616 9404 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6644 10103 6647
rect 11054 6644 11060 6656
rect 10091 6616 11060 6644
rect 10091 6613 10103 6616
rect 10045 6607 10103 6613
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11514 6604 11520 6656
rect 11572 6644 11578 6656
rect 11808 6644 11836 6684
rect 12250 6644 12256 6656
rect 11572 6616 11836 6644
rect 12211 6616 12256 6644
rect 11572 6604 11578 6616
rect 12250 6604 12256 6616
rect 12308 6604 12314 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12492 6616 12725 6644
rect 12492 6604 12498 6616
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 13372 6644 13400 6684
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 15378 6712 15384 6724
rect 15339 6684 15384 6712
rect 15378 6672 15384 6684
rect 15436 6672 15442 6724
rect 16758 6672 16764 6724
rect 16816 6712 16822 6724
rect 17773 6715 17831 6721
rect 17773 6712 17785 6715
rect 16816 6684 17785 6712
rect 16816 6672 16822 6684
rect 17773 6681 17785 6684
rect 17819 6681 17831 6715
rect 17880 6712 17908 6820
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 18279 6820 18460 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18340 6712 18368 6743
rect 17880 6684 18368 6712
rect 17773 6675 17831 6681
rect 14550 6644 14556 6656
rect 13372 6616 14556 6644
rect 12713 6607 12771 6613
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 15105 6647 15163 6653
rect 15105 6613 15117 6647
rect 15151 6644 15163 6647
rect 15286 6644 15292 6656
rect 15151 6616 15292 6644
rect 15151 6613 15163 6616
rect 15105 6607 15163 6613
rect 15286 6604 15292 6616
rect 15344 6644 15350 6656
rect 16574 6644 16580 6656
rect 15344 6616 16580 6644
rect 15344 6604 15350 6616
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16850 6644 16856 6656
rect 16811 6616 16856 6644
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17000 6616 17045 6644
rect 17000 6604 17006 6616
rect 17310 6604 17316 6656
rect 17368 6644 17374 6656
rect 18432 6644 18460 6820
rect 17368 6616 18460 6644
rect 17368 6604 17374 6616
rect 1104 6554 18860 6576
rect 1104 6502 3947 6554
rect 3999 6502 4011 6554
rect 4063 6502 4075 6554
rect 4127 6502 4139 6554
rect 4191 6502 9878 6554
rect 9930 6502 9942 6554
rect 9994 6502 10006 6554
rect 10058 6502 10070 6554
rect 10122 6502 15808 6554
rect 15860 6502 15872 6554
rect 15924 6502 15936 6554
rect 15988 6502 16000 6554
rect 16052 6502 18860 6554
rect 1104 6480 18860 6502
rect 3326 6440 3332 6452
rect 2983 6412 3332 6440
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 2682 6304 2688 6316
rect 2464 6276 2688 6304
rect 2464 6264 2470 6276
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 2983 6313 3011 6412
rect 3326 6400 3332 6412
rect 3384 6400 3390 6452
rect 3694 6400 3700 6452
rect 3752 6440 3758 6452
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 3752 6412 4629 6440
rect 3752 6400 3758 6412
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 6454 6440 6460 6452
rect 6415 6412 6460 6440
rect 4617 6403 4675 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6730 6400 6736 6452
rect 6788 6440 6794 6452
rect 7742 6440 7748 6452
rect 6788 6412 7748 6440
rect 6788 6400 6794 6412
rect 7742 6400 7748 6412
rect 7800 6440 7806 6452
rect 9861 6443 9919 6449
rect 7800 6412 8432 6440
rect 7800 6400 7806 6412
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 4798 6304 4804 6316
rect 4759 6276 4804 6304
rect 2961 6267 3019 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 4890 6264 4896 6316
rect 4948 6304 4954 6316
rect 8404 6313 8432 6412
rect 9861 6409 9873 6443
rect 9907 6440 9919 6443
rect 10410 6440 10416 6452
rect 9907 6412 10416 6440
rect 9907 6409 9919 6412
rect 9861 6403 9919 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 11882 6440 11888 6452
rect 11563 6412 11888 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12066 6400 12072 6452
rect 12124 6440 12130 6452
rect 12124 6412 12388 6440
rect 12124 6400 12130 6412
rect 12250 6372 12256 6384
rect 10520 6344 12256 6372
rect 10520 6313 10548 6344
rect 12250 6332 12256 6344
rect 12308 6332 12314 6384
rect 12360 6372 12388 6412
rect 12434 6400 12440 6452
rect 12492 6440 12498 6452
rect 15657 6443 15715 6449
rect 15657 6440 15669 6443
rect 12492 6412 15669 6440
rect 12492 6400 12498 6412
rect 15657 6409 15669 6412
rect 15703 6440 15715 6443
rect 17494 6440 17500 6452
rect 15703 6412 17500 6440
rect 15703 6409 15715 6412
rect 15657 6403 15715 6409
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 13078 6372 13084 6384
rect 12360 6344 13084 6372
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 15194 6372 15200 6384
rect 15155 6344 15200 6372
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 15286 6332 15292 6384
rect 15344 6372 15350 6384
rect 15381 6375 15439 6381
rect 15381 6372 15393 6375
rect 15344 6344 15393 6372
rect 15344 6332 15350 6344
rect 15381 6341 15393 6344
rect 15427 6341 15439 6375
rect 16390 6372 16396 6384
rect 16303 6344 16396 6372
rect 15381 6335 15439 6341
rect 5077 6307 5135 6313
rect 5077 6304 5089 6307
rect 4948 6276 5089 6304
rect 4948 6264 4954 6276
rect 5077 6273 5089 6276
rect 5123 6273 5135 6307
rect 8389 6307 8447 6313
rect 5077 6267 5135 6273
rect 6564 6276 6960 6304
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2501 6239 2559 6245
rect 1719 6208 2452 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 1946 6168 1952 6180
rect 1627 6140 1952 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 1946 6128 1952 6140
rect 2004 6128 2010 6180
rect 2424 6168 2452 6208
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 2590 6236 2596 6248
rect 2547 6208 2596 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 2590 6196 2596 6208
rect 2648 6196 2654 6248
rect 2700 6236 2728 6264
rect 3217 6239 3275 6245
rect 3217 6236 3229 6239
rect 2700 6208 3229 6236
rect 3217 6205 3229 6208
rect 3263 6205 3275 6239
rect 3217 6199 3275 6205
rect 4433 6239 4491 6245
rect 4433 6205 4445 6239
rect 4479 6236 4491 6239
rect 4982 6236 4988 6248
rect 4479 6208 4988 6236
rect 4479 6205 4491 6208
rect 4433 6199 4491 6205
rect 4982 6196 4988 6208
rect 5040 6196 5046 6248
rect 6564 6245 6592 6276
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 5276 6208 6561 6236
rect 5276 6168 5304 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 6730 6196 6736 6248
rect 6788 6236 6794 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6788 6208 6837 6236
rect 6788 6196 6794 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 6932 6236 6960 6276
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6273 10563 6307
rect 10505 6267 10563 6273
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11333 6307 11391 6313
rect 11333 6304 11345 6307
rect 11204 6276 11345 6304
rect 11204 6264 11210 6276
rect 11333 6273 11345 6276
rect 11379 6304 11391 6307
rect 11882 6304 11888 6316
rect 11379 6276 11888 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 11940 6276 12173 6304
rect 11940 6264 11946 6276
rect 12161 6273 12173 6276
rect 12207 6304 12219 6307
rect 13538 6304 13544 6316
rect 12207 6276 13544 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6304 13691 6307
rect 13679 6276 13952 6304
rect 13679 6273 13691 6276
rect 13633 6267 13691 6273
rect 11057 6239 11115 6245
rect 6932 6208 11008 6236
rect 6825 6199 6883 6205
rect 2424 6140 5304 6168
rect 5344 6171 5402 6177
rect 5344 6137 5356 6171
rect 5390 6168 5402 6171
rect 6638 6168 6644 6180
rect 5390 6140 6644 6168
rect 5390 6137 5402 6140
rect 5344 6131 5402 6137
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 7092 6171 7150 6177
rect 7092 6137 7104 6171
rect 7138 6168 7150 6171
rect 8294 6168 8300 6180
rect 7138 6140 8300 6168
rect 7138 6137 7150 6140
rect 7092 6131 7150 6137
rect 8294 6128 8300 6140
rect 8352 6128 8358 6180
rect 8656 6171 8714 6177
rect 8656 6137 8668 6171
rect 8702 6168 8714 6171
rect 9398 6168 9404 6180
rect 8702 6140 9404 6168
rect 8702 6137 8714 6140
rect 8656 6131 8714 6137
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 10229 6171 10287 6177
rect 10229 6137 10241 6171
rect 10275 6168 10287 6171
rect 10980 6168 11008 6208
rect 11057 6205 11069 6239
rect 11103 6236 11115 6239
rect 11514 6236 11520 6248
rect 11103 6208 11520 6236
rect 11103 6205 11115 6208
rect 11057 6199 11115 6205
rect 11514 6196 11520 6208
rect 11572 6196 11578 6248
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 12308 6208 12449 6236
rect 12308 6196 12314 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12802 6236 12808 6248
rect 12763 6208 12808 6236
rect 12437 6199 12495 6205
rect 12802 6196 12808 6208
rect 12860 6236 12866 6248
rect 13446 6236 13452 6248
rect 12860 6208 13452 6236
rect 12860 6196 12866 6208
rect 13446 6196 13452 6208
rect 13504 6196 13510 6248
rect 13722 6196 13728 6248
rect 13780 6236 13786 6248
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13780 6208 13829 6236
rect 13780 6196 13786 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13924 6236 13952 6276
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16316 6313 16344 6344
rect 16390 6332 16396 6344
rect 16448 6372 16454 6384
rect 16448 6344 17172 6372
rect 16448 6332 16454 6344
rect 16209 6307 16267 6313
rect 16209 6304 16221 6307
rect 16172 6276 16221 6304
rect 16172 6264 16178 6276
rect 16209 6273 16221 6276
rect 16255 6273 16267 6307
rect 16209 6267 16267 6273
rect 16301 6307 16359 6313
rect 16301 6273 16313 6307
rect 16347 6273 16359 6307
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 16301 6267 16359 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17144 6313 17172 6344
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6273 17187 6307
rect 17129 6267 17187 6273
rect 13924 6208 14127 6236
rect 13817 6199 13875 6205
rect 11149 6171 11207 6177
rect 11149 6168 11161 6171
rect 10275 6140 10732 6168
rect 10980 6140 11161 6168
rect 10275 6137 10287 6140
rect 10229 6131 10287 6137
rect 1854 6100 1860 6112
rect 1815 6072 1860 6100
rect 1854 6060 1860 6072
rect 1912 6060 1918 6112
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2593 6103 2651 6109
rect 2593 6069 2605 6103
rect 2639 6100 2651 6103
rect 3418 6100 3424 6112
rect 2639 6072 3424 6100
rect 2639 6069 2651 6072
rect 2593 6063 2651 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5718 6100 5724 6112
rect 4948 6072 5724 6100
rect 4948 6060 4954 6072
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 6656 6100 6684 6128
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 6656 6072 8217 6100
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9769 6103 9827 6109
rect 9769 6100 9781 6103
rect 9272 6072 9781 6100
rect 9272 6060 9278 6072
rect 9769 6069 9781 6072
rect 9815 6069 9827 6103
rect 10318 6100 10324 6112
rect 10279 6072 10324 6100
rect 9769 6063 9827 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10704 6109 10732 6140
rect 11149 6137 11161 6140
rect 11195 6168 11207 6171
rect 11790 6168 11796 6180
rect 11195 6140 11796 6168
rect 11195 6137 11207 6140
rect 11149 6131 11207 6137
rect 11790 6128 11796 6140
rect 11848 6128 11854 6180
rect 11977 6171 12035 6177
rect 11977 6137 11989 6171
rect 12023 6168 12035 6171
rect 12023 6140 13032 6168
rect 12023 6137 12035 6140
rect 11977 6131 12035 6137
rect 10689 6103 10747 6109
rect 10689 6069 10701 6103
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 13004 6109 13032 6140
rect 13078 6128 13084 6180
rect 13136 6128 13142 6180
rect 14099 6177 14127 6208
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 16942 6236 16948 6248
rect 14608 6208 16804 6236
rect 16903 6208 16948 6236
rect 14608 6196 14614 6208
rect 14084 6171 14142 6177
rect 14084 6137 14096 6171
rect 14130 6168 14142 6171
rect 14274 6168 14280 6180
rect 14130 6140 14280 6168
rect 14130 6137 14142 6140
rect 14084 6131 14142 6137
rect 14274 6128 14280 6140
rect 14332 6128 14338 6180
rect 14918 6128 14924 6180
rect 14976 6168 14982 6180
rect 15194 6168 15200 6180
rect 14976 6140 15200 6168
rect 14976 6128 14982 6140
rect 15194 6128 15200 6140
rect 15252 6128 15258 6180
rect 16117 6171 16175 6177
rect 16117 6137 16129 6171
rect 16163 6168 16175 6171
rect 16666 6168 16672 6180
rect 16163 6140 16672 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 16666 6128 16672 6140
rect 16724 6128 16730 6180
rect 16776 6168 16804 6208
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17589 6239 17647 6245
rect 17589 6236 17601 6239
rect 17420 6208 17601 6236
rect 17420 6177 17448 6208
rect 17589 6205 17601 6208
rect 17635 6205 17647 6239
rect 17589 6199 17647 6205
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 17920 6208 18061 6236
rect 17920 6196 17926 6208
rect 18049 6205 18061 6208
rect 18095 6236 18107 6239
rect 18417 6239 18475 6245
rect 18417 6236 18429 6239
rect 18095 6208 18429 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18417 6205 18429 6208
rect 18463 6205 18475 6239
rect 18417 6199 18475 6205
rect 17405 6171 17463 6177
rect 17405 6168 17417 6171
rect 16776 6140 17417 6168
rect 17405 6137 17417 6140
rect 17451 6137 17463 6171
rect 17405 6131 17463 6137
rect 11885 6103 11943 6109
rect 11885 6100 11897 6103
rect 11480 6072 11897 6100
rect 11480 6060 11486 6072
rect 11885 6069 11897 6072
rect 11931 6069 11943 6103
rect 11885 6063 11943 6069
rect 12989 6103 13047 6109
rect 12989 6069 13001 6103
rect 13035 6069 13047 6103
rect 13096 6100 13124 6128
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 13096 6072 13369 6100
rect 12989 6063 13047 6069
rect 13357 6069 13369 6072
rect 13403 6100 13415 6103
rect 14642 6100 14648 6112
rect 13403 6072 14648 6100
rect 13403 6069 13415 6072
rect 13357 6063 13415 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15746 6100 15752 6112
rect 15707 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16206 6060 16212 6112
rect 16264 6100 16270 6112
rect 16577 6103 16635 6109
rect 16577 6100 16589 6103
rect 16264 6072 16589 6100
rect 16264 6060 16270 6072
rect 16577 6069 16589 6072
rect 16623 6069 16635 6103
rect 17770 6100 17776 6112
rect 17731 6072 17776 6100
rect 16577 6063 16635 6069
rect 17770 6060 17776 6072
rect 17828 6060 17834 6112
rect 18230 6100 18236 6112
rect 18191 6072 18236 6100
rect 18230 6060 18236 6072
rect 18288 6060 18294 6112
rect 1104 6010 18860 6032
rect 1104 5958 6912 6010
rect 6964 5958 6976 6010
rect 7028 5958 7040 6010
rect 7092 5958 7104 6010
rect 7156 5958 12843 6010
rect 12895 5958 12907 6010
rect 12959 5958 12971 6010
rect 13023 5958 13035 6010
rect 13087 5958 18860 6010
rect 1104 5936 18860 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 1995 5868 2329 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 3145 5899 3203 5905
rect 3145 5896 3157 5899
rect 2317 5859 2375 5865
rect 2884 5868 3157 5896
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 1872 5624 1900 5723
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 2648 5732 2697 5760
rect 2648 5720 2654 5732
rect 2685 5729 2697 5732
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2406 5692 2412 5704
rect 2179 5664 2412 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2498 5652 2504 5704
rect 2556 5692 2562 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2556 5664 2789 5692
rect 2556 5652 2562 5664
rect 2777 5661 2789 5664
rect 2823 5661 2835 5695
rect 2777 5655 2835 5661
rect 2884 5624 2912 5868
rect 3145 5865 3157 5868
rect 3191 5865 3203 5899
rect 5902 5896 5908 5908
rect 5863 5868 5908 5896
rect 3145 5859 3203 5865
rect 5902 5856 5908 5868
rect 5960 5856 5966 5908
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 6365 5899 6423 5905
rect 6365 5896 6377 5899
rect 6043 5868 6377 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 6365 5865 6377 5868
rect 6411 5865 6423 5899
rect 6365 5859 6423 5865
rect 6472 5868 7052 5896
rect 3510 5828 3516 5840
rect 3471 5800 3516 5828
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 5350 5788 5356 5840
rect 5408 5828 5414 5840
rect 6472 5828 6500 5868
rect 5408 5800 6500 5828
rect 6825 5831 6883 5837
rect 5408 5788 5414 5800
rect 6825 5797 6837 5831
rect 6871 5828 6883 5831
rect 6914 5828 6920 5840
rect 6871 5800 6920 5828
rect 6871 5797 6883 5800
rect 6825 5791 6883 5797
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7024 5828 7052 5868
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 7377 5899 7435 5905
rect 7377 5896 7389 5899
rect 7340 5868 7389 5896
rect 7340 5856 7346 5868
rect 7377 5865 7389 5868
rect 7423 5865 7435 5899
rect 7377 5859 7435 5865
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 8168 5868 8217 5896
rect 8168 5856 8174 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 8205 5859 8263 5865
rect 9122 5856 9128 5908
rect 9180 5896 9186 5908
rect 10226 5896 10232 5908
rect 9180 5868 10232 5896
rect 9180 5856 9186 5868
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 10318 5856 10324 5908
rect 10376 5896 10382 5908
rect 11241 5899 11299 5905
rect 11241 5896 11253 5899
rect 10376 5868 11253 5896
rect 10376 5856 10382 5868
rect 11241 5865 11253 5868
rect 11287 5865 11299 5899
rect 11241 5859 11299 5865
rect 11422 5856 11428 5908
rect 11480 5896 11486 5908
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 11480 5868 12081 5896
rect 11480 5856 11486 5868
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13320 5868 13737 5896
rect 13320 5856 13326 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 14093 5899 14151 5905
rect 14093 5865 14105 5899
rect 14139 5896 14151 5899
rect 14553 5899 14611 5905
rect 14553 5896 14565 5899
rect 14139 5868 14565 5896
rect 14139 5865 14151 5868
rect 14093 5859 14151 5865
rect 14553 5865 14565 5868
rect 14599 5865 14611 5899
rect 14553 5859 14611 5865
rect 14921 5899 14979 5905
rect 14921 5865 14933 5899
rect 14967 5896 14979 5899
rect 15470 5896 15476 5908
rect 14967 5868 15476 5896
rect 14967 5865 14979 5868
rect 14921 5859 14979 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15746 5896 15752 5908
rect 15707 5868 15752 5896
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 8665 5831 8723 5837
rect 8665 5828 8677 5831
rect 7024 5800 7880 5828
rect 4338 5769 4344 5772
rect 4332 5760 4344 5769
rect 4299 5732 4344 5760
rect 4332 5723 4344 5732
rect 4338 5720 4344 5723
rect 4396 5720 4402 5772
rect 6733 5763 6791 5769
rect 6733 5729 6745 5763
rect 6779 5760 6791 5763
rect 7650 5760 7656 5772
rect 6779 5732 7656 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 7745 5763 7803 5769
rect 7745 5729 7757 5763
rect 7791 5729 7803 5763
rect 7852 5760 7880 5800
rect 8404 5800 8677 5828
rect 8404 5760 8432 5800
rect 8665 5797 8677 5800
rect 8711 5828 8723 5831
rect 9033 5831 9091 5837
rect 9033 5828 9045 5831
rect 8711 5800 9045 5828
rect 8711 5797 8723 5800
rect 8665 5791 8723 5797
rect 9033 5797 9045 5800
rect 9079 5828 9091 5831
rect 10410 5828 10416 5840
rect 9079 5800 10416 5828
rect 9079 5797 9091 5800
rect 9033 5791 9091 5797
rect 10410 5788 10416 5800
rect 10468 5788 10474 5840
rect 10594 5788 10600 5840
rect 10652 5828 10658 5840
rect 13538 5828 13544 5840
rect 10652 5800 13544 5828
rect 10652 5788 10658 5800
rect 13538 5788 13544 5800
rect 13596 5788 13602 5840
rect 13906 5788 13912 5840
rect 13964 5828 13970 5840
rect 14645 5831 14703 5837
rect 14645 5828 14657 5831
rect 13964 5800 14657 5828
rect 13964 5788 13970 5800
rect 14645 5797 14657 5800
rect 14691 5828 14703 5831
rect 15562 5828 15568 5840
rect 14691 5800 15568 5828
rect 14691 5797 14703 5800
rect 14645 5791 14703 5797
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 15657 5831 15715 5837
rect 15657 5797 15669 5831
rect 15703 5828 15715 5831
rect 16206 5828 16212 5840
rect 15703 5800 16212 5828
rect 15703 5797 15715 5800
rect 15657 5791 15715 5797
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 16660 5831 16718 5837
rect 16660 5797 16672 5831
rect 16706 5828 16718 5831
rect 16850 5828 16856 5840
rect 16706 5800 16856 5828
rect 16706 5797 16718 5800
rect 16660 5791 16718 5797
rect 16850 5788 16856 5800
rect 16908 5788 16914 5840
rect 17310 5788 17316 5840
rect 17368 5828 17374 5840
rect 17368 5800 18276 5828
rect 17368 5788 17374 5800
rect 8570 5760 8576 5772
rect 7852 5732 8432 5760
rect 8531 5732 8576 5760
rect 7745 5723 7803 5729
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5661 3019 5695
rect 3602 5692 3608 5704
rect 3563 5664 3608 5692
rect 2961 5655 3019 5661
rect 1872 5596 2912 5624
rect 2976 5624 3004 5655
rect 3602 5652 3608 5664
rect 3660 5652 3666 5704
rect 3786 5692 3792 5704
rect 3747 5664 3792 5692
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5661 4123 5695
rect 4065 5655 4123 5661
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5692 6239 5695
rect 6454 5692 6460 5704
rect 6227 5664 6460 5692
rect 6227 5661 6239 5664
rect 6181 5655 6239 5661
rect 3804 5624 3832 5652
rect 2976 5596 3832 5624
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 4080 5556 4108 5655
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6917 5695 6975 5701
rect 6917 5692 6929 5695
rect 6696 5664 6929 5692
rect 6696 5652 6702 5664
rect 6917 5661 6929 5664
rect 6963 5661 6975 5695
rect 6917 5655 6975 5661
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5692 7343 5695
rect 7374 5692 7380 5704
rect 7331 5664 7380 5692
rect 7331 5661 7343 5664
rect 7285 5655 7343 5661
rect 7374 5652 7380 5664
rect 7432 5692 7438 5704
rect 7760 5692 7788 5723
rect 8570 5720 8576 5732
rect 8628 5720 8634 5772
rect 10036 5763 10094 5769
rect 10036 5729 10048 5763
rect 10082 5760 10094 5763
rect 10318 5760 10324 5772
rect 10082 5732 10324 5760
rect 10082 5729 10094 5732
rect 10036 5723 10094 5729
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 11609 5763 11667 5769
rect 11609 5729 11621 5763
rect 11655 5760 11667 5763
rect 12342 5760 12348 5772
rect 11655 5732 12348 5760
rect 11655 5729 11667 5732
rect 11609 5723 11667 5729
rect 7432 5664 7788 5692
rect 7432 5652 7438 5664
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8021 5695 8079 5701
rect 7892 5664 7937 5692
rect 7892 5652 7898 5664
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 8294 5692 8300 5704
rect 8067 5664 8300 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8757 5695 8815 5701
rect 8757 5661 8769 5695
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 5074 5584 5080 5636
rect 5132 5624 5138 5636
rect 5537 5627 5595 5633
rect 5537 5624 5549 5627
rect 5132 5596 5549 5624
rect 5132 5584 5138 5596
rect 5537 5593 5549 5596
rect 5583 5593 5595 5627
rect 8312 5624 8340 5652
rect 8772 5624 8800 5655
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9217 5695 9275 5701
rect 9217 5692 9229 5695
rect 8904 5664 9229 5692
rect 8904 5652 8910 5664
rect 9217 5661 9229 5664
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 9769 5695 9827 5701
rect 9769 5692 9781 5695
rect 9732 5664 9781 5692
rect 9732 5652 9738 5664
rect 9769 5661 9781 5664
rect 9815 5661 9827 5695
rect 9769 5655 9827 5661
rect 11238 5652 11244 5704
rect 11296 5692 11302 5704
rect 11624 5692 11652 5723
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 12437 5763 12495 5769
rect 12437 5729 12449 5763
rect 12483 5760 12495 5763
rect 12526 5760 12532 5772
rect 12483 5732 12532 5760
rect 12483 5729 12495 5732
rect 12437 5723 12495 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12710 5720 12716 5772
rect 12768 5760 12774 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12768 5732 12909 5760
rect 12768 5720 12774 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 12989 5763 13047 5769
rect 12989 5729 13001 5763
rect 13035 5760 13047 5763
rect 13556 5760 13584 5788
rect 14185 5763 14243 5769
rect 14185 5760 14197 5763
rect 13035 5732 13400 5760
rect 13556 5732 14197 5760
rect 13035 5729 13047 5732
rect 12989 5723 13047 5729
rect 11296 5664 11652 5692
rect 11701 5695 11759 5701
rect 11296 5652 11302 5664
rect 11701 5661 11713 5695
rect 11747 5661 11759 5695
rect 11882 5692 11888 5704
rect 11843 5664 11888 5692
rect 11701 5655 11759 5661
rect 8312 5596 8800 5624
rect 5537 5587 5595 5593
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 9180 5596 9413 5624
rect 9180 5584 9186 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 11422 5584 11428 5636
rect 11480 5624 11486 5636
rect 11716 5624 11744 5655
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 12158 5652 12164 5704
rect 12216 5652 12222 5704
rect 13170 5692 13176 5704
rect 13131 5664 13176 5692
rect 13170 5652 13176 5664
rect 13228 5652 13234 5704
rect 13372 5692 13400 5732
rect 14185 5729 14197 5732
rect 14231 5729 14243 5763
rect 14185 5723 14243 5729
rect 14366 5720 14372 5772
rect 14424 5760 14430 5772
rect 14424 5732 14688 5760
rect 14424 5720 14430 5732
rect 13906 5692 13912 5704
rect 13372 5664 13912 5692
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 14660 5692 14688 5732
rect 14826 5720 14832 5772
rect 14884 5760 14890 5772
rect 15013 5763 15071 5769
rect 15013 5760 15025 5763
rect 14884 5732 15025 5760
rect 14884 5720 14890 5732
rect 15013 5729 15025 5732
rect 15059 5729 15071 5763
rect 15013 5723 15071 5729
rect 14734 5692 14740 5704
rect 14332 5664 14377 5692
rect 14660 5664 14740 5692
rect 14332 5652 14338 5664
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 15028 5692 15056 5723
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 16393 5763 16451 5769
rect 16393 5760 16405 5763
rect 15252 5732 16405 5760
rect 15252 5720 15258 5732
rect 16393 5729 16405 5732
rect 16439 5729 16451 5763
rect 17218 5760 17224 5772
rect 16393 5723 16451 5729
rect 16500 5732 17224 5760
rect 15562 5692 15568 5704
rect 15028 5664 15568 5692
rect 15562 5652 15568 5664
rect 15620 5652 15626 5704
rect 15654 5652 15660 5704
rect 15712 5692 15718 5704
rect 15841 5695 15899 5701
rect 15841 5692 15853 5695
rect 15712 5664 15853 5692
rect 15712 5652 15718 5664
rect 15841 5661 15853 5664
rect 15887 5661 15899 5695
rect 16114 5692 16120 5704
rect 16075 5664 16120 5692
rect 15841 5655 15899 5661
rect 16114 5652 16120 5664
rect 16172 5652 16178 5704
rect 16500 5692 16528 5732
rect 17218 5720 17224 5732
rect 17276 5720 17282 5772
rect 17494 5720 17500 5772
rect 17552 5760 17558 5772
rect 18248 5769 18276 5800
rect 17865 5763 17923 5769
rect 17865 5760 17877 5763
rect 17552 5732 17877 5760
rect 17552 5720 17558 5732
rect 17865 5729 17877 5732
rect 17911 5729 17923 5763
rect 17865 5723 17923 5729
rect 18233 5763 18291 5769
rect 18233 5729 18245 5763
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 16224 5664 16528 5692
rect 12176 5624 12204 5652
rect 13357 5627 13415 5633
rect 13357 5624 13369 5627
rect 11480 5596 13369 5624
rect 11480 5584 11486 5596
rect 13357 5593 13369 5596
rect 13403 5593 13415 5627
rect 13357 5587 13415 5593
rect 14553 5627 14611 5633
rect 14553 5593 14565 5627
rect 14599 5624 14611 5627
rect 16224 5624 16252 5664
rect 14599 5596 16252 5624
rect 14599 5593 14611 5596
rect 14553 5587 14611 5593
rect 4798 5556 4804 5568
rect 3384 5528 4804 5556
rect 3384 5516 3390 5528
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 5442 5556 5448 5568
rect 5403 5528 5448 5556
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 10410 5556 10416 5568
rect 6604 5528 10416 5556
rect 6604 5516 6610 5528
rect 10410 5516 10416 5528
rect 10468 5516 10474 5568
rect 11149 5559 11207 5565
rect 11149 5525 11161 5559
rect 11195 5556 11207 5559
rect 11238 5556 11244 5568
rect 11195 5528 11244 5556
rect 11195 5525 11207 5528
rect 11149 5519 11207 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 12250 5556 12256 5568
rect 12211 5528 12256 5556
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12526 5556 12532 5568
rect 12487 5528 12532 5556
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 17770 5556 17776 5568
rect 17731 5528 17776 5556
rect 17770 5516 17776 5528
rect 17828 5516 17834 5568
rect 18046 5556 18052 5568
rect 18007 5528 18052 5556
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 3947 5466
rect 3999 5414 4011 5466
rect 4063 5414 4075 5466
rect 4127 5414 4139 5466
rect 4191 5414 9878 5466
rect 9930 5414 9942 5466
rect 9994 5414 10006 5466
rect 10058 5414 10070 5466
rect 10122 5414 15808 5466
rect 15860 5414 15872 5466
rect 15924 5414 15936 5466
rect 15988 5414 16000 5466
rect 16052 5414 18860 5466
rect 1104 5392 18860 5414
rect 2498 5312 2504 5364
rect 2556 5352 2562 5364
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2556 5324 2605 5352
rect 2556 5312 2562 5324
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 3421 5355 3479 5361
rect 3421 5321 3433 5355
rect 3467 5352 3479 5355
rect 3602 5352 3608 5364
rect 3467 5324 3608 5352
rect 3467 5321 3479 5324
rect 3421 5315 3479 5321
rect 3602 5312 3608 5324
rect 3660 5312 3666 5364
rect 4338 5352 4344 5364
rect 4264 5324 4344 5352
rect 4264 5284 4292 5324
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 6178 5352 6184 5364
rect 4580 5324 6184 5352
rect 4580 5312 4586 5324
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6914 5352 6920 5364
rect 6875 5324 6920 5352
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 7745 5355 7803 5361
rect 7745 5352 7757 5355
rect 7708 5324 7757 5352
rect 7708 5312 7714 5324
rect 7745 5321 7757 5324
rect 7791 5321 7803 5355
rect 10318 5352 10324 5364
rect 10231 5324 10324 5352
rect 7745 5315 7803 5321
rect 10318 5312 10324 5324
rect 10376 5352 10382 5364
rect 11974 5352 11980 5364
rect 10376 5324 11980 5352
rect 10376 5312 10382 5324
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12342 5312 12348 5364
rect 12400 5352 12406 5364
rect 13906 5352 13912 5364
rect 12400 5324 13492 5352
rect 13867 5324 13912 5352
rect 12400 5312 12406 5324
rect 4430 5284 4436 5296
rect 2424 5256 4292 5284
rect 4391 5256 4436 5284
rect 1486 5176 1492 5228
rect 1544 5216 1550 5228
rect 2424 5225 2452 5256
rect 4430 5244 4436 5256
rect 4488 5244 4494 5296
rect 6638 5244 6644 5296
rect 6696 5244 6702 5296
rect 2225 5219 2283 5225
rect 2225 5216 2237 5219
rect 1544 5188 2237 5216
rect 1544 5176 1550 5188
rect 2225 5185 2237 5188
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2409 5219 2467 5225
rect 2409 5185 2421 5219
rect 2455 5185 2467 5219
rect 3234 5216 3240 5228
rect 3147 5188 3240 5216
rect 2409 5179 2467 5185
rect 3234 5176 3240 5188
rect 3292 5216 3298 5228
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3292 5188 3985 5216
rect 3292 5176 3298 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 6656 5216 6684 5244
rect 7374 5216 7380 5228
rect 6656 5188 6776 5216
rect 7335 5188 7380 5216
rect 3973 5179 4031 5185
rect 1394 5148 1400 5160
rect 1355 5120 1400 5148
rect 1394 5108 1400 5120
rect 1452 5108 1458 5160
rect 2130 5148 2136 5160
rect 2091 5120 2136 5148
rect 2130 5108 2136 5120
rect 2188 5108 2194 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 3326 5148 3332 5160
rect 2924 5120 3332 5148
rect 2924 5108 2930 5120
rect 3326 5108 3332 5120
rect 3384 5148 3390 5160
rect 3789 5151 3847 5157
rect 3789 5148 3801 5151
rect 3384 5120 3801 5148
rect 3384 5108 3390 5120
rect 3789 5117 3801 5120
rect 3835 5148 3847 5151
rect 4062 5148 4068 5160
rect 3835 5120 4068 5148
rect 3835 5117 3847 5120
rect 3789 5111 3847 5117
rect 4062 5108 4068 5120
rect 4120 5108 4126 5160
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5148 4307 5151
rect 4614 5148 4620 5160
rect 4295 5120 4620 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4724 5080 4752 5111
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 4976 5151 5034 5157
rect 4976 5117 4988 5151
rect 5022 5148 5034 5151
rect 5442 5148 5448 5160
rect 5022 5120 5448 5148
rect 5022 5117 5034 5120
rect 4976 5111 5034 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 6362 5148 6368 5160
rect 6323 5120 6368 5148
rect 6362 5108 6368 5120
rect 6420 5108 6426 5160
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 4212 5052 4752 5080
rect 5460 5080 5488 5108
rect 5626 5080 5632 5092
rect 5460 5052 5632 5080
rect 4212 5040 4218 5052
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 6656 5080 6684 5111
rect 6196 5052 6684 5080
rect 6748 5080 6776 5188
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 8294 5216 8300 5228
rect 7607 5188 8300 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 10870 5216 10876 5228
rect 10428 5188 10876 5216
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7340 5120 8217 5148
rect 7340 5108 7346 5120
rect 8205 5117 8217 5120
rect 8251 5148 8263 5151
rect 8846 5148 8852 5160
rect 8251 5120 8852 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 9214 5157 9220 5160
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5117 8999 5151
rect 9208 5148 9220 5157
rect 9175 5120 9220 5148
rect 8941 5111 8999 5117
rect 9208 5111 9220 5120
rect 9272 5148 9278 5160
rect 9582 5148 9588 5160
rect 9272 5120 9588 5148
rect 6748 5052 7328 5080
rect 6196 5024 6224 5052
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 5012 1823 5015
rect 1946 5012 1952 5024
rect 1811 4984 1952 5012
rect 1811 4981 1823 4984
rect 1765 4975 1823 4981
rect 1946 4972 1952 4984
rect 2004 4972 2010 5024
rect 2682 4972 2688 5024
rect 2740 5012 2746 5024
rect 2961 5015 3019 5021
rect 2961 5012 2973 5015
rect 2740 4984 2973 5012
rect 2740 4972 2746 4984
rect 2961 4981 2973 4984
rect 3007 4981 3019 5015
rect 2961 4975 3019 4981
rect 3053 5015 3111 5021
rect 3053 4981 3065 5015
rect 3099 5012 3111 5015
rect 3602 5012 3608 5024
rect 3099 4984 3608 5012
rect 3099 4981 3111 4984
rect 3053 4975 3111 4981
rect 3602 4972 3608 4984
rect 3660 4972 3666 5024
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 3881 5015 3939 5021
rect 3881 5012 3893 5015
rect 3752 4984 3893 5012
rect 3752 4972 3758 4984
rect 3881 4981 3893 4984
rect 3927 4981 3939 5015
rect 6086 5012 6092 5024
rect 6047 4984 6092 5012
rect 3881 4975 3939 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 6457 5015 6515 5021
rect 6236 4984 6281 5012
rect 6236 4972 6242 4984
rect 6457 4981 6469 5015
rect 6503 5012 6515 5015
rect 6730 5012 6736 5024
rect 6503 4984 6736 5012
rect 6503 4981 6515 4984
rect 6457 4975 6515 4981
rect 6730 4972 6736 4984
rect 6788 4972 6794 5024
rect 7300 5021 7328 5052
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8113 5083 8171 5089
rect 8113 5080 8125 5083
rect 7616 5052 8125 5080
rect 7616 5040 7622 5052
rect 8113 5049 8125 5052
rect 8159 5049 8171 5083
rect 8956 5080 8984 5111
rect 9214 5108 9220 5111
rect 9272 5108 9278 5120
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10428 5148 10456 5188
rect 10870 5176 10876 5188
rect 10928 5176 10934 5228
rect 12158 5176 12164 5228
rect 12216 5216 12222 5228
rect 12437 5219 12495 5225
rect 12437 5216 12449 5219
rect 12216 5188 12449 5216
rect 12216 5176 12222 5188
rect 12437 5185 12449 5188
rect 12483 5185 12495 5219
rect 13464 5216 13492 5324
rect 13906 5312 13912 5324
rect 13964 5312 13970 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 15010 5352 15016 5364
rect 14240 5324 15016 5352
rect 14240 5312 14246 5324
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17586 5352 17592 5364
rect 17184 5324 17592 5352
rect 17184 5312 17190 5324
rect 17586 5312 17592 5324
rect 17644 5352 17650 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 17644 5324 18429 5352
rect 17644 5312 17650 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 13538 5244 13544 5296
rect 13596 5284 13602 5296
rect 13817 5287 13875 5293
rect 13817 5284 13829 5287
rect 13596 5256 13829 5284
rect 13596 5244 13602 5256
rect 13817 5253 13829 5256
rect 13863 5253 13875 5287
rect 16298 5284 16304 5296
rect 13817 5247 13875 5253
rect 14099 5256 15424 5284
rect 14099 5216 14127 5256
rect 13464 5188 14127 5216
rect 12437 5179 12495 5185
rect 14366 5176 14372 5228
rect 14424 5216 14430 5228
rect 14461 5219 14519 5225
rect 14461 5216 14473 5219
rect 14424 5188 14473 5216
rect 14424 5176 14430 5188
rect 14461 5185 14473 5188
rect 14507 5185 14519 5219
rect 14461 5179 14519 5185
rect 9732 5120 10456 5148
rect 9732 5108 9738 5120
rect 9692 5080 9720 5108
rect 8956 5052 9720 5080
rect 8113 5043 8171 5049
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7926 5012 7932 5024
rect 7331 4984 7932 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 10134 5012 10140 5024
rect 9548 4984 10140 5012
rect 9548 4972 9554 4984
rect 10134 4972 10140 4984
rect 10192 4972 10198 5024
rect 10318 4972 10324 5024
rect 10376 5012 10382 5024
rect 10428 5021 10456 5120
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 11140 5151 11198 5157
rect 11140 5117 11152 5151
rect 11186 5148 11198 5151
rect 12342 5148 12348 5160
rect 11186 5120 12348 5148
rect 11186 5117 11198 5120
rect 11140 5111 11198 5117
rect 10612 5080 10640 5111
rect 12342 5108 12348 5120
rect 12400 5108 12406 5160
rect 12693 5151 12751 5157
rect 12693 5148 12705 5151
rect 12452 5120 12705 5148
rect 12158 5080 12164 5092
rect 10612 5052 12164 5080
rect 12158 5040 12164 5052
rect 12216 5040 12222 5092
rect 12452 5080 12480 5120
rect 12693 5117 12705 5120
rect 12739 5117 12751 5151
rect 14918 5148 14924 5160
rect 14879 5120 14924 5148
rect 12693 5111 12751 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 12268 5052 12480 5080
rect 12268 5024 12296 5052
rect 13722 5040 13728 5092
rect 13780 5080 13786 5092
rect 15396 5089 15424 5256
rect 16132 5256 16304 5284
rect 15562 5176 15568 5228
rect 15620 5216 15626 5228
rect 16132 5225 16160 5256
rect 16298 5244 16304 5256
rect 16356 5284 16362 5296
rect 17770 5284 17776 5296
rect 16356 5256 17776 5284
rect 16356 5244 16362 5256
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15620 5188 16129 5216
rect 15620 5176 15626 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16758 5216 16764 5228
rect 16719 5188 16764 5216
rect 16117 5179 16175 5185
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 16868 5225 16896 5256
rect 17770 5244 17776 5256
rect 17828 5244 17834 5296
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17678 5216 17684 5228
rect 17000 5188 17684 5216
rect 17000 5176 17006 5188
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 15470 5108 15476 5160
rect 15528 5148 15534 5160
rect 15933 5151 15991 5157
rect 15933 5148 15945 5151
rect 15528 5120 15945 5148
rect 15528 5108 15534 5120
rect 15933 5117 15945 5120
rect 15979 5117 15991 5151
rect 15933 5111 15991 5117
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17368 5120 18061 5148
rect 17368 5108 17374 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 15381 5083 15439 5089
rect 13780 5052 14780 5080
rect 13780 5040 13786 5052
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 10376 4984 10425 5012
rect 10376 4972 10382 4984
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 10413 4975 10471 4981
rect 10781 5015 10839 5021
rect 10781 4981 10793 5015
rect 10827 5012 10839 5015
rect 11146 5012 11152 5024
rect 10827 4984 11152 5012
rect 10827 4981 10839 4984
rect 10781 4975 10839 4981
rect 11146 4972 11152 4984
rect 11204 4972 11210 5024
rect 12250 5012 12256 5024
rect 12211 4984 12256 5012
rect 12250 4972 12256 4984
rect 12308 4972 12314 5024
rect 14182 4972 14188 5024
rect 14240 5012 14246 5024
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 14240 4984 14289 5012
rect 14240 4972 14246 4984
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14277 4975 14335 4981
rect 14369 5015 14427 5021
rect 14369 4981 14381 5015
rect 14415 5012 14427 5015
rect 14642 5012 14648 5024
rect 14415 4984 14648 5012
rect 14415 4981 14427 4984
rect 14369 4975 14427 4981
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 14752 5021 14780 5052
rect 15381 5049 15393 5083
rect 15427 5080 15439 5083
rect 16669 5083 16727 5089
rect 16669 5080 16681 5083
rect 15427 5052 16681 5080
rect 15427 5049 15439 5052
rect 15381 5043 15439 5049
rect 16669 5049 16681 5052
rect 16715 5080 16727 5083
rect 17954 5080 17960 5092
rect 16715 5052 17960 5080
rect 16715 5049 16727 5052
rect 16669 5043 16727 5049
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 14737 5015 14795 5021
rect 14737 4981 14749 5015
rect 14783 5012 14795 5015
rect 15194 5012 15200 5024
rect 14783 4984 15200 5012
rect 14783 4981 14795 4984
rect 14737 4975 14795 4981
rect 15194 4972 15200 4984
rect 15252 4972 15258 5024
rect 15470 5012 15476 5024
rect 15431 4984 15476 5012
rect 15470 4972 15476 4984
rect 15528 4972 15534 5024
rect 15654 4972 15660 5024
rect 15712 5012 15718 5024
rect 15841 5015 15899 5021
rect 15841 5012 15853 5015
rect 15712 4984 15853 5012
rect 15712 4972 15718 4984
rect 15841 4981 15853 4984
rect 15887 4981 15899 5015
rect 15841 4975 15899 4981
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16574 5012 16580 5024
rect 16347 4984 16580 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16574 4972 16580 4984
rect 16632 4972 16638 5024
rect 17126 5012 17132 5024
rect 17087 4984 17132 5012
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 17218 4972 17224 5024
rect 17276 5012 17282 5024
rect 17497 5015 17555 5021
rect 17497 5012 17509 5015
rect 17276 4984 17509 5012
rect 17276 4972 17282 4984
rect 17497 4981 17509 4984
rect 17543 4981 17555 5015
rect 17497 4975 17555 4981
rect 17586 4972 17592 5024
rect 17644 5012 17650 5024
rect 18230 5012 18236 5024
rect 17644 4984 17689 5012
rect 18191 4984 18236 5012
rect 17644 4972 17650 4984
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 6912 4922
rect 6964 4870 6976 4922
rect 7028 4870 7040 4922
rect 7092 4870 7104 4922
rect 7156 4870 12843 4922
rect 12895 4870 12907 4922
rect 12959 4870 12971 4922
rect 13023 4870 13035 4922
rect 13087 4870 18860 4922
rect 1104 4848 18860 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 1670 4808 1676 4820
rect 1627 4780 1676 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 1670 4768 1676 4780
rect 1728 4808 1734 4820
rect 3602 4808 3608 4820
rect 1728 4780 3608 4808
rect 1728 4768 1734 4780
rect 3602 4768 3608 4780
rect 3660 4768 3666 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3844 4780 3893 4808
rect 3844 4768 3850 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 6178 4808 6184 4820
rect 3881 4771 3939 4777
rect 4264 4780 6184 4808
rect 2768 4743 2826 4749
rect 1688 4712 2728 4740
rect 1688 4681 1716 4712
rect 1673 4675 1731 4681
rect 1673 4641 1685 4675
rect 1719 4641 1731 4675
rect 2038 4672 2044 4684
rect 1999 4644 2044 4672
rect 1673 4635 1731 4641
rect 2038 4632 2044 4644
rect 2096 4632 2102 4684
rect 2700 4672 2728 4712
rect 2768 4709 2780 4743
rect 2814 4740 2826 4743
rect 3234 4740 3240 4752
rect 2814 4712 3240 4740
rect 2814 4709 2826 4712
rect 2768 4703 2826 4709
rect 3234 4700 3240 4712
rect 3292 4700 3298 4752
rect 4264 4681 4292 4780
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 7101 4811 7159 4817
rect 7101 4777 7113 4811
rect 7147 4808 7159 4811
rect 7558 4808 7564 4820
rect 7147 4780 7564 4808
rect 7147 4777 7159 4780
rect 7101 4771 7159 4777
rect 7558 4768 7564 4780
rect 7616 4768 7622 4820
rect 8294 4768 8300 4820
rect 8352 4808 8358 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8352 4780 8585 4808
rect 8352 4768 8358 4780
rect 8573 4777 8585 4780
rect 8619 4777 8631 4811
rect 8573 4771 8631 4777
rect 9125 4811 9183 4817
rect 9125 4777 9137 4811
rect 9171 4808 9183 4811
rect 9766 4808 9772 4820
rect 9171 4780 9772 4808
rect 9171 4777 9183 4780
rect 9125 4771 9183 4777
rect 9766 4768 9772 4780
rect 9824 4768 9830 4820
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 10410 4808 10416 4820
rect 10367 4780 10416 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 10410 4768 10416 4780
rect 10468 4808 10474 4820
rect 10873 4811 10931 4817
rect 10873 4808 10885 4811
rect 10468 4780 10885 4808
rect 10468 4768 10474 4780
rect 10873 4777 10885 4780
rect 10919 4808 10931 4811
rect 11514 4808 11520 4820
rect 10919 4780 11520 4808
rect 10919 4777 10931 4780
rect 10873 4771 10931 4777
rect 11514 4768 11520 4780
rect 11572 4768 11578 4820
rect 11701 4811 11759 4817
rect 11701 4777 11713 4811
rect 11747 4808 11759 4811
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 11747 4780 12081 4808
rect 11747 4777 11759 4780
rect 11701 4771 11759 4777
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12069 4771 12127 4777
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 12897 4811 12955 4817
rect 12897 4808 12909 4811
rect 12768 4780 12909 4808
rect 12768 4768 12774 4780
rect 12897 4777 12909 4780
rect 12943 4777 12955 4811
rect 13354 4808 13360 4820
rect 13315 4780 13360 4808
rect 12897 4771 12955 4777
rect 13354 4768 13360 4780
rect 13412 4768 13418 4820
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 13504 4780 18000 4808
rect 13504 4768 13510 4780
rect 4522 4740 4528 4752
rect 4483 4712 4528 4740
rect 4522 4700 4528 4712
rect 4580 4700 4586 4752
rect 4614 4700 4620 4752
rect 4672 4740 4678 4752
rect 6549 4743 6607 4749
rect 6549 4740 6561 4743
rect 4672 4712 6561 4740
rect 4672 4700 4678 4712
rect 6549 4709 6561 4712
rect 6595 4709 6607 4743
rect 6549 4703 6607 4709
rect 7834 4700 7840 4752
rect 7892 4740 7898 4752
rect 10226 4740 10232 4752
rect 7892 4712 10232 4740
rect 7892 4700 7898 4712
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 11609 4743 11667 4749
rect 11609 4709 11621 4743
rect 11655 4740 11667 4743
rect 12526 4740 12532 4752
rect 11655 4712 12532 4740
rect 11655 4709 11667 4712
rect 11609 4703 11667 4709
rect 12526 4700 12532 4712
rect 12584 4700 12590 4752
rect 13265 4743 13323 4749
rect 13265 4709 13277 4743
rect 13311 4740 13323 4743
rect 14550 4740 14556 4752
rect 13311 4712 14556 4740
rect 13311 4709 13323 4712
rect 13265 4703 13323 4709
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 15562 4749 15568 4752
rect 15556 4740 15568 4749
rect 15523 4712 15568 4740
rect 15556 4703 15568 4712
rect 15562 4700 15568 4703
rect 15620 4700 15626 4752
rect 16942 4740 16948 4752
rect 16903 4712 16948 4740
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 17034 4700 17040 4752
rect 17092 4740 17098 4752
rect 17497 4743 17555 4749
rect 17497 4740 17509 4743
rect 17092 4712 17509 4740
rect 17092 4700 17098 4712
rect 17497 4709 17509 4712
rect 17543 4709 17555 4743
rect 17497 4703 17555 4709
rect 4249 4675 4307 4681
rect 2700 4644 4200 4672
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 2501 4607 2559 4613
rect 2501 4604 2513 4607
rect 1360 4576 2513 4604
rect 1360 4564 1366 4576
rect 2501 4573 2513 4576
rect 2547 4573 2559 4607
rect 2501 4567 2559 4573
rect 1854 4468 1860 4480
rect 1815 4440 1860 4468
rect 1854 4428 1860 4440
rect 1912 4428 1918 4480
rect 2222 4468 2228 4480
rect 2183 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 2516 4468 2544 4567
rect 4172 4536 4200 4644
rect 4249 4641 4261 4675
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 4338 4632 4344 4684
rect 4396 4672 4402 4684
rect 4801 4675 4859 4681
rect 4801 4672 4813 4675
rect 4396 4644 4813 4672
rect 4396 4632 4402 4644
rect 4801 4641 4813 4644
rect 4847 4641 4859 4675
rect 4801 4635 4859 4641
rect 4816 4604 4844 4635
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5350 4672 5356 4684
rect 5224 4644 5356 4672
rect 5224 4632 5230 4644
rect 5350 4632 5356 4644
rect 5408 4632 5414 4684
rect 5810 4672 5816 4684
rect 5771 4644 5816 4672
rect 5810 4632 5816 4644
rect 5868 4632 5874 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 7460 4675 7518 4681
rect 7460 4641 7472 4675
rect 7506 4672 7518 4675
rect 8202 4672 8208 4684
rect 7506 4644 8208 4672
rect 7506 4641 7518 4644
rect 7460 4635 7518 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9306 4672 9312 4684
rect 9263 4644 9312 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 9306 4632 9312 4644
rect 9364 4672 9370 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 9364 4644 9689 4672
rect 9364 4632 9370 4644
rect 9677 4641 9689 4644
rect 9723 4641 9735 4675
rect 9677 4635 9735 4641
rect 10134 4632 10140 4684
rect 10192 4672 10198 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10192 4644 10793 4672
rect 10192 4632 10198 4644
rect 10781 4641 10793 4644
rect 10827 4641 10839 4675
rect 10781 4635 10839 4641
rect 10888 4644 11468 4672
rect 5445 4607 5503 4613
rect 5445 4604 5457 4607
rect 4816 4576 5457 4604
rect 5445 4573 5457 4576
rect 5491 4573 5503 4607
rect 5626 4604 5632 4616
rect 5587 4576 5632 4604
rect 5445 4567 5503 4573
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6972 4576 7205 4604
rect 6972 4564 6978 4576
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8444 4576 9413 4604
rect 8444 4564 8450 4576
rect 9401 4573 9413 4576
rect 9447 4604 9459 4607
rect 10888 4604 10916 4644
rect 9447 4576 10916 4604
rect 11057 4607 11115 4613
rect 9447 4573 9459 4576
rect 9401 4567 9459 4573
rect 11057 4573 11069 4607
rect 11103 4604 11115 4607
rect 11330 4604 11336 4616
rect 11103 4576 11336 4604
rect 11103 4573 11115 4576
rect 11057 4567 11115 4573
rect 11330 4564 11336 4576
rect 11388 4564 11394 4616
rect 11440 4604 11468 4644
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 13981 4675 14039 4681
rect 13981 4672 13993 4675
rect 12492 4644 12537 4672
rect 13556 4644 13993 4672
rect 12492 4632 12498 4644
rect 11606 4604 11612 4616
rect 11440 4576 11612 4604
rect 11606 4564 11612 4576
rect 11664 4564 11670 4616
rect 11885 4607 11943 4613
rect 11885 4573 11897 4607
rect 11931 4604 11943 4607
rect 12250 4604 12256 4616
rect 11931 4576 12256 4604
rect 11931 4573 11943 4576
rect 11885 4567 11943 4573
rect 12250 4564 12256 4576
rect 12308 4564 12314 4616
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 13556 4613 13584 4644
rect 13981 4641 13993 4644
rect 14027 4672 14039 4675
rect 14274 4672 14280 4684
rect 14027 4644 14280 4672
rect 14027 4641 14039 4644
rect 13981 4635 14039 4641
rect 14274 4632 14280 4644
rect 14332 4632 14338 4684
rect 14458 4632 14464 4684
rect 14516 4672 14522 4684
rect 16761 4675 16819 4681
rect 16761 4672 16773 4675
rect 14516 4644 16773 4672
rect 14516 4632 14522 4644
rect 16761 4641 16773 4644
rect 16807 4672 16819 4675
rect 17310 4672 17316 4684
rect 16807 4644 17316 4672
rect 16807 4641 16819 4644
rect 16761 4635 16819 4641
rect 17310 4632 17316 4644
rect 17368 4632 17374 4684
rect 17972 4681 18000 4780
rect 17957 4675 18015 4681
rect 17957 4641 17969 4675
rect 18003 4672 18015 4675
rect 18325 4675 18383 4681
rect 18325 4672 18337 4675
rect 18003 4644 18337 4672
rect 18003 4641 18015 4644
rect 17957 4635 18015 4641
rect 18325 4641 18337 4644
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 12713 4607 12771 4613
rect 12713 4573 12725 4607
rect 12759 4573 12771 4607
rect 12713 4567 12771 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13722 4604 13728 4616
rect 13683 4576 13728 4604
rect 13541 4567 13599 4573
rect 6181 4539 6239 4545
rect 6181 4536 6193 4539
rect 4172 4508 6193 4536
rect 6181 4505 6193 4508
rect 6227 4536 6239 4539
rect 11146 4536 11152 4548
rect 6227 4508 7236 4536
rect 6227 4505 6239 4508
rect 6181 4499 6239 4505
rect 4065 4471 4123 4477
rect 4065 4468 4077 4471
rect 2516 4440 4077 4468
rect 4065 4437 4077 4440
rect 4111 4468 4123 4471
rect 4246 4468 4252 4480
rect 4111 4440 4252 4468
rect 4111 4437 4123 4440
rect 4065 4431 4123 4437
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4430 4468 4436 4480
rect 4391 4440 4436 4468
rect 4430 4428 4436 4440
rect 4488 4428 4494 4480
rect 4982 4468 4988 4480
rect 4943 4440 4988 4468
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5442 4428 5448 4480
rect 5500 4468 5506 4480
rect 5997 4471 6055 4477
rect 5997 4468 6009 4471
rect 5500 4440 6009 4468
rect 5500 4428 5506 4440
rect 5997 4437 6009 4440
rect 6043 4437 6055 4471
rect 6730 4468 6736 4480
rect 6691 4440 6736 4468
rect 5997 4431 6055 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 7208 4468 7236 4508
rect 8128 4508 11152 4536
rect 8128 4468 8156 4508
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 12342 4496 12348 4548
rect 12400 4536 12406 4548
rect 12728 4536 12756 4567
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 15289 4607 15347 4613
rect 15289 4604 15301 4607
rect 15252 4576 15301 4604
rect 15252 4564 15258 4576
rect 15289 4573 15301 4576
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 16942 4564 16948 4616
rect 17000 4604 17006 4616
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 17000 4576 17601 4604
rect 17000 4564 17006 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 17589 4567 17647 4573
rect 13170 4536 13176 4548
rect 12400 4508 13176 4536
rect 12400 4496 12406 4508
rect 13170 4496 13176 4508
rect 13228 4536 13234 4548
rect 17604 4536 17632 4567
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 17736 4576 17781 4604
rect 17736 4564 17742 4576
rect 18046 4536 18052 4548
rect 13228 4508 13492 4536
rect 17604 4508 18052 4536
rect 13228 4496 13234 4508
rect 8754 4468 8760 4480
rect 7208 4440 8156 4468
rect 8715 4440 8760 4468
rect 8754 4428 8760 4440
rect 8812 4428 8818 4480
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 9861 4471 9919 4477
rect 9861 4468 9873 4471
rect 9732 4440 9873 4468
rect 9732 4428 9738 4440
rect 9861 4437 9873 4440
rect 9907 4437 9919 4471
rect 9861 4431 9919 4437
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 10226 4468 10232 4480
rect 10183 4440 10232 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 10226 4428 10232 4440
rect 10284 4428 10290 4480
rect 10410 4468 10416 4480
rect 10371 4440 10416 4468
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 13354 4468 13360 4480
rect 11287 4440 13360 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13464 4468 13492 4508
rect 18046 4496 18052 4508
rect 18104 4496 18110 4548
rect 15105 4471 15163 4477
rect 15105 4468 15117 4471
rect 13464 4440 15117 4468
rect 15105 4437 15117 4440
rect 15151 4437 15163 4471
rect 16666 4468 16672 4480
rect 16627 4440 16672 4468
rect 15105 4431 15163 4437
rect 16666 4428 16672 4440
rect 16724 4428 16730 4480
rect 17129 4471 17187 4477
rect 17129 4437 17141 4471
rect 17175 4468 17187 4471
rect 17218 4468 17224 4480
rect 17175 4440 17224 4468
rect 17175 4437 17187 4440
rect 17129 4431 17187 4437
rect 17218 4428 17224 4440
rect 17276 4428 17282 4480
rect 17310 4428 17316 4480
rect 17368 4468 17374 4480
rect 17586 4468 17592 4480
rect 17368 4440 17592 4468
rect 17368 4428 17374 4440
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18141 4471 18199 4477
rect 18141 4468 18153 4471
rect 17920 4440 18153 4468
rect 17920 4428 17926 4440
rect 18141 4437 18153 4440
rect 18187 4437 18199 4471
rect 18141 4431 18199 4437
rect 1104 4378 18860 4400
rect 1104 4326 3947 4378
rect 3999 4326 4011 4378
rect 4063 4326 4075 4378
rect 4127 4326 4139 4378
rect 4191 4326 9878 4378
rect 9930 4326 9942 4378
rect 9994 4326 10006 4378
rect 10058 4326 10070 4378
rect 10122 4326 15808 4378
rect 15860 4326 15872 4378
rect 15924 4326 15936 4378
rect 15988 4326 16000 4378
rect 16052 4326 18860 4378
rect 1104 4304 18860 4326
rect 4522 4224 4528 4276
rect 4580 4264 4586 4276
rect 4798 4264 4804 4276
rect 4580 4236 4804 4264
rect 4580 4224 4586 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 6454 4264 6460 4276
rect 5776 4236 6460 4264
rect 5776 4224 5782 4236
rect 6454 4224 6460 4236
rect 6512 4224 6518 4276
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8202 4264 8208 4276
rect 7984 4236 8208 4264
rect 7984 4224 7990 4236
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10502 4264 10508 4276
rect 9732 4236 10508 4264
rect 9732 4224 9738 4236
rect 10502 4224 10508 4236
rect 10560 4264 10566 4276
rect 11514 4264 11520 4276
rect 10560 4236 11520 4264
rect 10560 4224 10566 4236
rect 11514 4224 11520 4236
rect 11572 4264 11578 4276
rect 12066 4264 12072 4276
rect 11572 4236 12072 4264
rect 11572 4224 11578 4236
rect 12066 4224 12072 4236
rect 12124 4264 12130 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 12124 4236 12173 4264
rect 12124 4224 12130 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 12434 4224 12440 4276
rect 12492 4264 12498 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 12492 4236 13737 4264
rect 12492 4224 12498 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 14090 4264 14096 4276
rect 13725 4227 13783 4233
rect 13832 4236 14096 4264
rect 1762 4156 1768 4208
rect 1820 4156 1826 4208
rect 3421 4199 3479 4205
rect 3421 4196 3433 4199
rect 3068 4168 3433 4196
rect 1780 4128 1808 4156
rect 1780 4100 1900 4128
rect 1489 4063 1547 4069
rect 1489 4029 1501 4063
rect 1535 4060 1547 4063
rect 1762 4060 1768 4072
rect 1535 4032 1768 4060
rect 1535 4029 1547 4032
rect 1489 4023 1547 4029
rect 1762 4020 1768 4032
rect 1820 4020 1826 4072
rect 1872 4069 1900 4100
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3068 4137 3096 4168
rect 3421 4165 3433 4168
rect 3467 4196 3479 4199
rect 6730 4196 6736 4208
rect 3467 4168 6736 4196
rect 3467 4165 3479 4168
rect 3421 4159 3479 4165
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 10137 4199 10195 4205
rect 10137 4165 10149 4199
rect 10183 4196 10195 4199
rect 10226 4196 10232 4208
rect 10183 4168 10232 4196
rect 10183 4165 10195 4168
rect 10137 4159 10195 4165
rect 10226 4156 10232 4168
rect 10284 4156 10290 4208
rect 11606 4196 11612 4208
rect 10796 4168 11612 4196
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 2832 4100 3065 4128
rect 2832 4088 2838 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3053 4091 3111 4097
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 4522 4128 4528 4140
rect 4483 4100 4528 4128
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 5040 4100 5181 4128
rect 5040 4088 5046 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5626 4128 5632 4140
rect 5399 4100 5632 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5626 4088 5632 4100
rect 5684 4128 5690 4140
rect 6086 4128 6092 4140
rect 5684 4100 6092 4128
rect 5684 4088 5690 4100
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10410 4088 10416 4140
rect 10468 4128 10474 4140
rect 10796 4137 10824 4168
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10468 4100 10609 4128
rect 10468 4088 10474 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 11422 4088 11428 4140
rect 11480 4088 11486 4140
rect 11532 4137 11560 4168
rect 11606 4156 11612 4168
rect 11664 4156 11670 4208
rect 13832 4196 13860 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 15010 4196 15016 4208
rect 11808 4168 13860 4196
rect 14016 4168 15016 4196
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4029 1915 4063
rect 1857 4023 1915 4029
rect 2225 4063 2283 4069
rect 2225 4029 2237 4063
rect 2271 4029 2283 4063
rect 2958 4060 2964 4072
rect 2919 4032 2964 4060
rect 2225 4023 2283 4029
rect 2240 3992 2268 4023
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 5442 4060 5448 4072
rect 4172 4032 5448 4060
rect 4172 3992 4200 4032
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 5592 4032 6837 4060
rect 5592 4020 5598 4032
rect 6825 4029 6837 4032
rect 6871 4060 6883 4063
rect 6914 4060 6920 4072
rect 6871 4032 6920 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 6914 4020 6920 4032
rect 6972 4060 6978 4072
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 6972 4032 8309 4060
rect 6972 4020 6978 4032
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 9674 4060 9680 4072
rect 8297 4023 8355 4029
rect 8404 4032 9680 4060
rect 2240 3964 4200 3992
rect 4249 3995 4307 4001
rect 4249 3961 4261 3995
rect 4295 3992 4307 3995
rect 4295 3964 5580 3992
rect 4295 3961 4307 3964
rect 4249 3955 4307 3961
rect 1670 3924 1676 3936
rect 1631 3896 1676 3924
rect 1670 3884 1676 3896
rect 1728 3884 1734 3936
rect 2038 3924 2044 3936
rect 1999 3896 2044 3924
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2406 3924 2412 3936
rect 2367 3896 2412 3924
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2590 3924 2596 3936
rect 2551 3896 2596 3924
rect 2590 3884 2596 3896
rect 2648 3884 2654 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4387 3896 4721 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 4798 3884 4804 3936
rect 4856 3924 4862 3936
rect 5552 3933 5580 3964
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 5905 3995 5963 4001
rect 5905 3992 5917 3995
rect 5868 3964 5917 3992
rect 5868 3952 5874 3964
rect 5905 3961 5917 3964
rect 5951 3992 5963 3995
rect 6638 3992 6644 4004
rect 5951 3964 6644 3992
rect 5951 3961 5963 3964
rect 5905 3955 5963 3961
rect 6638 3952 6644 3964
rect 6696 3952 6702 4004
rect 6730 3952 6736 4004
rect 6788 3992 6794 4004
rect 7070 3995 7128 4001
rect 7070 3992 7082 3995
rect 6788 3964 7082 3992
rect 6788 3952 6794 3964
rect 7070 3961 7082 3964
rect 7116 3961 7128 3995
rect 7070 3955 7128 3961
rect 7650 3952 7656 4004
rect 7708 3992 7714 4004
rect 8404 3992 8432 4032
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10318 4060 10324 4072
rect 9824 4032 10324 4060
rect 9824 4020 9830 4032
rect 10318 4020 10324 4032
rect 10376 4060 10382 4072
rect 11440 4060 11468 4088
rect 10376 4032 11468 4060
rect 10376 4020 10382 4032
rect 7708 3964 8432 3992
rect 8564 3995 8622 4001
rect 7708 3952 7714 3964
rect 8564 3961 8576 3995
rect 8610 3992 8622 3995
rect 9122 3992 9128 4004
rect 8610 3964 9128 3992
rect 8610 3961 8622 3964
rect 8564 3955 8622 3961
rect 9122 3952 9128 3964
rect 9180 3952 9186 4004
rect 11054 3992 11060 4004
rect 9223 3964 11060 3992
rect 5077 3927 5135 3933
rect 5077 3924 5089 3927
rect 4856 3896 5089 3924
rect 4856 3884 4862 3896
rect 5077 3893 5089 3896
rect 5123 3893 5135 3927
rect 5077 3887 5135 3893
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 6086 3924 6092 3936
rect 6043 3896 6092 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6270 3884 6276 3936
rect 6328 3924 6334 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6328 3896 6377 3924
rect 6328 3884 6334 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 6454 3884 6460 3936
rect 6512 3924 6518 3936
rect 9223 3924 9251 3964
rect 11054 3952 11060 3964
rect 11112 3952 11118 4004
rect 11146 3952 11152 4004
rect 11204 3992 11210 4004
rect 11425 3995 11483 4001
rect 11425 3992 11437 3995
rect 11204 3964 11437 3992
rect 11204 3952 11210 3964
rect 11425 3961 11437 3964
rect 11471 3992 11483 3995
rect 11808 3992 11836 4168
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 11940 4100 12449 4128
rect 11940 4088 11946 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 13262 4128 13268 4140
rect 12851 4100 13268 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13446 4128 13452 4140
rect 13407 4100 13452 4128
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13280 4060 13308 4088
rect 13357 4063 13415 4069
rect 13357 4060 13369 4063
rect 13280 4032 13369 4060
rect 13357 4029 13369 4032
rect 13403 4060 13415 4063
rect 14016 4060 14044 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 16666 4196 16672 4208
rect 16500 4168 16672 4196
rect 14274 4128 14280 4140
rect 14235 4100 14280 4128
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 15194 4088 15200 4140
rect 15252 4128 15258 4140
rect 15289 4131 15347 4137
rect 15289 4128 15301 4131
rect 15252 4100 15301 4128
rect 15252 4088 15258 4100
rect 15289 4097 15301 4100
rect 15335 4097 15347 4131
rect 15289 4091 15347 4097
rect 13403 4032 14044 4060
rect 14093 4063 14151 4069
rect 13403 4029 13415 4032
rect 13357 4023 13415 4029
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 14458 4060 14464 4072
rect 14139 4032 14464 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 14458 4020 14464 4032
rect 14516 4060 14522 4072
rect 14829 4063 14887 4069
rect 14829 4060 14841 4063
rect 14516 4032 14841 4060
rect 14516 4020 14522 4032
rect 14829 4029 14841 4032
rect 14875 4029 14887 4063
rect 14829 4023 14887 4029
rect 15556 4063 15614 4069
rect 15556 4029 15568 4063
rect 15602 4060 15614 4063
rect 16500 4060 16528 4168
rect 16666 4156 16672 4168
rect 16724 4156 16730 4208
rect 17770 4196 17776 4208
rect 17420 4168 17776 4196
rect 17034 4128 17040 4140
rect 15602 4032 16528 4060
rect 16592 4100 17040 4128
rect 15602 4029 15614 4032
rect 15556 4023 15614 4029
rect 11977 3995 12035 4001
rect 11977 3992 11989 3995
rect 11471 3964 11989 3992
rect 11471 3961 11483 3964
rect 11425 3955 11483 3961
rect 11977 3961 11989 3964
rect 12023 3961 12035 3995
rect 11977 3955 12035 3961
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 15013 3995 15071 4001
rect 15013 3992 15025 3995
rect 13596 3964 15025 3992
rect 13596 3952 13602 3964
rect 15013 3961 15025 3964
rect 15059 3961 15071 3995
rect 15013 3955 15071 3961
rect 6512 3896 9251 3924
rect 9677 3927 9735 3933
rect 6512 3884 6518 3896
rect 9677 3893 9689 3927
rect 9723 3924 9735 3927
rect 9950 3924 9956 3936
rect 9723 3896 9956 3924
rect 9723 3893 9735 3896
rect 9677 3887 9735 3893
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10091 3896 10517 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10505 3893 10517 3896
rect 10551 3924 10563 3927
rect 10686 3924 10692 3936
rect 10551 3896 10692 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10962 3924 10968 3936
rect 10923 3896 10968 3924
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11606 3924 11612 3936
rect 11379 3896 11612 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11606 3884 11612 3896
rect 11664 3924 11670 3936
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11664 3896 11805 3924
rect 11664 3884 11670 3896
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13170 3924 13176 3936
rect 12943 3896 13176 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 13265 3927 13323 3933
rect 13265 3893 13277 3927
rect 13311 3924 13323 3927
rect 13906 3924 13912 3936
rect 13311 3896 13912 3924
rect 13311 3893 13323 3896
rect 13265 3887 13323 3893
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 14182 3924 14188 3936
rect 14143 3896 14188 3924
rect 14182 3884 14188 3896
rect 14240 3884 14246 3936
rect 14734 3884 14740 3936
rect 14792 3924 14798 3936
rect 16592 3924 16620 4100
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17218 4128 17224 4140
rect 17179 4100 17224 4128
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17420 4137 17448 4168
rect 17770 4156 17776 4168
rect 17828 4156 17834 4208
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17405 4091 17463 4097
rect 16758 4020 16764 4072
rect 16816 4020 16822 4072
rect 17126 4060 17132 4072
rect 17087 4032 17132 4060
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4029 17647 4063
rect 18046 4060 18052 4072
rect 18007 4032 18052 4060
rect 17589 4023 17647 4029
rect 16776 3992 16804 4020
rect 16684 3964 16804 3992
rect 16684 3933 16712 3964
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17604 3992 17632 4023
rect 18046 4020 18052 4032
rect 18104 4060 18110 4072
rect 18417 4063 18475 4069
rect 18417 4060 18429 4063
rect 18104 4032 18429 4060
rect 18104 4020 18110 4032
rect 18417 4029 18429 4032
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 17000 3964 17632 3992
rect 17000 3952 17006 3964
rect 14792 3896 16620 3924
rect 16669 3927 16727 3933
rect 14792 3884 14798 3896
rect 16669 3893 16681 3927
rect 16715 3893 16727 3927
rect 16669 3887 16727 3893
rect 16761 3927 16819 3933
rect 16761 3893 16773 3927
rect 16807 3924 16819 3927
rect 16850 3924 16856 3936
rect 16807 3896 16856 3924
rect 16807 3893 16819 3896
rect 16761 3887 16819 3893
rect 16850 3884 16856 3896
rect 16908 3884 16914 3936
rect 17770 3924 17776 3936
rect 17731 3896 17776 3924
rect 17770 3884 17776 3896
rect 17828 3884 17834 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18233 3927 18291 3933
rect 18233 3924 18245 3927
rect 17920 3896 18245 3924
rect 17920 3884 17926 3896
rect 18233 3893 18245 3896
rect 18279 3893 18291 3927
rect 18233 3887 18291 3893
rect 1104 3834 18860 3856
rect 1104 3782 6912 3834
rect 6964 3782 6976 3834
rect 7028 3782 7040 3834
rect 7092 3782 7104 3834
rect 7156 3782 12843 3834
rect 12895 3782 12907 3834
rect 12959 3782 12971 3834
rect 13023 3782 13035 3834
rect 13087 3782 18860 3834
rect 1104 3760 18860 3782
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3234 3720 3240 3732
rect 2823 3692 3240 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3234 3680 3240 3692
rect 3292 3680 3298 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3878 3720 3884 3732
rect 3651 3692 3884 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4522 3680 4528 3732
rect 4580 3720 4586 3732
rect 5166 3720 5172 3732
rect 4580 3692 5172 3720
rect 4580 3680 4586 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 7285 3723 7343 3729
rect 5276 3692 5948 3720
rect 3694 3612 3700 3664
rect 3752 3652 3758 3664
rect 5276 3652 5304 3692
rect 3752 3624 5304 3652
rect 3752 3612 3758 3624
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 5782 3655 5840 3661
rect 5782 3652 5794 3655
rect 5500 3624 5794 3652
rect 5500 3612 5506 3624
rect 5782 3621 5794 3624
rect 5828 3621 5840 3655
rect 5920 3652 5948 3692
rect 7285 3689 7297 3723
rect 7331 3720 7343 3723
rect 7374 3720 7380 3732
rect 7331 3692 7380 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 8662 3720 8668 3732
rect 7484 3692 8668 3720
rect 7484 3652 7512 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 8754 3680 8760 3732
rect 8812 3720 8818 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 8812 3692 9137 3720
rect 8812 3680 8818 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 9217 3723 9275 3729
rect 9217 3689 9229 3723
rect 9263 3720 9275 3723
rect 10962 3720 10968 3732
rect 9263 3692 10968 3720
rect 9263 3689 9275 3692
rect 9217 3683 9275 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11054 3680 11060 3732
rect 11112 3720 11118 3732
rect 15933 3723 15991 3729
rect 11112 3692 15884 3720
rect 11112 3680 11118 3692
rect 7745 3655 7803 3661
rect 7745 3652 7757 3655
rect 5920 3624 7512 3652
rect 7576 3624 7757 3652
rect 5782 3615 5840 3621
rect 382 3544 388 3596
rect 440 3584 446 3596
rect 1653 3587 1711 3593
rect 1653 3584 1665 3587
rect 440 3556 1665 3584
rect 440 3544 446 3556
rect 1653 3553 1665 3556
rect 1699 3584 1711 3587
rect 2869 3587 2927 3593
rect 2869 3584 2881 3587
rect 1699 3556 2881 3584
rect 1699 3553 1711 3556
rect 1653 3547 1711 3553
rect 2869 3553 2881 3556
rect 2915 3553 2927 3587
rect 3510 3584 3516 3596
rect 3471 3556 3516 3584
rect 2869 3547 2927 3553
rect 3510 3544 3516 3556
rect 3568 3544 3574 3596
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4154 3584 4160 3596
rect 4111 3556 4160 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 4332 3587 4390 3593
rect 4332 3553 4344 3587
rect 4378 3584 4390 3587
rect 5626 3584 5632 3596
rect 4378 3556 5632 3584
rect 4378 3553 4390 3556
rect 4332 3547 4390 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 7193 3587 7251 3593
rect 7193 3584 7205 3587
rect 6604 3556 7205 3584
rect 6604 3544 6610 3556
rect 7193 3553 7205 3556
rect 7239 3584 7251 3587
rect 7576 3584 7604 3624
rect 7745 3621 7757 3624
rect 7791 3652 7803 3655
rect 8386 3652 8392 3664
rect 7791 3624 8392 3652
rect 7791 3621 7803 3624
rect 7745 3615 7803 3621
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 9306 3652 9312 3664
rect 8527 3624 9312 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 9306 3612 9312 3624
rect 9364 3612 9370 3664
rect 10686 3652 10692 3664
rect 9600 3624 10692 3652
rect 7239 3556 7604 3584
rect 7653 3587 7711 3593
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7653 3553 7665 3587
rect 7699 3584 7711 3587
rect 8205 3587 8263 3593
rect 7699 3556 8055 3584
rect 7699 3553 7711 3556
rect 7653 3547 7711 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 5534 3516 5540 3528
rect 5495 3488 5540 3516
rect 3789 3479 3847 3485
rect 3145 3383 3203 3389
rect 3145 3349 3157 3383
rect 3191 3380 3203 3383
rect 3418 3380 3424 3392
rect 3191 3352 3424 3380
rect 3191 3349 3203 3352
rect 3145 3343 3203 3349
rect 3418 3340 3424 3352
rect 3476 3340 3482 3392
rect 3804 3380 3832 3479
rect 5534 3476 5540 3488
rect 5592 3476 5598 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 7668 3516 7696 3547
rect 7926 3516 7932 3528
rect 7616 3488 7696 3516
rect 7887 3488 7932 3516
rect 7616 3476 7622 3488
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8027 3516 8055 3556
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 9030 3584 9036 3596
rect 8251 3556 9036 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 8938 3516 8944 3528
rect 8027 3488 8944 3516
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 9398 3516 9404 3528
rect 9311 3488 9404 3516
rect 9398 3476 9404 3488
rect 9456 3516 9462 3528
rect 9600 3516 9628 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 12802 3612 12808 3664
rect 12860 3652 12866 3664
rect 13164 3655 13222 3661
rect 13164 3652 13176 3655
rect 12860 3624 13176 3652
rect 12860 3612 12866 3624
rect 13164 3621 13176 3624
rect 13210 3652 13222 3655
rect 13446 3652 13452 3664
rect 13210 3624 13452 3652
rect 13210 3621 13222 3624
rect 13164 3615 13222 3621
rect 13446 3612 13452 3624
rect 13504 3612 13510 3664
rect 13906 3612 13912 3664
rect 13964 3652 13970 3664
rect 14369 3655 14427 3661
rect 14369 3652 14381 3655
rect 13964 3624 14381 3652
rect 13964 3612 13970 3624
rect 14369 3621 14381 3624
rect 14415 3621 14427 3655
rect 14369 3615 14427 3621
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 15381 3655 15439 3661
rect 15381 3652 15393 3655
rect 14792 3624 15393 3652
rect 14792 3612 14798 3624
rect 15381 3621 15393 3624
rect 15427 3621 15439 3655
rect 15856 3652 15884 3692
rect 15933 3689 15945 3723
rect 15979 3720 15991 3723
rect 16114 3720 16120 3732
rect 15979 3692 16120 3720
rect 15979 3689 15991 3692
rect 15933 3683 15991 3689
rect 16114 3680 16120 3692
rect 16172 3680 16178 3732
rect 16850 3720 16856 3732
rect 16811 3692 16856 3720
rect 16850 3680 16856 3692
rect 16908 3680 16914 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17313 3723 17371 3729
rect 17313 3720 17325 3723
rect 17000 3692 17325 3720
rect 17000 3680 17006 3692
rect 17313 3689 17325 3692
rect 17359 3689 17371 3723
rect 17494 3720 17500 3732
rect 17455 3692 17500 3720
rect 17313 3683 17371 3689
rect 17494 3680 17500 3692
rect 17552 3720 17558 3732
rect 17552 3692 18276 3720
rect 17552 3680 17558 3692
rect 15856 3624 16528 3652
rect 15381 3615 15439 3621
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9766 3584 9772 3596
rect 9723 3556 9772 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9766 3544 9772 3556
rect 9824 3544 9830 3596
rect 9950 3593 9956 3596
rect 9944 3584 9956 3593
rect 9863 3556 9956 3584
rect 9944 3547 9956 3556
rect 10008 3584 10014 3596
rect 10410 3584 10416 3596
rect 10008 3556 10416 3584
rect 9950 3544 9956 3547
rect 10008 3544 10014 3556
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 11681 3587 11739 3593
rect 11681 3584 11693 3587
rect 11256 3556 11693 3584
rect 11146 3516 11152 3528
rect 9456 3488 9628 3516
rect 11107 3488 11152 3516
rect 9456 3476 9462 3488
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5442 3448 5448 3460
rect 5224 3420 5448 3448
rect 5224 3408 5230 3420
rect 5442 3408 5448 3420
rect 5500 3408 5506 3460
rect 8846 3408 8852 3460
rect 8904 3448 8910 3460
rect 9674 3448 9680 3460
rect 8904 3420 9680 3448
rect 8904 3408 8910 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 11256 3448 11284 3556
rect 11681 3553 11693 3556
rect 11727 3553 11739 3587
rect 11681 3547 11739 3553
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3584 12955 3587
rect 13722 3584 13728 3596
rect 12943 3556 13728 3584
rect 12943 3553 12955 3556
rect 12897 3547 12955 3553
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14645 3587 14703 3593
rect 14645 3553 14657 3587
rect 14691 3584 14703 3587
rect 15930 3584 15936 3596
rect 14691 3556 15936 3584
rect 14691 3553 14703 3556
rect 14645 3547 14703 3553
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 16025 3587 16083 3593
rect 16025 3553 16037 3587
rect 16071 3584 16083 3587
rect 16206 3584 16212 3596
rect 16071 3556 16212 3584
rect 16071 3553 16083 3556
rect 16025 3547 16083 3553
rect 16206 3544 16212 3556
rect 16264 3544 16270 3596
rect 16500 3584 16528 3624
rect 16574 3612 16580 3664
rect 16632 3652 16638 3664
rect 16761 3655 16819 3661
rect 16761 3652 16773 3655
rect 16632 3624 16773 3652
rect 16632 3612 16638 3624
rect 16761 3621 16773 3624
rect 16807 3621 16819 3655
rect 18138 3652 18144 3664
rect 16761 3615 16819 3621
rect 17788 3624 18144 3652
rect 17788 3584 17816 3624
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18248 3593 18276 3692
rect 16500 3556 17816 3584
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3553 17923 3587
rect 17865 3547 17923 3553
rect 18233 3587 18291 3593
rect 18233 3553 18245 3587
rect 18279 3553 18291 3587
rect 18233 3547 18291 3553
rect 11422 3516 11428 3528
rect 11383 3488 11428 3516
rect 11422 3476 11428 3488
rect 11480 3476 11486 3528
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3516 14979 3519
rect 15654 3516 15660 3528
rect 14967 3488 15660 3516
rect 14967 3485 14979 3488
rect 14921 3479 14979 3485
rect 15654 3476 15660 3488
rect 15712 3476 15718 3528
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3516 16175 3519
rect 16298 3516 16304 3528
rect 16163 3488 16304 3516
rect 16163 3485 16175 3488
rect 16117 3479 16175 3485
rect 16298 3476 16304 3488
rect 16356 3476 16362 3528
rect 16666 3476 16672 3528
rect 16724 3516 16730 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16724 3488 16957 3516
rect 16724 3476 16730 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17773 3519 17831 3525
rect 17773 3485 17785 3519
rect 17819 3516 17831 3519
rect 17880 3516 17908 3547
rect 17819 3488 17908 3516
rect 17819 3485 17831 3488
rect 17773 3479 17831 3485
rect 12802 3448 12808 3460
rect 11072 3420 11284 3448
rect 12763 3420 12808 3448
rect 11072 3392 11100 3420
rect 12802 3408 12808 3420
rect 12860 3408 12866 3460
rect 15378 3408 15384 3460
rect 15436 3448 15442 3460
rect 17788 3448 17816 3479
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18690 3516 18696 3528
rect 18196 3488 18696 3516
rect 18196 3476 18202 3488
rect 18690 3476 18696 3488
rect 18748 3476 18754 3528
rect 15436 3420 17816 3448
rect 15436 3408 15442 3420
rect 6730 3380 6736 3392
rect 3804 3352 6736 3380
rect 6730 3340 6736 3352
rect 6788 3380 6794 3392
rect 6917 3383 6975 3389
rect 6917 3380 6929 3383
rect 6788 3352 6929 3380
rect 6788 3340 6794 3352
rect 6917 3349 6929 3352
rect 6963 3349 6975 3383
rect 6917 3343 6975 3349
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 8570 3380 8576 3392
rect 7064 3352 8576 3380
rect 7064 3340 7070 3352
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 9398 3380 9404 3392
rect 8803 3352 9404 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 11054 3380 11060 3392
rect 11015 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14274 3380 14280 3392
rect 13596 3352 14280 3380
rect 13596 3340 13602 3352
rect 14274 3340 14280 3352
rect 14332 3340 14338 3392
rect 15562 3380 15568 3392
rect 15523 3352 15568 3380
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 16393 3383 16451 3389
rect 16393 3349 16405 3383
rect 16439 3380 16451 3383
rect 16666 3380 16672 3392
rect 16439 3352 16672 3380
rect 16439 3349 16451 3352
rect 16393 3343 16451 3349
rect 16666 3340 16672 3352
rect 16724 3340 16730 3392
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 18414 3380 18420 3392
rect 18375 3352 18420 3380
rect 18414 3340 18420 3352
rect 18472 3340 18478 3392
rect 1104 3290 18860 3312
rect 1104 3238 3947 3290
rect 3999 3238 4011 3290
rect 4063 3238 4075 3290
rect 4127 3238 4139 3290
rect 4191 3238 9878 3290
rect 9930 3238 9942 3290
rect 9994 3238 10006 3290
rect 10058 3238 10070 3290
rect 10122 3238 15808 3290
rect 15860 3238 15872 3290
rect 15924 3238 15936 3290
rect 15988 3238 16000 3290
rect 16052 3238 18860 3290
rect 1104 3216 18860 3238
rect 2866 3176 2872 3188
rect 1780 3148 2872 3176
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 1486 2972 1492 2984
rect 1443 2944 1492 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 1486 2932 1492 2944
rect 1544 2932 1550 2984
rect 1780 2981 1808 3148
rect 2866 3136 2872 3148
rect 2924 3176 2930 3188
rect 2924 3148 3464 3176
rect 2924 3136 2930 3148
rect 3436 3108 3464 3148
rect 3510 3136 3516 3188
rect 3568 3176 3574 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 3568 3148 4261 3176
rect 3568 3136 3574 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 7650 3176 7656 3188
rect 5592 3148 7656 3176
rect 5592 3136 5598 3148
rect 7650 3136 7656 3148
rect 7708 3136 7714 3188
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3176 8263 3179
rect 8846 3176 8852 3188
rect 8251 3148 8852 3176
rect 8251 3145 8263 3148
rect 8205 3139 8263 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 9030 3176 9036 3188
rect 8991 3148 9036 3176
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 11054 3176 11060 3188
rect 9416 3148 11060 3176
rect 3786 3108 3792 3120
rect 3436 3080 3792 3108
rect 3786 3068 3792 3080
rect 3844 3068 3850 3120
rect 5718 3108 5724 3120
rect 5460 3080 5724 3108
rect 1854 3000 1860 3052
rect 1912 3040 1918 3052
rect 2774 3040 2780 3052
rect 1912 3012 2780 3040
rect 1912 3000 1918 3012
rect 2774 3000 2780 3012
rect 2832 3000 2838 3052
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3040 4951 3043
rect 5166 3040 5172 3052
rect 4939 3012 5172 3040
rect 4939 3009 4951 3012
rect 4893 3003 4951 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 1765 2975 1823 2981
rect 1765 2941 1777 2975
rect 1811 2941 1823 2975
rect 2130 2972 2136 2984
rect 2091 2944 2136 2972
rect 1765 2935 1823 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 2501 2975 2559 2981
rect 2501 2941 2513 2975
rect 2547 2941 2559 2975
rect 2501 2935 2559 2941
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2972 3019 2975
rect 3050 2972 3056 2984
rect 3007 2944 3056 2972
rect 3007 2941 3019 2944
rect 2961 2935 3019 2941
rect 2516 2904 2544 2935
rect 3050 2932 3056 2944
rect 3108 2932 3114 2984
rect 3326 2932 3332 2984
rect 3384 2972 3390 2984
rect 3513 2975 3571 2981
rect 3513 2972 3525 2975
rect 3384 2944 3525 2972
rect 3384 2932 3390 2944
rect 3513 2941 3525 2944
rect 3559 2941 3571 2975
rect 3513 2935 3571 2941
rect 3881 2975 3939 2981
rect 3881 2941 3893 2975
rect 3927 2972 3939 2975
rect 4798 2972 4804 2984
rect 3927 2944 4804 2972
rect 3927 2941 3939 2944
rect 3881 2935 3939 2941
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5460 2981 5488 3080
rect 5718 3068 5724 3080
rect 5776 3068 5782 3120
rect 6546 3068 6552 3120
rect 6604 3108 6610 3120
rect 7285 3111 7343 3117
rect 7285 3108 7297 3111
rect 6604 3080 7297 3108
rect 6604 3068 6610 3080
rect 7285 3077 7297 3080
rect 7331 3108 7343 3111
rect 8938 3108 8944 3120
rect 7331 3080 8944 3108
rect 7331 3077 7343 3080
rect 7285 3071 7343 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 5626 3040 5632 3052
rect 5587 3012 5632 3040
rect 5626 3000 5632 3012
rect 5684 3040 5690 3052
rect 6457 3043 6515 3049
rect 6457 3040 6469 3043
rect 5684 3012 6469 3040
rect 5684 3000 5690 3012
rect 6457 3009 6469 3012
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 8754 3040 8760 3052
rect 6696 3012 8760 3040
rect 6696 3000 6702 3012
rect 8754 3000 8760 3012
rect 8812 3000 8818 3052
rect 8849 3043 8907 3049
rect 8849 3009 8861 3043
rect 8895 3040 8907 3043
rect 9416 3040 9444 3148
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 12526 3136 12532 3188
rect 12584 3176 12590 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 12584 3148 12725 3176
rect 12584 3136 12590 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 15378 3176 15384 3188
rect 12713 3139 12771 3145
rect 13280 3148 15384 3176
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 9508 3080 10609 3108
rect 9508 3049 9536 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 10597 3071 10655 3077
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 10744 3080 11192 3108
rect 10744 3068 10750 3080
rect 8895 3012 9444 3040
rect 9493 3043 9551 3049
rect 8895 3009 8907 3012
rect 8849 3003 8907 3009
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 11164 3049 11192 3080
rect 11149 3043 11207 3049
rect 9640 3012 9685 3040
rect 10060 3012 10732 3040
rect 9640 3000 9646 3012
rect 5445 2975 5503 2981
rect 5445 2941 5457 2975
rect 5491 2941 5503 2975
rect 6270 2972 6276 2984
rect 6231 2944 6276 2972
rect 5445 2935 5503 2941
rect 6270 2932 6276 2944
rect 6328 2932 6334 2984
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6420 2944 6837 2972
rect 6420 2932 6426 2944
rect 6825 2941 6837 2944
rect 6871 2972 6883 2975
rect 7374 2972 7380 2984
rect 6871 2944 7380 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7650 2972 7656 2984
rect 7611 2944 7656 2972
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 7929 2975 7987 2981
rect 7929 2941 7941 2975
rect 7975 2972 7987 2975
rect 8478 2972 8484 2984
rect 7975 2944 8484 2972
rect 7975 2941 7987 2944
rect 7929 2935 7987 2941
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 9398 2972 9404 2984
rect 9359 2944 9404 2972
rect 9398 2932 9404 2944
rect 9456 2932 9462 2984
rect 10060 2981 10088 3012
rect 10045 2975 10103 2981
rect 10045 2972 10057 2975
rect 9508 2944 10057 2972
rect 3234 2904 3240 2916
rect 2516 2876 3096 2904
rect 3195 2876 3240 2904
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 1670 2796 1676 2848
rect 1728 2836 1734 2848
rect 1949 2839 2007 2845
rect 1949 2836 1961 2839
rect 1728 2808 1961 2836
rect 1728 2796 1734 2808
rect 1949 2805 1961 2808
rect 1995 2805 2007 2839
rect 2314 2836 2320 2848
rect 2275 2808 2320 2836
rect 1949 2799 2007 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 2682 2836 2688 2848
rect 2643 2808 2688 2836
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 3068 2836 3096 2876
rect 3234 2864 3240 2876
rect 3292 2864 3298 2916
rect 4522 2904 4528 2916
rect 3528 2876 4528 2904
rect 3528 2836 3556 2876
rect 4522 2864 4528 2876
rect 4580 2864 4586 2916
rect 4617 2907 4675 2913
rect 4617 2873 4629 2907
rect 4663 2904 4675 2907
rect 7558 2904 7564 2916
rect 4663 2876 5948 2904
rect 7519 2876 7564 2904
rect 4663 2873 4675 2876
rect 4617 2867 4675 2873
rect 3694 2836 3700 2848
rect 3068 2808 3556 2836
rect 3655 2808 3700 2836
rect 3694 2796 3700 2808
rect 3752 2796 3758 2848
rect 4062 2836 4068 2848
rect 4023 2808 4068 2836
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 5077 2839 5135 2845
rect 5077 2836 5089 2839
rect 4755 2808 5089 2836
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 5077 2805 5089 2808
rect 5123 2805 5135 2839
rect 5077 2799 5135 2805
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5920 2845 5948 2876
rect 7558 2864 7564 2876
rect 7616 2864 7622 2916
rect 8294 2864 8300 2916
rect 8352 2904 8358 2916
rect 8665 2907 8723 2913
rect 8665 2904 8677 2907
rect 8352 2876 8677 2904
rect 8352 2864 8358 2876
rect 8665 2873 8677 2876
rect 8711 2873 8723 2907
rect 8665 2867 8723 2873
rect 8754 2864 8760 2916
rect 8812 2904 8818 2916
rect 9508 2904 9536 2944
rect 10045 2941 10057 2944
rect 10091 2941 10103 2975
rect 10226 2972 10232 2984
rect 10139 2944 10232 2972
rect 10045 2935 10103 2941
rect 10226 2932 10232 2944
rect 10284 2972 10290 2984
rect 10594 2972 10600 2984
rect 10284 2944 10600 2972
rect 10284 2932 10290 2944
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10704 2972 10732 3012
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 11149 3003 11207 3009
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 12342 3040 12348 3052
rect 12084 3012 12348 3040
rect 10870 2972 10876 2984
rect 10704 2944 10876 2972
rect 10870 2932 10876 2944
rect 10928 2932 10934 2984
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 11020 2944 11069 2972
rect 11020 2932 11026 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 11793 2975 11851 2981
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 12084 2972 12112 3012
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 13170 3040 13176 3052
rect 13131 3012 13176 3040
rect 13170 3000 13176 3012
rect 13228 3000 13234 3052
rect 11839 2944 12112 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 13081 2975 13139 2981
rect 13081 2972 13093 2975
rect 12492 2944 13093 2972
rect 12492 2932 12498 2944
rect 13081 2941 13093 2944
rect 13127 2972 13139 2975
rect 13280 2972 13308 3148
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 17034 3136 17040 3188
rect 17092 3136 17098 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17368 3148 17417 3176
rect 17368 3136 17374 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17586 3176 17592 3188
rect 17547 3148 17592 3176
rect 17405 3139 17463 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 13998 3108 14004 3120
rect 13556 3080 14004 3108
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3040 13415 3043
rect 13446 3040 13452 3052
rect 13403 3012 13452 3040
rect 13403 3009 13415 3012
rect 13357 3003 13415 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13556 2981 13584 3080
rect 13998 3068 14004 3080
rect 14056 3068 14062 3120
rect 14734 3108 14740 3120
rect 14695 3080 14740 3108
rect 14734 3068 14740 3080
rect 14792 3068 14798 3120
rect 16574 3108 16580 3120
rect 16040 3080 16580 3108
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3009 13783 3043
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 13725 3003 13783 3009
rect 13127 2944 13308 2972
rect 13541 2975 13599 2981
rect 13127 2941 13139 2944
rect 13081 2935 13139 2941
rect 13541 2941 13553 2975
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 8812 2876 9536 2904
rect 9953 2907 10011 2913
rect 8812 2864 8818 2876
rect 9953 2873 9965 2907
rect 9999 2904 10011 2907
rect 10244 2904 10272 2932
rect 9999 2876 10272 2904
rect 9999 2873 10011 2876
rect 9953 2867 10011 2873
rect 10318 2864 10324 2916
rect 10376 2864 10382 2916
rect 10505 2907 10563 2913
rect 10505 2873 10517 2907
rect 10551 2904 10563 2907
rect 10686 2904 10692 2916
rect 10551 2876 10692 2904
rect 10551 2873 10563 2876
rect 10505 2867 10563 2873
rect 10686 2864 10692 2876
rect 10744 2864 10750 2916
rect 13262 2864 13268 2916
rect 13320 2904 13326 2916
rect 13740 2904 13768 3003
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3040 15163 3043
rect 15378 3040 15384 3052
rect 15151 3012 15384 3040
rect 15151 3009 15163 3012
rect 15105 3003 15163 3009
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 16040 3049 16068 3080
rect 16574 3068 16580 3080
rect 16632 3068 16638 3120
rect 17052 3108 17080 3136
rect 17773 3111 17831 3117
rect 17773 3108 17785 3111
rect 17052 3080 17785 3108
rect 17773 3077 17785 3080
rect 17819 3077 17831 3111
rect 17773 3071 17831 3077
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3009 16083 3043
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16025 3003 16083 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 16850 3040 16856 3052
rect 16811 3012 16856 3040
rect 16850 3000 16856 3012
rect 16908 3040 16914 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 16908 3012 17049 3040
rect 16908 3000 16914 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 14148 2944 14193 2972
rect 14148 2932 14154 2944
rect 14642 2932 14648 2984
rect 14700 2972 14706 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 14700 2944 15209 2972
rect 14700 2932 14706 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15562 2932 15568 2984
rect 15620 2972 15626 2984
rect 15749 2975 15807 2981
rect 15749 2972 15761 2975
rect 15620 2944 15761 2972
rect 15620 2932 15626 2944
rect 15749 2941 15761 2944
rect 15795 2941 15807 2975
rect 15749 2935 15807 2941
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 17221 2975 17279 2981
rect 17221 2972 17233 2975
rect 16264 2944 17233 2972
rect 16264 2932 16270 2944
rect 17221 2941 17233 2944
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17368 2944 18061 2972
rect 17368 2932 17374 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 13320 2876 13768 2904
rect 13320 2864 13326 2876
rect 14182 2864 14188 2916
rect 14240 2904 14246 2916
rect 14829 2907 14887 2913
rect 14829 2904 14841 2907
rect 14240 2876 14841 2904
rect 14240 2864 14246 2876
rect 14829 2873 14841 2876
rect 14875 2873 14887 2907
rect 16577 2907 16635 2913
rect 16577 2904 16589 2907
rect 14829 2867 14887 2873
rect 15396 2876 16589 2904
rect 5537 2839 5595 2845
rect 5537 2836 5549 2839
rect 5500 2808 5549 2836
rect 5500 2796 5506 2808
rect 5537 2805 5549 2808
rect 5583 2805 5595 2839
rect 5537 2799 5595 2805
rect 5905 2839 5963 2845
rect 5905 2805 5917 2839
rect 5951 2805 5963 2839
rect 5905 2799 5963 2805
rect 7101 2839 7159 2845
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 7282 2836 7288 2848
rect 7147 2808 7288 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 8573 2839 8631 2845
rect 8573 2805 8585 2839
rect 8619 2836 8631 2839
rect 9766 2836 9772 2848
rect 8619 2808 9772 2836
rect 8619 2805 8631 2808
rect 8573 2799 8631 2805
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 10229 2839 10287 2845
rect 10229 2836 10241 2839
rect 10192 2808 10241 2836
rect 10192 2796 10198 2808
rect 10229 2805 10241 2808
rect 10275 2805 10287 2839
rect 10336 2836 10364 2864
rect 10965 2839 11023 2845
rect 10965 2836 10977 2839
rect 10336 2808 10977 2836
rect 10229 2799 10287 2805
rect 10965 2805 10977 2808
rect 11011 2805 11023 2839
rect 11422 2836 11428 2848
rect 11383 2808 11428 2836
rect 10965 2799 11023 2805
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 12529 2839 12587 2845
rect 12529 2836 12541 2839
rect 11931 2808 12541 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 12529 2805 12541 2808
rect 12575 2836 12587 2839
rect 13630 2836 13636 2848
rect 12575 2808 13636 2836
rect 12575 2805 12587 2808
rect 12529 2799 12587 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 15396 2845 15424 2876
rect 16577 2873 16589 2876
rect 16623 2873 16635 2907
rect 16577 2867 16635 2873
rect 18325 2907 18383 2913
rect 18325 2873 18337 2907
rect 18371 2904 18383 2907
rect 19426 2904 19432 2916
rect 18371 2876 19432 2904
rect 18371 2873 18383 2876
rect 18325 2867 18383 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 15381 2839 15439 2845
rect 15381 2805 15393 2839
rect 15427 2805 15439 2839
rect 15381 2799 15439 2805
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 15841 2839 15899 2845
rect 15841 2836 15853 2839
rect 15528 2808 15853 2836
rect 15528 2796 15534 2808
rect 15841 2805 15853 2808
rect 15887 2805 15899 2839
rect 15841 2799 15899 2805
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16209 2839 16267 2845
rect 16209 2836 16221 2839
rect 16172 2808 16221 2836
rect 16172 2796 16178 2808
rect 16209 2805 16221 2808
rect 16255 2805 16267 2839
rect 16209 2799 16267 2805
rect 1104 2746 18860 2768
rect 1104 2694 6912 2746
rect 6964 2694 6976 2746
rect 7028 2694 7040 2746
rect 7092 2694 7104 2746
rect 7156 2694 12843 2746
rect 12895 2694 12907 2746
rect 12959 2694 12971 2746
rect 13023 2694 13035 2746
rect 13087 2694 18860 2746
rect 1104 2672 18860 2694
rect 1489 2635 1547 2641
rect 1489 2601 1501 2635
rect 1535 2632 1547 2635
rect 1854 2632 1860 2644
rect 1535 2604 1860 2632
rect 1535 2601 1547 2604
rect 1489 2595 1547 2601
rect 1854 2592 1860 2604
rect 1912 2592 1918 2644
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 4430 2632 4436 2644
rect 3568 2604 4436 2632
rect 3568 2592 3574 2604
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 5997 2635 6055 2641
rect 5997 2632 6009 2635
rect 5408 2604 6009 2632
rect 5408 2592 5414 2604
rect 5997 2601 6009 2604
rect 6043 2632 6055 2635
rect 6181 2635 6239 2641
rect 6181 2632 6193 2635
rect 6043 2604 6193 2632
rect 6043 2601 6055 2604
rect 5997 2595 6055 2601
rect 6181 2601 6193 2604
rect 6227 2601 6239 2635
rect 6181 2595 6239 2601
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8294 2632 8300 2644
rect 8067 2604 8300 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8389 2635 8447 2641
rect 8389 2601 8401 2635
rect 8435 2632 8447 2635
rect 8849 2635 8907 2641
rect 8849 2632 8861 2635
rect 8435 2604 8861 2632
rect 8435 2601 8447 2604
rect 8389 2595 8447 2601
rect 8849 2601 8861 2604
rect 8895 2601 8907 2635
rect 8849 2595 8907 2601
rect 8938 2592 8944 2644
rect 8996 2632 9002 2644
rect 9309 2635 9367 2641
rect 9309 2632 9321 2635
rect 8996 2604 9321 2632
rect 8996 2592 9002 2604
rect 9309 2601 9321 2604
rect 9355 2632 9367 2635
rect 10134 2632 10140 2644
rect 9355 2604 10140 2632
rect 9355 2601 9367 2604
rect 9309 2595 9367 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10686 2592 10692 2644
rect 10744 2632 10750 2644
rect 11054 2632 11060 2644
rect 10744 2604 11060 2632
rect 10744 2592 10750 2604
rect 11054 2592 11060 2604
rect 11112 2592 11118 2644
rect 11149 2635 11207 2641
rect 11149 2601 11161 2635
rect 11195 2632 11207 2635
rect 11330 2632 11336 2644
rect 11195 2604 11336 2632
rect 11195 2601 11207 2604
rect 11149 2595 11207 2601
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 11882 2632 11888 2644
rect 11572 2604 11888 2632
rect 11572 2592 11578 2604
rect 11882 2592 11888 2604
rect 11940 2632 11946 2644
rect 11977 2635 12035 2641
rect 11977 2632 11989 2635
rect 11940 2604 11989 2632
rect 11940 2592 11946 2604
rect 11977 2601 11989 2604
rect 12023 2601 12035 2635
rect 12989 2635 13047 2641
rect 12989 2632 13001 2635
rect 11977 2595 12035 2601
rect 12084 2604 13001 2632
rect 5074 2564 5080 2576
rect 4172 2536 5080 2564
rect 1118 2456 1124 2508
rect 1176 2496 1182 2508
rect 1581 2499 1639 2505
rect 1581 2496 1593 2499
rect 1176 2468 1593 2496
rect 1176 2456 1182 2468
rect 1581 2465 1593 2468
rect 1627 2465 1639 2499
rect 1946 2496 1952 2508
rect 1907 2468 1952 2496
rect 1581 2459 1639 2465
rect 1946 2456 1952 2468
rect 2004 2456 2010 2508
rect 2498 2496 2504 2508
rect 2459 2468 2504 2496
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 3418 2496 3424 2508
rect 3379 2468 3424 2496
rect 2869 2459 2927 2465
rect 2130 2428 2136 2440
rect 2091 2400 2136 2428
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 2685 2363 2743 2369
rect 2685 2329 2697 2363
rect 2731 2360 2743 2363
rect 2774 2360 2780 2372
rect 2731 2332 2780 2360
rect 2731 2329 2743 2332
rect 2685 2323 2743 2329
rect 2774 2320 2780 2332
rect 2832 2320 2838 2372
rect 2884 2360 2912 2459
rect 3418 2456 3424 2468
rect 3476 2456 3482 2508
rect 4172 2505 4200 2536
rect 5074 2524 5080 2536
rect 5132 2524 5138 2576
rect 5718 2524 5724 2576
rect 5776 2564 5782 2576
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 5776 2536 5825 2564
rect 5776 2524 5782 2536
rect 5813 2533 5825 2536
rect 5859 2533 5871 2567
rect 5813 2527 5871 2533
rect 8481 2567 8539 2573
rect 8481 2533 8493 2567
rect 8527 2564 8539 2567
rect 8662 2564 8668 2576
rect 8527 2536 8668 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 8662 2524 8668 2536
rect 8720 2524 8726 2576
rect 8754 2524 8760 2576
rect 8812 2564 8818 2576
rect 9217 2567 9275 2573
rect 9217 2564 9229 2567
rect 8812 2536 9229 2564
rect 8812 2524 8818 2536
rect 9217 2533 9229 2536
rect 9263 2533 9275 2567
rect 10226 2564 10232 2576
rect 10187 2536 10232 2564
rect 9217 2527 9275 2533
rect 10226 2524 10232 2536
rect 10284 2524 10290 2576
rect 10321 2567 10379 2573
rect 10321 2533 10333 2567
rect 10367 2564 10379 2567
rect 11422 2564 11428 2576
rect 10367 2536 11428 2564
rect 10367 2533 10379 2536
rect 10321 2527 10379 2533
rect 11422 2524 11428 2536
rect 11480 2524 11486 2576
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 12084 2564 12112 2604
rect 12989 2601 13001 2604
rect 13035 2601 13047 2635
rect 15194 2632 15200 2644
rect 15155 2604 15200 2632
rect 12989 2595 13047 2601
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 17037 2635 17095 2641
rect 17037 2601 17049 2635
rect 17083 2632 17095 2635
rect 17310 2632 17316 2644
rect 17083 2604 17316 2632
rect 17083 2601 17095 2604
rect 17037 2595 17095 2601
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 18138 2592 18144 2644
rect 18196 2632 18202 2644
rect 18417 2635 18475 2641
rect 18417 2632 18429 2635
rect 18196 2604 18429 2632
rect 18196 2592 18202 2604
rect 18417 2601 18429 2604
rect 18463 2601 18475 2635
rect 18417 2595 18475 2601
rect 11756 2536 12112 2564
rect 11756 2524 11762 2536
rect 12158 2524 12164 2576
rect 12216 2564 12222 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 12216 2536 14289 2564
rect 12216 2524 12222 2536
rect 14277 2533 14289 2536
rect 14323 2533 14335 2567
rect 14277 2527 14335 2533
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 17129 2567 17187 2573
rect 17129 2564 17141 2567
rect 15068 2536 17141 2564
rect 15068 2524 15074 2536
rect 17129 2533 17141 2536
rect 17175 2533 17187 2567
rect 17328 2564 17356 2592
rect 17328 2536 17724 2564
rect 17129 2527 17187 2533
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2465 4215 2499
rect 4706 2496 4712 2508
rect 4667 2468 4712 2496
rect 4157 2459 4215 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 5258 2496 5264 2508
rect 5219 2468 5264 2496
rect 5258 2456 5264 2468
rect 5316 2456 5322 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7374 2496 7380 2508
rect 6963 2468 7380 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7374 2456 7380 2468
rect 7432 2456 7438 2508
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 10778 2496 10784 2508
rect 7515 2468 10784 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11054 2456 11060 2508
rect 11112 2496 11118 2508
rect 11885 2499 11943 2505
rect 11885 2496 11897 2499
rect 11112 2468 11897 2496
rect 11112 2456 11118 2468
rect 11885 2465 11897 2468
rect 11931 2465 11943 2499
rect 11885 2459 11943 2465
rect 13354 2456 13360 2508
rect 13412 2496 13418 2508
rect 13449 2499 13507 2505
rect 13449 2496 13461 2499
rect 13412 2468 13461 2496
rect 13412 2456 13418 2468
rect 13449 2465 13461 2468
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 13814 2456 13820 2508
rect 13872 2496 13878 2508
rect 14001 2499 14059 2505
rect 14001 2496 14013 2499
rect 13872 2468 14013 2496
rect 13872 2456 13878 2468
rect 14001 2465 14013 2468
rect 14047 2465 14059 2499
rect 14001 2459 14059 2465
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2496 14611 2499
rect 15102 2496 15108 2508
rect 14599 2468 15108 2496
rect 14599 2465 14611 2468
rect 14553 2459 14611 2465
rect 15102 2456 15108 2468
rect 15160 2456 15166 2508
rect 15286 2456 15292 2508
rect 15344 2496 15350 2508
rect 15473 2499 15531 2505
rect 15473 2496 15485 2499
rect 15344 2468 15485 2496
rect 15344 2456 15350 2468
rect 15473 2465 15485 2468
rect 15519 2465 15531 2499
rect 17144 2496 17172 2527
rect 17696 2505 17724 2536
rect 17313 2499 17371 2505
rect 17313 2496 17325 2499
rect 17144 2468 17325 2496
rect 15473 2459 15531 2465
rect 17313 2465 17325 2468
rect 17359 2465 17371 2499
rect 17313 2459 17371 2465
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2465 17739 2499
rect 17681 2459 17739 2465
rect 3142 2388 3148 2440
rect 3200 2428 3206 2440
rect 3605 2431 3663 2437
rect 3605 2428 3617 2431
rect 3200 2400 3617 2428
rect 3200 2388 3206 2400
rect 3605 2397 3617 2400
rect 3651 2397 3663 2431
rect 3605 2391 3663 2397
rect 4246 2388 4252 2440
rect 4304 2428 4310 2440
rect 4341 2431 4399 2437
rect 4341 2428 4353 2431
rect 4304 2400 4353 2428
rect 4304 2388 4310 2400
rect 4341 2397 4353 2400
rect 4387 2397 4399 2431
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4341 2391 4399 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2428 5595 2431
rect 5810 2428 5816 2440
rect 5583 2400 5816 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6788 2400 7113 2428
rect 6788 2388 6794 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7616 2400 7665 2428
rect 7616 2388 7622 2400
rect 7653 2397 7665 2400
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 2884 2332 3740 2360
rect 1762 2292 1768 2304
rect 1723 2264 1768 2292
rect 1762 2252 1768 2264
rect 1820 2252 1826 2304
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 3329 2295 3387 2301
rect 3329 2261 3341 2295
rect 3375 2292 3387 2295
rect 3510 2292 3516 2304
rect 3375 2264 3516 2292
rect 3375 2261 3387 2264
rect 3329 2255 3387 2261
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 3712 2292 3740 2332
rect 3786 2320 3792 2372
rect 3844 2360 3850 2372
rect 6365 2363 6423 2369
rect 6365 2360 6377 2363
rect 3844 2332 6377 2360
rect 3844 2320 3850 2332
rect 6365 2329 6377 2332
rect 6411 2360 6423 2363
rect 7282 2360 7288 2372
rect 6411 2332 7288 2360
rect 6411 2329 6423 2332
rect 6365 2323 6423 2329
rect 7282 2320 7288 2332
rect 7340 2320 7346 2372
rect 8588 2360 8616 2391
rect 8754 2388 8760 2440
rect 8812 2428 8818 2440
rect 8812 2400 9076 2428
rect 8812 2388 8818 2400
rect 9048 2360 9076 2400
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 9180 2400 9413 2428
rect 9180 2388 9186 2400
rect 9401 2397 9413 2400
rect 9447 2428 9459 2431
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 9447 2400 10425 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 10413 2397 10425 2400
rect 10459 2428 10471 2431
rect 11238 2428 11244 2440
rect 10459 2400 11244 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 11238 2388 11244 2400
rect 11296 2428 11302 2440
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11296 2400 12081 2428
rect 11296 2388 11302 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12434 2428 12440 2440
rect 12395 2400 12440 2428
rect 12069 2391 12127 2397
rect 12434 2388 12440 2400
rect 12492 2388 12498 2440
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 8588 2332 8800 2360
rect 9048 2332 9873 2360
rect 6086 2292 6092 2304
rect 3712 2264 6092 2292
rect 6086 2252 6092 2264
rect 6144 2292 6150 2304
rect 6546 2292 6552 2304
rect 6144 2264 6552 2292
rect 6144 2252 6150 2264
rect 6546 2252 6552 2264
rect 6604 2252 6610 2304
rect 8772 2292 8800 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9861 2323 9919 2329
rect 10689 2363 10747 2369
rect 10689 2329 10701 2363
rect 10735 2360 10747 2363
rect 13096 2360 13124 2391
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 13630 2428 13636 2440
rect 13228 2400 13273 2428
rect 13591 2400 13636 2428
rect 13228 2388 13234 2400
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 10735 2332 13124 2360
rect 10735 2329 10747 2332
rect 10689 2323 10747 2329
rect 13906 2320 13912 2372
rect 13964 2360 13970 2372
rect 14752 2360 14780 2391
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 15657 2431 15715 2437
rect 15657 2428 15669 2431
rect 14884 2400 15669 2428
rect 14884 2388 14890 2400
rect 15657 2397 15669 2400
rect 15703 2397 15715 2431
rect 15657 2391 15715 2397
rect 17862 2388 17868 2440
rect 17920 2428 17926 2440
rect 17957 2431 18015 2437
rect 17957 2428 17969 2431
rect 17920 2400 17969 2428
rect 17920 2388 17926 2400
rect 17957 2397 17969 2400
rect 18003 2397 18015 2431
rect 17957 2391 18015 2397
rect 13964 2332 14780 2360
rect 13964 2320 13970 2332
rect 10410 2292 10416 2304
rect 8772 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 11517 2295 11575 2301
rect 11517 2261 11529 2295
rect 11563 2292 11575 2295
rect 11698 2292 11704 2304
rect 11563 2264 11704 2292
rect 11563 2261 11575 2264
rect 11517 2255 11575 2261
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 12124 2264 12633 2292
rect 12124 2252 12130 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 17494 2292 17500 2304
rect 17455 2264 17500 2292
rect 12621 2255 12679 2261
rect 17494 2252 17500 2264
rect 17552 2252 17558 2304
rect 1104 2202 18860 2224
rect 1104 2150 3947 2202
rect 3999 2150 4011 2202
rect 4063 2150 4075 2202
rect 4127 2150 4139 2202
rect 4191 2150 9878 2202
rect 9930 2150 9942 2202
rect 9994 2150 10006 2202
rect 10058 2150 10070 2202
rect 10122 2150 15808 2202
rect 15860 2150 15872 2202
rect 15924 2150 15936 2202
rect 15988 2150 16000 2202
rect 16052 2150 18860 2202
rect 1104 2128 18860 2150
rect 9766 2048 9772 2100
rect 9824 2088 9830 2100
rect 12066 2088 12072 2100
rect 9824 2060 12072 2088
rect 9824 2048 9830 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 10318 1436 10324 1488
rect 10376 1476 10382 1488
rect 14274 1476 14280 1488
rect 10376 1448 14280 1476
rect 10376 1436 10382 1448
rect 14274 1436 14280 1448
rect 14332 1436 14338 1488
rect 2590 1300 2596 1352
rect 2648 1340 2654 1352
rect 15194 1340 15200 1352
rect 2648 1312 15200 1340
rect 2648 1300 2654 1312
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
rect 15286 1272 15292 1284
rect 12360 1244 15292 1272
rect 3234 1164 3240 1216
rect 3292 1204 3298 1216
rect 12360 1204 12388 1244
rect 15286 1232 15292 1244
rect 15344 1232 15350 1284
rect 3292 1176 12388 1204
rect 3292 1164 3298 1176
rect 11238 1096 11244 1148
rect 11296 1136 11302 1148
rect 13630 1136 13636 1148
rect 11296 1108 13636 1136
rect 11296 1096 11302 1108
rect 13630 1096 13636 1108
rect 13688 1096 13694 1148
<< via1 >>
rect 4068 15172 4120 15224
rect 9404 15172 9456 15224
rect 6912 14662 6964 14714
rect 6976 14662 7028 14714
rect 7040 14662 7092 14714
rect 7104 14662 7156 14714
rect 12843 14662 12895 14714
rect 12907 14662 12959 14714
rect 12971 14662 13023 14714
rect 13035 14662 13087 14714
rect 1400 14603 1452 14612
rect 1400 14569 1409 14603
rect 1409 14569 1443 14603
rect 1443 14569 1452 14603
rect 1400 14560 1452 14569
rect 2044 14424 2096 14476
rect 2872 14424 2924 14476
rect 3700 14424 3752 14476
rect 1768 14399 1820 14408
rect 1768 14365 1777 14399
rect 1777 14365 1811 14399
rect 1811 14365 1820 14399
rect 1768 14356 1820 14365
rect 2320 14399 2372 14408
rect 2320 14365 2329 14399
rect 2329 14365 2363 14399
rect 2363 14365 2372 14399
rect 2320 14356 2372 14365
rect 1952 14288 2004 14340
rect 17316 14288 17368 14340
rect 3792 14220 3844 14272
rect 18052 14220 18104 14272
rect 3947 14118 3999 14170
rect 4011 14118 4063 14170
rect 4075 14118 4127 14170
rect 4139 14118 4191 14170
rect 9878 14118 9930 14170
rect 9942 14118 9994 14170
rect 10006 14118 10058 14170
rect 10070 14118 10122 14170
rect 15808 14118 15860 14170
rect 15872 14118 15924 14170
rect 15936 14118 15988 14170
rect 16000 14118 16052 14170
rect 2964 14016 3016 14068
rect 3792 14016 3844 14068
rect 5908 14016 5960 14068
rect 9404 14059 9456 14068
rect 9404 14025 9413 14059
rect 9413 14025 9447 14059
rect 9447 14025 9456 14059
rect 9404 14016 9456 14025
rect 17408 14016 17460 14068
rect 13912 13948 13964 14000
rect 1676 13880 1728 13932
rect 2780 13880 2832 13932
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 9680 13880 9732 13932
rect 9864 13923 9916 13932
rect 9864 13889 9873 13923
rect 9873 13889 9907 13923
rect 9907 13889 9916 13923
rect 9864 13880 9916 13889
rect 6092 13812 6144 13864
rect 9404 13812 9456 13864
rect 17868 13880 17920 13932
rect 17316 13812 17368 13864
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 17500 13676 17552 13728
rect 6912 13574 6964 13626
rect 6976 13574 7028 13626
rect 7040 13574 7092 13626
rect 7104 13574 7156 13626
rect 12843 13574 12895 13626
rect 12907 13574 12959 13626
rect 12971 13574 13023 13626
rect 13035 13574 13087 13626
rect 1492 13515 1544 13524
rect 1492 13481 1501 13515
rect 1501 13481 1535 13515
rect 1535 13481 1544 13515
rect 1492 13472 1544 13481
rect 17408 13515 17460 13524
rect 17408 13481 17417 13515
rect 17417 13481 17451 13515
rect 17451 13481 17460 13515
rect 17408 13472 17460 13481
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 2320 13311 2372 13320
rect 2320 13277 2329 13311
rect 2329 13277 2363 13311
rect 2363 13277 2372 13311
rect 2320 13268 2372 13277
rect 18052 13268 18104 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 3947 13030 3999 13082
rect 4011 13030 4063 13082
rect 4075 13030 4127 13082
rect 4139 13030 4191 13082
rect 9878 13030 9930 13082
rect 9942 13030 9994 13082
rect 10006 13030 10058 13082
rect 10070 13030 10122 13082
rect 15808 13030 15860 13082
rect 15872 13030 15924 13082
rect 15936 13030 15988 13082
rect 16000 13030 16052 13082
rect 9680 12928 9732 12980
rect 3976 12656 4028 12708
rect 5908 12656 5960 12708
rect 18604 12656 18656 12708
rect 9588 12588 9640 12640
rect 15752 12588 15804 12640
rect 6912 12486 6964 12538
rect 6976 12486 7028 12538
rect 7040 12486 7092 12538
rect 7104 12486 7156 12538
rect 12843 12486 12895 12538
rect 12907 12486 12959 12538
rect 12971 12486 13023 12538
rect 13035 12486 13087 12538
rect 6736 12384 6788 12436
rect 16948 12384 17000 12436
rect 9220 12316 9272 12368
rect 11060 12316 11112 12368
rect 3056 12248 3108 12300
rect 3700 12248 3752 12300
rect 10968 12248 11020 12300
rect 3424 12180 3476 12232
rect 10140 12180 10192 12232
rect 10324 12223 10376 12232
rect 10324 12189 10333 12223
rect 10333 12189 10367 12223
rect 10367 12189 10376 12223
rect 10324 12180 10376 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 10600 12180 10652 12232
rect 15752 12180 15804 12232
rect 3700 12112 3752 12164
rect 15200 12112 15252 12164
rect 7748 12044 7800 12096
rect 12072 12044 12124 12096
rect 3947 11942 3999 11994
rect 4011 11942 4063 11994
rect 4075 11942 4127 11994
rect 4139 11942 4191 11994
rect 9878 11942 9930 11994
rect 9942 11942 9994 11994
rect 10006 11942 10058 11994
rect 10070 11942 10122 11994
rect 15808 11942 15860 11994
rect 15872 11942 15924 11994
rect 15936 11942 15988 11994
rect 16000 11942 16052 11994
rect 3792 11840 3844 11892
rect 7932 11840 7984 11892
rect 10324 11883 10376 11892
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 10968 11840 11020 11892
rect 10048 11772 10100 11824
rect 3608 11704 3660 11756
rect 7564 11704 7616 11756
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 10784 11747 10836 11756
rect 7656 11704 7708 11713
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 10968 11747 11020 11756
rect 10968 11713 10977 11747
rect 10977 11713 11011 11747
rect 11011 11713 11020 11747
rect 12164 11840 12216 11892
rect 13912 11840 13964 11892
rect 10968 11704 11020 11713
rect 8116 11636 8168 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 10508 11636 10560 11688
rect 11612 11636 11664 11688
rect 17960 11840 18012 11892
rect 18144 11883 18196 11892
rect 18144 11849 18153 11883
rect 18153 11849 18187 11883
rect 18187 11849 18196 11883
rect 18144 11840 18196 11849
rect 18420 11883 18472 11892
rect 18420 11849 18429 11883
rect 18429 11849 18463 11883
rect 18463 11849 18472 11883
rect 18420 11840 18472 11849
rect 14464 11772 14516 11824
rect 16304 11772 16356 11824
rect 14372 11704 14424 11756
rect 18236 11704 18288 11756
rect 14924 11636 14976 11688
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 2044 11500 2096 11552
rect 2412 11543 2464 11552
rect 2412 11509 2421 11543
rect 2421 11509 2455 11543
rect 2455 11509 2464 11543
rect 7288 11568 7340 11620
rect 2412 11500 2464 11509
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 6736 11500 6788 11552
rect 7380 11500 7432 11552
rect 7748 11500 7800 11552
rect 10048 11568 10100 11620
rect 10140 11611 10192 11620
rect 10140 11577 10149 11611
rect 10149 11577 10183 11611
rect 10183 11577 10192 11611
rect 10140 11568 10192 11577
rect 15200 11568 15252 11620
rect 9772 11543 9824 11552
rect 9772 11509 9781 11543
rect 9781 11509 9815 11543
rect 9815 11509 9824 11543
rect 9772 11500 9824 11509
rect 10232 11500 10284 11552
rect 11244 11500 11296 11552
rect 11336 11500 11388 11552
rect 11704 11500 11756 11552
rect 15752 11500 15804 11552
rect 17684 11500 17736 11552
rect 6912 11398 6964 11450
rect 6976 11398 7028 11450
rect 7040 11398 7092 11450
rect 7104 11398 7156 11450
rect 12843 11398 12895 11450
rect 12907 11398 12959 11450
rect 12971 11398 13023 11450
rect 13035 11398 13087 11450
rect 2228 11296 2280 11348
rect 2504 11271 2556 11280
rect 2504 11237 2538 11271
rect 2538 11237 2556 11271
rect 2504 11228 2556 11237
rect 3700 11271 3752 11280
rect 3700 11237 3709 11271
rect 3709 11237 3743 11271
rect 3743 11237 3752 11271
rect 3700 11228 3752 11237
rect 6276 11296 6328 11348
rect 11336 11296 11388 11348
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 12072 11339 12124 11348
rect 12072 11305 12081 11339
rect 12081 11305 12115 11339
rect 12115 11305 12124 11339
rect 12072 11296 12124 11305
rect 12164 11296 12216 11348
rect 15568 11296 15620 11348
rect 15752 11296 15804 11348
rect 18420 11296 18472 11348
rect 6736 11160 6788 11212
rect 3792 11092 3844 11144
rect 6828 11092 6880 11144
rect 7380 11228 7432 11280
rect 10968 11228 11020 11280
rect 11796 11228 11848 11280
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 8024 11203 8076 11212
rect 8024 11169 8033 11203
rect 8033 11169 8067 11203
rect 8067 11169 8076 11203
rect 9220 11203 9272 11212
rect 8024 11160 8076 11169
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 11428 11160 11480 11212
rect 7656 11092 7708 11144
rect 8208 11092 8260 11144
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 11612 11092 11664 11144
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 3516 11024 3568 11076
rect 4804 11024 4856 11076
rect 7104 11024 7156 11076
rect 8300 11024 8352 11076
rect 1676 10999 1728 11008
rect 1676 10965 1685 10999
rect 1685 10965 1719 10999
rect 1719 10965 1728 10999
rect 1676 10956 1728 10965
rect 1860 10999 1912 11008
rect 1860 10965 1869 10999
rect 1869 10965 1903 10999
rect 1903 10965 1912 10999
rect 1860 10956 1912 10965
rect 2136 10999 2188 11008
rect 2136 10965 2145 10999
rect 2145 10965 2179 10999
rect 2179 10965 2188 10999
rect 2136 10956 2188 10965
rect 3608 10999 3660 11008
rect 3608 10965 3617 10999
rect 3617 10965 3651 10999
rect 3651 10965 3660 10999
rect 3608 10956 3660 10965
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 8116 10956 8168 11008
rect 8576 10956 8628 11008
rect 11520 10956 11572 11008
rect 12072 11024 12124 11076
rect 12348 11092 12400 11144
rect 13176 11228 13228 11280
rect 14464 11228 14516 11280
rect 12716 11024 12768 11076
rect 14188 11024 14240 11076
rect 16212 11228 16264 11280
rect 16948 11271 17000 11280
rect 16948 11237 16957 11271
rect 16957 11237 16991 11271
rect 16991 11237 17000 11271
rect 16948 11228 17000 11237
rect 17224 11271 17276 11280
rect 17224 11237 17233 11271
rect 17233 11237 17267 11271
rect 17267 11237 17276 11271
rect 17224 11228 17276 11237
rect 14924 11160 14976 11212
rect 15384 11160 15436 11212
rect 18144 11228 18196 11280
rect 17868 11203 17920 11212
rect 14464 10956 14516 11008
rect 15108 11092 15160 11144
rect 14832 11024 14884 11076
rect 15016 11067 15068 11076
rect 15016 11033 15025 11067
rect 15025 11033 15059 11067
rect 15059 11033 15068 11067
rect 15016 11024 15068 11033
rect 14924 10956 14976 11008
rect 17868 11169 17877 11203
rect 17877 11169 17911 11203
rect 17911 11169 17920 11203
rect 17868 11160 17920 11169
rect 16580 10956 16632 11008
rect 16856 11024 16908 11076
rect 17500 11067 17552 11076
rect 17500 11033 17509 11067
rect 17509 11033 17543 11067
rect 17543 11033 17552 11067
rect 17500 11024 17552 11033
rect 17132 10956 17184 11008
rect 3947 10854 3999 10906
rect 4011 10854 4063 10906
rect 4075 10854 4127 10906
rect 4139 10854 4191 10906
rect 9878 10854 9930 10906
rect 9942 10854 9994 10906
rect 10006 10854 10058 10906
rect 10070 10854 10122 10906
rect 15808 10854 15860 10906
rect 15872 10854 15924 10906
rect 15936 10854 15988 10906
rect 16000 10854 16052 10906
rect 2044 10752 2096 10804
rect 2412 10752 2464 10804
rect 4896 10752 4948 10804
rect 6368 10752 6420 10804
rect 7564 10752 7616 10804
rect 8484 10752 8536 10804
rect 1860 10659 1912 10668
rect 1860 10625 1869 10659
rect 1869 10625 1903 10659
rect 1903 10625 1912 10659
rect 1860 10616 1912 10625
rect 2504 10616 2556 10668
rect 2964 10616 3016 10668
rect 3608 10616 3660 10668
rect 3792 10616 3844 10668
rect 2136 10548 2188 10600
rect 4528 10548 4580 10600
rect 4712 10548 4764 10600
rect 6828 10684 6880 10736
rect 12164 10752 12216 10804
rect 12440 10752 12492 10804
rect 14924 10752 14976 10804
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 12256 10684 12308 10736
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 6276 10548 6328 10557
rect 10508 10616 10560 10668
rect 10968 10659 11020 10668
rect 10968 10625 10977 10659
rect 10977 10625 11011 10659
rect 11011 10625 11020 10659
rect 10968 10616 11020 10625
rect 11612 10616 11664 10668
rect 7104 10591 7156 10600
rect 7104 10557 7138 10591
rect 7138 10557 7156 10591
rect 3240 10480 3292 10532
rect 5080 10480 5132 10532
rect 6552 10480 6604 10532
rect 7104 10548 7156 10557
rect 8300 10548 8352 10600
rect 9864 10548 9916 10600
rect 11888 10548 11940 10600
rect 6920 10480 6972 10532
rect 8852 10480 8904 10532
rect 9680 10480 9732 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 2596 10412 2648 10464
rect 2780 10412 2832 10464
rect 4620 10412 4672 10464
rect 5356 10455 5408 10464
rect 5356 10421 5365 10455
rect 5365 10421 5399 10455
rect 5399 10421 5408 10455
rect 5356 10412 5408 10421
rect 12256 10523 12308 10532
rect 12256 10489 12265 10523
rect 12265 10489 12299 10523
rect 12299 10489 12308 10523
rect 12256 10480 12308 10489
rect 13268 10480 13320 10532
rect 17224 10752 17276 10804
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 17868 10616 17920 10668
rect 15108 10548 15160 10600
rect 14740 10480 14792 10532
rect 18144 10548 18196 10600
rect 16580 10480 16632 10532
rect 16672 10480 16724 10532
rect 10692 10455 10744 10464
rect 10692 10421 10701 10455
rect 10701 10421 10735 10455
rect 10735 10421 10744 10455
rect 10692 10412 10744 10421
rect 10784 10455 10836 10464
rect 10784 10421 10793 10455
rect 10793 10421 10827 10455
rect 10827 10421 10836 10455
rect 10784 10412 10836 10421
rect 11520 10412 11572 10464
rect 12072 10412 12124 10464
rect 15292 10455 15344 10464
rect 15292 10421 15301 10455
rect 15301 10421 15335 10455
rect 15335 10421 15344 10455
rect 15292 10412 15344 10421
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 16764 10412 16816 10464
rect 17224 10412 17276 10464
rect 17868 10412 17920 10464
rect 18420 10455 18472 10464
rect 18420 10421 18429 10455
rect 18429 10421 18463 10455
rect 18463 10421 18472 10455
rect 18420 10412 18472 10421
rect 6912 10310 6964 10362
rect 6976 10310 7028 10362
rect 7040 10310 7092 10362
rect 7104 10310 7156 10362
rect 12843 10310 12895 10362
rect 12907 10310 12959 10362
rect 12971 10310 13023 10362
rect 13035 10310 13087 10362
rect 1768 10208 1820 10260
rect 3240 10208 3292 10260
rect 4712 10251 4764 10260
rect 4712 10217 4721 10251
rect 4721 10217 4755 10251
rect 4755 10217 4764 10251
rect 4712 10208 4764 10217
rect 2044 10140 2096 10192
rect 2596 10140 2648 10192
rect 3700 10140 3752 10192
rect 4252 10140 4304 10192
rect 3516 10072 3568 10124
rect 4344 10072 4396 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2964 10004 3016 10056
rect 4436 10004 4488 10056
rect 4620 10072 4672 10124
rect 5540 10208 5592 10260
rect 9864 10251 9916 10260
rect 5448 10140 5500 10192
rect 6828 10140 6880 10192
rect 7564 10140 7616 10192
rect 8852 10140 8904 10192
rect 5540 10115 5592 10124
rect 5540 10081 5549 10115
rect 5549 10081 5583 10115
rect 5583 10081 5592 10115
rect 5540 10072 5592 10081
rect 6276 10072 6328 10124
rect 7472 10115 7524 10124
rect 7472 10081 7481 10115
rect 7481 10081 7515 10115
rect 7515 10081 7524 10115
rect 7472 10072 7524 10081
rect 7656 10072 7708 10124
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 4712 10004 4764 10056
rect 5080 10004 5132 10056
rect 5264 10004 5316 10056
rect 2688 9936 2740 9988
rect 3240 9936 3292 9988
rect 5356 9936 5408 9988
rect 6644 10004 6696 10056
rect 6552 9936 6604 9988
rect 2964 9868 3016 9920
rect 3424 9868 3476 9920
rect 5540 9868 5592 9920
rect 6736 9868 6788 9920
rect 9312 10004 9364 10056
rect 9864 10217 9873 10251
rect 9873 10217 9907 10251
rect 9907 10217 9916 10251
rect 9864 10208 9916 10217
rect 10692 10251 10744 10260
rect 10692 10217 10701 10251
rect 10701 10217 10735 10251
rect 10735 10217 10744 10251
rect 10692 10208 10744 10217
rect 11060 10251 11112 10260
rect 11060 10217 11069 10251
rect 11069 10217 11103 10251
rect 11103 10217 11112 10251
rect 11060 10208 11112 10217
rect 16212 10208 16264 10260
rect 16488 10208 16540 10260
rect 16764 10251 16816 10260
rect 16764 10217 16773 10251
rect 16773 10217 16807 10251
rect 16807 10217 16816 10251
rect 16764 10208 16816 10217
rect 17132 10251 17184 10260
rect 17132 10217 17141 10251
rect 17141 10217 17175 10251
rect 17175 10217 17184 10251
rect 17132 10208 17184 10217
rect 17960 10208 18012 10260
rect 18696 10208 18748 10260
rect 10048 10140 10100 10192
rect 11336 10072 11388 10124
rect 10048 10004 10100 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 9128 9936 9180 9988
rect 9496 9936 9548 9988
rect 9956 9936 10008 9988
rect 10968 9936 11020 9988
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 10232 9868 10284 9920
rect 10508 9868 10560 9920
rect 13084 10140 13136 10192
rect 16580 10140 16632 10192
rect 12164 10115 12216 10124
rect 12164 10081 12198 10115
rect 12198 10081 12216 10115
rect 12164 10072 12216 10081
rect 14556 10072 14608 10124
rect 16028 10072 16080 10124
rect 17776 10072 17828 10124
rect 18420 10072 18472 10124
rect 11888 10047 11940 10056
rect 11888 10013 11897 10047
rect 11897 10013 11931 10047
rect 11931 10013 11940 10047
rect 11888 10004 11940 10013
rect 14740 10047 14792 10056
rect 13360 9936 13412 9988
rect 13728 9936 13780 9988
rect 13268 9911 13320 9920
rect 13268 9877 13277 9911
rect 13277 9877 13311 9911
rect 13311 9877 13320 9911
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 15108 10004 15160 10056
rect 16580 9936 16632 9988
rect 13268 9868 13320 9877
rect 14004 9868 14056 9920
rect 15016 9911 15068 9920
rect 15016 9877 15025 9911
rect 15025 9877 15059 9911
rect 15059 9877 15068 9911
rect 15016 9868 15068 9877
rect 15660 9868 15712 9920
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 17592 9911 17644 9920
rect 17592 9877 17601 9911
rect 17601 9877 17635 9911
rect 17635 9877 17644 9911
rect 17592 9868 17644 9877
rect 17960 9868 18012 9920
rect 18236 9868 18288 9920
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 3947 9766 3999 9818
rect 4011 9766 4063 9818
rect 4075 9766 4127 9818
rect 4139 9766 4191 9818
rect 9878 9766 9930 9818
rect 9942 9766 9994 9818
rect 10006 9766 10058 9818
rect 10070 9766 10122 9818
rect 15808 9766 15860 9818
rect 15872 9766 15924 9818
rect 15936 9766 15988 9818
rect 16000 9766 16052 9818
rect 3792 9664 3844 9716
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 2964 9571 3016 9580
rect 2780 9528 2832 9537
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 5172 9664 5224 9716
rect 5264 9664 5316 9716
rect 6276 9707 6328 9716
rect 6276 9673 6285 9707
rect 6285 9673 6319 9707
rect 6319 9673 6328 9707
rect 6276 9664 6328 9673
rect 4344 9639 4396 9648
rect 4344 9605 4353 9639
rect 4353 9605 4387 9639
rect 4387 9605 4396 9639
rect 4344 9596 4396 9605
rect 4436 9596 4488 9648
rect 5816 9596 5868 9648
rect 7472 9664 7524 9716
rect 10324 9664 10376 9716
rect 10784 9664 10836 9716
rect 12164 9664 12216 9716
rect 13728 9707 13780 9716
rect 8208 9639 8260 9648
rect 4068 9528 4120 9580
rect 5080 9528 5132 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 1952 9460 2004 9512
rect 6276 9460 6328 9512
rect 6552 9460 6604 9512
rect 6920 9460 6972 9512
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 3240 9392 3292 9444
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2228 9324 2280 9333
rect 2412 9324 2464 9376
rect 3976 9367 4028 9376
rect 3976 9333 3985 9367
rect 3985 9333 4019 9367
rect 4019 9333 4028 9367
rect 4344 9392 4396 9444
rect 6000 9392 6052 9444
rect 6644 9392 6696 9444
rect 7380 9460 7432 9512
rect 8208 9605 8217 9639
rect 8217 9605 8251 9639
rect 8251 9605 8260 9639
rect 8208 9596 8260 9605
rect 9680 9639 9732 9648
rect 9680 9605 9689 9639
rect 9689 9605 9723 9639
rect 9723 9605 9732 9639
rect 9680 9596 9732 9605
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 10140 9528 10192 9580
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 13084 9596 13136 9648
rect 10968 9528 11020 9580
rect 13268 9528 13320 9580
rect 13728 9673 13737 9707
rect 13737 9673 13771 9707
rect 13771 9673 13780 9707
rect 13728 9664 13780 9673
rect 13820 9664 13872 9716
rect 14464 9664 14516 9716
rect 14740 9664 14792 9716
rect 15016 9664 15068 9716
rect 16120 9664 16172 9716
rect 17408 9664 17460 9716
rect 13912 9596 13964 9648
rect 14556 9639 14608 9648
rect 14556 9605 14565 9639
rect 14565 9605 14599 9639
rect 14599 9605 14608 9639
rect 14556 9596 14608 9605
rect 15200 9596 15252 9648
rect 16580 9596 16632 9648
rect 16672 9596 16724 9648
rect 15016 9528 15068 9580
rect 9404 9460 9456 9512
rect 9680 9392 9732 9444
rect 3976 9324 4028 9333
rect 4436 9324 4488 9376
rect 4620 9324 4672 9376
rect 4988 9324 5040 9376
rect 5264 9324 5316 9376
rect 5448 9324 5500 9376
rect 5816 9324 5868 9376
rect 9036 9324 9088 9376
rect 10600 9392 10652 9444
rect 10324 9324 10376 9376
rect 17684 9596 17736 9648
rect 15292 9528 15344 9580
rect 17316 9571 17368 9580
rect 17316 9537 17325 9571
rect 17325 9537 17359 9571
rect 17359 9537 17368 9571
rect 17316 9528 17368 9537
rect 17408 9528 17460 9580
rect 11060 9367 11112 9376
rect 11060 9333 11069 9367
rect 11069 9333 11103 9367
rect 11103 9333 11112 9367
rect 11060 9324 11112 9333
rect 11612 9324 11664 9376
rect 11888 9367 11940 9376
rect 11888 9333 11897 9367
rect 11897 9333 11931 9367
rect 11931 9333 11940 9367
rect 11888 9324 11940 9333
rect 12532 9324 12584 9376
rect 17776 9460 17828 9512
rect 18420 9460 18472 9512
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 13360 9324 13412 9376
rect 16764 9392 16816 9444
rect 16948 9392 17000 9444
rect 17316 9392 17368 9444
rect 17960 9392 18012 9444
rect 14096 9367 14148 9376
rect 14096 9333 14105 9367
rect 14105 9333 14139 9367
rect 14139 9333 14148 9367
rect 14096 9324 14148 9333
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14832 9324 14884 9376
rect 15936 9367 15988 9376
rect 15936 9333 15945 9367
rect 15945 9333 15979 9367
rect 15979 9333 15988 9367
rect 15936 9324 15988 9333
rect 16120 9324 16172 9376
rect 16304 9324 16356 9376
rect 17776 9367 17828 9376
rect 17776 9333 17785 9367
rect 17785 9333 17819 9367
rect 17819 9333 17828 9367
rect 17776 9324 17828 9333
rect 18236 9324 18288 9376
rect 6912 9222 6964 9274
rect 6976 9222 7028 9274
rect 7040 9222 7092 9274
rect 7104 9222 7156 9274
rect 12843 9222 12895 9274
rect 12907 9222 12959 9274
rect 12971 9222 13023 9274
rect 13035 9222 13087 9274
rect 1492 9120 1544 9172
rect 2412 9120 2464 9172
rect 4160 9120 4212 9172
rect 4988 9120 5040 9172
rect 5356 9120 5408 9172
rect 6000 9120 6052 9172
rect 6368 9120 6420 9172
rect 6736 9163 6788 9172
rect 6736 9129 6745 9163
rect 6745 9129 6779 9163
rect 6779 9129 6788 9163
rect 6736 9120 6788 9129
rect 9404 9163 9456 9172
rect 2964 9052 3016 9104
rect 3424 9095 3476 9104
rect 3424 9061 3433 9095
rect 3433 9061 3467 9095
rect 3467 9061 3476 9095
rect 3424 9052 3476 9061
rect 3976 9052 4028 9104
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 8024 9095 8076 9104
rect 8024 9061 8033 9095
rect 8033 9061 8067 9095
rect 8067 9061 8076 9095
rect 8024 9052 8076 9061
rect 10968 9120 11020 9172
rect 11428 9120 11480 9172
rect 11888 9120 11940 9172
rect 12072 9120 12124 9172
rect 9772 9052 9824 9104
rect 10232 9052 10284 9104
rect 12532 9052 12584 9104
rect 1400 8984 1452 9036
rect 2780 8984 2832 9036
rect 3792 8984 3844 9036
rect 5816 8984 5868 9036
rect 6184 8984 6236 9036
rect 7656 8984 7708 9036
rect 7932 9027 7984 9036
rect 7932 8993 7941 9027
rect 7941 8993 7975 9027
rect 7975 8993 7984 9027
rect 7932 8984 7984 8993
rect 8852 9027 8904 9036
rect 3148 8916 3200 8968
rect 3424 8916 3476 8968
rect 3700 8916 3752 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 4436 8916 4488 8968
rect 4620 8916 4672 8968
rect 7380 8916 7432 8968
rect 8208 8959 8260 8968
rect 8208 8925 8217 8959
rect 8217 8925 8251 8959
rect 8251 8925 8260 8959
rect 8208 8916 8260 8925
rect 8852 8993 8861 9027
rect 8861 8993 8895 9027
rect 8895 8993 8904 9027
rect 8852 8984 8904 8993
rect 8392 8916 8444 8968
rect 9588 8984 9640 9036
rect 10508 8984 10560 9036
rect 11152 8984 11204 9036
rect 9128 8959 9180 8968
rect 9128 8925 9137 8959
rect 9137 8925 9171 8959
rect 9171 8925 9180 8959
rect 9128 8916 9180 8925
rect 11520 8916 11572 8968
rect 2688 8848 2740 8900
rect 4068 8848 4120 8900
rect 4712 8848 4764 8900
rect 1124 8780 1176 8832
rect 3148 8823 3200 8832
rect 3148 8789 3157 8823
rect 3157 8789 3191 8823
rect 3191 8789 3200 8823
rect 3148 8780 3200 8789
rect 3608 8780 3660 8832
rect 4252 8780 4304 8832
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 8576 8780 8628 8832
rect 8852 8780 8904 8832
rect 9496 8780 9548 8832
rect 11336 8848 11388 8900
rect 13084 8984 13136 9036
rect 12164 8916 12216 8968
rect 13176 8848 13228 8900
rect 10876 8780 10928 8832
rect 10968 8780 11020 8832
rect 14832 9120 14884 9172
rect 15016 9163 15068 9172
rect 15016 9129 15025 9163
rect 15025 9129 15059 9163
rect 15059 9129 15068 9163
rect 15016 9120 15068 9129
rect 13820 9052 13872 9104
rect 14096 9052 14148 9104
rect 14280 9052 14332 9104
rect 14556 9052 14608 9104
rect 15936 9120 15988 9172
rect 16488 9120 16540 9172
rect 17592 9120 17644 9172
rect 15660 9095 15712 9104
rect 15660 9061 15694 9095
rect 15694 9061 15712 9095
rect 15660 9052 15712 9061
rect 17500 9052 17552 9104
rect 18420 9052 18472 9104
rect 17960 8984 18012 9036
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 14280 8780 14332 8832
rect 15108 8780 15160 8832
rect 17224 8916 17276 8968
rect 17868 8848 17920 8900
rect 16304 8780 16356 8832
rect 16580 8780 16632 8832
rect 16948 8823 17000 8832
rect 16948 8789 16957 8823
rect 16957 8789 16991 8823
rect 16991 8789 17000 8823
rect 16948 8780 17000 8789
rect 17592 8780 17644 8832
rect 3947 8678 3999 8730
rect 4011 8678 4063 8730
rect 4075 8678 4127 8730
rect 4139 8678 4191 8730
rect 9878 8678 9930 8730
rect 9942 8678 9994 8730
rect 10006 8678 10058 8730
rect 10070 8678 10122 8730
rect 15808 8678 15860 8730
rect 15872 8678 15924 8730
rect 15936 8678 15988 8730
rect 16000 8678 16052 8730
rect 2228 8576 2280 8628
rect 5816 8576 5868 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 7748 8576 7800 8628
rect 9680 8576 9732 8628
rect 10416 8576 10468 8628
rect 9404 8508 9456 8560
rect 11152 8576 11204 8628
rect 11612 8576 11664 8628
rect 11796 8576 11848 8628
rect 13268 8576 13320 8628
rect 14096 8619 14148 8628
rect 14096 8585 14105 8619
rect 14105 8585 14139 8619
rect 14139 8585 14148 8619
rect 14096 8576 14148 8585
rect 16120 8619 16172 8628
rect 16120 8585 16129 8619
rect 16129 8585 16163 8619
rect 16163 8585 16172 8619
rect 16120 8576 16172 8585
rect 12532 8508 12584 8560
rect 13360 8508 13412 8560
rect 17500 8576 17552 8628
rect 1400 8440 1452 8492
rect 9496 8440 9548 8492
rect 9864 8440 9916 8492
rect 3792 8372 3844 8424
rect 5908 8372 5960 8424
rect 6552 8372 6604 8424
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 9128 8372 9180 8424
rect 10324 8415 10376 8424
rect 10324 8381 10333 8415
rect 10333 8381 10367 8415
rect 10367 8381 10376 8415
rect 10324 8372 10376 8381
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 10600 8372 10652 8424
rect 11060 8372 11112 8424
rect 13176 8440 13228 8492
rect 13820 8483 13872 8492
rect 13820 8449 13829 8483
rect 13829 8449 13863 8483
rect 13863 8449 13872 8483
rect 13820 8440 13872 8449
rect 2688 8304 2740 8356
rect 4988 8304 5040 8356
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 7288 8304 7340 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3608 8236 3660 8288
rect 3792 8236 3844 8288
rect 4436 8279 4488 8288
rect 4436 8245 4445 8279
rect 4445 8245 4479 8279
rect 4479 8245 4488 8279
rect 4436 8236 4488 8245
rect 5724 8236 5776 8288
rect 7380 8236 7432 8288
rect 8852 8236 8904 8288
rect 10232 8304 10284 8356
rect 9680 8279 9732 8288
rect 9680 8245 9689 8279
rect 9689 8245 9723 8279
rect 9723 8245 9732 8279
rect 9680 8236 9732 8245
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 11336 8304 11388 8356
rect 12164 8236 12216 8288
rect 12256 8236 12308 8288
rect 12624 8236 12676 8288
rect 13176 8304 13228 8356
rect 13728 8304 13780 8356
rect 14280 8372 14332 8424
rect 15016 8372 15068 8424
rect 18788 8508 18840 8560
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 16580 8415 16632 8424
rect 16580 8381 16614 8415
rect 16614 8381 16632 8415
rect 16580 8372 16632 8381
rect 16856 8372 16908 8424
rect 14464 8304 14516 8356
rect 16672 8304 16724 8356
rect 13544 8279 13596 8288
rect 13544 8245 13553 8279
rect 13553 8245 13587 8279
rect 13587 8245 13596 8279
rect 13544 8236 13596 8245
rect 16396 8236 16448 8288
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 17960 8236 18012 8288
rect 18144 8236 18196 8288
rect 6912 8134 6964 8186
rect 6976 8134 7028 8186
rect 7040 8134 7092 8186
rect 7104 8134 7156 8186
rect 12843 8134 12895 8186
rect 12907 8134 12959 8186
rect 12971 8134 13023 8186
rect 13035 8134 13087 8186
rect 2780 8032 2832 8084
rect 3056 8075 3108 8084
rect 3056 8041 3065 8075
rect 3065 8041 3099 8075
rect 3099 8041 3108 8075
rect 3056 8032 3108 8041
rect 3884 8075 3936 8084
rect 3884 8041 3893 8075
rect 3893 8041 3927 8075
rect 3927 8041 3936 8075
rect 3884 8032 3936 8041
rect 4252 8032 4304 8084
rect 4896 8032 4948 8084
rect 7380 8075 7432 8084
rect 2412 7964 2464 8016
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 8024 8032 8076 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 10600 8032 10652 8084
rect 11796 8032 11848 8084
rect 5356 7964 5408 8016
rect 7196 7964 7248 8016
rect 2596 7896 2648 7948
rect 5908 7939 5960 7948
rect 2688 7828 2740 7880
rect 2872 7828 2924 7880
rect 4528 7871 4580 7880
rect 4528 7837 4537 7871
rect 4537 7837 4571 7871
rect 4571 7837 4580 7871
rect 4528 7828 4580 7837
rect 5908 7905 5917 7939
rect 5917 7905 5951 7939
rect 5951 7905 5960 7939
rect 5908 7896 5960 7905
rect 7380 7896 7432 7948
rect 2964 7760 3016 7812
rect 5172 7760 5224 7812
rect 5724 7828 5776 7880
rect 7104 7828 7156 7880
rect 10508 7964 10560 8016
rect 9312 7896 9364 7948
rect 9496 7896 9548 7948
rect 8576 7871 8628 7880
rect 8576 7837 8585 7871
rect 8585 7837 8619 7871
rect 8619 7837 8628 7871
rect 8760 7871 8812 7880
rect 8576 7828 8628 7837
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 12624 8032 12676 8084
rect 13912 8075 13964 8084
rect 13912 8041 13921 8075
rect 13921 8041 13955 8075
rect 13955 8041 13964 8075
rect 13912 8032 13964 8041
rect 14188 8032 14240 8084
rect 14740 8032 14792 8084
rect 16948 8032 17000 8084
rect 17500 8032 17552 8084
rect 12808 7964 12860 8016
rect 15384 7964 15436 8016
rect 16580 7964 16632 8016
rect 11888 7896 11940 7905
rect 13728 7896 13780 7948
rect 16856 7939 16908 7948
rect 7288 7803 7340 7812
rect 7288 7769 7297 7803
rect 7297 7769 7331 7803
rect 7331 7769 7340 7803
rect 7288 7760 7340 7769
rect 8208 7760 8260 7812
rect 11336 7828 11388 7880
rect 12164 7828 12216 7880
rect 13636 7828 13688 7880
rect 13912 7828 13964 7880
rect 13820 7803 13872 7812
rect 1676 7735 1728 7744
rect 1676 7701 1685 7735
rect 1685 7701 1719 7735
rect 1719 7701 1728 7735
rect 1676 7692 1728 7701
rect 2228 7692 2280 7744
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3608 7735 3660 7744
rect 3608 7701 3617 7735
rect 3617 7701 3651 7735
rect 3651 7701 3660 7735
rect 3608 7692 3660 7701
rect 4252 7692 4304 7744
rect 5632 7692 5684 7744
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 8484 7692 8536 7744
rect 8852 7692 8904 7744
rect 10324 7692 10376 7744
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 13820 7769 13829 7803
rect 13829 7769 13863 7803
rect 13863 7769 13872 7803
rect 15660 7828 15712 7880
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 18144 7939 18196 7948
rect 18144 7905 18153 7939
rect 18153 7905 18187 7939
rect 18187 7905 18196 7939
rect 18144 7896 18196 7905
rect 17684 7828 17736 7880
rect 13820 7760 13872 7769
rect 14740 7760 14792 7812
rect 16212 7760 16264 7812
rect 17500 7760 17552 7812
rect 14372 7692 14424 7744
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 15016 7735 15068 7744
rect 14832 7692 14884 7701
rect 15016 7701 15025 7735
rect 15025 7701 15059 7735
rect 15059 7701 15068 7735
rect 15016 7692 15068 7701
rect 15108 7692 15160 7744
rect 16580 7692 16632 7744
rect 17040 7692 17092 7744
rect 3947 7590 3999 7642
rect 4011 7590 4063 7642
rect 4075 7590 4127 7642
rect 4139 7590 4191 7642
rect 9878 7590 9930 7642
rect 9942 7590 9994 7642
rect 10006 7590 10058 7642
rect 10070 7590 10122 7642
rect 15808 7590 15860 7642
rect 15872 7590 15924 7642
rect 15936 7590 15988 7642
rect 16000 7590 16052 7642
rect 2412 7488 2464 7540
rect 4528 7488 4580 7540
rect 6000 7488 6052 7540
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2964 7420 3016 7472
rect 2872 7352 2924 7404
rect 3424 7352 3476 7404
rect 3792 7352 3844 7404
rect 4436 7420 4488 7472
rect 4804 7352 4856 7404
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5632 7352 5684 7404
rect 1400 7327 1452 7336
rect 1400 7293 1409 7327
rect 1409 7293 1443 7327
rect 1443 7293 1452 7327
rect 1400 7284 1452 7293
rect 2688 7284 2740 7336
rect 3608 7284 3660 7336
rect 4252 7284 4304 7336
rect 4436 7284 4488 7336
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 2872 7148 2924 7200
rect 3424 7148 3476 7200
rect 4344 7148 4396 7200
rect 7932 7488 7984 7540
rect 9588 7488 9640 7540
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 8760 7352 8812 7404
rect 9680 7352 9732 7404
rect 6736 7284 6788 7336
rect 7104 7284 7156 7336
rect 9404 7327 9456 7336
rect 9404 7293 9413 7327
rect 9413 7293 9447 7327
rect 9447 7293 9456 7327
rect 10324 7488 10376 7540
rect 11060 7488 11112 7540
rect 12808 7488 12860 7540
rect 10508 7420 10560 7472
rect 13544 7420 13596 7472
rect 15016 7488 15068 7540
rect 16856 7488 16908 7540
rect 18052 7488 18104 7540
rect 18512 7488 18564 7540
rect 10416 7352 10468 7404
rect 14280 7395 14332 7404
rect 9404 7284 9456 7293
rect 12256 7284 12308 7336
rect 14280 7361 14289 7395
rect 14289 7361 14323 7395
rect 14323 7361 14332 7395
rect 14280 7352 14332 7361
rect 16396 7352 16448 7404
rect 16580 7395 16632 7404
rect 16580 7361 16589 7395
rect 16589 7361 16623 7395
rect 16623 7361 16632 7395
rect 16580 7352 16632 7361
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 17500 7395 17552 7404
rect 16672 7352 16724 7361
rect 17500 7361 17509 7395
rect 17509 7361 17543 7395
rect 17543 7361 17552 7395
rect 17500 7352 17552 7361
rect 17960 7352 18012 7404
rect 18236 7352 18288 7404
rect 4896 7148 4948 7200
rect 5356 7148 5408 7200
rect 5632 7148 5684 7200
rect 7840 7216 7892 7268
rect 8392 7148 8444 7200
rect 8852 7148 8904 7200
rect 9588 7216 9640 7268
rect 10876 7216 10928 7268
rect 12164 7216 12216 7268
rect 13912 7284 13964 7336
rect 15384 7284 15436 7336
rect 16948 7284 17000 7336
rect 17868 7284 17920 7336
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 10324 7148 10376 7200
rect 10416 7148 10468 7200
rect 11888 7191 11940 7200
rect 11888 7157 11897 7191
rect 11897 7157 11931 7191
rect 11931 7157 11940 7191
rect 11888 7148 11940 7157
rect 12624 7148 12676 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 15936 7148 15988 7200
rect 16120 7191 16172 7200
rect 16120 7157 16129 7191
rect 16129 7157 16163 7191
rect 16163 7157 16172 7191
rect 16120 7148 16172 7157
rect 16212 7148 16264 7200
rect 16672 7148 16724 7200
rect 18236 7191 18288 7200
rect 18236 7157 18245 7191
rect 18245 7157 18279 7191
rect 18279 7157 18288 7191
rect 18236 7148 18288 7157
rect 6912 7046 6964 7098
rect 6976 7046 7028 7098
rect 7040 7046 7092 7098
rect 7104 7046 7156 7098
rect 12843 7046 12895 7098
rect 12907 7046 12959 7098
rect 12971 7046 13023 7098
rect 13035 7046 13087 7098
rect 18972 7055 19024 7064
rect 18972 7021 18981 7055
rect 18981 7021 19015 7055
rect 19015 7021 19024 7055
rect 18972 7012 19024 7021
rect 2688 6944 2740 6996
rect 3056 6944 3108 6996
rect 9404 6987 9456 6996
rect 1400 6876 1452 6928
rect 9404 6953 9413 6987
rect 9413 6953 9447 6987
rect 9447 6953 9456 6987
rect 9404 6944 9456 6953
rect 12348 6944 12400 6996
rect 12624 6944 12676 6996
rect 14372 6944 14424 6996
rect 14556 6944 14608 6996
rect 14740 6987 14792 6996
rect 14740 6953 14749 6987
rect 14749 6953 14783 6987
rect 14783 6953 14792 6987
rect 14740 6944 14792 6953
rect 15936 6944 15988 6996
rect 4804 6876 4856 6928
rect 1216 6740 1268 6792
rect 3424 6740 3476 6792
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 4252 6808 4304 6860
rect 5448 6876 5500 6928
rect 6736 6876 6788 6928
rect 6460 6808 6512 6860
rect 4344 6740 4396 6792
rect 4896 6783 4948 6792
rect 2596 6672 2648 6724
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 6644 6740 6696 6792
rect 7288 6783 7340 6792
rect 1400 6647 1452 6656
rect 1400 6613 1409 6647
rect 1409 6613 1443 6647
rect 1443 6613 1452 6647
rect 1400 6604 1452 6613
rect 2688 6604 2740 6656
rect 3056 6604 3108 6656
rect 5908 6672 5960 6724
rect 7288 6749 7297 6783
rect 7297 6749 7331 6783
rect 7331 6749 7340 6783
rect 7288 6740 7340 6749
rect 3424 6604 3476 6656
rect 4344 6604 4396 6656
rect 4620 6604 4672 6656
rect 5080 6604 5132 6656
rect 6368 6647 6420 6656
rect 6368 6613 6377 6647
rect 6377 6613 6411 6647
rect 6411 6613 6420 6647
rect 8024 6851 8076 6860
rect 8024 6817 8058 6851
rect 8058 6817 8076 6851
rect 10968 6876 11020 6928
rect 11060 6876 11112 6928
rect 11796 6876 11848 6928
rect 13544 6876 13596 6928
rect 13820 6876 13872 6928
rect 15016 6876 15068 6928
rect 15476 6876 15528 6928
rect 15660 6876 15712 6928
rect 10416 6851 10468 6860
rect 8024 6808 8076 6817
rect 10416 6817 10425 6851
rect 10425 6817 10459 6851
rect 10459 6817 10468 6851
rect 10416 6808 10468 6817
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 9772 6783 9824 6792
rect 9772 6749 9781 6783
rect 9781 6749 9815 6783
rect 9815 6749 9824 6783
rect 9772 6740 9824 6749
rect 10232 6740 10284 6792
rect 10600 6740 10652 6792
rect 11152 6851 11204 6860
rect 11152 6817 11186 6851
rect 11186 6817 11204 6851
rect 13268 6851 13320 6860
rect 11152 6808 11204 6817
rect 10876 6783 10928 6792
rect 10876 6749 10885 6783
rect 10885 6749 10919 6783
rect 10919 6749 10928 6783
rect 10876 6740 10928 6749
rect 13268 6817 13277 6851
rect 13277 6817 13311 6851
rect 13311 6817 13320 6851
rect 13268 6808 13320 6817
rect 15568 6808 15620 6860
rect 18696 6876 18748 6928
rect 16856 6808 16908 6860
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 10508 6672 10560 6724
rect 13912 6740 13964 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14924 6740 14976 6792
rect 16580 6740 16632 6792
rect 17316 6740 17368 6792
rect 17500 6783 17552 6792
rect 17500 6749 17509 6783
rect 17509 6749 17543 6783
rect 17543 6749 17552 6783
rect 17500 6740 17552 6749
rect 6368 6604 6420 6613
rect 8116 6604 8168 6656
rect 9404 6604 9456 6656
rect 11060 6604 11112 6656
rect 11520 6604 11572 6656
rect 12256 6647 12308 6656
rect 12256 6613 12265 6647
rect 12265 6613 12299 6647
rect 12299 6613 12308 6647
rect 12256 6604 12308 6613
rect 12440 6604 12492 6656
rect 15200 6672 15252 6724
rect 15384 6715 15436 6724
rect 15384 6681 15393 6715
rect 15393 6681 15427 6715
rect 15427 6681 15436 6715
rect 15384 6672 15436 6681
rect 16764 6672 16816 6724
rect 14556 6604 14608 6656
rect 15292 6604 15344 6656
rect 16580 6604 16632 6656
rect 16856 6647 16908 6656
rect 16856 6613 16865 6647
rect 16865 6613 16899 6647
rect 16899 6613 16908 6647
rect 16856 6604 16908 6613
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 17316 6604 17368 6656
rect 3947 6502 3999 6554
rect 4011 6502 4063 6554
rect 4075 6502 4127 6554
rect 4139 6502 4191 6554
rect 9878 6502 9930 6554
rect 9942 6502 9994 6554
rect 10006 6502 10058 6554
rect 10070 6502 10122 6554
rect 15808 6502 15860 6554
rect 15872 6502 15924 6554
rect 15936 6502 15988 6554
rect 16000 6502 16052 6554
rect 2412 6264 2464 6316
rect 2688 6307 2740 6316
rect 2688 6273 2697 6307
rect 2697 6273 2731 6307
rect 2731 6273 2740 6307
rect 2688 6264 2740 6273
rect 3332 6400 3384 6452
rect 3700 6400 3752 6452
rect 6460 6443 6512 6452
rect 6460 6409 6469 6443
rect 6469 6409 6503 6443
rect 6503 6409 6512 6443
rect 6460 6400 6512 6409
rect 6736 6400 6788 6452
rect 7748 6400 7800 6452
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 4896 6264 4948 6316
rect 10416 6400 10468 6452
rect 11888 6400 11940 6452
rect 12072 6400 12124 6452
rect 12256 6332 12308 6384
rect 12440 6400 12492 6452
rect 17500 6400 17552 6452
rect 13084 6332 13136 6384
rect 15200 6375 15252 6384
rect 15200 6341 15209 6375
rect 15209 6341 15243 6375
rect 15243 6341 15252 6375
rect 15200 6332 15252 6341
rect 15292 6332 15344 6384
rect 1952 6128 2004 6180
rect 2596 6196 2648 6248
rect 4988 6196 5040 6248
rect 6736 6196 6788 6248
rect 11152 6264 11204 6316
rect 11888 6264 11940 6316
rect 13544 6264 13596 6316
rect 6644 6128 6696 6180
rect 8300 6128 8352 6180
rect 9404 6128 9456 6180
rect 11520 6196 11572 6248
rect 12256 6196 12308 6248
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 13452 6239 13504 6248
rect 12808 6196 12860 6205
rect 13452 6205 13461 6239
rect 13461 6205 13495 6239
rect 13495 6205 13504 6239
rect 13452 6196 13504 6205
rect 13728 6196 13780 6248
rect 16120 6264 16172 6316
rect 16396 6332 16448 6384
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 1860 6103 1912 6112
rect 1860 6069 1869 6103
rect 1869 6069 1903 6103
rect 1903 6069 1912 6103
rect 1860 6060 1912 6069
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 3424 6060 3476 6112
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 4896 6060 4948 6112
rect 5724 6060 5776 6112
rect 9220 6060 9272 6112
rect 10324 6103 10376 6112
rect 10324 6069 10333 6103
rect 10333 6069 10367 6103
rect 10367 6069 10376 6103
rect 10324 6060 10376 6069
rect 11796 6128 11848 6180
rect 11428 6060 11480 6112
rect 13084 6128 13136 6180
rect 14556 6196 14608 6248
rect 16948 6239 17000 6248
rect 14280 6128 14332 6180
rect 14924 6128 14976 6180
rect 15200 6128 15252 6180
rect 16672 6128 16724 6180
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 17868 6196 17920 6248
rect 14648 6060 14700 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 16212 6060 16264 6112
rect 17776 6103 17828 6112
rect 17776 6069 17785 6103
rect 17785 6069 17819 6103
rect 17819 6069 17828 6103
rect 17776 6060 17828 6069
rect 18236 6103 18288 6112
rect 18236 6069 18245 6103
rect 18245 6069 18279 6103
rect 18279 6069 18288 6103
rect 18236 6060 18288 6069
rect 6912 5958 6964 6010
rect 6976 5958 7028 6010
rect 7040 5958 7092 6010
rect 7104 5958 7156 6010
rect 12843 5958 12895 6010
rect 12907 5958 12959 6010
rect 12971 5958 13023 6010
rect 13035 5958 13087 6010
rect 2596 5720 2648 5772
rect 2412 5652 2464 5704
rect 2504 5652 2556 5704
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 3516 5831 3568 5840
rect 3516 5797 3525 5831
rect 3525 5797 3559 5831
rect 3559 5797 3568 5831
rect 3516 5788 3568 5797
rect 5356 5788 5408 5840
rect 6920 5788 6972 5840
rect 7288 5856 7340 5908
rect 8116 5856 8168 5908
rect 9128 5856 9180 5908
rect 10232 5856 10284 5908
rect 10324 5856 10376 5908
rect 11428 5856 11480 5908
rect 13268 5856 13320 5908
rect 15476 5856 15528 5908
rect 15752 5899 15804 5908
rect 15752 5865 15761 5899
rect 15761 5865 15795 5899
rect 15795 5865 15804 5899
rect 15752 5856 15804 5865
rect 4344 5763 4396 5772
rect 4344 5729 4378 5763
rect 4378 5729 4396 5763
rect 4344 5720 4396 5729
rect 7656 5720 7708 5772
rect 10416 5788 10468 5840
rect 10600 5788 10652 5840
rect 13544 5831 13596 5840
rect 13544 5797 13553 5831
rect 13553 5797 13587 5831
rect 13587 5797 13596 5831
rect 13544 5788 13596 5797
rect 13912 5788 13964 5840
rect 15568 5788 15620 5840
rect 16212 5788 16264 5840
rect 16856 5788 16908 5840
rect 17316 5788 17368 5840
rect 8576 5763 8628 5772
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 3332 5516 3384 5568
rect 6460 5652 6512 5704
rect 6644 5652 6696 5704
rect 7380 5652 7432 5704
rect 8576 5729 8585 5763
rect 8585 5729 8619 5763
rect 8619 5729 8628 5763
rect 8576 5720 8628 5729
rect 10324 5720 10376 5772
rect 7840 5695 7892 5704
rect 7840 5661 7849 5695
rect 7849 5661 7883 5695
rect 7883 5661 7892 5695
rect 7840 5652 7892 5661
rect 8300 5652 8352 5704
rect 5080 5584 5132 5636
rect 8852 5652 8904 5704
rect 9680 5652 9732 5704
rect 11244 5652 11296 5704
rect 12348 5720 12400 5772
rect 12532 5720 12584 5772
rect 12716 5720 12768 5772
rect 11888 5695 11940 5704
rect 9128 5584 9180 5636
rect 11428 5584 11480 5636
rect 11888 5661 11897 5695
rect 11897 5661 11931 5695
rect 11931 5661 11940 5695
rect 11888 5652 11940 5661
rect 12164 5652 12216 5704
rect 13176 5695 13228 5704
rect 13176 5661 13185 5695
rect 13185 5661 13219 5695
rect 13219 5661 13228 5695
rect 13176 5652 13228 5661
rect 14372 5720 14424 5772
rect 13912 5652 13964 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14832 5720 14884 5772
rect 14280 5652 14332 5661
rect 14740 5652 14792 5704
rect 15200 5720 15252 5772
rect 15568 5652 15620 5704
rect 15660 5652 15712 5704
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 16120 5652 16172 5661
rect 17224 5720 17276 5772
rect 17500 5720 17552 5772
rect 4804 5516 4856 5568
rect 5448 5559 5500 5568
rect 5448 5525 5457 5559
rect 5457 5525 5491 5559
rect 5491 5525 5500 5559
rect 5448 5516 5500 5525
rect 6552 5516 6604 5568
rect 10416 5516 10468 5568
rect 11244 5516 11296 5568
rect 12256 5559 12308 5568
rect 12256 5525 12265 5559
rect 12265 5525 12299 5559
rect 12299 5525 12308 5559
rect 12256 5516 12308 5525
rect 12532 5559 12584 5568
rect 12532 5525 12541 5559
rect 12541 5525 12575 5559
rect 12575 5525 12584 5559
rect 12532 5516 12584 5525
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 17776 5559 17828 5568
rect 17776 5525 17785 5559
rect 17785 5525 17819 5559
rect 17819 5525 17828 5559
rect 17776 5516 17828 5525
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 3947 5414 3999 5466
rect 4011 5414 4063 5466
rect 4075 5414 4127 5466
rect 4139 5414 4191 5466
rect 9878 5414 9930 5466
rect 9942 5414 9994 5466
rect 10006 5414 10058 5466
rect 10070 5414 10122 5466
rect 15808 5414 15860 5466
rect 15872 5414 15924 5466
rect 15936 5414 15988 5466
rect 16000 5414 16052 5466
rect 2504 5312 2556 5364
rect 3608 5312 3660 5364
rect 4344 5312 4396 5364
rect 4528 5312 4580 5364
rect 6184 5312 6236 5364
rect 6920 5355 6972 5364
rect 6920 5321 6929 5355
rect 6929 5321 6963 5355
rect 6963 5321 6972 5355
rect 6920 5312 6972 5321
rect 7656 5312 7708 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 11980 5312 12032 5364
rect 12348 5312 12400 5364
rect 13912 5355 13964 5364
rect 4436 5287 4488 5296
rect 1492 5176 1544 5228
rect 4436 5253 4445 5287
rect 4445 5253 4479 5287
rect 4479 5253 4488 5287
rect 4436 5244 4488 5253
rect 6644 5244 6696 5296
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 7380 5219 7432 5228
rect 1400 5151 1452 5160
rect 1400 5117 1409 5151
rect 1409 5117 1443 5151
rect 1443 5117 1452 5151
rect 1400 5108 1452 5117
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 2872 5108 2924 5160
rect 3332 5108 3384 5160
rect 4068 5108 4120 5160
rect 4620 5108 4672 5160
rect 4160 5040 4212 5092
rect 4804 5108 4856 5160
rect 5448 5108 5500 5160
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 5632 5040 5684 5092
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 10876 5219 10928 5228
rect 7288 5108 7340 5160
rect 8852 5108 8904 5160
rect 9220 5151 9272 5160
rect 9220 5117 9254 5151
rect 9254 5117 9272 5151
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 1952 4972 2004 5024
rect 2688 4972 2740 5024
rect 3608 4972 3660 5024
rect 3700 4972 3752 5024
rect 6092 5015 6144 5024
rect 6092 4981 6101 5015
rect 6101 4981 6135 5015
rect 6135 4981 6144 5015
rect 6092 4972 6144 4981
rect 6184 5015 6236 5024
rect 6184 4981 6193 5015
rect 6193 4981 6227 5015
rect 6227 4981 6236 5015
rect 6184 4972 6236 4981
rect 6736 4972 6788 5024
rect 7564 5040 7616 5092
rect 9220 5108 9272 5117
rect 9588 5108 9640 5160
rect 9680 5108 9732 5160
rect 10876 5185 10885 5219
rect 10885 5185 10919 5219
rect 10919 5185 10928 5219
rect 10876 5176 10928 5185
rect 12164 5176 12216 5228
rect 13912 5321 13921 5355
rect 13921 5321 13955 5355
rect 13955 5321 13964 5355
rect 13912 5312 13964 5321
rect 14188 5312 14240 5364
rect 15016 5355 15068 5364
rect 15016 5321 15025 5355
rect 15025 5321 15059 5355
rect 15059 5321 15068 5355
rect 15016 5312 15068 5321
rect 17132 5312 17184 5364
rect 17592 5312 17644 5364
rect 13544 5244 13596 5296
rect 14372 5176 14424 5228
rect 7932 4972 7984 5024
rect 9496 4972 9548 5024
rect 10140 4972 10192 5024
rect 10324 4972 10376 5024
rect 12348 5108 12400 5160
rect 12164 5040 12216 5092
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 13728 5040 13780 5092
rect 15568 5176 15620 5228
rect 16304 5244 16356 5296
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 17776 5244 17828 5296
rect 16948 5176 17000 5228
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 15476 5108 15528 5160
rect 17316 5108 17368 5160
rect 11152 4972 11204 5024
rect 12256 5015 12308 5024
rect 12256 4981 12265 5015
rect 12265 4981 12299 5015
rect 12299 4981 12308 5015
rect 12256 4972 12308 4981
rect 14188 4972 14240 5024
rect 14648 4972 14700 5024
rect 17960 5040 18012 5092
rect 15200 4972 15252 5024
rect 15476 5015 15528 5024
rect 15476 4981 15485 5015
rect 15485 4981 15519 5015
rect 15519 4981 15528 5015
rect 15476 4972 15528 4981
rect 15660 4972 15712 5024
rect 16580 4972 16632 5024
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 17224 4972 17276 5024
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 18236 5015 18288 5024
rect 17592 4972 17644 4981
rect 18236 4981 18245 5015
rect 18245 4981 18279 5015
rect 18279 4981 18288 5015
rect 18236 4972 18288 4981
rect 6912 4870 6964 4922
rect 6976 4870 7028 4922
rect 7040 4870 7092 4922
rect 7104 4870 7156 4922
rect 12843 4870 12895 4922
rect 12907 4870 12959 4922
rect 12971 4870 13023 4922
rect 13035 4870 13087 4922
rect 1676 4768 1728 4820
rect 3608 4768 3660 4820
rect 3792 4768 3844 4820
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 3240 4700 3292 4752
rect 6184 4768 6236 4820
rect 7564 4768 7616 4820
rect 8300 4768 8352 4820
rect 9772 4768 9824 4820
rect 10416 4768 10468 4820
rect 11520 4768 11572 4820
rect 12716 4768 12768 4820
rect 13360 4811 13412 4820
rect 13360 4777 13369 4811
rect 13369 4777 13403 4811
rect 13403 4777 13412 4811
rect 13360 4768 13412 4777
rect 13452 4768 13504 4820
rect 4528 4743 4580 4752
rect 4528 4709 4537 4743
rect 4537 4709 4571 4743
rect 4571 4709 4580 4743
rect 4528 4700 4580 4709
rect 4620 4700 4672 4752
rect 7840 4700 7892 4752
rect 10232 4700 10284 4752
rect 12532 4700 12584 4752
rect 14556 4700 14608 4752
rect 15568 4743 15620 4752
rect 15568 4709 15602 4743
rect 15602 4709 15620 4743
rect 15568 4700 15620 4709
rect 16948 4743 17000 4752
rect 16948 4709 16957 4743
rect 16957 4709 16991 4743
rect 16991 4709 17000 4743
rect 16948 4700 17000 4709
rect 17040 4700 17092 4752
rect 1308 4564 1360 4616
rect 1860 4471 1912 4480
rect 1860 4437 1869 4471
rect 1869 4437 1903 4471
rect 1903 4437 1912 4471
rect 1860 4428 1912 4437
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 4344 4632 4396 4684
rect 5172 4632 5224 4684
rect 5356 4675 5408 4684
rect 5356 4641 5365 4675
rect 5365 4641 5399 4675
rect 5399 4641 5408 4675
rect 5356 4632 5408 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 8208 4632 8260 4684
rect 9312 4632 9364 4684
rect 10140 4632 10192 4684
rect 5632 4607 5684 4616
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 6920 4564 6972 4616
rect 8392 4564 8444 4616
rect 11336 4564 11388 4616
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 11612 4564 11664 4616
rect 12256 4564 12308 4616
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 14280 4632 14332 4684
rect 14464 4632 14516 4684
rect 17316 4632 17368 4684
rect 13728 4607 13780 4616
rect 4252 4428 4304 4480
rect 4436 4471 4488 4480
rect 4436 4437 4445 4471
rect 4445 4437 4479 4471
rect 4479 4437 4488 4471
rect 4436 4428 4488 4437
rect 4988 4471 5040 4480
rect 4988 4437 4997 4471
rect 4997 4437 5031 4471
rect 5031 4437 5040 4471
rect 4988 4428 5040 4437
rect 5448 4428 5500 4480
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 11152 4496 11204 4548
rect 12348 4496 12400 4548
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 15200 4564 15252 4616
rect 16948 4564 17000 4616
rect 13176 4496 13228 4548
rect 17684 4607 17736 4616
rect 17684 4573 17693 4607
rect 17693 4573 17727 4607
rect 17727 4573 17736 4607
rect 17684 4564 17736 4573
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 9680 4428 9732 4480
rect 10232 4428 10284 4480
rect 10416 4471 10468 4480
rect 10416 4437 10425 4471
rect 10425 4437 10459 4471
rect 10459 4437 10468 4471
rect 10416 4428 10468 4437
rect 13360 4428 13412 4480
rect 18052 4496 18104 4548
rect 16672 4471 16724 4480
rect 16672 4437 16681 4471
rect 16681 4437 16715 4471
rect 16715 4437 16724 4471
rect 16672 4428 16724 4437
rect 17224 4428 17276 4480
rect 17316 4428 17368 4480
rect 17592 4428 17644 4480
rect 17868 4428 17920 4480
rect 3947 4326 3999 4378
rect 4011 4326 4063 4378
rect 4075 4326 4127 4378
rect 4139 4326 4191 4378
rect 9878 4326 9930 4378
rect 9942 4326 9994 4378
rect 10006 4326 10058 4378
rect 10070 4326 10122 4378
rect 15808 4326 15860 4378
rect 15872 4326 15924 4378
rect 15936 4326 15988 4378
rect 16000 4326 16052 4378
rect 4528 4224 4580 4276
rect 4804 4224 4856 4276
rect 5724 4224 5776 4276
rect 6460 4224 6512 4276
rect 7932 4224 7984 4276
rect 8208 4267 8260 4276
rect 8208 4233 8217 4267
rect 8217 4233 8251 4267
rect 8251 4233 8260 4267
rect 8208 4224 8260 4233
rect 9680 4224 9732 4276
rect 10508 4224 10560 4276
rect 11520 4224 11572 4276
rect 12072 4224 12124 4276
rect 12440 4224 12492 4276
rect 1768 4156 1820 4208
rect 1768 4020 1820 4072
rect 2780 4088 2832 4140
rect 6736 4156 6788 4208
rect 10232 4156 10284 4208
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 4988 4088 5040 4140
rect 5632 4088 5684 4140
rect 6092 4131 6144 4140
rect 6092 4097 6101 4131
rect 6101 4097 6135 4131
rect 6135 4097 6144 4131
rect 6092 4088 6144 4097
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10416 4088 10468 4140
rect 11428 4088 11480 4140
rect 11612 4156 11664 4208
rect 14096 4224 14148 4276
rect 2964 4063 3016 4072
rect 2964 4029 2973 4063
rect 2973 4029 3007 4063
rect 3007 4029 3016 4063
rect 2964 4020 3016 4029
rect 5448 4020 5500 4072
rect 5540 4020 5592 4072
rect 6920 4020 6972 4072
rect 1676 3927 1728 3936
rect 1676 3893 1685 3927
rect 1685 3893 1719 3927
rect 1719 3893 1728 3927
rect 1676 3884 1728 3893
rect 2044 3927 2096 3936
rect 2044 3893 2053 3927
rect 2053 3893 2087 3927
rect 2087 3893 2096 3927
rect 2044 3884 2096 3893
rect 2412 3927 2464 3936
rect 2412 3893 2421 3927
rect 2421 3893 2455 3927
rect 2455 3893 2464 3927
rect 2412 3884 2464 3893
rect 2596 3927 2648 3936
rect 2596 3893 2605 3927
rect 2605 3893 2639 3927
rect 2639 3893 2648 3927
rect 2596 3884 2648 3893
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 4804 3884 4856 3936
rect 5816 3952 5868 4004
rect 6644 3952 6696 4004
rect 6736 3952 6788 4004
rect 7656 3952 7708 4004
rect 9680 4020 9732 4072
rect 9772 4020 9824 4072
rect 10324 4020 10376 4072
rect 9128 3952 9180 4004
rect 6092 3884 6144 3936
rect 6276 3884 6328 3936
rect 6460 3884 6512 3936
rect 11060 3952 11112 4004
rect 11152 3952 11204 4004
rect 11888 4088 11940 4140
rect 13268 4088 13320 4140
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 15016 4156 15068 4208
rect 14280 4131 14332 4140
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 15200 4088 15252 4140
rect 14464 4020 14516 4072
rect 16672 4156 16724 4208
rect 13544 3952 13596 4004
rect 9956 3884 10008 3936
rect 10692 3884 10744 3936
rect 10968 3927 11020 3936
rect 10968 3893 10977 3927
rect 10977 3893 11011 3927
rect 11011 3893 11020 3927
rect 10968 3884 11020 3893
rect 11612 3884 11664 3936
rect 13176 3884 13228 3936
rect 13912 3884 13964 3936
rect 14188 3927 14240 3936
rect 14188 3893 14197 3927
rect 14197 3893 14231 3927
rect 14231 3893 14240 3927
rect 14188 3884 14240 3893
rect 14740 3884 14792 3936
rect 17040 4088 17092 4140
rect 17224 4131 17276 4140
rect 17224 4097 17233 4131
rect 17233 4097 17267 4131
rect 17267 4097 17276 4131
rect 17224 4088 17276 4097
rect 17776 4156 17828 4208
rect 16764 4020 16816 4072
rect 17132 4063 17184 4072
rect 17132 4029 17141 4063
rect 17141 4029 17175 4063
rect 17175 4029 17184 4063
rect 17132 4020 17184 4029
rect 18052 4063 18104 4072
rect 16948 3952 17000 4004
rect 18052 4029 18061 4063
rect 18061 4029 18095 4063
rect 18095 4029 18104 4063
rect 18052 4020 18104 4029
rect 16856 3884 16908 3936
rect 17776 3927 17828 3936
rect 17776 3893 17785 3927
rect 17785 3893 17819 3927
rect 17819 3893 17828 3927
rect 17776 3884 17828 3893
rect 17868 3884 17920 3936
rect 6912 3782 6964 3834
rect 6976 3782 7028 3834
rect 7040 3782 7092 3834
rect 7104 3782 7156 3834
rect 12843 3782 12895 3834
rect 12907 3782 12959 3834
rect 12971 3782 13023 3834
rect 13035 3782 13087 3834
rect 3240 3680 3292 3732
rect 3884 3680 3936 3732
rect 4528 3680 4580 3732
rect 5172 3680 5224 3732
rect 3700 3612 3752 3664
rect 5448 3612 5500 3664
rect 7380 3680 7432 3732
rect 8668 3680 8720 3732
rect 8760 3680 8812 3732
rect 10968 3680 11020 3732
rect 11060 3680 11112 3732
rect 388 3544 440 3596
rect 3516 3587 3568 3596
rect 3516 3553 3525 3587
rect 3525 3553 3559 3587
rect 3559 3553 3568 3587
rect 3516 3544 3568 3553
rect 4160 3544 4212 3596
rect 5632 3544 5684 3596
rect 6552 3544 6604 3596
rect 8392 3612 8444 3664
rect 9312 3612 9364 3664
rect 1308 3476 1360 3528
rect 5540 3519 5592 3528
rect 3424 3340 3476 3392
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 7564 3476 7616 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9036 3544 9088 3596
rect 8944 3476 8996 3528
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 10692 3612 10744 3664
rect 12808 3612 12860 3664
rect 13452 3612 13504 3664
rect 13912 3612 13964 3664
rect 14740 3612 14792 3664
rect 16120 3680 16172 3732
rect 16856 3723 16908 3732
rect 16856 3689 16865 3723
rect 16865 3689 16899 3723
rect 16899 3689 16908 3723
rect 16856 3680 16908 3689
rect 16948 3680 17000 3732
rect 17500 3723 17552 3732
rect 17500 3689 17509 3723
rect 17509 3689 17543 3723
rect 17543 3689 17552 3723
rect 17500 3680 17552 3689
rect 9772 3544 9824 3596
rect 9956 3587 10008 3596
rect 9956 3553 9990 3587
rect 9990 3553 10008 3587
rect 9956 3544 10008 3553
rect 10416 3544 10468 3596
rect 11152 3519 11204 3528
rect 9404 3476 9456 3485
rect 11152 3485 11161 3519
rect 11161 3485 11195 3519
rect 11195 3485 11204 3519
rect 11152 3476 11204 3485
rect 5172 3408 5224 3460
rect 5448 3451 5500 3460
rect 5448 3417 5457 3451
rect 5457 3417 5491 3451
rect 5491 3417 5500 3451
rect 5448 3408 5500 3417
rect 8852 3408 8904 3460
rect 9680 3408 9732 3460
rect 13728 3544 13780 3596
rect 15936 3544 15988 3596
rect 16212 3544 16264 3596
rect 16580 3612 16632 3664
rect 18144 3612 18196 3664
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 15660 3476 15712 3528
rect 16304 3476 16356 3528
rect 16672 3476 16724 3528
rect 12808 3451 12860 3460
rect 12808 3417 12817 3451
rect 12817 3417 12851 3451
rect 12851 3417 12860 3451
rect 12808 3408 12860 3417
rect 15384 3408 15436 3460
rect 18144 3476 18196 3528
rect 18696 3476 18748 3528
rect 6736 3340 6788 3392
rect 7012 3340 7064 3392
rect 8576 3340 8628 3392
rect 9404 3340 9456 3392
rect 11060 3383 11112 3392
rect 11060 3349 11069 3383
rect 11069 3349 11103 3383
rect 11103 3349 11112 3383
rect 11060 3340 11112 3349
rect 13544 3340 13596 3392
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 16672 3340 16724 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 3947 3238 3999 3290
rect 4011 3238 4063 3290
rect 4075 3238 4127 3290
rect 4139 3238 4191 3290
rect 9878 3238 9930 3290
rect 9942 3238 9994 3290
rect 10006 3238 10058 3290
rect 10070 3238 10122 3290
rect 15808 3238 15860 3290
rect 15872 3238 15924 3290
rect 15936 3238 15988 3290
rect 16000 3238 16052 3290
rect 1492 2932 1544 2984
rect 2872 3136 2924 3188
rect 3516 3136 3568 3188
rect 5540 3136 5592 3188
rect 7656 3136 7708 3188
rect 8852 3136 8904 3188
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 3792 3068 3844 3120
rect 1860 3000 1912 3052
rect 2780 3000 2832 3052
rect 5172 3000 5224 3052
rect 2136 2975 2188 2984
rect 2136 2941 2145 2975
rect 2145 2941 2179 2975
rect 2179 2941 2188 2975
rect 2136 2932 2188 2941
rect 3056 2932 3108 2984
rect 3332 2932 3384 2984
rect 4804 2932 4856 2984
rect 5724 3068 5776 3120
rect 6552 3068 6604 3120
rect 8944 3068 8996 3120
rect 5632 3043 5684 3052
rect 5632 3009 5641 3043
rect 5641 3009 5675 3043
rect 5675 3009 5684 3043
rect 5632 3000 5684 3009
rect 6644 3000 6696 3052
rect 8760 3000 8812 3052
rect 11060 3136 11112 3188
rect 12532 3136 12584 3188
rect 10692 3068 10744 3120
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 9588 3000 9640 3009
rect 6276 2975 6328 2984
rect 6276 2941 6285 2975
rect 6285 2941 6319 2975
rect 6319 2941 6328 2975
rect 6276 2932 6328 2941
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 7380 2932 7432 2984
rect 7656 2975 7708 2984
rect 7656 2941 7665 2975
rect 7665 2941 7699 2975
rect 7699 2941 7708 2975
rect 7656 2932 7708 2941
rect 8484 2932 8536 2984
rect 9404 2975 9456 2984
rect 9404 2941 9413 2975
rect 9413 2941 9447 2975
rect 9447 2941 9456 2975
rect 9404 2932 9456 2941
rect 3240 2907 3292 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 1676 2796 1728 2848
rect 2320 2839 2372 2848
rect 2320 2805 2329 2839
rect 2329 2805 2363 2839
rect 2363 2805 2372 2839
rect 2320 2796 2372 2805
rect 2688 2839 2740 2848
rect 2688 2805 2697 2839
rect 2697 2805 2731 2839
rect 2731 2805 2740 2839
rect 2688 2796 2740 2805
rect 3240 2873 3249 2907
rect 3249 2873 3283 2907
rect 3283 2873 3292 2907
rect 3240 2864 3292 2873
rect 4528 2864 4580 2916
rect 7564 2907 7616 2916
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 4068 2839 4120 2848
rect 4068 2805 4077 2839
rect 4077 2805 4111 2839
rect 4111 2805 4120 2839
rect 4068 2796 4120 2805
rect 5448 2796 5500 2848
rect 7564 2873 7573 2907
rect 7573 2873 7607 2907
rect 7607 2873 7616 2907
rect 7564 2864 7616 2873
rect 8300 2864 8352 2916
rect 8760 2864 8812 2916
rect 10232 2932 10284 2984
rect 10600 2932 10652 2984
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 10876 2932 10928 2984
rect 10968 2932 11020 2984
rect 12348 3000 12400 3052
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 12440 2932 12492 2984
rect 15384 3136 15436 3188
rect 17040 3136 17092 3188
rect 17316 3136 17368 3188
rect 17592 3179 17644 3188
rect 17592 3145 17601 3179
rect 17601 3145 17635 3179
rect 17635 3145 17644 3179
rect 17592 3136 17644 3145
rect 13452 3000 13504 3052
rect 14004 3068 14056 3120
rect 14740 3111 14792 3120
rect 14740 3077 14749 3111
rect 14749 3077 14783 3111
rect 14783 3077 14792 3111
rect 14740 3068 14792 3077
rect 14280 3043 14332 3052
rect 10324 2864 10376 2916
rect 10692 2864 10744 2916
rect 13268 2864 13320 2916
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 15384 3000 15436 3052
rect 16580 3068 16632 3120
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 16856 3043 16908 3052
rect 16856 3009 16865 3043
rect 16865 3009 16899 3043
rect 16899 3009 16908 3043
rect 16856 3000 16908 3009
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14648 2932 14700 2984
rect 15568 2932 15620 2984
rect 16212 2932 16264 2984
rect 17316 2932 17368 2984
rect 14188 2864 14240 2916
rect 7288 2796 7340 2848
rect 9772 2796 9824 2848
rect 10140 2796 10192 2848
rect 11428 2839 11480 2848
rect 11428 2805 11437 2839
rect 11437 2805 11471 2839
rect 11471 2805 11480 2839
rect 11428 2796 11480 2805
rect 13636 2796 13688 2848
rect 19432 2864 19484 2916
rect 15476 2796 15528 2848
rect 16120 2796 16172 2848
rect 6912 2694 6964 2746
rect 6976 2694 7028 2746
rect 7040 2694 7092 2746
rect 7104 2694 7156 2746
rect 12843 2694 12895 2746
rect 12907 2694 12959 2746
rect 12971 2694 13023 2746
rect 13035 2694 13087 2746
rect 1860 2592 1912 2644
rect 3516 2592 3568 2644
rect 4436 2592 4488 2644
rect 5356 2592 5408 2644
rect 8300 2592 8352 2644
rect 8944 2592 8996 2644
rect 10140 2592 10192 2644
rect 10692 2592 10744 2644
rect 11060 2635 11112 2644
rect 11060 2601 11069 2635
rect 11069 2601 11103 2635
rect 11103 2601 11112 2635
rect 11060 2592 11112 2601
rect 11336 2592 11388 2644
rect 11520 2592 11572 2644
rect 11888 2592 11940 2644
rect 1124 2456 1176 2508
rect 1952 2499 2004 2508
rect 1952 2465 1961 2499
rect 1961 2465 1995 2499
rect 1995 2465 2004 2499
rect 1952 2456 2004 2465
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 3424 2499 3476 2508
rect 2136 2431 2188 2440
rect 2136 2397 2145 2431
rect 2145 2397 2179 2431
rect 2179 2397 2188 2431
rect 2136 2388 2188 2397
rect 2780 2320 2832 2372
rect 3424 2465 3433 2499
rect 3433 2465 3467 2499
rect 3467 2465 3476 2499
rect 3424 2456 3476 2465
rect 5080 2524 5132 2576
rect 5724 2524 5776 2576
rect 8668 2524 8720 2576
rect 8760 2524 8812 2576
rect 10232 2567 10284 2576
rect 10232 2533 10241 2567
rect 10241 2533 10275 2567
rect 10275 2533 10284 2567
rect 10232 2524 10284 2533
rect 11428 2524 11480 2576
rect 11704 2524 11756 2576
rect 15200 2635 15252 2644
rect 15200 2601 15209 2635
rect 15209 2601 15243 2635
rect 15243 2601 15252 2635
rect 15200 2592 15252 2601
rect 17316 2592 17368 2644
rect 18144 2592 18196 2644
rect 12164 2524 12216 2576
rect 15016 2524 15068 2576
rect 4712 2499 4764 2508
rect 4712 2465 4721 2499
rect 4721 2465 4755 2499
rect 4755 2465 4764 2499
rect 4712 2456 4764 2465
rect 5264 2499 5316 2508
rect 5264 2465 5273 2499
rect 5273 2465 5307 2499
rect 5307 2465 5316 2499
rect 5264 2456 5316 2465
rect 7380 2456 7432 2508
rect 10784 2456 10836 2508
rect 11060 2456 11112 2508
rect 13360 2456 13412 2508
rect 13820 2456 13872 2508
rect 15108 2456 15160 2508
rect 15292 2456 15344 2508
rect 3148 2388 3200 2440
rect 4252 2388 4304 2440
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5816 2388 5868 2440
rect 6736 2388 6788 2440
rect 7564 2388 7616 2440
rect 1768 2295 1820 2304
rect 1768 2261 1777 2295
rect 1777 2261 1811 2295
rect 1811 2261 1820 2295
rect 1768 2252 1820 2261
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 3516 2252 3568 2304
rect 3792 2320 3844 2372
rect 7288 2320 7340 2372
rect 8760 2388 8812 2440
rect 9128 2388 9180 2440
rect 11244 2431 11296 2440
rect 11244 2397 11253 2431
rect 11253 2397 11287 2431
rect 11287 2397 11296 2431
rect 11244 2388 11296 2397
rect 12440 2431 12492 2440
rect 12440 2397 12449 2431
rect 12449 2397 12483 2431
rect 12483 2397 12492 2431
rect 12440 2388 12492 2397
rect 6092 2252 6144 2304
rect 6552 2295 6604 2304
rect 6552 2261 6561 2295
rect 6561 2261 6595 2295
rect 6595 2261 6604 2295
rect 6552 2252 6604 2261
rect 13176 2431 13228 2440
rect 13176 2397 13185 2431
rect 13185 2397 13219 2431
rect 13219 2397 13228 2431
rect 13636 2431 13688 2440
rect 13176 2388 13228 2397
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 13912 2320 13964 2372
rect 14832 2388 14884 2440
rect 17868 2388 17920 2440
rect 10416 2252 10468 2304
rect 11704 2252 11756 2304
rect 12072 2252 12124 2304
rect 17500 2295 17552 2304
rect 17500 2261 17509 2295
rect 17509 2261 17543 2295
rect 17543 2261 17552 2295
rect 17500 2252 17552 2261
rect 3947 2150 3999 2202
rect 4011 2150 4063 2202
rect 4075 2150 4127 2202
rect 4139 2150 4191 2202
rect 9878 2150 9930 2202
rect 9942 2150 9994 2202
rect 10006 2150 10058 2202
rect 10070 2150 10122 2202
rect 15808 2150 15860 2202
rect 15872 2150 15924 2202
rect 15936 2150 15988 2202
rect 16000 2150 16052 2202
rect 9772 2048 9824 2100
rect 12072 2048 12124 2100
rect 10324 1436 10376 1488
rect 14280 1436 14332 1488
rect 2596 1300 2648 1352
rect 15200 1300 15252 1352
rect 3240 1164 3292 1216
rect 15292 1232 15344 1284
rect 11244 1096 11296 1148
rect 13636 1096 13688 1148
<< metal2 >>
rect 1950 16400 2006 17200
rect 4066 16960 4122 16969
rect 4066 16895 4122 16904
rect 2962 16688 3018 16697
rect 2962 16623 3018 16632
rect 1398 15600 1454 15609
rect 1398 15535 1454 15544
rect 1412 14618 1440 15535
rect 1674 15056 1730 15065
rect 1674 14991 1730 15000
rect 1400 14612 1452 14618
rect 1400 14554 1452 14560
rect 1688 13938 1716 14991
rect 1768 14408 1820 14414
rect 1766 14376 1768 14385
rect 1820 14376 1822 14385
rect 1964 14346 1992 16400
rect 2134 16280 2190 16289
rect 2134 16215 2190 16224
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1766 14311 1822 14320
rect 1952 14340 2004 14346
rect 1952 14282 2004 14288
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1504 13530 1532 13631
rect 1492 13524 1544 13530
rect 1492 13466 1544 13472
rect 2056 13394 2084 14418
rect 2148 13870 2176 16215
rect 2686 16008 2742 16017
rect 2686 15943 2742 15952
rect 2320 14408 2372 14414
rect 2320 14350 2372 14356
rect 2332 13977 2360 14350
rect 2318 13968 2374 13977
rect 2318 13903 2374 13912
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2320 13320 2372 13326
rect 1858 13288 1914 13297
rect 2320 13262 2372 13268
rect 1858 13223 1860 13232
rect 1912 13223 1914 13232
rect 1860 13194 1912 13200
rect 2134 13016 2190 13025
rect 2134 12951 2190 12960
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1674 11112 1730 11121
rect 1674 11047 1730 11056
rect 1688 11014 1716 11047
rect 1676 11008 1728 11014
rect 1676 10950 1728 10956
rect 1860 11008 1912 11014
rect 1860 10950 1912 10956
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9042 1440 9998
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1504 9178 1532 9318
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1124 8832 1176 8838
rect 1124 8774 1176 8780
rect 1136 5681 1164 8774
rect 1412 8498 1440 8978
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7342 1440 8230
rect 1400 7336 1452 7342
rect 1400 7278 1452 7284
rect 1306 7168 1362 7177
rect 1306 7103 1362 7112
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 1122 5672 1178 5681
rect 1122 5607 1178 5616
rect 388 3596 440 3602
rect 388 3538 440 3544
rect 400 800 428 3538
rect 1136 2514 1164 5607
rect 1228 4604 1256 6734
rect 1320 6644 1348 7103
rect 1412 6934 1440 7278
rect 1400 6928 1452 6934
rect 1400 6870 1452 6876
rect 1400 6656 1452 6662
rect 1320 6616 1400 6644
rect 1400 6598 1452 6604
rect 1412 5166 1440 6598
rect 1504 5930 1532 9114
rect 1688 8888 1716 10950
rect 1872 10674 1900 10950
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10266 1808 10406
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1964 9518 1992 11494
rect 2056 10810 2084 11494
rect 2148 11014 2176 12951
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10606 2176 10950
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 1952 9512 2004 9518
rect 1952 9454 2004 9460
rect 1688 8860 1808 8888
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6089 1624 7142
rect 1688 6769 1716 7686
rect 1674 6760 1730 6769
rect 1674 6695 1730 6704
rect 1582 6080 1638 6089
rect 1582 6015 1638 6024
rect 1504 5902 1624 5930
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1504 5234 1532 5510
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1400 5160 1452 5166
rect 1596 5114 1624 5902
rect 1400 5102 1452 5108
rect 1504 5086 1624 5114
rect 1308 4616 1360 4622
rect 1228 4576 1308 4604
rect 1308 4558 1360 4564
rect 1214 3632 1270 3641
rect 1214 3567 1270 3576
rect 1124 2508 1176 2514
rect 1124 2450 1176 2456
rect 1228 800 1256 3567
rect 1320 3534 1348 4558
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1504 2990 1532 5086
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4729 1624 4966
rect 1688 4826 1716 6695
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1780 4214 1808 8860
rect 1950 6216 2006 6225
rect 1950 6151 1952 6160
rect 2004 6151 2006 6160
rect 1952 6122 2004 6128
rect 1860 6112 1912 6118
rect 1860 6054 1912 6060
rect 1872 5137 1900 6054
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1860 4480 1912 4486
rect 1860 4422 1912 4428
rect 1768 4208 1820 4214
rect 1872 4185 1900 4422
rect 1768 4150 1820 4156
rect 1858 4176 1914 4185
rect 1858 4111 1914 4120
rect 1768 4072 1820 4078
rect 1768 4014 1820 4020
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 1688 3777 1716 3878
rect 1674 3768 1730 3777
rect 1674 3703 1730 3712
rect 1780 3346 1808 4014
rect 1780 3318 1900 3346
rect 1872 3058 1900 3318
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1676 2848 1728 2854
rect 1676 2790 1728 2796
rect 1596 2417 1624 2790
rect 1582 2408 1638 2417
rect 1582 2343 1638 2352
rect 386 0 442 800
rect 1214 0 1270 800
rect 1688 785 1716 2790
rect 1872 2650 1900 2994
rect 1860 2644 1912 2650
rect 1860 2586 1912 2592
rect 1964 2514 1992 4966
rect 2056 4729 2084 10134
rect 2240 9761 2268 11290
rect 2226 9752 2282 9761
rect 2226 9687 2282 9696
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2134 9208 2190 9217
rect 2134 9143 2190 9152
rect 2148 7721 2176 9143
rect 2240 8634 2268 9318
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2228 7744 2280 7750
rect 2134 7712 2190 7721
rect 2228 7686 2280 7692
rect 2134 7647 2190 7656
rect 2240 7410 2268 7686
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5166 2176 6054
rect 2226 5944 2282 5953
rect 2226 5879 2282 5888
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2042 4720 2098 4729
rect 2240 4672 2268 5879
rect 2042 4655 2044 4664
rect 2096 4655 2098 4664
rect 2044 4626 2096 4632
rect 2148 4644 2268 4672
rect 2056 4595 2084 4626
rect 2044 3936 2096 3942
rect 2044 3878 2096 3884
rect 2056 3097 2084 3878
rect 2042 3088 2098 3097
rect 2042 3023 2098 3032
rect 2148 2990 2176 4644
rect 2228 4480 2280 4486
rect 2226 4448 2228 4457
rect 2280 4448 2282 4457
rect 2226 4383 2282 4392
rect 2332 3380 2360 13262
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 10810 2452 11494
rect 2504 11280 2556 11286
rect 2504 11222 2556 11228
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2516 10674 2544 11222
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 10198 2636 10406
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2700 9994 2728 15943
rect 2870 15328 2926 15337
rect 2870 15263 2926 15272
rect 2778 14648 2834 14657
rect 2778 14583 2834 14592
rect 2792 13938 2820 14583
rect 2884 14482 2912 15263
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2976 14074 3004 16623
rect 4080 15230 4108 16895
rect 5906 16400 5962 17200
rect 9862 16400 9918 17200
rect 13910 16400 13966 17200
rect 16486 16960 16542 16969
rect 16486 16895 16542 16904
rect 15658 16552 15714 16561
rect 15658 16487 15714 16496
rect 4068 15224 4120 15230
rect 4068 15166 4120 15172
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 3712 12306 3740 14418
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 3804 14074 3832 14214
rect 3921 14172 4217 14192
rect 3977 14170 4001 14172
rect 4057 14170 4081 14172
rect 4137 14170 4161 14172
rect 3999 14118 4001 14170
rect 4063 14118 4075 14170
rect 4137 14118 4139 14170
rect 3977 14116 4001 14118
rect 4057 14116 4081 14118
rect 4137 14116 4161 14118
rect 3921 14096 4217 14116
rect 5920 14074 5948 16400
rect 9404 15224 9456 15230
rect 9404 15166 9456 15172
rect 6886 14716 7182 14736
rect 6942 14714 6966 14716
rect 7022 14714 7046 14716
rect 7102 14714 7126 14716
rect 6964 14662 6966 14714
rect 7028 14662 7040 14714
rect 7102 14662 7104 14714
rect 6942 14660 6966 14662
rect 7022 14660 7046 14662
rect 7102 14660 7126 14662
rect 6886 14640 7182 14660
rect 9416 14074 9444 15166
rect 9876 14396 9904 16400
rect 13450 15056 13506 15065
rect 13450 14991 13506 15000
rect 12817 14716 13113 14736
rect 12873 14714 12897 14716
rect 12953 14714 12977 14716
rect 13033 14714 13057 14716
rect 12895 14662 12897 14714
rect 12959 14662 12971 14714
rect 13033 14662 13035 14714
rect 12873 14660 12897 14662
rect 12953 14660 12977 14662
rect 13033 14660 13057 14662
rect 12817 14640 13113 14660
rect 9784 14368 9904 14396
rect 3792 14068 3844 14074
rect 3792 14010 3844 14016
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 9404 14068 9456 14074
rect 9404 14010 9456 14016
rect 9416 13870 9444 14010
rect 9784 13954 9812 14368
rect 9852 14172 10148 14192
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 9930 14118 9932 14170
rect 9994 14118 10006 14170
rect 10068 14118 10070 14170
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 9852 14096 10148 14116
rect 9784 13938 9904 13954
rect 9680 13932 9732 13938
rect 9784 13932 9916 13938
rect 9784 13926 9864 13932
rect 9680 13874 9732 13880
rect 9864 13874 9916 13880
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 3921 13084 4217 13104
rect 3977 13082 4001 13084
rect 4057 13082 4081 13084
rect 4137 13082 4161 13084
rect 3999 13030 4001 13082
rect 4063 13030 4075 13082
rect 4137 13030 4139 13082
rect 3977 13028 4001 13030
rect 4057 13028 4081 13030
rect 4137 13028 4161 13030
rect 3921 13008 4217 13028
rect 3974 12744 4030 12753
rect 3974 12679 3976 12688
rect 4028 12679 4030 12688
rect 5908 12708 5960 12714
rect 3976 12650 4028 12656
rect 5908 12650 5960 12656
rect 3790 12336 3846 12345
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3700 12300 3752 12306
rect 3790 12271 3846 12280
rect 3700 12242 3752 12248
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2792 9586 2820 10406
rect 2976 10062 3004 10610
rect 2964 10056 3016 10062
rect 2870 10024 2926 10033
rect 2964 9998 3016 10004
rect 2870 9959 2926 9968
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 9178 2452 9318
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2780 9036 2832 9042
rect 2780 8978 2832 8984
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8362 2728 8842
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2412 8016 2464 8022
rect 2412 7958 2464 7964
rect 2424 7546 2452 7958
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2424 7449 2452 7482
rect 2410 7440 2466 7449
rect 2410 7375 2466 7384
rect 2608 7290 2636 7890
rect 2700 7886 2728 8298
rect 2792 8090 2820 8978
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2884 7993 2912 9959
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2976 9586 3004 9862
rect 2964 9580 3016 9586
rect 2964 9522 3016 9528
rect 2976 9110 3004 9522
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 3068 9058 3096 12242
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3436 11665 3464 12174
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3514 12064 3570 12073
rect 3514 11999 3570 12008
rect 3422 11656 3478 11665
rect 3422 11591 3478 11600
rect 3330 11384 3386 11393
rect 3330 11319 3386 11328
rect 3240 10532 3292 10538
rect 3240 10474 3292 10480
rect 3252 10266 3280 10474
rect 3240 10260 3292 10266
rect 3240 10202 3292 10208
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3252 9625 3280 9930
rect 3238 9616 3294 9625
rect 3238 9551 3294 9560
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 3068 9030 3188 9058
rect 3160 8974 3188 9030
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2870 7984 2926 7993
rect 2870 7919 2926 7928
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2872 7880 2924 7886
rect 2872 7822 2924 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2700 7342 2728 7686
rect 2778 7440 2834 7449
rect 2884 7410 2912 7822
rect 2976 7818 3004 8230
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2964 7812 3016 7818
rect 2964 7754 3016 7760
rect 2976 7478 3004 7754
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2778 7375 2834 7384
rect 2872 7404 2924 7410
rect 2516 7262 2636 7290
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 5710 2452 6258
rect 2516 5930 2544 7262
rect 2688 6996 2740 7002
rect 2688 6938 2740 6944
rect 2700 6905 2728 6938
rect 2686 6896 2742 6905
rect 2686 6831 2742 6840
rect 2596 6724 2648 6730
rect 2596 6666 2648 6672
rect 2608 6254 2636 6666
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6322 2728 6598
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2596 6248 2648 6254
rect 2596 6190 2648 6196
rect 2516 5902 2728 5930
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2516 5370 2544 5646
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2608 3942 2636 5714
rect 2700 5030 2728 5902
rect 2688 5024 2740 5030
rect 2688 4966 2740 4972
rect 2700 4593 2728 4966
rect 2686 4584 2742 4593
rect 2686 4519 2742 4528
rect 2792 4146 2820 7375
rect 2872 7346 2924 7352
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2884 5166 2912 7142
rect 3068 7002 3096 8026
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2962 6896 3018 6905
rect 2962 6831 3018 6840
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2976 4078 3004 6831
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3068 5386 3096 6598
rect 3160 5953 3188 8774
rect 3146 5944 3202 5953
rect 3146 5879 3202 5888
rect 3252 5817 3280 9386
rect 3344 8265 3372 11319
rect 3528 11082 3556 11999
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3620 11014 3648 11698
rect 3712 11286 3740 12106
rect 3804 11898 3832 12271
rect 3921 11996 4217 12016
rect 3977 11994 4001 11996
rect 4057 11994 4081 11996
rect 4137 11994 4161 11996
rect 3999 11942 4001 11994
rect 4063 11942 4075 11994
rect 4137 11942 4139 11994
rect 3977 11940 4001 11942
rect 4057 11940 4081 11942
rect 4137 11940 4161 11942
rect 3921 11920 4217 11940
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3700 11280 3752 11286
rect 3700 11222 3752 11228
rect 3608 11008 3660 11014
rect 3422 10976 3478 10985
rect 3608 10950 3660 10956
rect 3422 10911 3478 10920
rect 3436 9926 3464 10911
rect 3620 10674 3648 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 10124 3568 10130
rect 3620 10112 3648 10610
rect 3712 10198 3740 11222
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10674 3832 11086
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 3921 10908 4217 10928
rect 3977 10906 4001 10908
rect 4057 10906 4081 10908
rect 4137 10906 4161 10908
rect 3999 10854 4001 10906
rect 4063 10854 4075 10906
rect 4137 10854 4139 10906
rect 3977 10852 4001 10854
rect 4057 10852 4081 10854
rect 4137 10852 4161 10854
rect 3921 10832 4217 10852
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3568 10084 3648 10112
rect 3516 10066 3568 10072
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3804 9722 3832 10610
rect 4264 10198 4292 10950
rect 4526 10704 4582 10713
rect 4526 10639 4582 10648
rect 4540 10606 4568 10639
rect 4528 10600 4580 10606
rect 4528 10542 4580 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4252 10192 4304 10198
rect 4252 10134 4304 10140
rect 4632 10130 4660 10406
rect 4724 10266 4752 10542
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 3921 9820 4217 9840
rect 3977 9818 4001 9820
rect 4057 9818 4081 9820
rect 4137 9818 4161 9820
rect 3999 9766 4001 9818
rect 4063 9766 4075 9818
rect 4137 9766 4139 9818
rect 3977 9764 4001 9766
rect 4057 9764 4081 9766
rect 4137 9764 4161 9766
rect 3921 9744 4217 9764
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3514 9616 3570 9625
rect 3514 9551 3570 9560
rect 3424 9104 3476 9110
rect 3422 9072 3424 9081
rect 3476 9072 3478 9081
rect 3422 9007 3478 9016
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3330 8256 3386 8265
rect 3330 8191 3386 8200
rect 3436 8106 3464 8910
rect 3344 8078 3464 8106
rect 3344 7018 3372 8078
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3436 7206 3464 7346
rect 3424 7200 3476 7206
rect 3424 7142 3476 7148
rect 3344 6990 3464 7018
rect 3436 6798 3464 6990
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3238 5808 3294 5817
rect 3238 5743 3294 5752
rect 3344 5574 3372 6394
rect 3436 6118 3464 6598
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3528 5930 3556 9551
rect 3804 9042 3832 9658
rect 4356 9654 4384 10066
rect 4436 10056 4488 10062
rect 4434 10024 4436 10033
rect 4712 10056 4764 10062
rect 4488 10024 4490 10033
rect 4712 9998 4764 10004
rect 4434 9959 4490 9968
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4618 9616 4674 9625
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3988 9110 4016 9318
rect 3976 9104 4028 9110
rect 3976 9046 4028 9052
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8294 3648 8774
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3606 8120 3662 8129
rect 3606 8055 3662 8064
rect 3620 7750 3648 8055
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3620 7342 3648 7686
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3620 6338 3648 7278
rect 3712 7041 3740 8910
rect 3804 8430 3832 8978
rect 4080 8906 4108 9522
rect 4344 9444 4396 9450
rect 4344 9386 4396 9392
rect 4250 9344 4306 9353
rect 4250 9279 4306 9288
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4172 8974 4200 9114
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4264 8838 4292 9279
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 3921 8732 4217 8752
rect 3977 8730 4001 8732
rect 4057 8730 4081 8732
rect 4137 8730 4161 8732
rect 3999 8678 4001 8730
rect 4063 8678 4075 8730
rect 4137 8678 4139 8730
rect 3977 8676 4001 8678
rect 4057 8676 4081 8678
rect 4137 8676 4161 8678
rect 3921 8656 4217 8676
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3792 8288 3844 8294
rect 3792 8230 3844 8236
rect 3882 8256 3938 8265
rect 3804 7410 3832 8230
rect 3882 8191 3938 8200
rect 3896 8090 3924 8191
rect 4264 8090 4292 8774
rect 3884 8084 3936 8090
rect 3884 8026 3936 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 3921 7644 4217 7664
rect 3977 7642 4001 7644
rect 4057 7642 4081 7644
rect 4137 7642 4161 7644
rect 3999 7590 4001 7642
rect 4063 7590 4075 7642
rect 4137 7590 4139 7642
rect 3977 7588 4001 7590
rect 4057 7588 4081 7590
rect 4137 7588 4161 7590
rect 3921 7568 4217 7588
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 4264 7342 4292 7686
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4356 7206 4384 9386
rect 4448 9382 4476 9590
rect 4618 9551 4674 9560
rect 4632 9382 4660 9551
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4620 9376 4672 9382
rect 4724 9353 4752 9998
rect 4816 9489 4844 11018
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4802 9480 4858 9489
rect 4802 9415 4858 9424
rect 4620 9318 4672 9324
rect 4710 9344 4766 9353
rect 4632 8974 4660 9318
rect 4710 9279 4766 9288
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4448 8412 4476 8910
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4448 8384 4568 8412
rect 4436 8288 4488 8294
rect 4436 8230 4488 8236
rect 4448 7478 4476 8230
rect 4540 7993 4568 8384
rect 4526 7984 4582 7993
rect 4526 7919 4582 7928
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4540 7546 4568 7822
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 3698 7032 3754 7041
rect 3698 6967 3754 6976
rect 4158 7032 4214 7041
rect 4448 6984 4476 7278
rect 4158 6967 4214 6976
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3698 6488 3754 6497
rect 3698 6423 3700 6432
rect 3752 6423 3754 6432
rect 3700 6394 3752 6400
rect 3620 6310 3740 6338
rect 3436 5902 3556 5930
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3068 5358 3188 5386
rect 2964 4072 3016 4078
rect 2884 4032 2964 4060
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2424 3505 2452 3878
rect 2410 3496 2466 3505
rect 2410 3431 2466 3440
rect 2332 3352 2636 3380
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2148 2689 2176 2926
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2134 2680 2190 2689
rect 2134 2615 2190 2624
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 1768 2304 1820 2310
rect 1768 2246 1820 2252
rect 1780 2145 1808 2246
rect 1766 2136 1822 2145
rect 1766 2071 1822 2080
rect 2148 800 2176 2382
rect 2332 1873 2360 2790
rect 2502 2544 2558 2553
rect 2502 2479 2504 2488
rect 2556 2479 2558 2488
rect 2504 2450 2556 2456
rect 2318 1864 2374 1873
rect 2318 1799 2374 1808
rect 2608 1358 2636 3352
rect 2884 3194 2912 4032
rect 2964 4014 3016 4020
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2778 3088 2834 3097
rect 2778 3023 2780 3032
rect 2832 3023 2834 3032
rect 2780 2994 2832 3000
rect 3056 2984 3108 2990
rect 3054 2952 3056 2961
rect 3160 2972 3188 5358
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3252 4758 3280 5170
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3252 4146 3280 4694
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3738 3280 4082
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3344 2990 3372 5102
rect 3436 4049 3464 5902
rect 3516 5840 3568 5846
rect 3514 5808 3516 5817
rect 3568 5808 3570 5817
rect 3514 5743 3570 5752
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3620 5370 3648 5646
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3712 5030 3740 6310
rect 3804 5710 3832 6734
rect 4172 6644 4200 6967
rect 4264 6956 4476 6984
rect 4264 6866 4292 6956
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4356 6662 4384 6734
rect 4632 6662 4660 8774
rect 4344 6656 4396 6662
rect 4172 6616 4292 6644
rect 3921 6556 4217 6576
rect 3977 6554 4001 6556
rect 4057 6554 4081 6556
rect 4137 6554 4161 6556
rect 3999 6502 4001 6554
rect 4063 6502 4075 6554
rect 4137 6502 4139 6554
rect 3977 6500 4001 6502
rect 4057 6500 4081 6502
rect 4137 6500 4161 6502
rect 3921 6480 4217 6500
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3608 5024 3660 5030
rect 3608 4966 3660 4972
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3620 4826 3648 4966
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 3620 4185 3648 4762
rect 3606 4176 3662 4185
rect 3606 4111 3662 4120
rect 3422 4040 3478 4049
rect 3422 3975 3478 3984
rect 3712 3942 3740 4966
rect 3804 4826 3832 5646
rect 3921 5468 4217 5488
rect 3977 5466 4001 5468
rect 4057 5466 4081 5468
rect 4137 5466 4161 5468
rect 3999 5414 4001 5466
rect 4063 5414 4075 5466
rect 4137 5414 4139 5466
rect 3977 5412 4001 5414
rect 4057 5412 4081 5414
rect 4137 5412 4161 5414
rect 3921 5392 4217 5412
rect 4068 5160 4120 5166
rect 4066 5128 4068 5137
rect 4120 5128 4122 5137
rect 4066 5063 4122 5072
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 4172 4468 4200 5034
rect 4264 4672 4292 6616
rect 4344 6598 4396 6604
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4356 5778 4384 6054
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5370 4384 5714
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4436 5296 4488 5302
rect 4434 5264 4436 5273
rect 4488 5264 4490 5273
rect 4434 5199 4490 5208
rect 4540 4758 4568 5306
rect 4632 5166 4660 6598
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4632 4758 4660 5102
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4344 4684 4396 4690
rect 4264 4644 4344 4672
rect 4344 4626 4396 4632
rect 4252 4480 4304 4486
rect 4172 4440 4252 4468
rect 4436 4480 4488 4486
rect 4252 4422 4304 4428
rect 4434 4448 4436 4457
rect 4488 4448 4490 4457
rect 3921 4380 4217 4400
rect 3977 4378 4001 4380
rect 4057 4378 4081 4380
rect 4137 4378 4161 4380
rect 3999 4326 4001 4378
rect 4063 4326 4075 4378
rect 4137 4326 4139 4378
rect 3977 4324 4001 4326
rect 4057 4324 4081 4326
rect 4137 4324 4161 4326
rect 3921 4304 4217 4324
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3712 3670 3740 3878
rect 3896 3738 3924 3878
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3700 3664 3752 3670
rect 3700 3606 3752 3612
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 4160 3596 4212 3602
rect 4264 3584 4292 4422
rect 4434 4383 4490 4392
rect 4212 3556 4292 3584
rect 4160 3538 4212 3544
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3108 2952 3188 2972
rect 3110 2944 3188 2952
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3054 2887 3110 2896
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2596 1352 2648 1358
rect 2596 1294 2648 1300
rect 1674 776 1730 785
rect 1674 711 1730 720
rect 2134 0 2190 800
rect 2700 513 2728 2790
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2780 2372 2832 2378
rect 2780 2314 2832 2320
rect 2686 504 2742 513
rect 2686 439 2742 448
rect 2792 241 2820 2314
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 1193 3096 2246
rect 3054 1184 3110 1193
rect 3054 1119 3110 1128
rect 3160 1034 3188 2382
rect 3252 1222 3280 2858
rect 3436 2514 3464 3334
rect 3528 3194 3556 3538
rect 3921 3292 4217 3312
rect 3977 3290 4001 3292
rect 4057 3290 4081 3292
rect 4137 3290 4161 3292
rect 3999 3238 4001 3290
rect 4063 3238 4075 3290
rect 4137 3238 4139 3290
rect 3977 3236 4001 3238
rect 4057 3236 4081 3238
rect 4137 3236 4161 3238
rect 3921 3216 4217 3236
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3528 2553 3556 2586
rect 3514 2544 3570 2553
rect 3424 2508 3476 2514
rect 3514 2479 3570 2488
rect 3424 2450 3476 2456
rect 3528 2310 3556 2479
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3712 1465 3740 2790
rect 3804 2378 3832 3062
rect 4068 2848 4120 2854
rect 4066 2816 4068 2825
rect 4120 2816 4122 2825
rect 4066 2751 4122 2760
rect 4448 2650 4476 4383
rect 4540 4282 4568 4694
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4540 3738 4568 4082
rect 4528 3732 4580 3738
rect 4528 3674 4580 3680
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4540 2825 4568 2858
rect 4526 2816 4582 2825
rect 4526 2751 4582 2760
rect 4436 2644 4488 2650
rect 4436 2586 4488 2592
rect 4724 2514 4752 8842
rect 4816 7410 4844 9415
rect 4908 8344 4936 10746
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10062 5120 10474
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5538 10432 5594 10441
rect 5080 10056 5132 10062
rect 5264 10056 5316 10062
rect 5080 9998 5132 10004
rect 5184 10016 5264 10044
rect 5092 9586 5120 9998
rect 5184 9722 5212 10016
rect 5368 10033 5396 10406
rect 5538 10367 5594 10376
rect 5552 10266 5580 10367
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5264 9998 5316 10004
rect 5354 10024 5410 10033
rect 5354 9959 5356 9968
rect 5408 9959 5410 9968
rect 5356 9930 5408 9936
rect 5368 9899 5396 9930
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5276 9625 5304 9658
rect 5262 9616 5318 9625
rect 5080 9580 5132 9586
rect 5262 9551 5318 9560
rect 5080 9522 5132 9528
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9178 5028 9318
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4988 8356 5040 8362
rect 4908 8316 4988 8344
rect 4988 8298 5040 8304
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4908 7857 4936 8026
rect 4894 7848 4950 7857
rect 4894 7783 4950 7792
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4896 7200 4948 7206
rect 4894 7168 4896 7177
rect 4948 7168 4950 7177
rect 4894 7103 4950 7112
rect 4804 6928 4856 6934
rect 4804 6870 4856 6876
rect 4816 6322 4844 6870
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6322 4936 6734
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 6202 4936 6258
rect 5000 6254 5028 8298
rect 5092 6662 5120 9522
rect 5460 9466 5488 10134
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9926 5580 10066
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5368 9438 5488 9466
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7410 5212 7754
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5170 7304 5226 7313
rect 5170 7239 5226 7248
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 4816 6174 4936 6202
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 4816 5574 4844 6174
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4816 5166 4844 5510
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4816 3942 4844 4218
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4804 2984 4856 2990
rect 4908 2972 4936 6054
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 5000 4146 5028 4422
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4856 2944 4936 2972
rect 4804 2926 4856 2932
rect 5092 2582 5120 5578
rect 5184 4690 5212 7239
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5184 3466 5212 3674
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5184 3058 5212 3402
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5080 2576 5132 2582
rect 5080 2518 5132 2524
rect 5276 2514 5304 9318
rect 5368 9178 5396 9438
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5356 8016 5408 8022
rect 5356 7958 5408 7964
rect 5368 7206 5396 7958
rect 5460 7585 5488 9318
rect 5446 7576 5502 7585
rect 5446 7511 5502 7520
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 5846 5396 7142
rect 5448 6928 5500 6934
rect 5448 6870 5500 6876
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 5460 5692 5488 6870
rect 5368 5664 5488 5692
rect 5368 5012 5396 5664
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 5166 5488 5510
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5368 4984 5488 5012
rect 5356 4684 5408 4690
rect 5356 4626 5408 4632
rect 5368 2825 5396 4626
rect 5460 4486 5488 4984
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4078 5488 4422
rect 5552 4264 5580 9862
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5736 9058 5764 9522
rect 5828 9382 5856 9590
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5736 9042 5856 9058
rect 5736 9036 5868 9042
rect 5736 9030 5816 9036
rect 5816 8978 5868 8984
rect 5828 8634 5856 8978
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 8514 5948 12650
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6012 9178 6040 9386
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5920 8486 6040 8514
rect 5908 8424 5960 8430
rect 5814 8392 5870 8401
rect 5908 8366 5960 8372
rect 5814 8327 5870 8336
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 7886 5764 8230
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 7410 5672 7686
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5630 7304 5686 7313
rect 5630 7239 5686 7248
rect 5644 7206 5672 7239
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5736 6118 5764 7822
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5644 4622 5672 5034
rect 5828 4690 5856 8327
rect 5920 7954 5948 8366
rect 5908 7948 5960 7954
rect 5908 7890 5960 7896
rect 6012 7546 6040 8486
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6104 6984 6132 13806
rect 6886 13628 7182 13648
rect 6942 13626 6966 13628
rect 7022 13626 7046 13628
rect 7102 13626 7126 13628
rect 6964 13574 6966 13626
rect 7028 13574 7040 13626
rect 7102 13574 7104 13626
rect 6942 13572 6966 13574
rect 7022 13572 7046 13574
rect 7102 13572 7126 13574
rect 6886 13552 7182 13572
rect 9692 12986 9720 13874
rect 12162 13832 12218 13841
rect 12162 13767 12218 13776
rect 9852 13084 10148 13104
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 9930 13030 9932 13082
rect 9994 13030 10006 13082
rect 10068 13030 10070 13082
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 9852 13008 10148 13028
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 6886 12540 7182 12560
rect 6942 12538 6966 12540
rect 7022 12538 7046 12540
rect 7102 12538 7126 12540
rect 6964 12486 6966 12538
rect 7028 12486 7040 12538
rect 7102 12486 7104 12538
rect 6942 12484 6966 12486
rect 7022 12484 7046 12486
rect 7102 12484 7126 12486
rect 6886 12464 7182 12484
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6748 11558 6776 12378
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7288 11620 7340 11626
rect 7288 11562 7340 11568
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 6288 10606 6316 11290
rect 6380 10810 6408 11494
rect 6748 11218 6776 11494
rect 6886 11452 7182 11472
rect 6942 11450 6966 11452
rect 7022 11450 7046 11452
rect 7102 11450 7126 11452
rect 6964 11398 6966 11450
rect 7028 11398 7040 11450
rect 7102 11398 7104 11450
rect 6942 11396 6966 11398
rect 7022 11396 7046 11398
rect 7102 11396 7126 11398
rect 6886 11376 7182 11396
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6840 10742 6868 11086
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9722 6316 10066
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6196 9042 6224 9143
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6196 8634 6224 8978
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6012 6956 6132 6984
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5920 5914 5948 6666
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5724 4276 5776 4282
rect 5552 4236 5724 4264
rect 5724 4218 5776 4224
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5460 3466 5488 3606
rect 5552 3534 5580 4014
rect 5644 3602 5672 4082
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5540 3188 5592 3194
rect 5460 3148 5540 3176
rect 5460 2854 5488 3148
rect 5540 3130 5592 3136
rect 5644 3058 5672 3538
rect 5736 3126 5764 4218
rect 5828 4010 5856 4626
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 6012 3505 6040 6956
rect 6196 5370 6224 8570
rect 6288 6644 6316 9454
rect 6380 9178 6408 10610
rect 6552 10532 6604 10538
rect 6840 10520 6868 10678
rect 7116 10606 7144 11018
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 6920 10532 6972 10538
rect 6840 10492 6920 10520
rect 6552 10474 6604 10480
rect 6920 10474 6972 10480
rect 6564 9994 6592 10474
rect 6886 10364 7182 10384
rect 6942 10362 6966 10364
rect 7022 10362 7046 10364
rect 7102 10362 7126 10364
rect 6964 10310 6966 10362
rect 7028 10310 7040 10362
rect 7102 10310 7104 10362
rect 6942 10308 6966 10310
rect 7022 10308 7046 10310
rect 7102 10308 7126 10310
rect 6886 10288 7182 10308
rect 6828 10192 6880 10198
rect 6880 10152 6960 10180
rect 6828 10134 6880 10140
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6552 9988 6604 9994
rect 6552 9930 6604 9936
rect 6564 9518 6592 9930
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6564 8430 6592 9454
rect 6656 9450 6684 9998
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6748 9178 6776 9862
rect 6932 9518 6960 10152
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 6886 9276 7182 9296
rect 6942 9274 6966 9276
rect 7022 9274 7046 9276
rect 7102 9274 7126 9276
rect 6964 9222 6966 9274
rect 7028 9222 7040 9274
rect 7102 9222 7104 9274
rect 6942 9220 6966 9222
rect 7022 9220 7046 9222
rect 7102 9220 7126 9222
rect 6886 9200 7182 9220
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7300 8786 7328 11562
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7392 11286 7420 11494
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7576 10810 7604 11698
rect 7668 11150 7696 11698
rect 7760 11558 7788 12038
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7576 10198 7604 10746
rect 7564 10192 7616 10198
rect 7564 10134 7616 10140
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7656 10124 7708 10130
rect 7656 10066 7708 10072
rect 7484 9722 7512 10066
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 8974 7420 9454
rect 7668 9042 7696 10066
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7562 8936 7618 8945
rect 7562 8871 7618 8880
rect 7300 8758 7512 8786
rect 6552 8424 6604 8430
rect 6366 8392 6422 8401
rect 6552 8366 6604 8372
rect 6366 8327 6368 8336
rect 6420 8327 6422 8336
rect 7288 8356 7340 8362
rect 6368 8298 6420 8304
rect 7288 8298 7340 8304
rect 6886 8188 7182 8208
rect 6942 8186 6966 8188
rect 7022 8186 7046 8188
rect 7102 8186 7126 8188
rect 6964 8134 6966 8186
rect 7028 8134 7040 8186
rect 7102 8134 7104 8186
rect 6942 8132 6966 8134
rect 7022 8132 7046 8134
rect 7102 8132 7126 8134
rect 6886 8112 7182 8132
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7104 7880 7156 7886
rect 6550 7848 6606 7857
rect 7104 7822 7156 7828
rect 6550 7783 6606 7792
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6368 6656 6420 6662
rect 6288 6616 6368 6644
rect 6368 6598 6420 6604
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6380 5166 6408 6598
rect 6472 6458 6500 6802
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 5710 6500 6394
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6564 5574 6592 7783
rect 7116 7342 7144 7822
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7208 7290 7236 7958
rect 7300 7818 7328 8298
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 8090 7420 8230
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7288 7812 7340 7818
rect 7288 7754 7340 7760
rect 7392 7410 7420 7890
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 6748 6934 6776 7278
rect 7208 7262 7420 7290
rect 7392 7177 7420 7262
rect 7378 7168 7434 7177
rect 6886 7100 7182 7120
rect 7378 7103 7434 7112
rect 6942 7098 6966 7100
rect 7022 7098 7046 7100
rect 7102 7098 7126 7100
rect 6964 7046 6966 7098
rect 7028 7046 7040 7098
rect 7102 7046 7104 7098
rect 6942 7044 6966 7046
rect 7022 7044 7046 7046
rect 7102 7044 7126 7046
rect 6886 7024 7182 7044
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 6656 6186 6684 6734
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6748 6254 6776 6394
rect 6736 6248 6788 6254
rect 6736 6190 6788 6196
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6656 5710 6684 6122
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6644 5296 6696 5302
rect 6644 5238 6696 5244
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6104 4146 6132 4966
rect 6196 4826 6224 4966
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 6366 4720 6422 4729
rect 6366 4655 6368 4664
rect 6420 4655 6422 4664
rect 6368 4626 6420 4632
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 5998 3496 6054 3505
rect 5998 3431 6054 3440
rect 5724 3120 5776 3126
rect 5724 3062 5776 3068
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5448 2848 5500 2854
rect 5354 2816 5410 2825
rect 5448 2790 5500 2796
rect 5354 2751 5410 2760
rect 5368 2650 5396 2751
rect 5460 2689 5488 2790
rect 5446 2680 5502 2689
rect 5356 2644 5408 2650
rect 5446 2615 5502 2624
rect 5356 2586 5408 2592
rect 5736 2582 5764 3062
rect 5724 2576 5776 2582
rect 5724 2518 5776 2524
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 3921 2204 4217 2224
rect 3977 2202 4001 2204
rect 4057 2202 4081 2204
rect 4137 2202 4161 2204
rect 3999 2150 4001 2202
rect 4063 2150 4075 2202
rect 4137 2150 4139 2202
rect 3977 2148 4001 2150
rect 4057 2148 4081 2150
rect 4137 2148 4161 2150
rect 3921 2128 4217 2148
rect 3698 1456 3754 1465
rect 4264 1442 4292 2382
rect 3698 1391 3754 1400
rect 3988 1414 4292 1442
rect 3240 1216 3292 1222
rect 3240 1158 3292 1164
rect 3068 1006 3188 1034
rect 3068 800 3096 1006
rect 3988 800 4016 1414
rect 4908 800 4936 2382
rect 5828 800 5856 2382
rect 6104 2310 6132 3878
rect 6288 2990 6316 3878
rect 6380 2990 6408 4626
rect 6656 4468 6684 5238
rect 6748 5030 6776 6190
rect 6886 6012 7182 6032
rect 6942 6010 6966 6012
rect 7022 6010 7046 6012
rect 7102 6010 7126 6012
rect 6964 5958 6966 6010
rect 7028 5958 7040 6010
rect 7102 5958 7104 6010
rect 6942 5956 6966 5958
rect 7022 5956 7046 5958
rect 7102 5956 7126 5958
rect 6886 5936 7182 5956
rect 7300 5914 7328 6734
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6932 5370 6960 5782
rect 7392 5710 7420 7103
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6748 4808 6776 4966
rect 6886 4924 7182 4944
rect 6942 4922 6966 4924
rect 7022 4922 7046 4924
rect 7102 4922 7126 4924
rect 6964 4870 6966 4922
rect 7028 4870 7040 4922
rect 7102 4870 7104 4922
rect 6942 4868 6966 4870
rect 7022 4868 7046 4870
rect 7102 4868 7126 4870
rect 6886 4848 7182 4868
rect 6748 4780 6960 4808
rect 6932 4622 6960 4780
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6736 4480 6788 4486
rect 6656 4440 6736 4468
rect 6736 4422 6788 4428
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6472 3942 6500 4218
rect 6748 4214 6776 4422
rect 6736 4208 6788 4214
rect 6550 4176 6606 4185
rect 6736 4150 6788 4156
rect 6550 4111 6606 4120
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6564 3602 6592 4111
rect 6932 4078 6960 4558
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6552 3120 6604 3126
rect 6552 3062 6604 3068
rect 6276 2984 6328 2990
rect 6276 2926 6328 2932
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6564 2310 6592 3062
rect 6656 3058 6684 3946
rect 6748 3398 6776 3946
rect 6886 3836 7182 3856
rect 6942 3834 6966 3836
rect 7022 3834 7046 3836
rect 7102 3834 7126 3836
rect 6964 3782 6966 3834
rect 7028 3782 7040 3834
rect 7102 3782 7104 3834
rect 6942 3780 6966 3782
rect 7022 3780 7046 3782
rect 7102 3780 7126 3782
rect 6886 3760 7182 3780
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3097 7052 3334
rect 7010 3088 7066 3097
rect 6644 3052 6696 3058
rect 7010 3023 7066 3032
rect 6644 2994 6696 3000
rect 7300 2854 7328 5102
rect 7392 3738 7420 5170
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7288 2848 7340 2854
rect 7392 2825 7420 2926
rect 7288 2790 7340 2796
rect 7378 2816 7434 2825
rect 6886 2748 7182 2768
rect 6942 2746 6966 2748
rect 7022 2746 7046 2748
rect 7102 2746 7126 2748
rect 6964 2694 6966 2746
rect 7028 2694 7040 2746
rect 7102 2694 7104 2746
rect 6942 2692 6966 2694
rect 7022 2692 7046 2694
rect 7102 2692 7126 2694
rect 6886 2672 7182 2692
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6552 2304 6604 2310
rect 6552 2246 6604 2252
rect 6748 800 6776 2382
rect 7300 2378 7328 2790
rect 7378 2751 7434 2760
rect 7380 2508 7432 2514
rect 7484 2496 7512 8758
rect 7576 5098 7604 8871
rect 7760 8634 7788 11494
rect 7944 11218 7972 11834
rect 8116 11688 8168 11694
rect 8116 11630 8168 11636
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 11121 8064 11154
rect 8022 11112 8078 11121
rect 8022 11047 8078 11056
rect 8128 11014 8156 11630
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8298 11112 8354 11121
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8220 9654 8248 11086
rect 8298 11047 8300 11056
rect 8352 11047 8354 11056
rect 8300 11018 8352 11024
rect 8300 10600 8352 10606
rect 8404 10588 8432 11630
rect 9232 11218 9260 12310
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 8944 11144 8996 11150
rect 8942 11112 8944 11121
rect 8996 11112 8998 11121
rect 8942 11047 8998 11056
rect 8576 11008 8628 11014
rect 8576 10950 8628 10956
rect 8588 10849 8616 10950
rect 8574 10840 8630 10849
rect 8484 10804 8536 10810
rect 8574 10775 8630 10784
rect 8484 10746 8536 10752
rect 8496 10713 8524 10746
rect 8482 10704 8538 10713
rect 8482 10639 8538 10648
rect 8352 10560 8432 10588
rect 8300 10542 8352 10548
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8312 9518 8340 10542
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8864 10198 8892 10474
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9312 10056 9364 10062
rect 9310 10024 9312 10033
rect 9364 10024 9366 10033
rect 9128 9988 9180 9994
rect 9508 9994 9536 10066
rect 9310 9959 9366 9968
rect 9496 9988 9548 9994
rect 9128 9930 9180 9936
rect 9496 9930 9548 9936
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7944 7546 7972 8978
rect 8036 8090 8064 9046
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 8024 8084 8076 8090
rect 8024 8026 8076 8032
rect 8220 7818 8248 8910
rect 8312 8430 8340 9454
rect 9048 9382 9076 9862
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6458 7788 6734
rect 7748 6452 7800 6458
rect 7748 6394 7800 6400
rect 7852 6225 7880 7210
rect 8036 6984 8064 7686
rect 8404 7392 8432 8910
rect 8864 8838 8892 8978
rect 9140 8974 9168 9930
rect 9600 9738 9628 12582
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10140 12232 10192 12238
rect 10324 12232 10376 12238
rect 10192 12192 10272 12220
rect 10140 12174 10192 12180
rect 9852 11996 10148 12016
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 9930 11942 9932 11994
rect 9994 11942 10006 11994
rect 10068 11942 10070 11994
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 9852 11920 10148 11940
rect 10048 11824 10100 11830
rect 10100 11784 10180 11812
rect 10048 11766 10100 11772
rect 10046 11656 10102 11665
rect 10152 11626 10180 11784
rect 10046 11591 10048 11600
rect 10100 11591 10102 11600
rect 10140 11620 10192 11626
rect 10048 11562 10100 11568
rect 10140 11562 10192 11568
rect 10244 11558 10272 12192
rect 10324 12174 10376 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10336 11898 10364 12174
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10520 11694 10548 12174
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9784 11121 9812 11494
rect 10232 11144 10284 11150
rect 9770 11112 9826 11121
rect 10232 11086 10284 11092
rect 9770 11047 9826 11056
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9324 9710 9628 9738
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8852 8832 8904 8838
rect 8904 8792 8984 8820
rect 8852 8774 8904 8780
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8496 7750 8524 8026
rect 8588 7886 8616 8774
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8772 7410 8800 7822
rect 8864 7750 8892 8230
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8760 7404 8812 7410
rect 8404 7364 8524 7392
rect 8390 7304 8446 7313
rect 8390 7239 8446 7248
rect 8404 7206 8432 7239
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 7944 6956 8064 6984
rect 7838 6216 7894 6225
rect 7838 6151 7894 6160
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7668 5370 7696 5714
rect 7840 5704 7892 5710
rect 7838 5672 7840 5681
rect 7892 5672 7894 5681
rect 7838 5607 7894 5616
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7576 4826 7604 5034
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7852 4758 7880 5607
rect 7944 5030 7972 6956
rect 8024 6860 8076 6866
rect 8076 6820 8432 6848
rect 8024 6802 8076 6808
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 5914 8156 6598
rect 8300 6180 8352 6186
rect 8300 6122 8352 6128
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8312 5710 8340 6122
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8312 5234 8340 5646
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 8312 4826 8340 5170
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7562 4448 7618 4457
rect 7562 4383 7618 4392
rect 7576 3534 7604 4383
rect 8220 4282 8248 4626
rect 8404 4622 8432 6820
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 7656 4004 7708 4010
rect 7656 3946 7708 3952
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7576 2922 7604 3470
rect 7668 3194 7696 3946
rect 7944 3534 7972 4218
rect 8496 3754 8524 7364
rect 8760 7346 8812 7352
rect 8864 7206 8892 7686
rect 8852 7200 8904 7206
rect 8852 7142 8904 7148
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8588 5234 8616 5714
rect 8864 5710 8892 7142
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8864 5166 8892 5646
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8404 3726 8524 3754
rect 8404 3670 8432 3726
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8588 3398 8616 3839
rect 8666 3768 8722 3777
rect 8772 3738 8800 4422
rect 8666 3703 8668 3712
rect 8720 3703 8722 3712
rect 8760 3732 8812 3738
rect 8668 3674 8720 3680
rect 8760 3674 8812 3680
rect 8956 3534 8984 8792
rect 9140 8430 9168 8910
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9324 7954 9352 9710
rect 9692 9654 9720 10474
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9416 9178 9444 9454
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9402 8936 9458 8945
rect 9402 8871 9458 8880
rect 9416 8566 9444 8871
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9404 8560 9456 8566
rect 9404 8502 9456 8508
rect 9508 8498 9536 8774
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9600 8265 9628 8978
rect 9692 8634 9720 9386
rect 9784 9110 9812 11047
rect 9852 10908 10148 10928
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 9930 10854 9932 10906
rect 9994 10854 10006 10906
rect 10068 10854 10070 10906
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 9852 10832 10148 10852
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9876 10266 9904 10542
rect 9864 10260 9916 10266
rect 9864 10202 9916 10208
rect 10048 10192 10100 10198
rect 9954 10160 10010 10169
rect 10048 10134 10100 10140
rect 9954 10095 10010 10104
rect 9968 9994 9996 10095
rect 10060 10062 10088 10134
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 9956 9988 10008 9994
rect 9956 9930 10008 9936
rect 10244 9926 10272 11086
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10520 10062 10548 10610
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 9852 9820 10148 9840
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 9930 9766 9932 9818
rect 9994 9766 10006 9818
rect 10068 9766 10070 9818
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 9852 9744 10148 9764
rect 10336 9722 10364 9998
rect 10508 9920 10560 9926
rect 10508 9862 10560 9868
rect 10324 9716 10376 9722
rect 10324 9658 10376 9664
rect 10322 9616 10378 9625
rect 10140 9580 10192 9586
rect 10192 9540 10272 9568
rect 10322 9551 10324 9560
rect 10140 9522 10192 9528
rect 10244 9364 10272 9540
rect 10376 9551 10378 9560
rect 10324 9522 10376 9528
rect 10324 9376 10376 9382
rect 10244 9336 10324 9364
rect 10324 9318 10376 9324
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 9852 8732 10148 8752
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 9930 8678 9932 8730
rect 9994 8678 10006 8730
rect 10068 8678 10070 8730
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 9852 8656 10148 8676
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9876 8294 9904 8434
rect 10244 8362 10272 9046
rect 10336 8430 10364 9318
rect 10520 9042 10548 9862
rect 10612 9450 10640 12174
rect 10980 11898 11008 12242
rect 11072 12209 11100 12310
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 10968 11892 11020 11898
rect 10968 11834 11020 11840
rect 10782 11792 10838 11801
rect 11978 11792 12034 11801
rect 10782 11727 10784 11736
rect 10836 11727 10838 11736
rect 10968 11756 11020 11762
rect 10784 11698 10836 11704
rect 11978 11727 12034 11736
rect 10968 11698 11020 11704
rect 10980 11286 11008 11698
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11702 11656 11758 11665
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11336 11552 11388 11558
rect 11336 11494 11388 11500
rect 10968 11280 11020 11286
rect 10874 11248 10930 11257
rect 10968 11222 11020 11228
rect 10874 11183 10930 11192
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10704 10266 10732 10406
rect 10692 10260 10744 10266
rect 10692 10202 10744 10208
rect 10796 9722 10824 10406
rect 10784 9716 10836 9722
rect 10784 9658 10836 9664
rect 10600 9444 10652 9450
rect 10600 9386 10652 9392
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 9680 8288 9732 8294
rect 9586 8256 9642 8265
rect 9680 8230 9732 8236
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 9586 8191 9642 8200
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9496 7948 9548 7954
rect 9496 7890 9548 7896
rect 9404 7336 9456 7342
rect 9404 7278 9456 7284
rect 9416 7002 9444 7278
rect 9404 6996 9456 7002
rect 9324 6956 9404 6984
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9140 5642 9168 5850
rect 9128 5636 9180 5642
rect 9128 5578 9180 5584
rect 9140 5137 9168 5578
rect 9232 5166 9260 6054
rect 9220 5160 9272 5166
rect 9126 5128 9182 5137
rect 9220 5102 9272 5108
rect 9126 5063 9182 5072
rect 9324 4690 9352 6956
rect 9404 6938 9456 6944
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6186 9444 6598
rect 9404 6180 9456 6186
rect 9404 6122 9456 6128
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8864 3194 8892 3402
rect 9048 3194 9076 3538
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8944 3120 8996 3126
rect 7654 3088 7710 3097
rect 8944 3062 8996 3068
rect 7654 3023 7710 3032
rect 8760 3052 8812 3058
rect 7668 2990 7696 3023
rect 8760 2994 8812 3000
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 7564 2916 7616 2922
rect 7564 2858 7616 2864
rect 8300 2916 8352 2922
rect 8300 2858 8352 2864
rect 8312 2650 8340 2858
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 7432 2468 7512 2496
rect 7380 2450 7432 2456
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7576 800 7604 2382
rect 8496 800 8524 2926
rect 8772 2922 8800 2994
rect 8760 2916 8812 2922
rect 8760 2858 8812 2864
rect 8772 2582 8800 2858
rect 8956 2650 8984 3062
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8668 2576 8720 2582
rect 8668 2518 8720 2524
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 8680 2428 8708 2518
rect 9140 2446 9168 3946
rect 9312 3664 9364 3670
rect 9312 3606 9364 3612
rect 8760 2440 8812 2446
rect 8680 2400 8760 2428
rect 8760 2382 8812 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9324 1850 9352 3606
rect 9416 3534 9444 6122
rect 9508 5030 9536 7890
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9600 7274 9628 7482
rect 9692 7410 9720 8230
rect 9876 7993 9904 8230
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 9852 7644 10148 7664
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 9930 7590 9932 7642
rect 9994 7590 10006 7642
rect 10068 7590 10070 7642
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 9852 7568 10148 7588
rect 10336 7546 10364 7686
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 10428 7410 10456 8570
rect 10520 8430 10548 8978
rect 10888 8922 10916 11183
rect 10980 10674 11008 11222
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 11058 10568 11114 10577
rect 11058 10503 11114 10512
rect 11072 10266 11100 10503
rect 11060 10260 11112 10266
rect 11060 10202 11112 10208
rect 11150 10160 11206 10169
rect 11150 10095 11206 10104
rect 11164 10062 11192 10095
rect 11152 10056 11204 10062
rect 11058 10024 11114 10033
rect 10968 9988 11020 9994
rect 11152 9998 11204 10004
rect 11058 9959 11114 9968
rect 10968 9930 11020 9936
rect 10980 9586 11008 9930
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11072 9382 11100 9959
rect 11164 9897 11192 9998
rect 11150 9888 11206 9897
rect 11150 9823 11206 9832
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10796 8894 10916 8922
rect 10598 8800 10654 8809
rect 10598 8735 10654 8744
rect 10612 8430 10640 8735
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10612 8090 10640 8366
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10520 7585 10548 7958
rect 10506 7576 10562 7585
rect 10796 7562 10824 8894
rect 10980 8838 11008 9114
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10506 7511 10562 7520
rect 10612 7534 10824 7562
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 9588 7268 9640 7274
rect 9588 7210 9640 7216
rect 10324 7200 10376 7206
rect 10324 7142 10376 7148
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10336 6905 10364 7142
rect 10428 7041 10456 7142
rect 10414 7032 10470 7041
rect 10414 6967 10470 6976
rect 10322 6896 10378 6905
rect 10520 6866 10548 7414
rect 10322 6831 10378 6840
rect 10416 6860 10468 6866
rect 10416 6802 10468 6808
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9692 5166 9720 5646
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9416 2990 9444 3334
rect 9600 3058 9628 5102
rect 9784 4826 9812 6734
rect 9852 6556 10148 6576
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 9930 6502 9932 6554
rect 9994 6502 10006 6554
rect 10068 6502 10070 6554
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 9852 6480 10148 6500
rect 10244 5914 10272 6734
rect 10428 6458 10456 6802
rect 10612 6798 10640 7534
rect 10690 7440 10746 7449
rect 10690 7375 10746 7384
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10336 5914 10364 6054
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 9852 5468 10148 5488
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 9930 5414 9932 5466
rect 9994 5414 10006 5466
rect 10068 5414 10070 5466
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 9852 5392 10148 5412
rect 10244 5352 10272 5850
rect 10416 5840 10468 5846
rect 10414 5808 10416 5817
rect 10468 5808 10470 5817
rect 10324 5772 10376 5778
rect 10414 5743 10470 5752
rect 10324 5714 10376 5720
rect 10336 5370 10364 5714
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 9876 5324 10272 5352
rect 10324 5364 10376 5370
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4706 9904 5324
rect 10324 5306 10376 5312
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 9784 4678 9904 4706
rect 10152 4690 10180 4966
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10140 4684 10192 4690
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 4282 9720 4422
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9692 4078 9720 4218
rect 9784 4162 9812 4678
rect 10140 4626 10192 4632
rect 10244 4486 10272 4694
rect 10232 4480 10284 4486
rect 10230 4448 10232 4457
rect 10284 4448 10286 4457
rect 9852 4380 10148 4400
rect 10230 4383 10286 4392
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 9930 4326 9932 4378
rect 9994 4326 10006 4378
rect 10068 4326 10070 4378
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 9852 4304 10148 4324
rect 10232 4208 10284 4214
rect 9784 4146 9904 4162
rect 10232 4150 10284 4156
rect 9784 4140 9916 4146
rect 9784 4134 9864 4140
rect 9864 4082 9916 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3602 9812 4014
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9968 3602 9996 3878
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9404 2984 9456 2990
rect 9404 2926 9456 2932
rect 9692 2553 9720 3402
rect 9852 3292 10148 3312
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 9930 3238 9932 3290
rect 9994 3238 10006 3290
rect 10068 3238 10070 3290
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 9852 3216 10148 3236
rect 10244 3074 10272 4150
rect 10336 4078 10364 4966
rect 10428 4826 10456 5510
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10428 4146 10456 4422
rect 10520 4282 10548 6666
rect 10600 5840 10652 5846
rect 10600 5782 10652 5788
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10244 3046 10364 3074
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9678 2544 9734 2553
rect 9678 2479 9734 2488
rect 9784 2106 9812 2790
rect 10152 2650 10180 2790
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10152 2417 10180 2586
rect 10244 2582 10272 2926
rect 10336 2922 10364 3046
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 10138 2408 10194 2417
rect 10138 2343 10194 2352
rect 10428 2310 10456 3538
rect 10506 3224 10562 3233
rect 10506 3159 10562 3168
rect 10520 2961 10548 3159
rect 10612 2990 10640 5782
rect 10704 3942 10732 7375
rect 10888 7274 10916 8774
rect 11164 8634 11192 8978
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11060 8424 11112 8430
rect 10980 8384 11060 8412
rect 10980 7750 11008 8384
rect 11060 8366 11112 8372
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10782 7032 10838 7041
rect 10782 6967 10838 6976
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10704 3126 10732 3606
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10600 2984 10652 2990
rect 10506 2952 10562 2961
rect 10600 2926 10652 2932
rect 10506 2887 10562 2896
rect 10692 2916 10744 2922
rect 10692 2858 10744 2864
rect 10704 2650 10732 2858
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10796 2514 10824 6967
rect 10980 6934 11008 7686
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11072 6934 11100 7482
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 11060 6928 11112 6934
rect 11060 6870 11112 6876
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10888 5234 10916 6734
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10966 6352 11022 6361
rect 10966 6287 11022 6296
rect 10876 5228 10928 5234
rect 10876 5170 10928 5176
rect 10980 5114 11008 6287
rect 10888 5086 11008 5114
rect 10888 2990 10916 5086
rect 11072 4593 11100 6598
rect 11164 6322 11192 6802
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11256 5710 11284 11494
rect 11348 11354 11376 11494
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11428 11212 11480 11218
rect 11428 11154 11480 11160
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9058 11376 10066
rect 11440 9178 11468 11154
rect 11624 11150 11652 11630
rect 11702 11591 11758 11600
rect 11716 11558 11744 11591
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10470 11560 10950
rect 11624 10674 11652 11086
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11348 9030 11468 9058
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11348 8362 11376 8842
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7886 11376 8298
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11244 5704 11296 5710
rect 11164 5664 11244 5692
rect 11164 5030 11192 5664
rect 11244 5646 11296 5652
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11058 4584 11114 4593
rect 11058 4519 11114 4528
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4010 11192 4490
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 11152 4004 11204 4010
rect 11152 3946 11204 3952
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3738 11008 3878
rect 11072 3738 11100 3946
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11060 3732 11112 3738
rect 11060 3674 11112 3680
rect 11072 3482 11100 3674
rect 10980 3454 11100 3482
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 10980 3074 11008 3454
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3194 11100 3334
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10980 3046 11100 3074
rect 10876 2984 10928 2990
rect 10968 2984 11020 2990
rect 10876 2926 10928 2932
rect 10966 2952 10968 2961
rect 11020 2952 11022 2961
rect 10966 2887 11022 2896
rect 11072 2650 11100 3046
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11164 2530 11192 3470
rect 11072 2514 11192 2530
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 11060 2508 11192 2514
rect 11112 2502 11192 2508
rect 11060 2450 11112 2456
rect 11256 2446 11284 5510
rect 11348 4622 11376 7822
rect 11440 6644 11468 9030
rect 11520 8968 11572 8974
rect 11624 8945 11652 9318
rect 11520 8910 11572 8916
rect 11610 8936 11666 8945
rect 11532 8809 11560 8910
rect 11610 8871 11666 8880
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 11520 6656 11572 6662
rect 11440 6616 11520 6644
rect 11440 6118 11468 6616
rect 11520 6598 11572 6604
rect 11520 6248 11572 6254
rect 11518 6216 11520 6225
rect 11572 6216 11574 6225
rect 11518 6151 11574 6160
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11440 5914 11468 6054
rect 11428 5908 11480 5914
rect 11428 5850 11480 5856
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11336 4616 11388 4622
rect 11336 4558 11388 4564
rect 11440 4468 11468 5578
rect 11518 5264 11574 5273
rect 11518 5199 11574 5208
rect 11532 4826 11560 5199
rect 11520 4820 11572 4826
rect 11520 4762 11572 4768
rect 11624 4622 11652 8570
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11348 4440 11468 4468
rect 11348 3913 11376 4440
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11334 3904 11390 3913
rect 11334 3839 11390 3848
rect 11440 3534 11468 4082
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11532 3210 11560 4218
rect 11624 4214 11652 4558
rect 11612 4208 11664 4214
rect 11612 4150 11664 4156
rect 11612 3936 11664 3942
rect 11610 3904 11612 3913
rect 11664 3904 11666 3913
rect 11610 3839 11666 3848
rect 11348 3182 11560 3210
rect 11348 2650 11376 3182
rect 11716 3097 11744 11290
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11808 8634 11836 11222
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 10062 11928 10542
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11900 9178 11928 9318
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11992 8480 12020 11727
rect 12084 11354 12112 12038
rect 12176 11898 12204 13767
rect 12817 13628 13113 13648
rect 12873 13626 12897 13628
rect 12953 13626 12977 13628
rect 13033 13626 13057 13628
rect 12895 13574 12897 13626
rect 12959 13574 12971 13626
rect 13033 13574 13035 13626
rect 12873 13572 12897 13574
rect 12953 13572 12977 13574
rect 13033 13572 13057 13574
rect 12817 13552 13113 13572
rect 12817 12540 13113 12560
rect 12873 12538 12897 12540
rect 12953 12538 12977 12540
rect 13033 12538 13057 12540
rect 12895 12486 12897 12538
rect 12959 12486 12971 12538
rect 13033 12486 13035 12538
rect 12873 12484 12897 12486
rect 12953 12484 12977 12486
rect 13033 12484 13057 12486
rect 12817 12464 13113 12484
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12176 11801 12204 11834
rect 12162 11792 12218 11801
rect 12162 11727 12218 11736
rect 12817 11452 13113 11472
rect 12873 11450 12897 11452
rect 12953 11450 12977 11452
rect 13033 11450 13057 11452
rect 12895 11398 12897 11450
rect 12959 11398 12971 11450
rect 13033 11398 13035 11450
rect 12873 11396 12897 11398
rect 12953 11396 12977 11398
rect 13033 11396 13057 11398
rect 12817 11376 13113 11396
rect 12072 11348 12124 11354
rect 12072 11290 12124 11296
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12176 11257 12204 11290
rect 13176 11280 13228 11286
rect 12162 11248 12218 11257
rect 13176 11222 13228 11228
rect 12162 11183 12218 11192
rect 12164 11144 12216 11150
rect 12070 11112 12126 11121
rect 12348 11144 12400 11150
rect 12164 11086 12216 11092
rect 12254 11112 12310 11121
rect 12070 11047 12072 11056
rect 12124 11047 12126 11056
rect 12072 11018 12124 11024
rect 12176 10810 12204 11086
rect 12348 11086 12400 11092
rect 12438 11112 12494 11121
rect 12254 11047 12310 11056
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10742 12296 11047
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12256 10532 12308 10538
rect 12256 10474 12308 10480
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12084 9178 12112 10406
rect 12164 10124 12216 10130
rect 12164 10066 12216 10072
rect 12176 9722 12204 10066
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11900 8452 12020 8480
rect 11794 8120 11850 8129
rect 11900 8106 11928 8452
rect 11900 8078 12020 8106
rect 11794 8055 11796 8064
rect 11848 8055 11850 8064
rect 11796 8026 11848 8032
rect 11886 7984 11942 7993
rect 11886 7919 11888 7928
rect 11940 7919 11942 7928
rect 11888 7890 11940 7896
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11808 6186 11836 6870
rect 11900 6458 11928 7142
rect 11992 7018 12020 8078
rect 12084 7449 12112 9114
rect 12176 8974 12204 9658
rect 12164 8968 12216 8974
rect 12268 8945 12296 10474
rect 12164 8910 12216 8916
rect 12254 8936 12310 8945
rect 12254 8871 12310 8880
rect 12164 8288 12216 8294
rect 12256 8288 12308 8294
rect 12164 8230 12216 8236
rect 12254 8256 12256 8265
rect 12308 8256 12310 8265
rect 12176 7886 12204 8230
rect 12254 8191 12310 8200
rect 12360 8129 12388 11086
rect 12438 11047 12494 11056
rect 12716 11076 12768 11082
rect 12452 10810 12480 11047
rect 12716 11018 12768 11024
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12544 9382 12572 9823
rect 12532 9376 12584 9382
rect 12452 9336 12532 9364
rect 12346 8120 12402 8129
rect 12346 8055 12402 8064
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12070 7440 12126 7449
rect 12070 7375 12126 7384
rect 12176 7274 12204 7822
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 11992 6990 12204 7018
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 11888 6316 11940 6322
rect 11888 6258 11940 6264
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11900 5710 11928 6258
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11702 3088 11758 3097
rect 11702 3023 11758 3032
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11518 2816 11574 2825
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11440 2582 11468 2790
rect 11518 2751 11574 2760
rect 11532 2650 11560 2751
rect 11900 2650 11928 4082
rect 11992 3058 12020 5306
rect 12084 4282 12112 6394
rect 12176 5710 12204 6990
rect 12268 6662 12296 7278
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12256 6656 12308 6662
rect 12256 6598 12308 6604
rect 12268 6390 12296 6598
rect 12360 6497 12388 6938
rect 12452 6769 12480 9336
rect 12532 9318 12584 9324
rect 12532 9104 12584 9110
rect 12532 9046 12584 9052
rect 12544 8673 12572 9046
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12452 6662 12480 6695
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12346 6488 12402 6497
rect 12346 6423 12402 6432
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12256 6384 12308 6390
rect 12256 6326 12308 6332
rect 12256 6248 12308 6254
rect 12254 6216 12256 6225
rect 12308 6216 12310 6225
rect 12254 6151 12310 6160
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12256 5568 12308 5574
rect 12254 5536 12256 5545
rect 12308 5536 12310 5545
rect 12254 5471 12310 5480
rect 12162 5400 12218 5409
rect 12162 5335 12218 5344
rect 12176 5234 12204 5335
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12268 5114 12296 5471
rect 12360 5370 12388 5714
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5273 12480 6394
rect 12544 5778 12572 8502
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12636 8090 12664 8230
rect 12624 8084 12676 8090
rect 12624 8026 12676 8032
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12636 7002 12664 7142
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12728 5896 12756 11018
rect 12817 10364 13113 10384
rect 12873 10362 12897 10364
rect 12953 10362 12977 10364
rect 13033 10362 13057 10364
rect 12895 10310 12897 10362
rect 12959 10310 12971 10362
rect 13033 10310 13035 10362
rect 12873 10308 12897 10310
rect 12953 10308 12977 10310
rect 13033 10308 13057 10310
rect 12817 10288 13113 10308
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13096 9654 13124 10134
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12817 9276 13113 9296
rect 12873 9274 12897 9276
rect 12953 9274 12977 9276
rect 13033 9274 13057 9276
rect 12895 9222 12897 9274
rect 12959 9222 12971 9274
rect 13033 9222 13035 9274
rect 12873 9220 12897 9222
rect 12953 9220 12977 9222
rect 13033 9220 13057 9222
rect 12817 9200 13113 9220
rect 13084 9036 13136 9042
rect 13188 9024 13216 11222
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 9926 13308 10474
rect 13360 9988 13412 9994
rect 13360 9930 13412 9936
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13280 9586 13308 9862
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13372 9382 13400 9930
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13136 8996 13216 9024
rect 13084 8978 13136 8984
rect 13096 8537 13124 8978
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 13082 8528 13138 8537
rect 13188 8498 13216 8842
rect 13280 8634 13308 9318
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13372 8566 13400 9318
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13082 8463 13138 8472
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 12817 8188 13113 8208
rect 12873 8186 12897 8188
rect 12953 8186 12977 8188
rect 13033 8186 13057 8188
rect 12895 8134 12897 8186
rect 12959 8134 12971 8186
rect 13033 8134 13035 8186
rect 12873 8132 12897 8134
rect 12953 8132 12977 8134
rect 13033 8132 13057 8134
rect 12817 8112 13113 8132
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12820 7546 12848 7958
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12817 7100 13113 7120
rect 12873 7098 12897 7100
rect 12953 7098 12977 7100
rect 13033 7098 13057 7100
rect 12895 7046 12897 7098
rect 12959 7046 12971 7098
rect 13033 7046 13035 7098
rect 12873 7044 12897 7046
rect 12953 7044 12977 7046
rect 13033 7044 13057 7046
rect 12817 7024 13113 7044
rect 13084 6384 13136 6390
rect 12806 6352 12862 6361
rect 13084 6326 13136 6332
rect 12806 6287 12862 6296
rect 12820 6254 12848 6287
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 13096 6186 13124 6326
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12817 6012 13113 6032
rect 12873 6010 12897 6012
rect 12953 6010 12977 6012
rect 13033 6010 13057 6012
rect 12895 5958 12897 6010
rect 12959 5958 12971 6010
rect 13033 5958 13035 6010
rect 12873 5956 12897 5958
rect 12953 5956 12977 5958
rect 13033 5956 13057 5958
rect 12817 5936 13113 5956
rect 12636 5868 12756 5896
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12438 5264 12494 5273
rect 12438 5199 12494 5208
rect 12176 5098 12296 5114
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12164 5092 12296 5098
rect 12216 5086 12296 5092
rect 12164 5034 12216 5040
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 4622 12296 4966
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12360 4554 12388 5102
rect 12544 4758 12572 5510
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12452 4282 12480 4626
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12438 4176 12494 4185
rect 12438 4111 12494 4120
rect 12452 3777 12480 4111
rect 12438 3768 12494 3777
rect 12438 3703 12494 3712
rect 12346 3224 12402 3233
rect 12544 3194 12572 4558
rect 12346 3159 12402 3168
rect 12532 3188 12584 3194
rect 12360 3058 12388 3159
rect 12532 3130 12584 3136
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12440 2984 12492 2990
rect 12636 2961 12664 5868
rect 13188 5794 13216 8298
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13280 5914 13308 6802
rect 13464 6338 13492 14991
rect 13924 14006 13952 16400
rect 15014 15736 15070 15745
rect 15014 15671 15070 15680
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 13924 11898 13952 13942
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 13728 9988 13780 9994
rect 13728 9930 13780 9936
rect 13740 9722 13768 9930
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 13728 9716 13780 9722
rect 13728 9658 13780 9664
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13832 9194 13860 9658
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 13740 9166 13860 9194
rect 13634 8800 13690 8809
rect 13634 8735 13690 8744
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 7993 13584 8230
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 13556 7478 13584 7919
rect 13648 7886 13676 8735
rect 13740 8673 13768 9166
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13726 8664 13782 8673
rect 13726 8599 13782 8608
rect 13832 8498 13860 9046
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13740 7954 13768 8298
rect 13728 7948 13780 7954
rect 13728 7890 13780 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13832 7818 13860 8434
rect 13924 8090 13952 9590
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13544 7472 13596 7478
rect 13544 7414 13596 7420
rect 13556 6934 13584 7414
rect 13924 7342 13952 7822
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13544 6928 13596 6934
rect 13544 6870 13596 6876
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13634 6760 13690 6769
rect 13372 6310 13492 6338
rect 13556 6322 13584 6734
rect 13634 6695 13690 6704
rect 13544 6316 13596 6322
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13372 5817 13400 6310
rect 13544 6258 13596 6264
rect 13452 6248 13504 6254
rect 13452 6190 13504 6196
rect 13358 5808 13414 5817
rect 12716 5772 12768 5778
rect 13188 5766 13308 5794
rect 12716 5714 12768 5720
rect 12728 4826 12756 5714
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12817 4924 13113 4944
rect 12873 4922 12897 4924
rect 12953 4922 12977 4924
rect 13033 4922 13057 4924
rect 12895 4870 12897 4922
rect 12959 4870 12971 4922
rect 13033 4870 13035 4922
rect 12873 4868 12897 4870
rect 12953 4868 12977 4870
rect 13033 4868 13057 4870
rect 12817 4848 13113 4868
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 13188 4554 13216 5646
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13280 4146 13308 5766
rect 13358 5743 13414 5752
rect 13372 4826 13400 5743
rect 13464 4826 13492 6190
rect 13542 5944 13598 5953
rect 13542 5879 13598 5888
rect 13556 5846 13584 5879
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13542 5672 13598 5681
rect 13542 5607 13598 5616
rect 13556 5302 13584 5607
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13372 4570 13400 4762
rect 13648 4729 13676 6695
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13740 5409 13768 6190
rect 13726 5400 13782 5409
rect 13726 5335 13782 5344
rect 13740 5098 13768 5335
rect 13728 5092 13780 5098
rect 13728 5034 13780 5040
rect 13634 4720 13690 4729
rect 13634 4655 13690 4664
rect 13372 4542 13492 4570
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12817 3836 13113 3856
rect 12873 3834 12897 3836
rect 12953 3834 12977 3836
rect 13033 3834 13057 3836
rect 12895 3782 12897 3834
rect 12959 3782 12971 3834
rect 13033 3782 13035 3834
rect 12873 3780 12897 3782
rect 12953 3780 12977 3782
rect 13033 3780 13057 3782
rect 12817 3760 13113 3780
rect 12808 3664 12860 3670
rect 12808 3606 12860 3612
rect 12820 3466 12848 3606
rect 12808 3460 12860 3466
rect 12808 3402 12860 3408
rect 13188 3058 13216 3878
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12440 2926 12492 2932
rect 12622 2952 12678 2961
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11428 2576 11480 2582
rect 11428 2518 11480 2524
rect 11704 2576 11756 2582
rect 11704 2518 11756 2524
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11716 2310 11744 2518
rect 10416 2304 10468 2310
rect 10414 2272 10416 2281
rect 11704 2304 11756 2310
rect 10468 2272 10470 2281
rect 9852 2204 10148 2224
rect 11704 2246 11756 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 10414 2207 10470 2216
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 9930 2150 9932 2202
rect 9994 2150 10006 2202
rect 10068 2150 10070 2202
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 9852 2128 10148 2148
rect 12084 2106 12112 2246
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 9324 1822 9444 1850
rect 9416 800 9444 1822
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10336 800 10364 1430
rect 11244 1148 11296 1154
rect 11244 1090 11296 1096
rect 11256 800 11284 1090
rect 12176 800 12204 2518
rect 12452 2446 12480 2926
rect 12622 2887 12678 2896
rect 13268 2916 13320 2922
rect 13268 2858 13320 2864
rect 12817 2748 13113 2768
rect 12873 2746 12897 2748
rect 12953 2746 12977 2748
rect 13033 2746 13057 2748
rect 12895 2694 12897 2746
rect 12959 2694 12971 2746
rect 13033 2694 13035 2746
rect 12873 2692 12897 2694
rect 12953 2692 12977 2694
rect 13033 2692 13057 2694
rect 12817 2672 13113 2692
rect 12440 2440 12492 2446
rect 12440 2382 12492 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 13188 2281 13216 2382
rect 13174 2272 13230 2281
rect 13174 2207 13230 2216
rect 13280 1442 13308 2858
rect 13372 2514 13400 4422
rect 13464 4264 13492 4542
rect 13464 4236 13584 4264
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13464 3670 13492 4082
rect 13556 4010 13584 4236
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13452 3664 13504 3670
rect 13452 3606 13504 3612
rect 13544 3392 13596 3398
rect 13464 3340 13544 3346
rect 13464 3334 13596 3340
rect 13464 3318 13584 3334
rect 13464 3058 13492 3318
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13648 2854 13676 4655
rect 13740 4622 13768 5034
rect 13832 4842 13860 6870
rect 13912 6792 13964 6798
rect 13910 6760 13912 6769
rect 13964 6760 13966 6769
rect 13910 6695 13966 6704
rect 13910 6488 13966 6497
rect 13910 6423 13966 6432
rect 13924 5846 13952 6423
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13924 5370 13952 5646
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13832 4814 13952 4842
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13818 4584 13874 4593
rect 13740 3602 13768 4558
rect 13818 4519 13874 4528
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 13832 2514 13860 4519
rect 13924 3942 13952 4814
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13924 3670 13952 3878
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 14016 3126 14044 9862
rect 14094 9480 14150 9489
rect 14094 9415 14150 9424
rect 14108 9382 14136 9415
rect 14200 9382 14228 11018
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14188 9376 14240 9382
rect 14188 9318 14240 9324
rect 14108 9110 14136 9318
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14108 8634 14136 9046
rect 14096 8628 14148 8634
rect 14096 8570 14148 8576
rect 14200 8514 14228 9318
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14292 8945 14320 9046
rect 14278 8936 14334 8945
rect 14278 8871 14334 8880
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 14108 8486 14228 8514
rect 14108 4282 14136 8486
rect 14292 8430 14320 8774
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14200 5522 14228 8026
rect 14292 7410 14320 8366
rect 14384 7750 14412 11698
rect 14476 11286 14504 11766
rect 14924 11688 14976 11694
rect 14646 11656 14702 11665
rect 14924 11630 14976 11636
rect 14646 11591 14702 11600
rect 14464 11280 14516 11286
rect 14464 11222 14516 11228
rect 14464 11008 14516 11014
rect 14464 10950 14516 10956
rect 14476 9722 14504 10950
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14568 9654 14596 10066
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14372 6996 14424 7002
rect 14372 6938 14424 6944
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14292 6186 14320 6734
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14292 5710 14320 6122
rect 14384 5778 14412 6938
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14280 5704 14332 5710
rect 14278 5672 14280 5681
rect 14332 5672 14334 5681
rect 14278 5607 14334 5616
rect 14200 5494 14320 5522
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14200 5273 14228 5306
rect 14186 5264 14242 5273
rect 14186 5199 14242 5208
rect 14200 5030 14228 5199
rect 14188 5024 14240 5030
rect 14188 4966 14240 4972
rect 14292 4842 14320 5494
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14200 4814 14320 4842
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14200 3942 14228 4814
rect 14280 4684 14332 4690
rect 14384 4672 14412 5170
rect 14476 4690 14504 8298
rect 14568 7002 14596 9046
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 6254 14596 6598
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14660 6118 14688 11591
rect 14936 11218 14964 11630
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 15028 11082 15056 15671
rect 15474 15464 15530 15473
rect 15474 15399 15530 15408
rect 15198 14648 15254 14657
rect 15198 14583 15254 14592
rect 15212 12170 15240 14583
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 14832 11076 14884 11082
rect 14832 11018 14884 11024
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14740 10532 14792 10538
rect 14740 10474 14792 10480
rect 14752 10062 14780 10474
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14752 8090 14780 9658
rect 14844 9382 14872 11018
rect 14924 11008 14976 11014
rect 14924 10950 14976 10956
rect 14936 10810 14964 10950
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14832 9376 14884 9382
rect 14832 9318 14884 9324
rect 14844 9178 14872 9318
rect 14832 9172 14884 9178
rect 14832 9114 14884 9120
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14752 7818 14780 8026
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14738 7576 14794 7585
rect 14738 7511 14794 7520
rect 14752 7002 14780 7511
rect 14844 7313 14872 7686
rect 14830 7304 14886 7313
rect 14830 7239 14886 7248
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14936 6882 14964 10746
rect 15120 10606 15148 11086
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10062 15148 10542
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15016 9920 15068 9926
rect 15014 9888 15016 9897
rect 15068 9888 15070 9897
rect 15014 9823 15070 9832
rect 15028 9722 15056 9823
rect 15016 9716 15068 9722
rect 15016 9658 15068 9664
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15028 9178 15056 9522
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 15120 8838 15148 9998
rect 15212 9654 15240 11562
rect 15384 11212 15436 11218
rect 15304 11172 15384 11200
rect 15304 10470 15332 11172
rect 15384 11154 15436 11160
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 9648 15252 9654
rect 15200 9590 15252 9596
rect 15304 9586 15332 10406
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15028 7750 15056 8366
rect 15396 8022 15424 10406
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15108 7744 15160 7750
rect 15108 7686 15160 7692
rect 15016 7540 15068 7546
rect 15016 7482 15068 7488
rect 15028 6934 15056 7482
rect 14844 6854 14964 6882
rect 15016 6928 15068 6934
rect 15016 6870 15068 6876
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14844 5778 14872 6854
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 15014 6760 15070 6769
rect 14936 6186 14964 6734
rect 15014 6695 15070 6704
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14832 5772 14884 5778
rect 14832 5714 14884 5720
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14556 4752 14608 4758
rect 14556 4694 14608 4700
rect 14332 4644 14412 4672
rect 14464 4684 14516 4690
rect 14280 4626 14332 4632
rect 14464 4626 14516 4632
rect 14292 4146 14320 4626
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14108 2553 14136 2926
rect 14200 2922 14228 3878
rect 14292 3398 14320 4082
rect 14476 4078 14504 4626
rect 14568 4146 14596 4694
rect 14660 4457 14688 4966
rect 14646 4448 14702 4457
rect 14646 4383 14702 4392
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14188 2916 14240 2922
rect 14188 2858 14240 2864
rect 14094 2544 14150 2553
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13820 2508 13872 2514
rect 14094 2479 14150 2488
rect 13820 2450 13872 2456
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13096 1414 13308 1442
rect 13096 800 13124 1414
rect 13648 1154 13676 2382
rect 13912 2372 13964 2378
rect 13912 2314 13964 2320
rect 13636 1148 13688 1154
rect 13636 1090 13688 1096
rect 13924 800 13952 2314
rect 14292 1494 14320 2994
rect 14660 2990 14688 4383
rect 14752 3942 14780 5646
rect 14922 5536 14978 5545
rect 14922 5471 14978 5480
rect 14936 5166 14964 5471
rect 15028 5370 15056 6695
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14740 3936 14792 3942
rect 14740 3878 14792 3884
rect 14752 3670 14780 3878
rect 14740 3664 14792 3670
rect 14740 3606 14792 3612
rect 14752 3233 14780 3606
rect 14738 3224 14794 3233
rect 14738 3159 14794 3168
rect 14752 3126 14780 3159
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 15028 2582 15056 4150
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 15120 2514 15148 7686
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15396 6730 15424 7278
rect 15488 6934 15516 15399
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15580 11257 15608 11290
rect 15566 11248 15622 11257
rect 15566 11183 15622 11192
rect 15672 11132 15700 16487
rect 16210 14240 16266 14249
rect 15782 14172 16078 14192
rect 16210 14175 16266 14184
rect 15838 14170 15862 14172
rect 15918 14170 15942 14172
rect 15998 14170 16022 14172
rect 15860 14118 15862 14170
rect 15924 14118 15936 14170
rect 15998 14118 16000 14170
rect 15838 14116 15862 14118
rect 15918 14116 15942 14118
rect 15998 14116 16022 14118
rect 15782 14096 16078 14116
rect 15782 13084 16078 13104
rect 15838 13082 15862 13084
rect 15918 13082 15942 13084
rect 15998 13082 16022 13084
rect 15860 13030 15862 13082
rect 15924 13030 15936 13082
rect 15998 13030 16000 13082
rect 15838 13028 15862 13030
rect 15918 13028 15942 13030
rect 15998 13028 16022 13030
rect 15782 13008 16078 13028
rect 15750 12744 15806 12753
rect 15750 12679 15806 12688
rect 15764 12646 15792 12679
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15750 12336 15806 12345
rect 15750 12271 15806 12280
rect 15764 12238 15792 12271
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15782 11996 16078 12016
rect 15838 11994 15862 11996
rect 15918 11994 15942 11996
rect 15998 11994 16022 11996
rect 15860 11942 15862 11994
rect 15924 11942 15936 11994
rect 15998 11942 16000 11994
rect 15838 11940 15862 11942
rect 15918 11940 15942 11942
rect 15998 11940 16022 11942
rect 15782 11920 16078 11940
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11354 15792 11494
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 16224 11286 16252 14175
rect 16394 13560 16450 13569
rect 16394 13495 16450 13504
rect 16302 11928 16358 11937
rect 16302 11863 16358 11872
rect 16316 11830 16344 11863
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 15580 11104 15700 11132
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15384 6724 15436 6730
rect 15384 6666 15436 6672
rect 15212 6390 15240 6666
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6390 15332 6598
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 6180 15252 6186
rect 15200 6122 15252 6128
rect 15212 5778 15240 6122
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5030 15240 5714
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15200 5024 15252 5030
rect 15200 4966 15252 4972
rect 15212 4622 15240 4966
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15212 4146 15240 4558
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15198 3088 15254 3097
rect 15198 3023 15254 3032
rect 15212 2650 15240 3023
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15304 2514 15332 5510
rect 15396 3466 15424 6666
rect 15488 5914 15516 6870
rect 15580 6866 15608 11104
rect 15782 10908 16078 10928
rect 15838 10906 15862 10908
rect 15918 10906 15942 10908
rect 15998 10906 16022 10908
rect 15860 10854 15862 10906
rect 15924 10854 15936 10906
rect 15998 10854 16000 10906
rect 15838 10852 15862 10854
rect 15918 10852 15942 10854
rect 15998 10852 16022 10854
rect 15782 10832 16078 10852
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16040 10130 16068 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15672 9110 15700 9862
rect 15782 9820 16078 9840
rect 15838 9818 15862 9820
rect 15918 9818 15942 9820
rect 15998 9818 16022 9820
rect 15860 9766 15862 9818
rect 15924 9766 15936 9818
rect 15998 9766 16000 9818
rect 15838 9764 15862 9766
rect 15918 9764 15942 9766
rect 15998 9764 16022 9766
rect 15782 9744 16078 9764
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16132 9382 16160 9658
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15948 9178 15976 9318
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15672 7886 15700 9046
rect 16118 8936 16174 8945
rect 16118 8871 16174 8880
rect 15782 8732 16078 8752
rect 15838 8730 15862 8732
rect 15918 8730 15942 8732
rect 15998 8730 16022 8732
rect 15860 8678 15862 8730
rect 15924 8678 15936 8730
rect 15998 8678 16000 8730
rect 15838 8676 15862 8678
rect 15918 8676 15942 8678
rect 15998 8676 16022 8678
rect 15782 8656 16078 8676
rect 16132 8634 16160 8871
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16224 8378 16252 10202
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 16316 8838 16344 9318
rect 16304 8832 16356 8838
rect 16304 8774 16356 8780
rect 16316 8498 16344 8774
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16302 8392 16358 8401
rect 16224 8350 16302 8378
rect 16408 8378 16436 13495
rect 16500 10266 16528 16895
rect 17866 16400 17922 17200
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17328 13870 17356 14282
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17420 13530 17448 14010
rect 17880 13938 17908 16400
rect 18418 16144 18474 16153
rect 18418 16079 18474 16088
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 18064 13870 18092 14214
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16960 11286 16988 12378
rect 17512 11676 17540 13670
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17420 11648 17540 11676
rect 16948 11280 17000 11286
rect 16948 11222 17000 11228
rect 17224 11280 17276 11286
rect 17276 11240 17356 11268
rect 17224 11222 17276 11228
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10538 16620 10950
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16672 10532 16724 10538
rect 16672 10474 16724 10480
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16592 10198 16620 10474
rect 16580 10192 16632 10198
rect 16580 10134 16632 10140
rect 16486 10024 16542 10033
rect 16486 9959 16542 9968
rect 16580 9988 16632 9994
rect 16500 9178 16528 9959
rect 16580 9930 16632 9936
rect 16592 9654 16620 9930
rect 16684 9654 16712 10474
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16776 10266 16804 10406
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16580 9648 16632 9654
rect 16580 9590 16632 9596
rect 16672 9648 16724 9654
rect 16868 9625 16896 11018
rect 16672 9590 16724 9596
rect 16854 9616 16910 9625
rect 16854 9551 16910 9560
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16488 9172 16540 9178
rect 16488 9114 16540 9120
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16592 8430 16620 8774
rect 16580 8424 16632 8430
rect 16408 8350 16528 8378
rect 16580 8366 16632 8372
rect 16302 8327 16358 8336
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 15782 7644 16078 7664
rect 15838 7642 15862 7644
rect 15918 7642 15942 7644
rect 15998 7642 16022 7644
rect 15860 7590 15862 7642
rect 15924 7590 15936 7642
rect 15998 7590 16000 7642
rect 15838 7588 15862 7590
rect 15918 7588 15942 7590
rect 15998 7588 16022 7590
rect 15782 7568 16078 7588
rect 16224 7206 16252 7754
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15672 6934 15700 7142
rect 15948 7002 15976 7142
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15660 6928 15712 6934
rect 15660 6870 15712 6876
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15488 5166 15516 5850
rect 15580 5846 15608 6802
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15672 5710 15700 6870
rect 15782 6556 16078 6576
rect 15838 6554 15862 6556
rect 15918 6554 15942 6556
rect 15998 6554 16022 6556
rect 15860 6502 15862 6554
rect 15924 6502 15936 6554
rect 15998 6502 16000 6554
rect 15838 6500 15862 6502
rect 15918 6500 15942 6502
rect 15998 6500 16022 6502
rect 15782 6480 16078 6500
rect 16132 6322 16160 7142
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 15764 5914 15792 6054
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 16224 5846 16252 6054
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 16120 5704 16172 5710
rect 16316 5658 16344 8327
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 7410 16436 8230
rect 16500 7857 16528 8350
rect 16592 8022 16620 8366
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16486 7848 16542 7857
rect 16486 7783 16542 7792
rect 16580 7744 16632 7750
rect 16580 7686 16632 7692
rect 16592 7410 16620 7686
rect 16684 7410 16712 8298
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16408 6390 16436 7346
rect 16776 7290 16804 9386
rect 16868 8430 16896 9551
rect 16960 9450 16988 11222
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17144 10266 17172 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17236 10470 17264 10746
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16960 8090 16988 8774
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16856 7948 16908 7954
rect 17052 7936 17080 9687
rect 17144 9081 17172 10202
rect 17130 9072 17186 9081
rect 17130 9007 17186 9016
rect 16908 7908 17080 7936
rect 16856 7890 16908 7896
rect 16868 7546 16896 7890
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16592 7262 16804 7290
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16592 6798 16620 7262
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 16592 6662 16620 6734
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16684 6186 16712 7142
rect 16960 6905 16988 7278
rect 16946 6896 17002 6905
rect 16856 6860 16908 6866
rect 16946 6831 17002 6840
rect 16856 6802 16908 6808
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16672 6180 16724 6186
rect 16672 6122 16724 6128
rect 16120 5646 16172 5652
rect 15580 5352 15608 5646
rect 15782 5468 16078 5488
rect 15838 5466 15862 5468
rect 15918 5466 15942 5468
rect 15998 5466 16022 5468
rect 15860 5414 15862 5466
rect 15924 5414 15936 5466
rect 15998 5414 16000 5466
rect 15838 5412 15862 5414
rect 15918 5412 15942 5414
rect 15998 5412 16022 5414
rect 15782 5392 16078 5412
rect 15580 5324 15700 5352
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15384 3460 15436 3466
rect 15384 3402 15436 3408
rect 15396 3194 15424 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15382 3088 15438 3097
rect 15382 3023 15384 3032
rect 15436 3023 15438 3032
rect 15384 2994 15436 3000
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15292 2508 15344 2514
rect 15292 2450 15344 2456
rect 14832 2440 14884 2446
rect 15396 2417 15424 2994
rect 15488 2854 15516 4966
rect 15580 4758 15608 5170
rect 15672 5030 15700 5324
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15568 4752 15620 4758
rect 15568 4694 15620 4700
rect 15782 4380 16078 4400
rect 15838 4378 15862 4380
rect 15918 4378 15942 4380
rect 15998 4378 16022 4380
rect 15860 4326 15862 4378
rect 15924 4326 15936 4378
rect 15998 4326 16000 4378
rect 15838 4324 15862 4326
rect 15918 4324 15942 4326
rect 15998 4324 16022 4326
rect 15782 4304 16078 4324
rect 16132 3738 16160 5646
rect 16224 5630 16344 5658
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16224 3602 16252 5630
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 16212 3596 16264 3602
rect 16212 3538 16264 3544
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15948 3482 15976 3538
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15580 2990 15608 3334
rect 15568 2984 15620 2990
rect 15568 2926 15620 2932
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 14832 2382 14884 2388
rect 15382 2408 15438 2417
rect 14280 1488 14332 1494
rect 14280 1430 14332 1436
rect 14844 800 14872 2382
rect 15382 2343 15438 2352
rect 15672 1850 15700 3470
rect 15948 3454 16160 3482
rect 15782 3292 16078 3312
rect 15838 3290 15862 3292
rect 15918 3290 15942 3292
rect 15998 3290 16022 3292
rect 15860 3238 15862 3290
rect 15924 3238 15936 3290
rect 15998 3238 16000 3290
rect 15838 3236 15862 3238
rect 15918 3236 15942 3238
rect 15998 3236 16022 3238
rect 15782 3216 16078 3236
rect 16132 2854 16160 3454
rect 16224 2990 16252 3538
rect 16316 3534 16344 5238
rect 16776 5234 16804 6666
rect 16868 6662 16896 6802
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16868 5846 16896 6598
rect 16960 6254 16988 6598
rect 17052 6322 17080 7686
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16764 5228 16816 5234
rect 16868 5216 16896 5782
rect 17144 5370 17172 9007
rect 17236 8974 17264 10406
rect 17328 10169 17356 11240
rect 17314 10160 17370 10169
rect 17314 10095 17370 10104
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17328 9586 17356 9998
rect 17420 9722 17448 11648
rect 17684 11552 17736 11558
rect 17684 11494 17736 11500
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17328 8650 17356 9386
rect 17236 8622 17356 8650
rect 17236 5778 17264 8622
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 6662 17356 6734
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17328 5846 17356 6598
rect 17316 5840 17368 5846
rect 17316 5782 17368 5788
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16948 5228 17000 5234
rect 16868 5188 16948 5216
rect 16764 5170 16816 5176
rect 16948 5170 17000 5176
rect 17236 5030 17264 5714
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 16580 5024 16632 5030
rect 16580 4966 16632 4972
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17224 5024 17276 5030
rect 17224 4966 17276 4972
rect 16592 3670 16620 4966
rect 16948 4752 17000 4758
rect 16946 4720 16948 4729
rect 17040 4752 17092 4758
rect 17000 4720 17002 4729
rect 17040 4694 17092 4700
rect 16946 4655 17002 4664
rect 16960 4622 16988 4655
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 16672 4480 16724 4486
rect 16672 4422 16724 4428
rect 16684 4214 16712 4422
rect 16672 4208 16724 4214
rect 16672 4150 16724 4156
rect 16946 4176 17002 4185
rect 16580 3664 16632 3670
rect 16580 3606 16632 3612
rect 16684 3534 16712 4150
rect 17052 4146 17080 4694
rect 16946 4111 17002 4120
rect 17040 4140 17092 4146
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 16776 3641 16804 4014
rect 16960 4010 16988 4111
rect 17040 4082 17092 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16856 3936 16908 3942
rect 16856 3878 16908 3884
rect 16868 3738 16896 3878
rect 16960 3738 16988 3946
rect 16856 3732 16908 3738
rect 16856 3674 16908 3680
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16762 3632 16818 3641
rect 16818 3590 16896 3618
rect 16762 3567 16818 3576
rect 16304 3528 16356 3534
rect 16672 3528 16724 3534
rect 16304 3470 16356 3476
rect 16486 3496 16542 3505
rect 16486 3431 16542 3440
rect 16592 3476 16672 3482
rect 16592 3470 16724 3476
rect 16592 3454 16712 3470
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 16500 2938 16528 3431
rect 16592 3126 16620 3454
rect 16672 3392 16724 3398
rect 16672 3334 16724 3340
rect 16580 3120 16632 3126
rect 16580 3062 16632 3068
rect 16684 3058 16712 3334
rect 16868 3058 16896 3590
rect 17052 3194 17080 4082
rect 17144 4078 17172 4966
rect 17236 4570 17264 4966
rect 17328 4690 17356 5102
rect 17316 4684 17368 4690
rect 17316 4626 17368 4632
rect 17236 4542 17356 4570
rect 17328 4486 17356 4542
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17236 4146 17264 4422
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17314 4040 17370 4049
rect 17314 3975 17370 3984
rect 17328 3194 17356 3975
rect 17040 3188 17092 3194
rect 17040 3130 17092 3136
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 17328 2990 17356 3130
rect 17316 2984 17368 2990
rect 16500 2910 16712 2938
rect 17420 2972 17448 9522
rect 17512 9110 17540 11018
rect 17696 10441 17724 11494
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10674 17908 11154
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17868 10464 17920 10470
rect 17682 10432 17738 10441
rect 17868 10406 17920 10412
rect 17682 10367 17738 10376
rect 17776 10124 17828 10130
rect 17776 10066 17828 10072
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 9178 17632 9862
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 9104 17552 9110
rect 17500 9046 17552 9052
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17512 8090 17540 8570
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 7410 17540 7754
rect 17604 7449 17632 8774
rect 17696 8129 17724 9590
rect 17788 9518 17816 10066
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17776 9376 17828 9382
rect 17880 9353 17908 10406
rect 17972 10266 18000 11834
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17972 9450 18000 9862
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17776 9318 17828 9324
rect 17866 9344 17922 9353
rect 17788 8537 17816 9318
rect 17866 9279 17922 9288
rect 17960 9036 18012 9042
rect 17960 8978 18012 8984
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17774 8528 17830 8537
rect 17774 8463 17830 8472
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17682 8120 17738 8129
rect 17682 8055 17738 8064
rect 17684 7880 17736 7886
rect 17682 7848 17684 7857
rect 17736 7848 17738 7857
rect 17682 7783 17738 7792
rect 17590 7440 17646 7449
rect 17500 7404 17552 7410
rect 17590 7375 17646 7384
rect 17500 7346 17552 7352
rect 17512 6798 17540 7346
rect 17500 6792 17552 6798
rect 17788 6769 17816 8230
rect 17880 7857 17908 8842
rect 17972 8294 18000 8978
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 18064 7546 18092 13262
rect 18142 13152 18198 13161
rect 18142 13087 18198 13096
rect 18156 12209 18184 13087
rect 18142 12200 18198 12209
rect 18142 12135 18198 12144
rect 18156 11898 18184 12135
rect 18144 11892 18196 11898
rect 18144 11834 18196 11840
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18156 10606 18184 11222
rect 18248 10849 18276 11698
rect 18234 10840 18290 10849
rect 18234 10775 18290 10784
rect 18144 10600 18196 10606
rect 18248 10577 18276 10775
rect 18144 10542 18196 10548
rect 18234 10568 18290 10577
rect 18234 10503 18290 10512
rect 18248 9926 18276 10503
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 9042 18276 9318
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18144 8288 18196 8294
rect 18144 8230 18196 8236
rect 18156 7954 18184 8230
rect 18144 7948 18196 7954
rect 18144 7890 18196 7896
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17868 7336 17920 7342
rect 17868 7278 17920 7284
rect 17500 6734 17552 6740
rect 17774 6760 17830 6769
rect 17774 6695 17830 6704
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17512 5778 17540 6394
rect 17880 6254 17908 7278
rect 17868 6248 17920 6254
rect 17774 6216 17830 6225
rect 17868 6190 17920 6196
rect 17774 6151 17830 6160
rect 17788 6118 17816 6151
rect 17776 6112 17828 6118
rect 17776 6054 17828 6060
rect 17500 5772 17552 5778
rect 17500 5714 17552 5720
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17604 5030 17632 5306
rect 17788 5302 17816 5510
rect 17776 5296 17828 5302
rect 17776 5238 17828 5244
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 5024 17644 5030
rect 17512 4984 17592 5012
rect 17512 3738 17540 4984
rect 17592 4966 17644 4972
rect 17696 4622 17724 5170
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17604 3194 17632 4422
rect 17788 4214 17816 5238
rect 17972 5098 18000 7346
rect 18052 7336 18104 7342
rect 18050 7304 18052 7313
rect 18104 7304 18106 7313
rect 18050 7239 18106 7248
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 5137 18092 5510
rect 18050 5128 18106 5137
rect 17960 5092 18012 5098
rect 18050 5063 18106 5072
rect 17960 5034 18012 5040
rect 18052 4548 18104 4554
rect 18052 4490 18104 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 4208 17828 4214
rect 17776 4150 17828 4156
rect 17880 4049 17908 4422
rect 18064 4078 18092 4490
rect 18052 4072 18104 4078
rect 17866 4040 17922 4049
rect 18052 4014 18104 4020
rect 17866 3975 17922 3984
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17788 3641 17816 3878
rect 17774 3632 17830 3641
rect 17774 3567 17830 3576
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17604 3097 17632 3130
rect 17590 3088 17646 3097
rect 17590 3023 17646 3032
rect 17420 2944 17632 2972
rect 17316 2926 17368 2932
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15782 2204 16078 2224
rect 15838 2202 15862 2204
rect 15918 2202 15942 2204
rect 15998 2202 16022 2204
rect 15860 2150 15862 2202
rect 15924 2150 15936 2202
rect 15998 2150 16000 2202
rect 15838 2148 15862 2150
rect 15918 2148 15942 2150
rect 15998 2148 16022 2150
rect 15782 2128 16078 2148
rect 15672 1822 15792 1850
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 800
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15212 513 15240 1294
rect 15292 1284 15344 1290
rect 15292 1226 15344 1232
rect 15198 504 15254 513
rect 15198 439 15254 448
rect 15304 241 15332 1226
rect 15764 800 15792 1822
rect 16684 800 16712 2910
rect 17328 2650 17356 2926
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17512 2145 17540 2246
rect 17498 2136 17554 2145
rect 17498 2071 17554 2080
rect 17604 800 17632 2944
rect 17880 2553 17908 3878
rect 18156 3670 18184 7890
rect 18248 7410 18276 8978
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 6633 18276 7142
rect 18234 6624 18290 6633
rect 18234 6559 18290 6568
rect 18236 6112 18288 6118
rect 18236 6054 18288 6060
rect 18248 5953 18276 6054
rect 18234 5944 18290 5953
rect 18234 5879 18290 5888
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4321 18276 4966
rect 18234 4312 18290 4321
rect 18234 4247 18290 4256
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 2825 18092 3334
rect 18050 2816 18106 2825
rect 18050 2751 18106 2760
rect 18156 2650 18184 3470
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 17866 2544 17922 2553
rect 17866 2479 17922 2488
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17880 921 17908 2382
rect 18340 1737 18368 13806
rect 18432 11898 18460 16079
rect 18604 12708 18656 12714
rect 18604 12650 18656 12656
rect 18420 11892 18472 11898
rect 18420 11834 18472 11840
rect 18432 11354 18460 11834
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18432 10130 18460 10406
rect 18420 10124 18472 10130
rect 18420 10066 18472 10072
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9518 18460 9862
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 18432 9110 18460 9454
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18512 7540 18564 7546
rect 18512 7482 18564 7488
rect 18420 5568 18472 5574
rect 18418 5536 18420 5545
rect 18472 5536 18474 5545
rect 18418 5471 18474 5480
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 3233 18460 3334
rect 18418 3224 18474 3233
rect 18418 3159 18474 3168
rect 18326 1728 18382 1737
rect 18326 1663 18382 1672
rect 17866 912 17922 921
rect 17866 847 17922 856
rect 18524 800 18552 7482
rect 18616 1329 18644 12650
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18708 6934 18736 10202
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 18708 3534 18736 6870
rect 18800 4729 18828 8502
rect 18972 7064 19024 7070
rect 18970 7032 18972 7041
rect 19024 7032 19026 7041
rect 18970 6967 19026 6976
rect 18786 4720 18842 4729
rect 18786 4655 18842 4664
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 18602 1320 18658 1329
rect 18602 1255 18658 1264
rect 19444 800 19472 2858
rect 15290 232 15346 241
rect 15290 167 15346 176
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 4066 16904 4122 16960
rect 2962 16632 3018 16688
rect 1398 15544 1454 15600
rect 1674 15000 1730 15056
rect 1766 14356 1768 14376
rect 1768 14356 1820 14376
rect 1820 14356 1822 14376
rect 1766 14320 1822 14356
rect 2134 16224 2190 16280
rect 1490 13640 1546 13696
rect 2686 15952 2742 16008
rect 2318 13912 2374 13968
rect 1858 13252 1914 13288
rect 1858 13232 1860 13252
rect 1860 13232 1912 13252
rect 1912 13232 1914 13252
rect 2134 12960 2190 13016
rect 1674 11056 1730 11112
rect 1306 7112 1362 7168
rect 1122 5616 1178 5672
rect 1674 6704 1730 6760
rect 1582 6024 1638 6080
rect 1214 3576 1270 3632
rect 1582 4664 1638 4720
rect 1950 6180 2006 6216
rect 1950 6160 1952 6180
rect 1952 6160 2004 6180
rect 2004 6160 2006 6180
rect 1858 5072 1914 5128
rect 1858 4120 1914 4176
rect 1674 3712 1730 3768
rect 1582 2352 1638 2408
rect 2226 9696 2282 9752
rect 2134 9152 2190 9208
rect 2134 7656 2190 7712
rect 2226 5888 2282 5944
rect 2042 4684 2098 4720
rect 2042 4664 2044 4684
rect 2044 4664 2096 4684
rect 2096 4664 2098 4684
rect 2042 3032 2098 3088
rect 2226 4428 2228 4448
rect 2228 4428 2280 4448
rect 2280 4428 2282 4448
rect 2226 4392 2282 4428
rect 2870 15272 2926 15328
rect 2778 14592 2834 14648
rect 16486 16904 16542 16960
rect 15658 16496 15714 16552
rect 3921 14170 3977 14172
rect 4001 14170 4057 14172
rect 4081 14170 4137 14172
rect 4161 14170 4217 14172
rect 3921 14118 3947 14170
rect 3947 14118 3977 14170
rect 4001 14118 4011 14170
rect 4011 14118 4057 14170
rect 4081 14118 4127 14170
rect 4127 14118 4137 14170
rect 4161 14118 4191 14170
rect 4191 14118 4217 14170
rect 3921 14116 3977 14118
rect 4001 14116 4057 14118
rect 4081 14116 4137 14118
rect 4161 14116 4217 14118
rect 6886 14714 6942 14716
rect 6966 14714 7022 14716
rect 7046 14714 7102 14716
rect 7126 14714 7182 14716
rect 6886 14662 6912 14714
rect 6912 14662 6942 14714
rect 6966 14662 6976 14714
rect 6976 14662 7022 14714
rect 7046 14662 7092 14714
rect 7092 14662 7102 14714
rect 7126 14662 7156 14714
rect 7156 14662 7182 14714
rect 6886 14660 6942 14662
rect 6966 14660 7022 14662
rect 7046 14660 7102 14662
rect 7126 14660 7182 14662
rect 13450 15000 13506 15056
rect 12817 14714 12873 14716
rect 12897 14714 12953 14716
rect 12977 14714 13033 14716
rect 13057 14714 13113 14716
rect 12817 14662 12843 14714
rect 12843 14662 12873 14714
rect 12897 14662 12907 14714
rect 12907 14662 12953 14714
rect 12977 14662 13023 14714
rect 13023 14662 13033 14714
rect 13057 14662 13087 14714
rect 13087 14662 13113 14714
rect 12817 14660 12873 14662
rect 12897 14660 12953 14662
rect 12977 14660 13033 14662
rect 13057 14660 13113 14662
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9878 14170
rect 9878 14118 9908 14170
rect 9932 14118 9942 14170
rect 9942 14118 9988 14170
rect 10012 14118 10058 14170
rect 10058 14118 10068 14170
rect 10092 14118 10122 14170
rect 10122 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 3921 13082 3977 13084
rect 4001 13082 4057 13084
rect 4081 13082 4137 13084
rect 4161 13082 4217 13084
rect 3921 13030 3947 13082
rect 3947 13030 3977 13082
rect 4001 13030 4011 13082
rect 4011 13030 4057 13082
rect 4081 13030 4127 13082
rect 4127 13030 4137 13082
rect 4161 13030 4191 13082
rect 4191 13030 4217 13082
rect 3921 13028 3977 13030
rect 4001 13028 4057 13030
rect 4081 13028 4137 13030
rect 4161 13028 4217 13030
rect 3974 12708 4030 12744
rect 3974 12688 3976 12708
rect 3976 12688 4028 12708
rect 4028 12688 4030 12708
rect 3790 12280 3846 12336
rect 2870 9968 2926 10024
rect 2410 7384 2466 7440
rect 3514 12008 3570 12064
rect 3422 11600 3478 11656
rect 3330 11328 3386 11384
rect 3238 9560 3294 9616
rect 2870 7928 2926 7984
rect 2778 7384 2834 7440
rect 2686 6840 2742 6896
rect 2686 4528 2742 4584
rect 2962 6840 3018 6896
rect 3146 5888 3202 5944
rect 3921 11994 3977 11996
rect 4001 11994 4057 11996
rect 4081 11994 4137 11996
rect 4161 11994 4217 11996
rect 3921 11942 3947 11994
rect 3947 11942 3977 11994
rect 4001 11942 4011 11994
rect 4011 11942 4057 11994
rect 4081 11942 4127 11994
rect 4127 11942 4137 11994
rect 4161 11942 4191 11994
rect 4191 11942 4217 11994
rect 3921 11940 3977 11942
rect 4001 11940 4057 11942
rect 4081 11940 4137 11942
rect 4161 11940 4217 11942
rect 3422 10920 3478 10976
rect 3921 10906 3977 10908
rect 4001 10906 4057 10908
rect 4081 10906 4137 10908
rect 4161 10906 4217 10908
rect 3921 10854 3947 10906
rect 3947 10854 3977 10906
rect 4001 10854 4011 10906
rect 4011 10854 4057 10906
rect 4081 10854 4127 10906
rect 4127 10854 4137 10906
rect 4161 10854 4191 10906
rect 4191 10854 4217 10906
rect 3921 10852 3977 10854
rect 4001 10852 4057 10854
rect 4081 10852 4137 10854
rect 4161 10852 4217 10854
rect 4526 10648 4582 10704
rect 3921 9818 3977 9820
rect 4001 9818 4057 9820
rect 4081 9818 4137 9820
rect 4161 9818 4217 9820
rect 3921 9766 3947 9818
rect 3947 9766 3977 9818
rect 4001 9766 4011 9818
rect 4011 9766 4057 9818
rect 4081 9766 4127 9818
rect 4127 9766 4137 9818
rect 4161 9766 4191 9818
rect 4191 9766 4217 9818
rect 3921 9764 3977 9766
rect 4001 9764 4057 9766
rect 4081 9764 4137 9766
rect 4161 9764 4217 9766
rect 3514 9560 3570 9616
rect 3422 9052 3424 9072
rect 3424 9052 3476 9072
rect 3476 9052 3478 9072
rect 3422 9016 3478 9052
rect 3330 8200 3386 8256
rect 3238 5752 3294 5808
rect 4434 10004 4436 10024
rect 4436 10004 4488 10024
rect 4488 10004 4490 10024
rect 4434 9968 4490 10004
rect 3606 8064 3662 8120
rect 4250 9288 4306 9344
rect 3921 8730 3977 8732
rect 4001 8730 4057 8732
rect 4081 8730 4137 8732
rect 4161 8730 4217 8732
rect 3921 8678 3947 8730
rect 3947 8678 3977 8730
rect 4001 8678 4011 8730
rect 4011 8678 4057 8730
rect 4081 8678 4127 8730
rect 4127 8678 4137 8730
rect 4161 8678 4191 8730
rect 4191 8678 4217 8730
rect 3921 8676 3977 8678
rect 4001 8676 4057 8678
rect 4081 8676 4137 8678
rect 4161 8676 4217 8678
rect 3882 8200 3938 8256
rect 3921 7642 3977 7644
rect 4001 7642 4057 7644
rect 4081 7642 4137 7644
rect 4161 7642 4217 7644
rect 3921 7590 3947 7642
rect 3947 7590 3977 7642
rect 4001 7590 4011 7642
rect 4011 7590 4057 7642
rect 4081 7590 4127 7642
rect 4127 7590 4137 7642
rect 4161 7590 4191 7642
rect 4191 7590 4217 7642
rect 3921 7588 3977 7590
rect 4001 7588 4057 7590
rect 4081 7588 4137 7590
rect 4161 7588 4217 7590
rect 4618 9560 4674 9616
rect 4802 9424 4858 9480
rect 4710 9288 4766 9344
rect 4526 7928 4582 7984
rect 3698 6976 3754 7032
rect 4158 6976 4214 7032
rect 3698 6452 3754 6488
rect 3698 6432 3700 6452
rect 3700 6432 3752 6452
rect 3752 6432 3754 6452
rect 2410 3440 2466 3496
rect 2134 2624 2190 2680
rect 1766 2080 1822 2136
rect 2502 2508 2558 2544
rect 2502 2488 2504 2508
rect 2504 2488 2556 2508
rect 2556 2488 2558 2508
rect 2318 1808 2374 1864
rect 2778 3052 2834 3088
rect 2778 3032 2780 3052
rect 2780 3032 2832 3052
rect 2832 3032 2834 3052
rect 3514 5788 3516 5808
rect 3516 5788 3568 5808
rect 3568 5788 3570 5808
rect 3514 5752 3570 5788
rect 3921 6554 3977 6556
rect 4001 6554 4057 6556
rect 4081 6554 4137 6556
rect 4161 6554 4217 6556
rect 3921 6502 3947 6554
rect 3947 6502 3977 6554
rect 4001 6502 4011 6554
rect 4011 6502 4057 6554
rect 4081 6502 4127 6554
rect 4127 6502 4137 6554
rect 4161 6502 4191 6554
rect 4191 6502 4217 6554
rect 3921 6500 3977 6502
rect 4001 6500 4057 6502
rect 4081 6500 4137 6502
rect 4161 6500 4217 6502
rect 3606 4120 3662 4176
rect 3422 3984 3478 4040
rect 3921 5466 3977 5468
rect 4001 5466 4057 5468
rect 4081 5466 4137 5468
rect 4161 5466 4217 5468
rect 3921 5414 3947 5466
rect 3947 5414 3977 5466
rect 4001 5414 4011 5466
rect 4011 5414 4057 5466
rect 4081 5414 4127 5466
rect 4127 5414 4137 5466
rect 4161 5414 4191 5466
rect 4191 5414 4217 5466
rect 3921 5412 3977 5414
rect 4001 5412 4057 5414
rect 4081 5412 4137 5414
rect 4161 5412 4217 5414
rect 4066 5108 4068 5128
rect 4068 5108 4120 5128
rect 4120 5108 4122 5128
rect 4066 5072 4122 5108
rect 4434 5244 4436 5264
rect 4436 5244 4488 5264
rect 4488 5244 4490 5264
rect 4434 5208 4490 5244
rect 4434 4428 4436 4448
rect 4436 4428 4488 4448
rect 4488 4428 4490 4448
rect 3921 4378 3977 4380
rect 4001 4378 4057 4380
rect 4081 4378 4137 4380
rect 4161 4378 4217 4380
rect 3921 4326 3947 4378
rect 3947 4326 3977 4378
rect 4001 4326 4011 4378
rect 4011 4326 4057 4378
rect 4081 4326 4127 4378
rect 4127 4326 4137 4378
rect 4161 4326 4191 4378
rect 4191 4326 4217 4378
rect 3921 4324 3977 4326
rect 4001 4324 4057 4326
rect 4081 4324 4137 4326
rect 4161 4324 4217 4326
rect 4434 4392 4490 4428
rect 3054 2932 3056 2952
rect 3056 2932 3108 2952
rect 3108 2932 3110 2952
rect 3054 2896 3110 2932
rect 1674 720 1730 776
rect 2686 448 2742 504
rect 3054 1128 3110 1184
rect 3921 3290 3977 3292
rect 4001 3290 4057 3292
rect 4081 3290 4137 3292
rect 4161 3290 4217 3292
rect 3921 3238 3947 3290
rect 3947 3238 3977 3290
rect 4001 3238 4011 3290
rect 4011 3238 4057 3290
rect 4081 3238 4127 3290
rect 4127 3238 4137 3290
rect 4161 3238 4191 3290
rect 4191 3238 4217 3290
rect 3921 3236 3977 3238
rect 4001 3236 4057 3238
rect 4081 3236 4137 3238
rect 4161 3236 4217 3238
rect 3514 2488 3570 2544
rect 4066 2796 4068 2816
rect 4068 2796 4120 2816
rect 4120 2796 4122 2816
rect 4066 2760 4122 2796
rect 4526 2760 4582 2816
rect 5538 10376 5594 10432
rect 5354 9988 5410 10024
rect 5354 9968 5356 9988
rect 5356 9968 5408 9988
rect 5408 9968 5410 9988
rect 5262 9560 5318 9616
rect 4894 7792 4950 7848
rect 4894 7148 4896 7168
rect 4896 7148 4948 7168
rect 4948 7148 4950 7168
rect 4894 7112 4950 7148
rect 5170 7248 5226 7304
rect 5446 7520 5502 7576
rect 5814 8336 5870 8392
rect 5630 7248 5686 7304
rect 6886 13626 6942 13628
rect 6966 13626 7022 13628
rect 7046 13626 7102 13628
rect 7126 13626 7182 13628
rect 6886 13574 6912 13626
rect 6912 13574 6942 13626
rect 6966 13574 6976 13626
rect 6976 13574 7022 13626
rect 7046 13574 7092 13626
rect 7092 13574 7102 13626
rect 7126 13574 7156 13626
rect 7156 13574 7182 13626
rect 6886 13572 6942 13574
rect 6966 13572 7022 13574
rect 7046 13572 7102 13574
rect 7126 13572 7182 13574
rect 12162 13776 12218 13832
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9878 13082
rect 9878 13030 9908 13082
rect 9932 13030 9942 13082
rect 9942 13030 9988 13082
rect 10012 13030 10058 13082
rect 10058 13030 10068 13082
rect 10092 13030 10122 13082
rect 10122 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 6886 12538 6942 12540
rect 6966 12538 7022 12540
rect 7046 12538 7102 12540
rect 7126 12538 7182 12540
rect 6886 12486 6912 12538
rect 6912 12486 6942 12538
rect 6966 12486 6976 12538
rect 6976 12486 7022 12538
rect 7046 12486 7092 12538
rect 7092 12486 7102 12538
rect 7126 12486 7156 12538
rect 7156 12486 7182 12538
rect 6886 12484 6942 12486
rect 6966 12484 7022 12486
rect 7046 12484 7102 12486
rect 7126 12484 7182 12486
rect 6886 11450 6942 11452
rect 6966 11450 7022 11452
rect 7046 11450 7102 11452
rect 7126 11450 7182 11452
rect 6886 11398 6912 11450
rect 6912 11398 6942 11450
rect 6966 11398 6976 11450
rect 6976 11398 7022 11450
rect 7046 11398 7092 11450
rect 7092 11398 7102 11450
rect 7126 11398 7156 11450
rect 7156 11398 7182 11450
rect 6886 11396 6942 11398
rect 6966 11396 7022 11398
rect 7046 11396 7102 11398
rect 7126 11396 7182 11398
rect 6182 9152 6238 9208
rect 6886 10362 6942 10364
rect 6966 10362 7022 10364
rect 7046 10362 7102 10364
rect 7126 10362 7182 10364
rect 6886 10310 6912 10362
rect 6912 10310 6942 10362
rect 6966 10310 6976 10362
rect 6976 10310 7022 10362
rect 7046 10310 7092 10362
rect 7092 10310 7102 10362
rect 7126 10310 7156 10362
rect 7156 10310 7182 10362
rect 6886 10308 6942 10310
rect 6966 10308 7022 10310
rect 7046 10308 7102 10310
rect 7126 10308 7182 10310
rect 6886 9274 6942 9276
rect 6966 9274 7022 9276
rect 7046 9274 7102 9276
rect 7126 9274 7182 9276
rect 6886 9222 6912 9274
rect 6912 9222 6942 9274
rect 6966 9222 6976 9274
rect 6976 9222 7022 9274
rect 7046 9222 7092 9274
rect 7092 9222 7102 9274
rect 7126 9222 7156 9274
rect 7156 9222 7182 9274
rect 6886 9220 6942 9222
rect 6966 9220 7022 9222
rect 7046 9220 7102 9222
rect 7126 9220 7182 9222
rect 7562 8880 7618 8936
rect 6366 8356 6422 8392
rect 6366 8336 6368 8356
rect 6368 8336 6420 8356
rect 6420 8336 6422 8356
rect 6886 8186 6942 8188
rect 6966 8186 7022 8188
rect 7046 8186 7102 8188
rect 7126 8186 7182 8188
rect 6886 8134 6912 8186
rect 6912 8134 6942 8186
rect 6966 8134 6976 8186
rect 6976 8134 7022 8186
rect 7046 8134 7092 8186
rect 7092 8134 7102 8186
rect 7126 8134 7156 8186
rect 7156 8134 7182 8186
rect 6886 8132 6942 8134
rect 6966 8132 7022 8134
rect 7046 8132 7102 8134
rect 7126 8132 7182 8134
rect 6550 7792 6606 7848
rect 7378 7112 7434 7168
rect 6886 7098 6942 7100
rect 6966 7098 7022 7100
rect 7046 7098 7102 7100
rect 7126 7098 7182 7100
rect 6886 7046 6912 7098
rect 6912 7046 6942 7098
rect 6966 7046 6976 7098
rect 6976 7046 7022 7098
rect 7046 7046 7092 7098
rect 7092 7046 7102 7098
rect 7126 7046 7156 7098
rect 7156 7046 7182 7098
rect 6886 7044 6942 7046
rect 6966 7044 7022 7046
rect 7046 7044 7102 7046
rect 7126 7044 7182 7046
rect 6366 4684 6422 4720
rect 6366 4664 6368 4684
rect 6368 4664 6420 4684
rect 6420 4664 6422 4684
rect 5998 3440 6054 3496
rect 5354 2760 5410 2816
rect 5446 2624 5502 2680
rect 3921 2202 3977 2204
rect 4001 2202 4057 2204
rect 4081 2202 4137 2204
rect 4161 2202 4217 2204
rect 3921 2150 3947 2202
rect 3947 2150 3977 2202
rect 4001 2150 4011 2202
rect 4011 2150 4057 2202
rect 4081 2150 4127 2202
rect 4127 2150 4137 2202
rect 4161 2150 4191 2202
rect 4191 2150 4217 2202
rect 3921 2148 3977 2150
rect 4001 2148 4057 2150
rect 4081 2148 4137 2150
rect 4161 2148 4217 2150
rect 3698 1400 3754 1456
rect 6886 6010 6942 6012
rect 6966 6010 7022 6012
rect 7046 6010 7102 6012
rect 7126 6010 7182 6012
rect 6886 5958 6912 6010
rect 6912 5958 6942 6010
rect 6966 5958 6976 6010
rect 6976 5958 7022 6010
rect 7046 5958 7092 6010
rect 7092 5958 7102 6010
rect 7126 5958 7156 6010
rect 7156 5958 7182 6010
rect 6886 5956 6942 5958
rect 6966 5956 7022 5958
rect 7046 5956 7102 5958
rect 7126 5956 7182 5958
rect 6886 4922 6942 4924
rect 6966 4922 7022 4924
rect 7046 4922 7102 4924
rect 7126 4922 7182 4924
rect 6886 4870 6912 4922
rect 6912 4870 6942 4922
rect 6966 4870 6976 4922
rect 6976 4870 7022 4922
rect 7046 4870 7092 4922
rect 7092 4870 7102 4922
rect 7126 4870 7156 4922
rect 7156 4870 7182 4922
rect 6886 4868 6942 4870
rect 6966 4868 7022 4870
rect 7046 4868 7102 4870
rect 7126 4868 7182 4870
rect 6550 4120 6606 4176
rect 6886 3834 6942 3836
rect 6966 3834 7022 3836
rect 7046 3834 7102 3836
rect 7126 3834 7182 3836
rect 6886 3782 6912 3834
rect 6912 3782 6942 3834
rect 6966 3782 6976 3834
rect 6976 3782 7022 3834
rect 7046 3782 7092 3834
rect 7092 3782 7102 3834
rect 7126 3782 7156 3834
rect 7156 3782 7182 3834
rect 6886 3780 6942 3782
rect 6966 3780 7022 3782
rect 7046 3780 7102 3782
rect 7126 3780 7182 3782
rect 7010 3032 7066 3088
rect 6886 2746 6942 2748
rect 6966 2746 7022 2748
rect 7046 2746 7102 2748
rect 7126 2746 7182 2748
rect 6886 2694 6912 2746
rect 6912 2694 6942 2746
rect 6966 2694 6976 2746
rect 6976 2694 7022 2746
rect 7046 2694 7092 2746
rect 7092 2694 7102 2746
rect 7126 2694 7156 2746
rect 7156 2694 7182 2746
rect 6886 2692 6942 2694
rect 6966 2692 7022 2694
rect 7046 2692 7102 2694
rect 7126 2692 7182 2694
rect 7378 2760 7434 2816
rect 8022 11056 8078 11112
rect 8298 11076 8354 11112
rect 8298 11056 8300 11076
rect 8300 11056 8352 11076
rect 8352 11056 8354 11076
rect 8942 11092 8944 11112
rect 8944 11092 8996 11112
rect 8996 11092 8998 11112
rect 8942 11056 8998 11092
rect 8574 10784 8630 10840
rect 8482 10648 8538 10704
rect 9310 10004 9312 10024
rect 9312 10004 9364 10024
rect 9364 10004 9366 10024
rect 9310 9968 9366 10004
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9878 11994
rect 9878 11942 9908 11994
rect 9932 11942 9942 11994
rect 9942 11942 9988 11994
rect 10012 11942 10058 11994
rect 10058 11942 10068 11994
rect 10092 11942 10122 11994
rect 10122 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10046 11620 10102 11656
rect 10046 11600 10048 11620
rect 10048 11600 10100 11620
rect 10100 11600 10102 11620
rect 9770 11056 9826 11112
rect 8390 7248 8446 7304
rect 7838 6160 7894 6216
rect 7838 5652 7840 5672
rect 7840 5652 7892 5672
rect 7892 5652 7894 5672
rect 7838 5616 7894 5652
rect 7562 4392 7618 4448
rect 8574 3848 8630 3904
rect 8666 3732 8722 3768
rect 8666 3712 8668 3732
rect 8668 3712 8720 3732
rect 8720 3712 8722 3732
rect 9402 8880 9458 8936
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9878 10906
rect 9878 10854 9908 10906
rect 9932 10854 9942 10906
rect 9942 10854 9988 10906
rect 10012 10854 10058 10906
rect 10058 10854 10068 10906
rect 10092 10854 10122 10906
rect 10122 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9954 10104 10010 10160
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9878 9818
rect 9878 9766 9908 9818
rect 9932 9766 9942 9818
rect 9942 9766 9988 9818
rect 10012 9766 10058 9818
rect 10058 9766 10068 9818
rect 10092 9766 10122 9818
rect 10122 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10322 9580 10378 9616
rect 10322 9560 10324 9580
rect 10324 9560 10376 9580
rect 10376 9560 10378 9580
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9878 8730
rect 9878 8678 9908 8730
rect 9932 8678 9942 8730
rect 9942 8678 9988 8730
rect 10012 8678 10058 8730
rect 10058 8678 10068 8730
rect 10092 8678 10122 8730
rect 10122 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 11058 12144 11114 12200
rect 10782 11756 10838 11792
rect 10782 11736 10784 11756
rect 10784 11736 10836 11756
rect 10836 11736 10838 11756
rect 11978 11736 12034 11792
rect 10874 11192 10930 11248
rect 9586 8200 9642 8256
rect 9126 5072 9182 5128
rect 7654 3032 7710 3088
rect 9862 7928 9918 7984
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9878 7642
rect 9878 7590 9908 7642
rect 9932 7590 9942 7642
rect 9942 7590 9988 7642
rect 10012 7590 10058 7642
rect 10058 7590 10068 7642
rect 10092 7590 10122 7642
rect 10122 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 11058 10512 11114 10568
rect 11150 10104 11206 10160
rect 11058 9968 11114 10024
rect 11150 9832 11206 9888
rect 10598 8744 10654 8800
rect 10506 7520 10562 7576
rect 10414 6976 10470 7032
rect 10322 6840 10378 6896
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9878 6554
rect 9878 6502 9908 6554
rect 9932 6502 9942 6554
rect 9942 6502 9988 6554
rect 10012 6502 10058 6554
rect 10058 6502 10068 6554
rect 10092 6502 10122 6554
rect 10122 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10690 7384 10746 7440
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9878 5466
rect 9878 5414 9908 5466
rect 9932 5414 9942 5466
rect 9942 5414 9988 5466
rect 10012 5414 10058 5466
rect 10058 5414 10068 5466
rect 10092 5414 10122 5466
rect 10122 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10414 5788 10416 5808
rect 10416 5788 10468 5808
rect 10468 5788 10470 5808
rect 10414 5752 10470 5788
rect 10230 4428 10232 4448
rect 10232 4428 10284 4448
rect 10284 4428 10286 4448
rect 10230 4392 10286 4428
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9878 4378
rect 9878 4326 9908 4378
rect 9932 4326 9942 4378
rect 9942 4326 9988 4378
rect 10012 4326 10058 4378
rect 10058 4326 10068 4378
rect 10092 4326 10122 4378
rect 10122 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9878 3290
rect 9878 3238 9908 3290
rect 9932 3238 9942 3290
rect 9942 3238 9988 3290
rect 10012 3238 10058 3290
rect 10058 3238 10068 3290
rect 10092 3238 10122 3290
rect 10122 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 9678 2488 9734 2544
rect 10138 2352 10194 2408
rect 10506 3168 10562 3224
rect 10782 6976 10838 7032
rect 10506 2896 10562 2952
rect 10966 6296 11022 6352
rect 11702 11600 11758 11656
rect 11058 4528 11114 4584
rect 10966 2932 10968 2952
rect 10968 2932 11020 2952
rect 11020 2932 11022 2952
rect 10966 2896 11022 2932
rect 11610 8880 11666 8936
rect 11518 8744 11574 8800
rect 11518 6196 11520 6216
rect 11520 6196 11572 6216
rect 11572 6196 11574 6216
rect 11518 6160 11574 6196
rect 11518 5208 11574 5264
rect 11334 3848 11390 3904
rect 11610 3884 11612 3904
rect 11612 3884 11664 3904
rect 11664 3884 11666 3904
rect 11610 3848 11666 3884
rect 12817 13626 12873 13628
rect 12897 13626 12953 13628
rect 12977 13626 13033 13628
rect 13057 13626 13113 13628
rect 12817 13574 12843 13626
rect 12843 13574 12873 13626
rect 12897 13574 12907 13626
rect 12907 13574 12953 13626
rect 12977 13574 13023 13626
rect 13023 13574 13033 13626
rect 13057 13574 13087 13626
rect 13087 13574 13113 13626
rect 12817 13572 12873 13574
rect 12897 13572 12953 13574
rect 12977 13572 13033 13574
rect 13057 13572 13113 13574
rect 12817 12538 12873 12540
rect 12897 12538 12953 12540
rect 12977 12538 13033 12540
rect 13057 12538 13113 12540
rect 12817 12486 12843 12538
rect 12843 12486 12873 12538
rect 12897 12486 12907 12538
rect 12907 12486 12953 12538
rect 12977 12486 13023 12538
rect 13023 12486 13033 12538
rect 13057 12486 13087 12538
rect 13087 12486 13113 12538
rect 12817 12484 12873 12486
rect 12897 12484 12953 12486
rect 12977 12484 13033 12486
rect 13057 12484 13113 12486
rect 12162 11736 12218 11792
rect 12817 11450 12873 11452
rect 12897 11450 12953 11452
rect 12977 11450 13033 11452
rect 13057 11450 13113 11452
rect 12817 11398 12843 11450
rect 12843 11398 12873 11450
rect 12897 11398 12907 11450
rect 12907 11398 12953 11450
rect 12977 11398 13023 11450
rect 13023 11398 13033 11450
rect 13057 11398 13087 11450
rect 13087 11398 13113 11450
rect 12817 11396 12873 11398
rect 12897 11396 12953 11398
rect 12977 11396 13033 11398
rect 13057 11396 13113 11398
rect 12162 11192 12218 11248
rect 12070 11076 12126 11112
rect 12070 11056 12072 11076
rect 12072 11056 12124 11076
rect 12124 11056 12126 11076
rect 12254 11056 12310 11112
rect 11794 8084 11850 8120
rect 11794 8064 11796 8084
rect 11796 8064 11848 8084
rect 11848 8064 11850 8084
rect 11886 7948 11942 7984
rect 11886 7928 11888 7948
rect 11888 7928 11940 7948
rect 11940 7928 11942 7948
rect 12254 8880 12310 8936
rect 12254 8236 12256 8256
rect 12256 8236 12308 8256
rect 12308 8236 12310 8256
rect 12254 8200 12310 8236
rect 12438 11056 12494 11112
rect 12530 9832 12586 9888
rect 12346 8064 12402 8120
rect 12070 7384 12126 7440
rect 11702 3032 11758 3088
rect 11518 2760 11574 2816
rect 12530 8608 12586 8664
rect 12438 6704 12494 6760
rect 12346 6432 12402 6488
rect 12254 6196 12256 6216
rect 12256 6196 12308 6216
rect 12308 6196 12310 6216
rect 12254 6160 12310 6196
rect 12254 5516 12256 5536
rect 12256 5516 12308 5536
rect 12308 5516 12310 5536
rect 12254 5480 12310 5516
rect 12162 5344 12218 5400
rect 12817 10362 12873 10364
rect 12897 10362 12953 10364
rect 12977 10362 13033 10364
rect 13057 10362 13113 10364
rect 12817 10310 12843 10362
rect 12843 10310 12873 10362
rect 12897 10310 12907 10362
rect 12907 10310 12953 10362
rect 12977 10310 13023 10362
rect 13023 10310 13033 10362
rect 13057 10310 13087 10362
rect 13087 10310 13113 10362
rect 12817 10308 12873 10310
rect 12897 10308 12953 10310
rect 12977 10308 13033 10310
rect 13057 10308 13113 10310
rect 12817 9274 12873 9276
rect 12897 9274 12953 9276
rect 12977 9274 13033 9276
rect 13057 9274 13113 9276
rect 12817 9222 12843 9274
rect 12843 9222 12873 9274
rect 12897 9222 12907 9274
rect 12907 9222 12953 9274
rect 12977 9222 13023 9274
rect 13023 9222 13033 9274
rect 13057 9222 13087 9274
rect 13087 9222 13113 9274
rect 12817 9220 12873 9222
rect 12897 9220 12953 9222
rect 12977 9220 13033 9222
rect 13057 9220 13113 9222
rect 13082 8472 13138 8528
rect 12817 8186 12873 8188
rect 12897 8186 12953 8188
rect 12977 8186 13033 8188
rect 13057 8186 13113 8188
rect 12817 8134 12843 8186
rect 12843 8134 12873 8186
rect 12897 8134 12907 8186
rect 12907 8134 12953 8186
rect 12977 8134 13023 8186
rect 13023 8134 13033 8186
rect 13057 8134 13087 8186
rect 13087 8134 13113 8186
rect 12817 8132 12873 8134
rect 12897 8132 12953 8134
rect 12977 8132 13033 8134
rect 13057 8132 13113 8134
rect 12817 7098 12873 7100
rect 12897 7098 12953 7100
rect 12977 7098 13033 7100
rect 13057 7098 13113 7100
rect 12817 7046 12843 7098
rect 12843 7046 12873 7098
rect 12897 7046 12907 7098
rect 12907 7046 12953 7098
rect 12977 7046 13023 7098
rect 13023 7046 13033 7098
rect 13057 7046 13087 7098
rect 13087 7046 13113 7098
rect 12817 7044 12873 7046
rect 12897 7044 12953 7046
rect 12977 7044 13033 7046
rect 13057 7044 13113 7046
rect 12806 6296 12862 6352
rect 12817 6010 12873 6012
rect 12897 6010 12953 6012
rect 12977 6010 13033 6012
rect 13057 6010 13113 6012
rect 12817 5958 12843 6010
rect 12843 5958 12873 6010
rect 12897 5958 12907 6010
rect 12907 5958 12953 6010
rect 12977 5958 13023 6010
rect 13023 5958 13033 6010
rect 13057 5958 13087 6010
rect 13087 5958 13113 6010
rect 12817 5956 12873 5958
rect 12897 5956 12953 5958
rect 12977 5956 13033 5958
rect 13057 5956 13113 5958
rect 12438 5208 12494 5264
rect 12438 4120 12494 4176
rect 12438 3712 12494 3768
rect 12346 3168 12402 3224
rect 15014 15680 15070 15736
rect 13634 8744 13690 8800
rect 13542 7928 13598 7984
rect 13726 8608 13782 8664
rect 13634 6704 13690 6760
rect 12817 4922 12873 4924
rect 12897 4922 12953 4924
rect 12977 4922 13033 4924
rect 13057 4922 13113 4924
rect 12817 4870 12843 4922
rect 12843 4870 12873 4922
rect 12897 4870 12907 4922
rect 12907 4870 12953 4922
rect 12977 4870 13023 4922
rect 13023 4870 13033 4922
rect 13057 4870 13087 4922
rect 13087 4870 13113 4922
rect 12817 4868 12873 4870
rect 12897 4868 12953 4870
rect 12977 4868 13033 4870
rect 13057 4868 13113 4870
rect 13358 5752 13414 5808
rect 13542 5888 13598 5944
rect 13542 5616 13598 5672
rect 13726 5344 13782 5400
rect 13634 4664 13690 4720
rect 12817 3834 12873 3836
rect 12897 3834 12953 3836
rect 12977 3834 13033 3836
rect 13057 3834 13113 3836
rect 12817 3782 12843 3834
rect 12843 3782 12873 3834
rect 12897 3782 12907 3834
rect 12907 3782 12953 3834
rect 12977 3782 13023 3834
rect 13023 3782 13033 3834
rect 13057 3782 13087 3834
rect 13087 3782 13113 3834
rect 12817 3780 12873 3782
rect 12897 3780 12953 3782
rect 12977 3780 13033 3782
rect 13057 3780 13113 3782
rect 10414 2252 10416 2272
rect 10416 2252 10468 2272
rect 10468 2252 10470 2272
rect 10414 2216 10470 2252
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9878 2202
rect 9878 2150 9908 2202
rect 9932 2150 9942 2202
rect 9942 2150 9988 2202
rect 10012 2150 10058 2202
rect 10058 2150 10068 2202
rect 10092 2150 10122 2202
rect 10122 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 12622 2896 12678 2952
rect 12817 2746 12873 2748
rect 12897 2746 12953 2748
rect 12977 2746 13033 2748
rect 13057 2746 13113 2748
rect 12817 2694 12843 2746
rect 12843 2694 12873 2746
rect 12897 2694 12907 2746
rect 12907 2694 12953 2746
rect 12977 2694 13023 2746
rect 13023 2694 13033 2746
rect 13057 2694 13087 2746
rect 13087 2694 13113 2746
rect 12817 2692 12873 2694
rect 12897 2692 12953 2694
rect 12977 2692 13033 2694
rect 13057 2692 13113 2694
rect 13174 2216 13230 2272
rect 13910 6740 13912 6760
rect 13912 6740 13964 6760
rect 13964 6740 13966 6760
rect 13910 6704 13966 6740
rect 13910 6432 13966 6488
rect 13818 4528 13874 4584
rect 14094 9424 14150 9480
rect 14278 8880 14334 8936
rect 14646 11600 14702 11656
rect 14278 5652 14280 5672
rect 14280 5652 14332 5672
rect 14332 5652 14334 5672
rect 14278 5616 14334 5652
rect 14186 5208 14242 5264
rect 15474 15408 15530 15464
rect 15198 14592 15254 14648
rect 14738 7520 14794 7576
rect 14830 7248 14886 7304
rect 15014 9868 15016 9888
rect 15016 9868 15068 9888
rect 15068 9868 15070 9888
rect 15014 9832 15070 9868
rect 15014 6704 15070 6760
rect 14646 4392 14702 4448
rect 14094 2488 14150 2544
rect 14922 5480 14978 5536
rect 14738 3168 14794 3224
rect 15566 11192 15622 11248
rect 16210 14184 16266 14240
rect 15782 14170 15838 14172
rect 15862 14170 15918 14172
rect 15942 14170 15998 14172
rect 16022 14170 16078 14172
rect 15782 14118 15808 14170
rect 15808 14118 15838 14170
rect 15862 14118 15872 14170
rect 15872 14118 15918 14170
rect 15942 14118 15988 14170
rect 15988 14118 15998 14170
rect 16022 14118 16052 14170
rect 16052 14118 16078 14170
rect 15782 14116 15838 14118
rect 15862 14116 15918 14118
rect 15942 14116 15998 14118
rect 16022 14116 16078 14118
rect 15782 13082 15838 13084
rect 15862 13082 15918 13084
rect 15942 13082 15998 13084
rect 16022 13082 16078 13084
rect 15782 13030 15808 13082
rect 15808 13030 15838 13082
rect 15862 13030 15872 13082
rect 15872 13030 15918 13082
rect 15942 13030 15988 13082
rect 15988 13030 15998 13082
rect 16022 13030 16052 13082
rect 16052 13030 16078 13082
rect 15782 13028 15838 13030
rect 15862 13028 15918 13030
rect 15942 13028 15998 13030
rect 16022 13028 16078 13030
rect 15750 12688 15806 12744
rect 15750 12280 15806 12336
rect 15782 11994 15838 11996
rect 15862 11994 15918 11996
rect 15942 11994 15998 11996
rect 16022 11994 16078 11996
rect 15782 11942 15808 11994
rect 15808 11942 15838 11994
rect 15862 11942 15872 11994
rect 15872 11942 15918 11994
rect 15942 11942 15988 11994
rect 15988 11942 15998 11994
rect 16022 11942 16052 11994
rect 16052 11942 16078 11994
rect 15782 11940 15838 11942
rect 15862 11940 15918 11942
rect 15942 11940 15998 11942
rect 16022 11940 16078 11942
rect 16394 13504 16450 13560
rect 16302 11872 16358 11928
rect 15198 3032 15254 3088
rect 15782 10906 15838 10908
rect 15862 10906 15918 10908
rect 15942 10906 15998 10908
rect 16022 10906 16078 10908
rect 15782 10854 15808 10906
rect 15808 10854 15838 10906
rect 15862 10854 15872 10906
rect 15872 10854 15918 10906
rect 15942 10854 15988 10906
rect 15988 10854 15998 10906
rect 16022 10854 16052 10906
rect 16052 10854 16078 10906
rect 15782 10852 15838 10854
rect 15862 10852 15918 10854
rect 15942 10852 15998 10854
rect 16022 10852 16078 10854
rect 15782 9818 15838 9820
rect 15862 9818 15918 9820
rect 15942 9818 15998 9820
rect 16022 9818 16078 9820
rect 15782 9766 15808 9818
rect 15808 9766 15838 9818
rect 15862 9766 15872 9818
rect 15872 9766 15918 9818
rect 15942 9766 15988 9818
rect 15988 9766 15998 9818
rect 16022 9766 16052 9818
rect 16052 9766 16078 9818
rect 15782 9764 15838 9766
rect 15862 9764 15918 9766
rect 15942 9764 15998 9766
rect 16022 9764 16078 9766
rect 16118 8880 16174 8936
rect 15782 8730 15838 8732
rect 15862 8730 15918 8732
rect 15942 8730 15998 8732
rect 16022 8730 16078 8732
rect 15782 8678 15808 8730
rect 15808 8678 15838 8730
rect 15862 8678 15872 8730
rect 15872 8678 15918 8730
rect 15942 8678 15988 8730
rect 15988 8678 15998 8730
rect 16022 8678 16052 8730
rect 16052 8678 16078 8730
rect 15782 8676 15838 8678
rect 15862 8676 15918 8678
rect 15942 8676 15998 8678
rect 16022 8676 16078 8678
rect 16302 8336 16358 8392
rect 18418 16088 18474 16144
rect 16486 9968 16542 10024
rect 16854 9560 16910 9616
rect 15782 7642 15838 7644
rect 15862 7642 15918 7644
rect 15942 7642 15998 7644
rect 16022 7642 16078 7644
rect 15782 7590 15808 7642
rect 15808 7590 15838 7642
rect 15862 7590 15872 7642
rect 15872 7590 15918 7642
rect 15942 7590 15988 7642
rect 15988 7590 15998 7642
rect 16022 7590 16052 7642
rect 16052 7590 16078 7642
rect 15782 7588 15838 7590
rect 15862 7588 15918 7590
rect 15942 7588 15998 7590
rect 16022 7588 16078 7590
rect 15782 6554 15838 6556
rect 15862 6554 15918 6556
rect 15942 6554 15998 6556
rect 16022 6554 16078 6556
rect 15782 6502 15808 6554
rect 15808 6502 15838 6554
rect 15862 6502 15872 6554
rect 15872 6502 15918 6554
rect 15942 6502 15988 6554
rect 15988 6502 15998 6554
rect 16022 6502 16052 6554
rect 16052 6502 16078 6554
rect 15782 6500 15838 6502
rect 15862 6500 15918 6502
rect 15942 6500 15998 6502
rect 16022 6500 16078 6502
rect 16486 7792 16542 7848
rect 17038 9696 17094 9752
rect 17130 9016 17186 9072
rect 16946 6840 17002 6896
rect 15782 5466 15838 5468
rect 15862 5466 15918 5468
rect 15942 5466 15998 5468
rect 16022 5466 16078 5468
rect 15782 5414 15808 5466
rect 15808 5414 15838 5466
rect 15862 5414 15872 5466
rect 15872 5414 15918 5466
rect 15942 5414 15988 5466
rect 15988 5414 15998 5466
rect 16022 5414 16052 5466
rect 16052 5414 16078 5466
rect 15782 5412 15838 5414
rect 15862 5412 15918 5414
rect 15942 5412 15998 5414
rect 16022 5412 16078 5414
rect 15382 3052 15438 3088
rect 15382 3032 15384 3052
rect 15384 3032 15436 3052
rect 15436 3032 15438 3052
rect 15782 4378 15838 4380
rect 15862 4378 15918 4380
rect 15942 4378 15998 4380
rect 16022 4378 16078 4380
rect 15782 4326 15808 4378
rect 15808 4326 15838 4378
rect 15862 4326 15872 4378
rect 15872 4326 15918 4378
rect 15942 4326 15988 4378
rect 15988 4326 15998 4378
rect 16022 4326 16052 4378
rect 16052 4326 16078 4378
rect 15782 4324 15838 4326
rect 15862 4324 15918 4326
rect 15942 4324 15998 4326
rect 16022 4324 16078 4326
rect 15382 2352 15438 2408
rect 15782 3290 15838 3292
rect 15862 3290 15918 3292
rect 15942 3290 15998 3292
rect 16022 3290 16078 3292
rect 15782 3238 15808 3290
rect 15808 3238 15838 3290
rect 15862 3238 15872 3290
rect 15872 3238 15918 3290
rect 15942 3238 15988 3290
rect 15988 3238 15998 3290
rect 16022 3238 16052 3290
rect 16052 3238 16078 3290
rect 15782 3236 15838 3238
rect 15862 3236 15918 3238
rect 15942 3236 15998 3238
rect 16022 3236 16078 3238
rect 17314 10104 17370 10160
rect 16946 4700 16948 4720
rect 16948 4700 17000 4720
rect 17000 4700 17002 4720
rect 16946 4664 17002 4700
rect 16946 4120 17002 4176
rect 16762 3576 16818 3632
rect 16486 3440 16542 3496
rect 17314 3984 17370 4040
rect 17682 10376 17738 10432
rect 17866 9288 17922 9344
rect 17774 8472 17830 8528
rect 17682 8064 17738 8120
rect 17682 7828 17684 7848
rect 17684 7828 17736 7848
rect 17736 7828 17738 7848
rect 17682 7792 17738 7828
rect 17590 7384 17646 7440
rect 17866 7792 17922 7848
rect 18142 13096 18198 13152
rect 18142 12144 18198 12200
rect 18234 10784 18290 10840
rect 18234 10512 18290 10568
rect 17774 6704 17830 6760
rect 17774 6160 17830 6216
rect 18050 7284 18052 7304
rect 18052 7284 18104 7304
rect 18104 7284 18106 7304
rect 18050 7248 18106 7284
rect 18050 5072 18106 5128
rect 17866 3984 17922 4040
rect 17774 3576 17830 3632
rect 17590 3032 17646 3088
rect 15782 2202 15838 2204
rect 15862 2202 15918 2204
rect 15942 2202 15998 2204
rect 16022 2202 16078 2204
rect 15782 2150 15808 2202
rect 15808 2150 15838 2202
rect 15862 2150 15872 2202
rect 15872 2150 15918 2202
rect 15942 2150 15988 2202
rect 15988 2150 15998 2202
rect 16022 2150 16052 2202
rect 16052 2150 16078 2202
rect 15782 2148 15838 2150
rect 15862 2148 15918 2150
rect 15942 2148 15998 2150
rect 16022 2148 16078 2150
rect 2778 176 2834 232
rect 15198 448 15254 504
rect 17498 2080 17554 2136
rect 18234 6568 18290 6624
rect 18234 5888 18290 5944
rect 18234 4256 18290 4312
rect 18050 2760 18106 2816
rect 17866 2488 17922 2544
rect 18418 5516 18420 5536
rect 18420 5516 18472 5536
rect 18472 5516 18474 5536
rect 18418 5480 18474 5516
rect 18418 3168 18474 3224
rect 18326 1672 18382 1728
rect 17866 856 17922 912
rect 18970 7012 18972 7032
rect 18972 7012 19024 7032
rect 19024 7012 19026 7032
rect 18970 6976 19026 7012
rect 18786 4664 18842 4720
rect 18602 1264 18658 1320
rect 15290 176 15346 232
<< metal3 >>
rect 0 16962 800 16992
rect 4061 16962 4127 16965
rect 0 16960 4127 16962
rect 0 16904 4066 16960
rect 4122 16904 4127 16960
rect 0 16902 4127 16904
rect 0 16872 800 16902
rect 4061 16899 4127 16902
rect 16481 16962 16547 16965
rect 19200 16962 20000 16992
rect 16481 16960 20000 16962
rect 16481 16904 16486 16960
rect 16542 16904 20000 16960
rect 16481 16902 20000 16904
rect 16481 16899 16547 16902
rect 19200 16872 20000 16902
rect 0 16690 800 16720
rect 2957 16690 3023 16693
rect 0 16688 3023 16690
rect 0 16632 2962 16688
rect 3018 16632 3023 16688
rect 0 16630 3023 16632
rect 0 16600 800 16630
rect 2957 16627 3023 16630
rect 15653 16554 15719 16557
rect 19200 16554 20000 16584
rect 15653 16552 20000 16554
rect 15653 16496 15658 16552
rect 15714 16496 20000 16552
rect 15653 16494 20000 16496
rect 15653 16491 15719 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 2129 16282 2195 16285
rect 0 16280 2195 16282
rect 0 16224 2134 16280
rect 2190 16224 2195 16280
rect 0 16222 2195 16224
rect 0 16192 800 16222
rect 2129 16219 2195 16222
rect 18413 16146 18479 16149
rect 19200 16146 20000 16176
rect 18413 16144 20000 16146
rect 18413 16088 18418 16144
rect 18474 16088 20000 16144
rect 18413 16086 20000 16088
rect 18413 16083 18479 16086
rect 19200 16056 20000 16086
rect 0 16010 800 16040
rect 2681 16010 2747 16013
rect 0 16008 2747 16010
rect 0 15952 2686 16008
rect 2742 15952 2747 16008
rect 0 15950 2747 15952
rect 0 15920 800 15950
rect 2681 15947 2747 15950
rect 15009 15738 15075 15741
rect 19200 15738 20000 15768
rect 15009 15736 20000 15738
rect 15009 15680 15014 15736
rect 15070 15680 20000 15736
rect 15009 15678 20000 15680
rect 15009 15675 15075 15678
rect 19200 15648 20000 15678
rect 0 15602 800 15632
rect 1393 15602 1459 15605
rect 0 15600 1459 15602
rect 0 15544 1398 15600
rect 1454 15544 1459 15600
rect 0 15542 1459 15544
rect 0 15512 800 15542
rect 1393 15539 1459 15542
rect 15469 15466 15535 15469
rect 19200 15466 20000 15496
rect 15469 15464 20000 15466
rect 15469 15408 15474 15464
rect 15530 15408 20000 15464
rect 15469 15406 20000 15408
rect 15469 15403 15535 15406
rect 19200 15376 20000 15406
rect 0 15330 800 15360
rect 2865 15330 2931 15333
rect 0 15328 2931 15330
rect 0 15272 2870 15328
rect 2926 15272 2931 15328
rect 0 15270 2931 15272
rect 0 15240 800 15270
rect 2865 15267 2931 15270
rect 0 15058 800 15088
rect 1669 15058 1735 15061
rect 0 15056 1735 15058
rect 0 15000 1674 15056
rect 1730 15000 1735 15056
rect 0 14998 1735 15000
rect 0 14968 800 14998
rect 1669 14995 1735 14998
rect 13445 15058 13511 15061
rect 19200 15058 20000 15088
rect 13445 15056 20000 15058
rect 13445 15000 13450 15056
rect 13506 15000 20000 15056
rect 13445 14998 20000 15000
rect 13445 14995 13511 14998
rect 19200 14968 20000 14998
rect 6874 14720 7194 14721
rect 0 14650 800 14680
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7194 14720
rect 6874 14655 7194 14656
rect 12805 14720 13125 14721
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 14655 13125 14656
rect 2773 14650 2839 14653
rect 0 14648 2839 14650
rect 0 14592 2778 14648
rect 2834 14592 2839 14648
rect 0 14590 2839 14592
rect 0 14560 800 14590
rect 2773 14587 2839 14590
rect 15193 14650 15259 14653
rect 19200 14650 20000 14680
rect 15193 14648 20000 14650
rect 15193 14592 15198 14648
rect 15254 14592 20000 14648
rect 15193 14590 20000 14592
rect 15193 14587 15259 14590
rect 19200 14560 20000 14590
rect 0 14378 800 14408
rect 1761 14378 1827 14381
rect 0 14376 1827 14378
rect 0 14320 1766 14376
rect 1822 14320 1827 14376
rect 0 14318 1827 14320
rect 0 14288 800 14318
rect 1761 14315 1827 14318
rect 16205 14242 16271 14245
rect 19200 14242 20000 14272
rect 16205 14240 20000 14242
rect 16205 14184 16210 14240
rect 16266 14184 20000 14240
rect 16205 14182 20000 14184
rect 16205 14179 16271 14182
rect 3909 14176 4229 14177
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 14111 4229 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 15770 14176 16090 14177
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16090 14176
rect 19200 14152 20000 14182
rect 15770 14111 16090 14112
rect 0 13970 800 14000
rect 2313 13970 2379 13973
rect 0 13968 2379 13970
rect 0 13912 2318 13968
rect 2374 13912 2379 13968
rect 0 13910 2379 13912
rect 0 13880 800 13910
rect 2313 13907 2379 13910
rect 12157 13834 12223 13837
rect 19200 13834 20000 13864
rect 12157 13832 20000 13834
rect 12157 13776 12162 13832
rect 12218 13776 20000 13832
rect 12157 13774 20000 13776
rect 12157 13771 12223 13774
rect 19200 13744 20000 13774
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 6874 13632 7194 13633
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7194 13632
rect 6874 13567 7194 13568
rect 12805 13632 13125 13633
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 13567 13125 13568
rect 16389 13562 16455 13565
rect 19200 13562 20000 13592
rect 16389 13560 20000 13562
rect 16389 13504 16394 13560
rect 16450 13504 20000 13560
rect 16389 13502 20000 13504
rect 16389 13499 16455 13502
rect 19200 13472 20000 13502
rect 0 13290 800 13320
rect 1853 13290 1919 13293
rect 0 13288 1919 13290
rect 0 13232 1858 13288
rect 1914 13232 1919 13288
rect 0 13230 1919 13232
rect 0 13200 800 13230
rect 1853 13227 1919 13230
rect 18137 13154 18203 13157
rect 19200 13154 20000 13184
rect 18137 13152 20000 13154
rect 18137 13096 18142 13152
rect 18198 13096 20000 13152
rect 18137 13094 20000 13096
rect 18137 13091 18203 13094
rect 3909 13088 4229 13089
rect 0 13018 800 13048
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 13023 4229 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 15770 13088 16090 13089
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16090 13088
rect 19200 13064 20000 13094
rect 15770 13023 16090 13024
rect 2129 13018 2195 13021
rect 0 13016 2195 13018
rect 0 12960 2134 13016
rect 2190 12960 2195 13016
rect 0 12958 2195 12960
rect 0 12928 800 12958
rect 2129 12955 2195 12958
rect 0 12746 800 12776
rect 3969 12746 4035 12749
rect 0 12744 4035 12746
rect 0 12688 3974 12744
rect 4030 12688 4035 12744
rect 0 12686 4035 12688
rect 0 12656 800 12686
rect 3969 12683 4035 12686
rect 15745 12746 15811 12749
rect 19200 12746 20000 12776
rect 15745 12744 20000 12746
rect 15745 12688 15750 12744
rect 15806 12688 20000 12744
rect 15745 12686 20000 12688
rect 15745 12683 15811 12686
rect 19200 12656 20000 12686
rect 6874 12544 7194 12545
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7194 12544
rect 6874 12479 7194 12480
rect 12805 12544 13125 12545
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 12479 13125 12480
rect 0 12338 800 12368
rect 3785 12338 3851 12341
rect 0 12336 3851 12338
rect 0 12280 3790 12336
rect 3846 12280 3851 12336
rect 0 12278 3851 12280
rect 0 12248 800 12278
rect 3785 12275 3851 12278
rect 15745 12338 15811 12341
rect 19200 12338 20000 12368
rect 15745 12336 20000 12338
rect 15745 12280 15750 12336
rect 15806 12280 20000 12336
rect 15745 12278 20000 12280
rect 15745 12275 15811 12278
rect 19200 12248 20000 12278
rect 11053 12202 11119 12205
rect 18137 12202 18203 12205
rect 11053 12200 18203 12202
rect 11053 12144 11058 12200
rect 11114 12144 18142 12200
rect 18198 12144 18203 12200
rect 11053 12142 18203 12144
rect 11053 12139 11119 12142
rect 18137 12139 18203 12142
rect 0 12066 800 12096
rect 3509 12066 3575 12069
rect 0 12064 3575 12066
rect 0 12008 3514 12064
rect 3570 12008 3575 12064
rect 0 12006 3575 12008
rect 0 11976 800 12006
rect 3509 12003 3575 12006
rect 3909 12000 4229 12001
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 11935 4229 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 15770 12000 16090 12001
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16090 12000
rect 15770 11935 16090 11936
rect 16297 11930 16363 11933
rect 19200 11930 20000 11960
rect 16297 11928 20000 11930
rect 16297 11872 16302 11928
rect 16358 11872 20000 11928
rect 16297 11870 20000 11872
rect 16297 11867 16363 11870
rect 19200 11840 20000 11870
rect 10777 11794 10843 11797
rect 11973 11794 12039 11797
rect 12157 11794 12223 11797
rect 10777 11792 12223 11794
rect 10777 11736 10782 11792
rect 10838 11736 11978 11792
rect 12034 11736 12162 11792
rect 12218 11736 12223 11792
rect 10777 11734 12223 11736
rect 10777 11731 10843 11734
rect 11973 11731 12039 11734
rect 12157 11731 12223 11734
rect 0 11658 800 11688
rect 3417 11658 3483 11661
rect 0 11656 3483 11658
rect 0 11600 3422 11656
rect 3478 11600 3483 11656
rect 0 11598 3483 11600
rect 0 11568 800 11598
rect 3417 11595 3483 11598
rect 10041 11658 10107 11661
rect 11697 11658 11763 11661
rect 10041 11656 11763 11658
rect 10041 11600 10046 11656
rect 10102 11600 11702 11656
rect 11758 11600 11763 11656
rect 10041 11598 11763 11600
rect 10041 11595 10107 11598
rect 11697 11595 11763 11598
rect 14641 11658 14707 11661
rect 19200 11658 20000 11688
rect 14641 11656 20000 11658
rect 14641 11600 14646 11656
rect 14702 11600 20000 11656
rect 14641 11598 20000 11600
rect 14641 11595 14707 11598
rect 19200 11568 20000 11598
rect 6874 11456 7194 11457
rect 0 11386 800 11416
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7194 11456
rect 6874 11391 7194 11392
rect 12805 11456 13125 11457
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 11391 13125 11392
rect 3325 11386 3391 11389
rect 0 11384 3391 11386
rect 0 11328 3330 11384
rect 3386 11328 3391 11384
rect 0 11326 3391 11328
rect 0 11296 800 11326
rect 3325 11323 3391 11326
rect 10869 11250 10935 11253
rect 12157 11250 12223 11253
rect 10869 11248 12223 11250
rect 10869 11192 10874 11248
rect 10930 11192 12162 11248
rect 12218 11192 12223 11248
rect 10869 11190 12223 11192
rect 10869 11187 10935 11190
rect 12157 11187 12223 11190
rect 15561 11250 15627 11253
rect 19200 11250 20000 11280
rect 15561 11248 20000 11250
rect 15561 11192 15566 11248
rect 15622 11192 20000 11248
rect 15561 11190 20000 11192
rect 15561 11187 15627 11190
rect 19200 11160 20000 11190
rect 1669 11114 1735 11117
rect 8017 11114 8083 11117
rect 1669 11112 8083 11114
rect 1669 11056 1674 11112
rect 1730 11056 8022 11112
rect 8078 11056 8083 11112
rect 1669 11054 8083 11056
rect 1669 11051 1735 11054
rect 8017 11051 8083 11054
rect 8293 11114 8359 11117
rect 8937 11114 9003 11117
rect 8293 11112 9003 11114
rect 8293 11056 8298 11112
rect 8354 11056 8942 11112
rect 8998 11056 9003 11112
rect 8293 11054 9003 11056
rect 8293 11051 8359 11054
rect 8937 11051 9003 11054
rect 9765 11114 9831 11117
rect 12065 11114 12131 11117
rect 9765 11112 12131 11114
rect 9765 11056 9770 11112
rect 9826 11056 12070 11112
rect 12126 11056 12131 11112
rect 9765 11054 12131 11056
rect 9765 11051 9831 11054
rect 12065 11051 12131 11054
rect 12249 11114 12315 11117
rect 12433 11114 12499 11117
rect 12249 11112 12499 11114
rect 12249 11056 12254 11112
rect 12310 11056 12438 11112
rect 12494 11056 12499 11112
rect 12249 11054 12499 11056
rect 12249 11051 12315 11054
rect 12433 11051 12499 11054
rect 0 10978 800 11008
rect 3417 10978 3483 10981
rect 0 10976 3483 10978
rect 0 10920 3422 10976
rect 3478 10920 3483 10976
rect 0 10918 3483 10920
rect 0 10888 800 10918
rect 3417 10915 3483 10918
rect 3909 10912 4229 10913
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 10847 4229 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 15770 10912 16090 10913
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16090 10912
rect 15770 10847 16090 10848
rect 8569 10842 8635 10845
rect 4340 10840 8635 10842
rect 4340 10784 8574 10840
rect 8630 10784 8635 10840
rect 4340 10782 8635 10784
rect 0 10706 800 10736
rect 4340 10706 4400 10782
rect 8569 10779 8635 10782
rect 18229 10842 18295 10845
rect 19200 10842 20000 10872
rect 18229 10840 20000 10842
rect 18229 10784 18234 10840
rect 18290 10784 20000 10840
rect 18229 10782 20000 10784
rect 18229 10779 18295 10782
rect 19200 10752 20000 10782
rect 0 10646 4400 10706
rect 4521 10706 4587 10709
rect 8477 10706 8543 10709
rect 4521 10704 8543 10706
rect 4521 10648 4526 10704
rect 4582 10648 8482 10704
rect 8538 10648 8543 10704
rect 4521 10646 8543 10648
rect 0 10616 800 10646
rect 4521 10643 4587 10646
rect 8477 10643 8543 10646
rect 11053 10570 11119 10573
rect 18229 10570 18295 10573
rect 11053 10568 18295 10570
rect 11053 10512 11058 10568
rect 11114 10512 18234 10568
rect 18290 10512 18295 10568
rect 11053 10510 18295 10512
rect 11053 10507 11119 10510
rect 18229 10507 18295 10510
rect 0 10434 800 10464
rect 5533 10434 5599 10437
rect 0 10432 5599 10434
rect 0 10376 5538 10432
rect 5594 10376 5599 10432
rect 0 10374 5599 10376
rect 0 10344 800 10374
rect 5533 10371 5599 10374
rect 17677 10434 17743 10437
rect 19200 10434 20000 10464
rect 17677 10432 20000 10434
rect 17677 10376 17682 10432
rect 17738 10376 20000 10432
rect 17677 10374 20000 10376
rect 17677 10371 17743 10374
rect 6874 10368 7194 10369
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7194 10368
rect 6874 10303 7194 10304
rect 12805 10368 13125 10369
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 19200 10344 20000 10374
rect 12805 10303 13125 10304
rect 9949 10162 10015 10165
rect 11145 10162 11211 10165
rect 9949 10160 11211 10162
rect 9949 10104 9954 10160
rect 10010 10104 11150 10160
rect 11206 10104 11211 10160
rect 9949 10102 11211 10104
rect 9949 10099 10015 10102
rect 11145 10099 11211 10102
rect 17309 10162 17375 10165
rect 17309 10160 17418 10162
rect 17309 10104 17314 10160
rect 17370 10104 17418 10160
rect 17309 10099 17418 10104
rect 0 10026 800 10056
rect 2865 10026 2931 10029
rect 0 10024 2931 10026
rect 0 9968 2870 10024
rect 2926 9968 2931 10024
rect 0 9966 2931 9968
rect 0 9936 800 9966
rect 2865 9963 2931 9966
rect 4429 10026 4495 10029
rect 5349 10026 5415 10029
rect 4429 10024 5415 10026
rect 4429 9968 4434 10024
rect 4490 9968 5354 10024
rect 5410 9968 5415 10024
rect 4429 9966 5415 9968
rect 4429 9963 4495 9966
rect 5349 9963 5415 9966
rect 9305 10026 9371 10029
rect 11053 10026 11119 10029
rect 9305 10024 11119 10026
rect 9305 9968 9310 10024
rect 9366 9968 11058 10024
rect 11114 9968 11119 10024
rect 9305 9966 11119 9968
rect 9305 9963 9371 9966
rect 11053 9963 11119 9966
rect 16481 10026 16547 10029
rect 17358 10026 17418 10099
rect 19200 10026 20000 10056
rect 16481 10024 20000 10026
rect 16481 9968 16486 10024
rect 16542 9968 20000 10024
rect 16481 9966 20000 9968
rect 16481 9963 16547 9966
rect 19200 9936 20000 9966
rect 11145 9890 11211 9893
rect 12382 9890 12388 9892
rect 11145 9888 12388 9890
rect 11145 9832 11150 9888
rect 11206 9832 12388 9888
rect 11145 9830 12388 9832
rect 11145 9827 11211 9830
rect 12382 9828 12388 9830
rect 12452 9828 12458 9892
rect 12525 9890 12591 9893
rect 15009 9890 15075 9893
rect 12525 9888 15075 9890
rect 12525 9832 12530 9888
rect 12586 9832 15014 9888
rect 15070 9832 15075 9888
rect 12525 9830 15075 9832
rect 12525 9827 12591 9830
rect 15009 9827 15075 9830
rect 3909 9824 4229 9825
rect 0 9754 800 9784
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 9759 4229 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 15770 9824 16090 9825
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16090 9824
rect 15770 9759 16090 9760
rect 2221 9754 2287 9757
rect 0 9752 2287 9754
rect 0 9696 2226 9752
rect 2282 9696 2287 9752
rect 0 9694 2287 9696
rect 0 9664 800 9694
rect 2221 9691 2287 9694
rect 17033 9754 17099 9757
rect 19200 9754 20000 9784
rect 17033 9752 20000 9754
rect 17033 9696 17038 9752
rect 17094 9696 20000 9752
rect 17033 9694 20000 9696
rect 17033 9691 17099 9694
rect 19200 9664 20000 9694
rect 3233 9618 3299 9621
rect 3509 9618 3575 9621
rect 3233 9616 3575 9618
rect 3233 9560 3238 9616
rect 3294 9560 3514 9616
rect 3570 9560 3575 9616
rect 3233 9558 3575 9560
rect 3233 9555 3299 9558
rect 3509 9555 3575 9558
rect 4613 9618 4679 9621
rect 5257 9618 5323 9621
rect 4613 9616 5323 9618
rect 4613 9560 4618 9616
rect 4674 9560 5262 9616
rect 5318 9560 5323 9616
rect 4613 9558 5323 9560
rect 4613 9555 4679 9558
rect 5257 9555 5323 9558
rect 10317 9618 10383 9621
rect 16849 9618 16915 9621
rect 10317 9616 16915 9618
rect 10317 9560 10322 9616
rect 10378 9560 16854 9616
rect 16910 9560 16915 9616
rect 10317 9558 16915 9560
rect 10317 9555 10383 9558
rect 16849 9555 16915 9558
rect 4797 9482 4863 9485
rect 14089 9482 14155 9485
rect 4797 9480 14155 9482
rect 4797 9424 4802 9480
rect 4858 9424 14094 9480
rect 14150 9424 14155 9480
rect 4797 9422 14155 9424
rect 4797 9419 4863 9422
rect 14089 9419 14155 9422
rect 0 9346 800 9376
rect 4245 9346 4311 9349
rect 0 9344 4311 9346
rect 0 9288 4250 9344
rect 4306 9288 4311 9344
rect 0 9286 4311 9288
rect 0 9256 800 9286
rect 4245 9283 4311 9286
rect 4705 9344 4771 9349
rect 4705 9288 4710 9344
rect 4766 9288 4771 9344
rect 4705 9283 4771 9288
rect 17861 9346 17927 9349
rect 19200 9346 20000 9376
rect 17861 9344 20000 9346
rect 17861 9288 17866 9344
rect 17922 9288 20000 9344
rect 17861 9286 20000 9288
rect 17861 9283 17927 9286
rect 2129 9210 2195 9213
rect 4708 9210 4768 9283
rect 6874 9280 7194 9281
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7194 9280
rect 6874 9215 7194 9216
rect 12805 9280 13125 9281
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 19200 9256 20000 9286
rect 12805 9215 13125 9216
rect 6177 9210 6243 9213
rect 2129 9208 6243 9210
rect 2129 9152 2134 9208
rect 2190 9152 6182 9208
rect 6238 9152 6243 9208
rect 2129 9150 6243 9152
rect 2129 9147 2195 9150
rect 6177 9147 6243 9150
rect 0 9074 800 9104
rect 3417 9074 3483 9077
rect 0 9072 3483 9074
rect 0 9016 3422 9072
rect 3478 9016 3483 9072
rect 0 9014 3483 9016
rect 0 8984 800 9014
rect 3417 9011 3483 9014
rect 12382 9012 12388 9076
rect 12452 9074 12458 9076
rect 13486 9074 13492 9076
rect 12452 9014 13492 9074
rect 12452 9012 12458 9014
rect 13486 9012 13492 9014
rect 13556 9074 13562 9076
rect 17125 9074 17191 9077
rect 13556 9072 17191 9074
rect 13556 9016 17130 9072
rect 17186 9016 17191 9072
rect 13556 9014 17191 9016
rect 13556 9012 13562 9014
rect 17125 9011 17191 9014
rect 7557 8938 7623 8941
rect 9397 8938 9463 8941
rect 3742 8936 9463 8938
rect 3742 8880 7562 8936
rect 7618 8880 9402 8936
rect 9458 8880 9463 8936
rect 3742 8878 9463 8880
rect 0 8802 800 8832
rect 3742 8802 3802 8878
rect 7557 8875 7623 8878
rect 9397 8875 9463 8878
rect 11605 8938 11671 8941
rect 12249 8938 12315 8941
rect 14273 8938 14339 8941
rect 11605 8936 14339 8938
rect 11605 8880 11610 8936
rect 11666 8880 12254 8936
rect 12310 8880 14278 8936
rect 14334 8880 14339 8936
rect 11605 8878 14339 8880
rect 11605 8875 11671 8878
rect 12249 8875 12315 8878
rect 14273 8875 14339 8878
rect 16113 8938 16179 8941
rect 19200 8938 20000 8968
rect 16113 8936 20000 8938
rect 16113 8880 16118 8936
rect 16174 8880 20000 8936
rect 16113 8878 20000 8880
rect 16113 8875 16179 8878
rect 19200 8848 20000 8878
rect 0 8742 3802 8802
rect 10593 8802 10659 8805
rect 11513 8802 11579 8805
rect 13629 8802 13695 8805
rect 10593 8800 13695 8802
rect 10593 8744 10598 8800
rect 10654 8744 11518 8800
rect 11574 8744 13634 8800
rect 13690 8744 13695 8800
rect 10593 8742 13695 8744
rect 0 8712 800 8742
rect 10593 8739 10659 8742
rect 11513 8739 11579 8742
rect 13629 8739 13695 8742
rect 3909 8736 4229 8737
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3909 8671 4229 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 15770 8736 16090 8737
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16090 8736
rect 15770 8671 16090 8672
rect 12525 8666 12591 8669
rect 13721 8666 13787 8669
rect 12525 8664 13787 8666
rect 12525 8608 12530 8664
rect 12586 8608 13726 8664
rect 13782 8608 13787 8664
rect 12525 8606 13787 8608
rect 12525 8603 12591 8606
rect 13721 8603 13787 8606
rect 13077 8530 13143 8533
rect 13302 8530 13308 8532
rect 13077 8528 13308 8530
rect 13077 8472 13082 8528
rect 13138 8472 13308 8528
rect 13077 8470 13308 8472
rect 13077 8467 13143 8470
rect 13302 8468 13308 8470
rect 13372 8468 13378 8532
rect 17769 8530 17835 8533
rect 19200 8530 20000 8560
rect 17769 8528 20000 8530
rect 17769 8472 17774 8528
rect 17830 8472 20000 8528
rect 17769 8470 20000 8472
rect 17769 8467 17835 8470
rect 19200 8440 20000 8470
rect 0 8394 800 8424
rect 5809 8394 5875 8397
rect 0 8392 5875 8394
rect 0 8336 5814 8392
rect 5870 8336 5875 8392
rect 0 8334 5875 8336
rect 0 8304 800 8334
rect 5809 8331 5875 8334
rect 6361 8394 6427 8397
rect 16297 8394 16363 8397
rect 6361 8392 16363 8394
rect 6361 8336 6366 8392
rect 6422 8336 16302 8392
rect 16358 8336 16363 8392
rect 6361 8334 16363 8336
rect 6361 8331 6427 8334
rect 16297 8331 16363 8334
rect 3325 8258 3391 8261
rect 3877 8258 3943 8261
rect 3325 8256 3943 8258
rect 3325 8200 3330 8256
rect 3386 8200 3882 8256
rect 3938 8200 3943 8256
rect 3325 8198 3943 8200
rect 3325 8195 3391 8198
rect 3877 8195 3943 8198
rect 9581 8258 9647 8261
rect 12249 8258 12315 8261
rect 9581 8256 12315 8258
rect 9581 8200 9586 8256
rect 9642 8200 12254 8256
rect 12310 8200 12315 8256
rect 9581 8198 12315 8200
rect 9581 8195 9647 8198
rect 12249 8195 12315 8198
rect 6874 8192 7194 8193
rect 0 8122 800 8152
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7194 8192
rect 6874 8127 7194 8128
rect 12805 8192 13125 8193
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 12805 8127 13125 8128
rect 3601 8122 3667 8125
rect 0 8120 3667 8122
rect 0 8064 3606 8120
rect 3662 8064 3667 8120
rect 0 8062 3667 8064
rect 0 8032 800 8062
rect 3601 8059 3667 8062
rect 11789 8122 11855 8125
rect 12341 8122 12407 8125
rect 11789 8120 12407 8122
rect 11789 8064 11794 8120
rect 11850 8064 12346 8120
rect 12402 8064 12407 8120
rect 11789 8062 12407 8064
rect 11789 8059 11855 8062
rect 12341 8059 12407 8062
rect 17677 8122 17743 8125
rect 19200 8122 20000 8152
rect 17677 8120 20000 8122
rect 17677 8064 17682 8120
rect 17738 8064 20000 8120
rect 17677 8062 20000 8064
rect 17677 8059 17743 8062
rect 19200 8032 20000 8062
rect 2865 7986 2931 7989
rect 3366 7986 3372 7988
rect 2865 7984 3372 7986
rect 2865 7928 2870 7984
rect 2926 7928 3372 7984
rect 2865 7926 3372 7928
rect 2865 7923 2931 7926
rect 3366 7924 3372 7926
rect 3436 7924 3442 7988
rect 4521 7986 4587 7989
rect 9857 7986 9923 7989
rect 11881 7986 11947 7989
rect 13537 7986 13603 7989
rect 4521 7984 4722 7986
rect 4521 7928 4526 7984
rect 4582 7928 4722 7984
rect 4521 7926 4722 7928
rect 4521 7923 4587 7926
rect 0 7714 800 7744
rect 2129 7714 2195 7717
rect 0 7712 2195 7714
rect 0 7656 2134 7712
rect 2190 7656 2195 7712
rect 0 7654 2195 7656
rect 0 7624 800 7654
rect 2129 7651 2195 7654
rect 3909 7648 4229 7649
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 7583 4229 7584
rect 0 7442 800 7472
rect 2405 7442 2471 7445
rect 2773 7442 2839 7445
rect 0 7440 2839 7442
rect 0 7384 2410 7440
rect 2466 7384 2778 7440
rect 2834 7384 2839 7440
rect 0 7382 2839 7384
rect 0 7352 800 7382
rect 2405 7379 2471 7382
rect 2773 7379 2839 7382
rect 4662 7306 4722 7926
rect 9857 7984 13603 7986
rect 9857 7928 9862 7984
rect 9918 7928 11886 7984
rect 11942 7928 13542 7984
rect 13598 7928 13603 7984
rect 9857 7926 13603 7928
rect 9857 7923 9923 7926
rect 11881 7923 11947 7926
rect 13537 7923 13603 7926
rect 4889 7850 4955 7853
rect 6545 7850 6611 7853
rect 16481 7850 16547 7853
rect 17677 7850 17743 7853
rect 4889 7848 6611 7850
rect 4889 7792 4894 7848
rect 4950 7792 6550 7848
rect 6606 7792 6611 7848
rect 4889 7790 6611 7792
rect 4889 7787 4955 7790
rect 6545 7787 6611 7790
rect 14736 7848 17743 7850
rect 14736 7792 16486 7848
rect 16542 7792 17682 7848
rect 17738 7792 17743 7848
rect 14736 7790 17743 7792
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 14736 7581 14796 7790
rect 16481 7787 16547 7790
rect 17677 7787 17743 7790
rect 17861 7850 17927 7853
rect 19200 7850 20000 7880
rect 17861 7848 20000 7850
rect 17861 7792 17866 7848
rect 17922 7792 20000 7848
rect 17861 7790 20000 7792
rect 17861 7787 17927 7790
rect 19200 7760 20000 7790
rect 15770 7648 16090 7649
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16090 7648
rect 15770 7583 16090 7584
rect 5441 7578 5507 7581
rect 10501 7578 10567 7581
rect 14733 7578 14799 7581
rect 5441 7576 5642 7578
rect 5441 7520 5446 7576
rect 5502 7520 5642 7576
rect 5441 7518 5642 7520
rect 5441 7515 5507 7518
rect 5582 7309 5642 7518
rect 10501 7576 14799 7578
rect 10501 7520 10506 7576
rect 10562 7520 14738 7576
rect 14794 7520 14799 7576
rect 10501 7518 14799 7520
rect 10501 7515 10567 7518
rect 14733 7515 14799 7518
rect 10685 7442 10751 7445
rect 12065 7442 12131 7445
rect 17585 7442 17651 7445
rect 19200 7442 20000 7472
rect 10685 7440 17418 7442
rect 10685 7384 10690 7440
rect 10746 7384 12070 7440
rect 12126 7384 17418 7440
rect 10685 7382 17418 7384
rect 10685 7379 10751 7382
rect 12065 7379 12131 7382
rect 5165 7306 5231 7309
rect 4662 7304 5231 7306
rect 4662 7248 5170 7304
rect 5226 7248 5231 7304
rect 4662 7246 5231 7248
rect 5582 7304 5691 7309
rect 5582 7248 5630 7304
rect 5686 7248 5691 7304
rect 5582 7246 5691 7248
rect 5165 7243 5231 7246
rect 5625 7243 5691 7246
rect 8385 7306 8451 7309
rect 11462 7306 11468 7308
rect 8385 7304 11468 7306
rect 8385 7248 8390 7304
rect 8446 7248 11468 7304
rect 8385 7246 11468 7248
rect 8385 7243 8451 7246
rect 11462 7244 11468 7246
rect 11532 7306 11538 7308
rect 14825 7306 14891 7309
rect 11532 7304 14891 7306
rect 11532 7248 14830 7304
rect 14886 7248 14891 7304
rect 11532 7246 14891 7248
rect 17358 7306 17418 7382
rect 17585 7440 20000 7442
rect 17585 7384 17590 7440
rect 17646 7384 20000 7440
rect 17585 7382 20000 7384
rect 17585 7379 17651 7382
rect 19200 7352 20000 7382
rect 18045 7306 18111 7309
rect 17358 7304 18111 7306
rect 17358 7248 18050 7304
rect 18106 7248 18111 7304
rect 17358 7246 18111 7248
rect 11532 7244 11538 7246
rect 14825 7243 14891 7246
rect 18045 7243 18111 7246
rect 1301 7170 1367 7173
rect 4889 7170 4955 7173
rect 1301 7168 4955 7170
rect 1301 7112 1306 7168
rect 1362 7112 4894 7168
rect 4950 7112 4955 7168
rect 1301 7110 4955 7112
rect 1301 7107 1367 7110
rect 4889 7107 4955 7110
rect 7373 7170 7439 7173
rect 12566 7170 12572 7172
rect 7373 7168 12572 7170
rect 7373 7112 7378 7168
rect 7434 7112 12572 7168
rect 7373 7110 12572 7112
rect 7373 7107 7439 7110
rect 12566 7108 12572 7110
rect 12636 7108 12642 7172
rect 6874 7104 7194 7105
rect 0 7034 800 7064
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7194 7104
rect 6874 7039 7194 7040
rect 12805 7104 13125 7105
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 7039 13125 7040
rect 3693 7034 3759 7037
rect 4153 7034 4219 7037
rect 0 7032 4219 7034
rect 0 6976 3698 7032
rect 3754 6976 4158 7032
rect 4214 6976 4219 7032
rect 0 6974 4219 6976
rect 0 6944 800 6974
rect 3693 6971 3759 6974
rect 4153 6971 4219 6974
rect 10409 7034 10475 7037
rect 10777 7034 10843 7037
rect 10409 7032 10843 7034
rect 10409 6976 10414 7032
rect 10470 6976 10782 7032
rect 10838 6976 10843 7032
rect 10409 6974 10843 6976
rect 10409 6971 10475 6974
rect 10777 6971 10843 6974
rect 18965 7034 19031 7037
rect 19200 7034 20000 7064
rect 18965 7032 20000 7034
rect 18965 6976 18970 7032
rect 19026 6976 20000 7032
rect 18965 6974 20000 6976
rect 18965 6971 19031 6974
rect 19200 6944 20000 6974
rect 2681 6898 2747 6901
rect 2957 6898 3023 6901
rect 2681 6896 3023 6898
rect 2681 6840 2686 6896
rect 2742 6840 2962 6896
rect 3018 6840 3023 6896
rect 2681 6838 3023 6840
rect 2681 6835 2747 6838
rect 2957 6835 3023 6838
rect 10317 6898 10383 6901
rect 16941 6898 17007 6901
rect 10317 6896 17007 6898
rect 10317 6840 10322 6896
rect 10378 6840 16946 6896
rect 17002 6840 17007 6896
rect 10317 6838 17007 6840
rect 10317 6835 10383 6838
rect 16941 6835 17007 6838
rect 0 6762 800 6792
rect 1669 6762 1735 6765
rect 0 6760 1735 6762
rect 0 6704 1674 6760
rect 1730 6704 1735 6760
rect 0 6702 1735 6704
rect 0 6672 800 6702
rect 1669 6699 1735 6702
rect 12433 6762 12499 6765
rect 13629 6762 13695 6765
rect 13905 6762 13971 6765
rect 12433 6760 13971 6762
rect 12433 6704 12438 6760
rect 12494 6704 13634 6760
rect 13690 6704 13910 6760
rect 13966 6704 13971 6760
rect 12433 6702 13971 6704
rect 12433 6699 12499 6702
rect 13629 6699 13695 6702
rect 13905 6699 13971 6702
rect 15009 6762 15075 6765
rect 17769 6762 17835 6765
rect 15009 6760 17835 6762
rect 15009 6704 15014 6760
rect 15070 6704 17774 6760
rect 17830 6704 17835 6760
rect 15009 6702 17835 6704
rect 15009 6699 15075 6702
rect 17769 6699 17835 6702
rect 18229 6626 18295 6629
rect 19200 6626 20000 6656
rect 18229 6624 20000 6626
rect 18229 6568 18234 6624
rect 18290 6568 20000 6624
rect 18229 6566 20000 6568
rect 18229 6563 18295 6566
rect 3909 6560 4229 6561
rect 0 6490 800 6520
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3909 6495 4229 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 15770 6560 16090 6561
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16090 6560
rect 19200 6536 20000 6566
rect 15770 6495 16090 6496
rect 3693 6490 3759 6493
rect 0 6488 3759 6490
rect 0 6432 3698 6488
rect 3754 6432 3759 6488
rect 0 6430 3759 6432
rect 0 6400 800 6430
rect 3693 6427 3759 6430
rect 12341 6490 12407 6493
rect 13905 6490 13971 6493
rect 12341 6488 13971 6490
rect 12341 6432 12346 6488
rect 12402 6432 13910 6488
rect 13966 6432 13971 6488
rect 12341 6430 13971 6432
rect 12341 6427 12407 6430
rect 13905 6427 13971 6430
rect 10961 6354 11027 6357
rect 12801 6354 12867 6357
rect 10961 6352 12867 6354
rect 10961 6296 10966 6352
rect 11022 6296 12806 6352
rect 12862 6296 12867 6352
rect 10961 6294 12867 6296
rect 10961 6291 11027 6294
rect 12801 6291 12867 6294
rect 1945 6218 2011 6221
rect 3366 6218 3372 6220
rect 1945 6216 3372 6218
rect 1945 6160 1950 6216
rect 2006 6160 3372 6216
rect 1945 6158 3372 6160
rect 1945 6155 2011 6158
rect 3366 6156 3372 6158
rect 3436 6218 3442 6220
rect 7833 6218 7899 6221
rect 3436 6216 7899 6218
rect 3436 6160 7838 6216
rect 7894 6160 7899 6216
rect 3436 6158 7899 6160
rect 3436 6156 3442 6158
rect 7833 6155 7899 6158
rect 11513 6218 11579 6221
rect 12249 6218 12315 6221
rect 11513 6216 12315 6218
rect 11513 6160 11518 6216
rect 11574 6160 12254 6216
rect 12310 6160 12315 6216
rect 11513 6158 12315 6160
rect 11513 6155 11579 6158
rect 12249 6155 12315 6158
rect 17769 6218 17835 6221
rect 19200 6218 20000 6248
rect 17769 6216 20000 6218
rect 17769 6160 17774 6216
rect 17830 6160 20000 6216
rect 17769 6158 20000 6160
rect 17769 6155 17835 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 1577 6082 1643 6085
rect 0 6080 1643 6082
rect 0 6024 1582 6080
rect 1638 6024 1643 6080
rect 0 6022 1643 6024
rect 0 5992 800 6022
rect 1577 6019 1643 6022
rect 6874 6016 7194 6017
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7194 6016
rect 6874 5951 7194 5952
rect 12805 6016 13125 6017
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12805 5951 13125 5952
rect 2221 5946 2287 5949
rect 3141 5946 3207 5949
rect 13537 5948 13603 5949
rect 2221 5944 3207 5946
rect 2221 5888 2226 5944
rect 2282 5888 3146 5944
rect 3202 5888 3207 5944
rect 2221 5886 3207 5888
rect 2221 5883 2287 5886
rect 3141 5883 3207 5886
rect 13486 5884 13492 5948
rect 13556 5946 13603 5948
rect 18229 5946 18295 5949
rect 19200 5946 20000 5976
rect 13556 5944 13648 5946
rect 13598 5888 13648 5944
rect 13556 5886 13648 5888
rect 18229 5944 20000 5946
rect 18229 5888 18234 5944
rect 18290 5888 20000 5944
rect 18229 5886 20000 5888
rect 13556 5884 13603 5886
rect 13537 5883 13603 5884
rect 18229 5883 18295 5886
rect 19200 5856 20000 5886
rect 0 5810 800 5840
rect 3233 5810 3299 5813
rect 0 5808 3299 5810
rect 0 5752 3238 5808
rect 3294 5752 3299 5808
rect 0 5750 3299 5752
rect 0 5720 800 5750
rect 3233 5747 3299 5750
rect 3366 5748 3372 5812
rect 3436 5810 3442 5812
rect 3509 5810 3575 5813
rect 3436 5808 3575 5810
rect 3436 5752 3514 5808
rect 3570 5752 3575 5808
rect 3436 5750 3575 5752
rect 3436 5748 3442 5750
rect 3509 5747 3575 5750
rect 10409 5810 10475 5813
rect 13353 5810 13419 5813
rect 10409 5808 13419 5810
rect 10409 5752 10414 5808
rect 10470 5752 13358 5808
rect 13414 5752 13419 5808
rect 10409 5750 13419 5752
rect 10409 5747 10475 5750
rect 13353 5747 13419 5750
rect 1117 5674 1183 5677
rect 7833 5674 7899 5677
rect 1117 5672 7899 5674
rect 1117 5616 1122 5672
rect 1178 5616 7838 5672
rect 7894 5616 7899 5672
rect 1117 5614 7899 5616
rect 1117 5611 1183 5614
rect 7833 5611 7899 5614
rect 13537 5674 13603 5677
rect 14273 5674 14339 5677
rect 13537 5672 14339 5674
rect 13537 5616 13542 5672
rect 13598 5616 14278 5672
rect 14334 5616 14339 5672
rect 13537 5614 14339 5616
rect 13537 5611 13603 5614
rect 14273 5611 14339 5614
rect 12249 5538 12315 5541
rect 14917 5538 14983 5541
rect 12249 5536 14983 5538
rect 12249 5480 12254 5536
rect 12310 5480 14922 5536
rect 14978 5480 14983 5536
rect 12249 5478 14983 5480
rect 12249 5475 12315 5478
rect 14917 5475 14983 5478
rect 18413 5538 18479 5541
rect 19200 5538 20000 5568
rect 18413 5536 20000 5538
rect 18413 5480 18418 5536
rect 18474 5480 20000 5536
rect 18413 5478 20000 5480
rect 18413 5475 18479 5478
rect 3909 5472 4229 5473
rect 0 5402 800 5432
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 5407 4229 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 15770 5472 16090 5473
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16090 5472
rect 19200 5448 20000 5478
rect 15770 5407 16090 5408
rect 12157 5402 12223 5405
rect 13721 5402 13787 5405
rect 0 5342 3618 5402
rect 0 5312 800 5342
rect 3558 5266 3618 5342
rect 12157 5400 13787 5402
rect 12157 5344 12162 5400
rect 12218 5344 13726 5400
rect 13782 5344 13787 5400
rect 12157 5342 13787 5344
rect 12157 5339 12223 5342
rect 13721 5339 13787 5342
rect 4429 5266 4495 5269
rect 3558 5264 4495 5266
rect 3558 5208 4434 5264
rect 4490 5208 4495 5264
rect 3558 5206 4495 5208
rect 4429 5203 4495 5206
rect 11513 5266 11579 5269
rect 12433 5266 12499 5269
rect 11513 5264 12499 5266
rect 11513 5208 11518 5264
rect 11574 5208 12438 5264
rect 12494 5208 12499 5264
rect 11513 5206 12499 5208
rect 11513 5203 11579 5206
rect 12433 5203 12499 5206
rect 12566 5204 12572 5268
rect 12636 5266 12642 5268
rect 14181 5266 14247 5269
rect 12636 5264 14247 5266
rect 12636 5208 14186 5264
rect 14242 5208 14247 5264
rect 12636 5206 14247 5208
rect 12636 5204 12642 5206
rect 14181 5203 14247 5206
rect 0 5130 800 5160
rect 1853 5130 1919 5133
rect 0 5128 1919 5130
rect 0 5072 1858 5128
rect 1914 5072 1919 5128
rect 0 5070 1919 5072
rect 0 5040 800 5070
rect 1853 5067 1919 5070
rect 4061 5130 4127 5133
rect 9121 5130 9187 5133
rect 4061 5128 9187 5130
rect 4061 5072 4066 5128
rect 4122 5072 9126 5128
rect 9182 5072 9187 5128
rect 4061 5070 9187 5072
rect 4061 5067 4127 5070
rect 9121 5067 9187 5070
rect 18045 5130 18111 5133
rect 19200 5130 20000 5160
rect 18045 5128 20000 5130
rect 18045 5072 18050 5128
rect 18106 5072 20000 5128
rect 18045 5070 20000 5072
rect 18045 5067 18111 5070
rect 19200 5040 20000 5070
rect 6874 4928 7194 4929
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7194 4928
rect 6874 4863 7194 4864
rect 12805 4928 13125 4929
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 12805 4863 13125 4864
rect 0 4722 800 4752
rect 1577 4722 1643 4725
rect 0 4720 1643 4722
rect 0 4664 1582 4720
rect 1638 4664 1643 4720
rect 0 4662 1643 4664
rect 0 4632 800 4662
rect 1577 4659 1643 4662
rect 2037 4722 2103 4725
rect 6361 4722 6427 4725
rect 2037 4720 6427 4722
rect 2037 4664 2042 4720
rect 2098 4664 6366 4720
rect 6422 4664 6427 4720
rect 2037 4662 6427 4664
rect 2037 4659 2103 4662
rect 6361 4659 6427 4662
rect 13629 4722 13695 4725
rect 16941 4722 17007 4725
rect 13629 4720 17007 4722
rect 13629 4664 13634 4720
rect 13690 4664 16946 4720
rect 17002 4664 17007 4720
rect 13629 4662 17007 4664
rect 13629 4659 13695 4662
rect 16941 4659 17007 4662
rect 18781 4722 18847 4725
rect 19200 4722 20000 4752
rect 18781 4720 20000 4722
rect 18781 4664 18786 4720
rect 18842 4664 20000 4720
rect 18781 4662 20000 4664
rect 18781 4659 18847 4662
rect 19200 4632 20000 4662
rect 2681 4586 2747 4589
rect 11053 4586 11119 4589
rect 13813 4586 13879 4589
rect 2681 4584 4492 4586
rect 2681 4528 2686 4584
rect 2742 4528 4492 4584
rect 2681 4526 4492 4528
rect 2681 4523 2747 4526
rect 0 4450 800 4480
rect 4432 4453 4492 4526
rect 11053 4584 13879 4586
rect 11053 4528 11058 4584
rect 11114 4528 13818 4584
rect 13874 4528 13879 4584
rect 11053 4526 13879 4528
rect 11053 4523 11119 4526
rect 13813 4523 13879 4526
rect 2221 4450 2287 4453
rect 0 4448 2287 4450
rect 0 4392 2226 4448
rect 2282 4392 2287 4448
rect 0 4390 2287 4392
rect 0 4360 800 4390
rect 2221 4387 2287 4390
rect 4429 4450 4495 4453
rect 7557 4450 7623 4453
rect 4429 4448 7623 4450
rect 4429 4392 4434 4448
rect 4490 4392 7562 4448
rect 7618 4392 7623 4448
rect 4429 4390 7623 4392
rect 4429 4387 4495 4390
rect 7557 4387 7623 4390
rect 10225 4450 10291 4453
rect 13302 4450 13308 4452
rect 10225 4448 13308 4450
rect 10225 4392 10230 4448
rect 10286 4392 13308 4448
rect 10225 4390 13308 4392
rect 10225 4387 10291 4390
rect 13302 4388 13308 4390
rect 13372 4450 13378 4452
rect 14641 4450 14707 4453
rect 13372 4448 14707 4450
rect 13372 4392 14646 4448
rect 14702 4392 14707 4448
rect 13372 4390 14707 4392
rect 13372 4388 13378 4390
rect 14641 4387 14707 4390
rect 3909 4384 4229 4385
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 4319 4229 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 15770 4384 16090 4385
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16090 4384
rect 15770 4319 16090 4320
rect 18229 4314 18295 4317
rect 19200 4314 20000 4344
rect 18229 4312 20000 4314
rect 18229 4256 18234 4312
rect 18290 4256 20000 4312
rect 18229 4254 20000 4256
rect 18229 4251 18295 4254
rect 19200 4224 20000 4254
rect 0 4178 800 4208
rect 1853 4178 1919 4181
rect 0 4176 1919 4178
rect 0 4120 1858 4176
rect 1914 4120 1919 4176
rect 0 4118 1919 4120
rect 0 4088 800 4118
rect 1853 4115 1919 4118
rect 3601 4178 3667 4181
rect 6545 4178 6611 4181
rect 3601 4176 6611 4178
rect 3601 4120 3606 4176
rect 3662 4120 6550 4176
rect 6606 4120 6611 4176
rect 3601 4118 6611 4120
rect 3601 4115 3667 4118
rect 6545 4115 6611 4118
rect 12433 4178 12499 4181
rect 16941 4178 17007 4181
rect 12433 4176 17007 4178
rect 12433 4120 12438 4176
rect 12494 4120 16946 4176
rect 17002 4120 17007 4176
rect 12433 4118 17007 4120
rect 12433 4115 12499 4118
rect 16941 4115 17007 4118
rect 3417 4042 3483 4045
rect 17309 4042 17375 4045
rect 3417 4040 17375 4042
rect 3417 3984 3422 4040
rect 3478 3984 17314 4040
rect 17370 3984 17375 4040
rect 3417 3982 17375 3984
rect 3417 3979 3483 3982
rect 17309 3979 17375 3982
rect 17861 4042 17927 4045
rect 19200 4042 20000 4072
rect 17861 4040 20000 4042
rect 17861 3984 17866 4040
rect 17922 3984 20000 4040
rect 17861 3982 20000 3984
rect 17861 3979 17927 3982
rect 19200 3952 20000 3982
rect 8569 3906 8635 3909
rect 11329 3906 11395 3909
rect 8569 3904 11395 3906
rect 8569 3848 8574 3904
rect 8630 3848 11334 3904
rect 11390 3848 11395 3904
rect 8569 3846 11395 3848
rect 8569 3843 8635 3846
rect 11329 3843 11395 3846
rect 11462 3844 11468 3908
rect 11532 3906 11538 3908
rect 11605 3906 11671 3909
rect 11532 3904 11671 3906
rect 11532 3848 11610 3904
rect 11666 3848 11671 3904
rect 11532 3846 11671 3848
rect 11532 3844 11538 3846
rect 11605 3843 11671 3846
rect 6874 3840 7194 3841
rect 0 3770 800 3800
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7194 3840
rect 6874 3775 7194 3776
rect 12805 3840 13125 3841
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 3775 13125 3776
rect 1669 3770 1735 3773
rect 0 3768 1735 3770
rect 0 3712 1674 3768
rect 1730 3712 1735 3768
rect 0 3710 1735 3712
rect 0 3680 800 3710
rect 1669 3707 1735 3710
rect 8661 3770 8727 3773
rect 12433 3770 12499 3773
rect 8661 3768 12499 3770
rect 8661 3712 8666 3768
rect 8722 3712 12438 3768
rect 12494 3712 12499 3768
rect 8661 3710 12499 3712
rect 8661 3707 8727 3710
rect 12433 3707 12499 3710
rect 1209 3634 1275 3637
rect 16757 3634 16823 3637
rect 1209 3632 16823 3634
rect 1209 3576 1214 3632
rect 1270 3576 16762 3632
rect 16818 3576 16823 3632
rect 1209 3574 16823 3576
rect 1209 3571 1275 3574
rect 16757 3571 16823 3574
rect 17769 3634 17835 3637
rect 19200 3634 20000 3664
rect 17769 3632 20000 3634
rect 17769 3576 17774 3632
rect 17830 3576 20000 3632
rect 17769 3574 20000 3576
rect 17769 3571 17835 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 2405 3498 2471 3501
rect 0 3496 2471 3498
rect 0 3440 2410 3496
rect 2466 3440 2471 3496
rect 0 3438 2471 3440
rect 0 3408 800 3438
rect 2405 3435 2471 3438
rect 5993 3498 6059 3501
rect 16481 3498 16547 3501
rect 5993 3496 16547 3498
rect 5993 3440 5998 3496
rect 6054 3440 16486 3496
rect 16542 3440 16547 3496
rect 5993 3438 16547 3440
rect 5993 3435 6059 3438
rect 16481 3435 16547 3438
rect 3909 3296 4229 3297
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 3231 4229 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 15770 3296 16090 3297
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16090 3296
rect 15770 3231 16090 3232
rect 10501 3226 10567 3229
rect 12341 3226 12407 3229
rect 14733 3226 14799 3229
rect 10501 3224 11898 3226
rect 10501 3168 10506 3224
rect 10562 3168 11898 3224
rect 10501 3166 11898 3168
rect 10501 3163 10567 3166
rect 0 3090 800 3120
rect 2037 3090 2103 3093
rect 0 3088 2103 3090
rect 0 3032 2042 3088
rect 2098 3032 2103 3088
rect 0 3030 2103 3032
rect 0 3000 800 3030
rect 2037 3027 2103 3030
rect 2773 3090 2839 3093
rect 7005 3090 7071 3093
rect 2773 3088 7071 3090
rect 2773 3032 2778 3088
rect 2834 3032 7010 3088
rect 7066 3032 7071 3088
rect 2773 3030 7071 3032
rect 2773 3027 2839 3030
rect 7005 3027 7071 3030
rect 7649 3090 7715 3093
rect 11697 3090 11763 3093
rect 7649 3088 11763 3090
rect 7649 3032 7654 3088
rect 7710 3032 11702 3088
rect 11758 3032 11763 3088
rect 7649 3030 11763 3032
rect 11838 3090 11898 3166
rect 12341 3224 14799 3226
rect 12341 3168 12346 3224
rect 12402 3168 14738 3224
rect 14794 3168 14799 3224
rect 12341 3166 14799 3168
rect 12341 3163 12407 3166
rect 14733 3163 14799 3166
rect 18413 3226 18479 3229
rect 19200 3226 20000 3256
rect 18413 3224 20000 3226
rect 18413 3168 18418 3224
rect 18474 3168 20000 3224
rect 18413 3166 20000 3168
rect 18413 3163 18479 3166
rect 19200 3136 20000 3166
rect 15193 3090 15259 3093
rect 11838 3088 15259 3090
rect 11838 3032 15198 3088
rect 15254 3032 15259 3088
rect 11838 3030 15259 3032
rect 7649 3027 7715 3030
rect 11697 3027 11763 3030
rect 15193 3027 15259 3030
rect 15377 3090 15443 3093
rect 17585 3090 17651 3093
rect 15377 3088 17651 3090
rect 15377 3032 15382 3088
rect 15438 3032 17590 3088
rect 17646 3032 17651 3088
rect 15377 3030 17651 3032
rect 15377 3027 15443 3030
rect 17585 3027 17651 3030
rect 3049 2954 3115 2957
rect 10501 2954 10567 2957
rect 3049 2952 10567 2954
rect 3049 2896 3054 2952
rect 3110 2896 10506 2952
rect 10562 2896 10567 2952
rect 3049 2894 10567 2896
rect 3049 2891 3115 2894
rect 10501 2891 10567 2894
rect 10961 2954 11027 2957
rect 12617 2954 12683 2957
rect 10961 2952 12683 2954
rect 10961 2896 10966 2952
rect 11022 2896 12622 2952
rect 12678 2896 12683 2952
rect 10961 2894 12683 2896
rect 10961 2891 11027 2894
rect 12617 2891 12683 2894
rect 0 2818 800 2848
rect 4061 2818 4127 2821
rect 0 2816 4127 2818
rect 0 2760 4066 2816
rect 4122 2760 4127 2816
rect 0 2758 4127 2760
rect 0 2728 800 2758
rect 4061 2755 4127 2758
rect 4521 2818 4587 2821
rect 5349 2818 5415 2821
rect 4521 2816 5415 2818
rect 4521 2760 4526 2816
rect 4582 2760 5354 2816
rect 5410 2760 5415 2816
rect 4521 2758 5415 2760
rect 4521 2755 4587 2758
rect 5349 2755 5415 2758
rect 7373 2818 7439 2821
rect 11513 2818 11579 2821
rect 7373 2816 11579 2818
rect 7373 2760 7378 2816
rect 7434 2760 11518 2816
rect 11574 2760 11579 2816
rect 7373 2758 11579 2760
rect 7373 2755 7439 2758
rect 11513 2755 11579 2758
rect 18045 2818 18111 2821
rect 19200 2818 20000 2848
rect 18045 2816 20000 2818
rect 18045 2760 18050 2816
rect 18106 2760 20000 2816
rect 18045 2758 20000 2760
rect 18045 2755 18111 2758
rect 6874 2752 7194 2753
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7194 2752
rect 6874 2687 7194 2688
rect 12805 2752 13125 2753
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 19200 2728 20000 2758
rect 12805 2687 13125 2688
rect 2129 2682 2195 2685
rect 5441 2682 5507 2685
rect 2129 2680 5507 2682
rect 2129 2624 2134 2680
rect 2190 2624 5446 2680
rect 5502 2624 5507 2680
rect 2129 2622 5507 2624
rect 2129 2619 2195 2622
rect 5441 2619 5507 2622
rect 2497 2546 2563 2549
rect 3509 2546 3575 2549
rect 2497 2544 3575 2546
rect 2497 2488 2502 2544
rect 2558 2488 3514 2544
rect 3570 2488 3575 2544
rect 2497 2486 3575 2488
rect 2497 2483 2563 2486
rect 3509 2483 3575 2486
rect 9673 2546 9739 2549
rect 14089 2546 14155 2549
rect 9673 2544 14155 2546
rect 9673 2488 9678 2544
rect 9734 2488 14094 2544
rect 14150 2488 14155 2544
rect 9673 2486 14155 2488
rect 9673 2483 9739 2486
rect 14089 2483 14155 2486
rect 17861 2546 17927 2549
rect 17861 2544 18154 2546
rect 17861 2488 17866 2544
rect 17922 2488 18154 2544
rect 17861 2486 18154 2488
rect 17861 2483 17927 2486
rect 0 2410 800 2440
rect 1577 2410 1643 2413
rect 0 2408 1643 2410
rect 0 2352 1582 2408
rect 1638 2352 1643 2408
rect 0 2350 1643 2352
rect 0 2320 800 2350
rect 1577 2347 1643 2350
rect 10133 2410 10199 2413
rect 15377 2410 15443 2413
rect 10133 2408 15443 2410
rect 10133 2352 10138 2408
rect 10194 2352 15382 2408
rect 15438 2352 15443 2408
rect 10133 2350 15443 2352
rect 18094 2410 18154 2486
rect 19200 2410 20000 2440
rect 18094 2350 20000 2410
rect 10133 2347 10199 2350
rect 15377 2347 15443 2350
rect 19200 2320 20000 2350
rect 10409 2274 10475 2277
rect 13169 2274 13235 2277
rect 10409 2272 13235 2274
rect 10409 2216 10414 2272
rect 10470 2216 13174 2272
rect 13230 2216 13235 2272
rect 10409 2214 13235 2216
rect 10409 2211 10475 2214
rect 13169 2211 13235 2214
rect 3909 2208 4229 2209
rect 0 2138 800 2168
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2143 4229 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 15770 2208 16090 2209
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16090 2208
rect 15770 2143 16090 2144
rect 1761 2138 1827 2141
rect 0 2136 1827 2138
rect 0 2080 1766 2136
rect 1822 2080 1827 2136
rect 0 2078 1827 2080
rect 0 2048 800 2078
rect 1761 2075 1827 2078
rect 17493 2138 17559 2141
rect 19200 2138 20000 2168
rect 17493 2136 20000 2138
rect 17493 2080 17498 2136
rect 17554 2080 20000 2136
rect 17493 2078 20000 2080
rect 17493 2075 17559 2078
rect 19200 2048 20000 2078
rect 0 1866 800 1896
rect 2313 1866 2379 1869
rect 0 1864 2379 1866
rect 0 1808 2318 1864
rect 2374 1808 2379 1864
rect 0 1806 2379 1808
rect 0 1776 800 1806
rect 2313 1803 2379 1806
rect 18321 1730 18387 1733
rect 19200 1730 20000 1760
rect 18321 1728 20000 1730
rect 18321 1672 18326 1728
rect 18382 1672 20000 1728
rect 18321 1670 20000 1672
rect 18321 1667 18387 1670
rect 19200 1640 20000 1670
rect 0 1458 800 1488
rect 3693 1458 3759 1461
rect 0 1456 3759 1458
rect 0 1400 3698 1456
rect 3754 1400 3759 1456
rect 0 1398 3759 1400
rect 0 1368 800 1398
rect 3693 1395 3759 1398
rect 18597 1322 18663 1325
rect 19200 1322 20000 1352
rect 18597 1320 20000 1322
rect 18597 1264 18602 1320
rect 18658 1264 20000 1320
rect 18597 1262 20000 1264
rect 18597 1259 18663 1262
rect 19200 1232 20000 1262
rect 0 1186 800 1216
rect 3049 1186 3115 1189
rect 0 1184 3115 1186
rect 0 1128 3054 1184
rect 3110 1128 3115 1184
rect 0 1126 3115 1128
rect 0 1096 800 1126
rect 3049 1123 3115 1126
rect 17861 914 17927 917
rect 19200 914 20000 944
rect 17861 912 20000 914
rect 17861 856 17866 912
rect 17922 856 20000 912
rect 17861 854 20000 856
rect 17861 851 17927 854
rect 19200 824 20000 854
rect 0 778 800 808
rect 1669 778 1735 781
rect 0 776 1735 778
rect 0 720 1674 776
rect 1730 720 1735 776
rect 0 718 1735 720
rect 0 688 800 718
rect 1669 715 1735 718
rect 0 506 800 536
rect 2681 506 2747 509
rect 0 504 2747 506
rect 0 448 2686 504
rect 2742 448 2747 504
rect 0 446 2747 448
rect 0 416 800 446
rect 2681 443 2747 446
rect 15193 506 15259 509
rect 19200 506 20000 536
rect 15193 504 20000 506
rect 15193 448 15198 504
rect 15254 448 20000 504
rect 15193 446 20000 448
rect 15193 443 15259 446
rect 19200 416 20000 446
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
rect 15285 234 15351 237
rect 19200 234 20000 264
rect 15285 232 20000 234
rect 15285 176 15290 232
rect 15346 176 20000 232
rect 15285 174 20000 176
rect 15285 171 15351 174
rect 19200 144 20000 174
<< via3 >>
rect 6882 14716 6946 14720
rect 6882 14660 6886 14716
rect 6886 14660 6942 14716
rect 6942 14660 6946 14716
rect 6882 14656 6946 14660
rect 6962 14716 7026 14720
rect 6962 14660 6966 14716
rect 6966 14660 7022 14716
rect 7022 14660 7026 14716
rect 6962 14656 7026 14660
rect 7042 14716 7106 14720
rect 7042 14660 7046 14716
rect 7046 14660 7102 14716
rect 7102 14660 7106 14716
rect 7042 14656 7106 14660
rect 7122 14716 7186 14720
rect 7122 14660 7126 14716
rect 7126 14660 7182 14716
rect 7182 14660 7186 14716
rect 7122 14656 7186 14660
rect 12813 14716 12877 14720
rect 12813 14660 12817 14716
rect 12817 14660 12873 14716
rect 12873 14660 12877 14716
rect 12813 14656 12877 14660
rect 12893 14716 12957 14720
rect 12893 14660 12897 14716
rect 12897 14660 12953 14716
rect 12953 14660 12957 14716
rect 12893 14656 12957 14660
rect 12973 14716 13037 14720
rect 12973 14660 12977 14716
rect 12977 14660 13033 14716
rect 13033 14660 13037 14716
rect 12973 14656 13037 14660
rect 13053 14716 13117 14720
rect 13053 14660 13057 14716
rect 13057 14660 13113 14716
rect 13113 14660 13117 14716
rect 13053 14656 13117 14660
rect 3917 14172 3981 14176
rect 3917 14116 3921 14172
rect 3921 14116 3977 14172
rect 3977 14116 3981 14172
rect 3917 14112 3981 14116
rect 3997 14172 4061 14176
rect 3997 14116 4001 14172
rect 4001 14116 4057 14172
rect 4057 14116 4061 14172
rect 3997 14112 4061 14116
rect 4077 14172 4141 14176
rect 4077 14116 4081 14172
rect 4081 14116 4137 14172
rect 4137 14116 4141 14172
rect 4077 14112 4141 14116
rect 4157 14172 4221 14176
rect 4157 14116 4161 14172
rect 4161 14116 4217 14172
rect 4217 14116 4221 14172
rect 4157 14112 4221 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 15778 14172 15842 14176
rect 15778 14116 15782 14172
rect 15782 14116 15838 14172
rect 15838 14116 15842 14172
rect 15778 14112 15842 14116
rect 15858 14172 15922 14176
rect 15858 14116 15862 14172
rect 15862 14116 15918 14172
rect 15918 14116 15922 14172
rect 15858 14112 15922 14116
rect 15938 14172 16002 14176
rect 15938 14116 15942 14172
rect 15942 14116 15998 14172
rect 15998 14116 16002 14172
rect 15938 14112 16002 14116
rect 16018 14172 16082 14176
rect 16018 14116 16022 14172
rect 16022 14116 16078 14172
rect 16078 14116 16082 14172
rect 16018 14112 16082 14116
rect 6882 13628 6946 13632
rect 6882 13572 6886 13628
rect 6886 13572 6942 13628
rect 6942 13572 6946 13628
rect 6882 13568 6946 13572
rect 6962 13628 7026 13632
rect 6962 13572 6966 13628
rect 6966 13572 7022 13628
rect 7022 13572 7026 13628
rect 6962 13568 7026 13572
rect 7042 13628 7106 13632
rect 7042 13572 7046 13628
rect 7046 13572 7102 13628
rect 7102 13572 7106 13628
rect 7042 13568 7106 13572
rect 7122 13628 7186 13632
rect 7122 13572 7126 13628
rect 7126 13572 7182 13628
rect 7182 13572 7186 13628
rect 7122 13568 7186 13572
rect 12813 13628 12877 13632
rect 12813 13572 12817 13628
rect 12817 13572 12873 13628
rect 12873 13572 12877 13628
rect 12813 13568 12877 13572
rect 12893 13628 12957 13632
rect 12893 13572 12897 13628
rect 12897 13572 12953 13628
rect 12953 13572 12957 13628
rect 12893 13568 12957 13572
rect 12973 13628 13037 13632
rect 12973 13572 12977 13628
rect 12977 13572 13033 13628
rect 13033 13572 13037 13628
rect 12973 13568 13037 13572
rect 13053 13628 13117 13632
rect 13053 13572 13057 13628
rect 13057 13572 13113 13628
rect 13113 13572 13117 13628
rect 13053 13568 13117 13572
rect 3917 13084 3981 13088
rect 3917 13028 3921 13084
rect 3921 13028 3977 13084
rect 3977 13028 3981 13084
rect 3917 13024 3981 13028
rect 3997 13084 4061 13088
rect 3997 13028 4001 13084
rect 4001 13028 4057 13084
rect 4057 13028 4061 13084
rect 3997 13024 4061 13028
rect 4077 13084 4141 13088
rect 4077 13028 4081 13084
rect 4081 13028 4137 13084
rect 4137 13028 4141 13084
rect 4077 13024 4141 13028
rect 4157 13084 4221 13088
rect 4157 13028 4161 13084
rect 4161 13028 4217 13084
rect 4217 13028 4221 13084
rect 4157 13024 4221 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 15778 13084 15842 13088
rect 15778 13028 15782 13084
rect 15782 13028 15838 13084
rect 15838 13028 15842 13084
rect 15778 13024 15842 13028
rect 15858 13084 15922 13088
rect 15858 13028 15862 13084
rect 15862 13028 15918 13084
rect 15918 13028 15922 13084
rect 15858 13024 15922 13028
rect 15938 13084 16002 13088
rect 15938 13028 15942 13084
rect 15942 13028 15998 13084
rect 15998 13028 16002 13084
rect 15938 13024 16002 13028
rect 16018 13084 16082 13088
rect 16018 13028 16022 13084
rect 16022 13028 16078 13084
rect 16078 13028 16082 13084
rect 16018 13024 16082 13028
rect 6882 12540 6946 12544
rect 6882 12484 6886 12540
rect 6886 12484 6942 12540
rect 6942 12484 6946 12540
rect 6882 12480 6946 12484
rect 6962 12540 7026 12544
rect 6962 12484 6966 12540
rect 6966 12484 7022 12540
rect 7022 12484 7026 12540
rect 6962 12480 7026 12484
rect 7042 12540 7106 12544
rect 7042 12484 7046 12540
rect 7046 12484 7102 12540
rect 7102 12484 7106 12540
rect 7042 12480 7106 12484
rect 7122 12540 7186 12544
rect 7122 12484 7126 12540
rect 7126 12484 7182 12540
rect 7182 12484 7186 12540
rect 7122 12480 7186 12484
rect 12813 12540 12877 12544
rect 12813 12484 12817 12540
rect 12817 12484 12873 12540
rect 12873 12484 12877 12540
rect 12813 12480 12877 12484
rect 12893 12540 12957 12544
rect 12893 12484 12897 12540
rect 12897 12484 12953 12540
rect 12953 12484 12957 12540
rect 12893 12480 12957 12484
rect 12973 12540 13037 12544
rect 12973 12484 12977 12540
rect 12977 12484 13033 12540
rect 13033 12484 13037 12540
rect 12973 12480 13037 12484
rect 13053 12540 13117 12544
rect 13053 12484 13057 12540
rect 13057 12484 13113 12540
rect 13113 12484 13117 12540
rect 13053 12480 13117 12484
rect 3917 11996 3981 12000
rect 3917 11940 3921 11996
rect 3921 11940 3977 11996
rect 3977 11940 3981 11996
rect 3917 11936 3981 11940
rect 3997 11996 4061 12000
rect 3997 11940 4001 11996
rect 4001 11940 4057 11996
rect 4057 11940 4061 11996
rect 3997 11936 4061 11940
rect 4077 11996 4141 12000
rect 4077 11940 4081 11996
rect 4081 11940 4137 11996
rect 4137 11940 4141 11996
rect 4077 11936 4141 11940
rect 4157 11996 4221 12000
rect 4157 11940 4161 11996
rect 4161 11940 4217 11996
rect 4217 11940 4221 11996
rect 4157 11936 4221 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 15778 11996 15842 12000
rect 15778 11940 15782 11996
rect 15782 11940 15838 11996
rect 15838 11940 15842 11996
rect 15778 11936 15842 11940
rect 15858 11996 15922 12000
rect 15858 11940 15862 11996
rect 15862 11940 15918 11996
rect 15918 11940 15922 11996
rect 15858 11936 15922 11940
rect 15938 11996 16002 12000
rect 15938 11940 15942 11996
rect 15942 11940 15998 11996
rect 15998 11940 16002 11996
rect 15938 11936 16002 11940
rect 16018 11996 16082 12000
rect 16018 11940 16022 11996
rect 16022 11940 16078 11996
rect 16078 11940 16082 11996
rect 16018 11936 16082 11940
rect 6882 11452 6946 11456
rect 6882 11396 6886 11452
rect 6886 11396 6942 11452
rect 6942 11396 6946 11452
rect 6882 11392 6946 11396
rect 6962 11452 7026 11456
rect 6962 11396 6966 11452
rect 6966 11396 7022 11452
rect 7022 11396 7026 11452
rect 6962 11392 7026 11396
rect 7042 11452 7106 11456
rect 7042 11396 7046 11452
rect 7046 11396 7102 11452
rect 7102 11396 7106 11452
rect 7042 11392 7106 11396
rect 7122 11452 7186 11456
rect 7122 11396 7126 11452
rect 7126 11396 7182 11452
rect 7182 11396 7186 11452
rect 7122 11392 7186 11396
rect 12813 11452 12877 11456
rect 12813 11396 12817 11452
rect 12817 11396 12873 11452
rect 12873 11396 12877 11452
rect 12813 11392 12877 11396
rect 12893 11452 12957 11456
rect 12893 11396 12897 11452
rect 12897 11396 12953 11452
rect 12953 11396 12957 11452
rect 12893 11392 12957 11396
rect 12973 11452 13037 11456
rect 12973 11396 12977 11452
rect 12977 11396 13033 11452
rect 13033 11396 13037 11452
rect 12973 11392 13037 11396
rect 13053 11452 13117 11456
rect 13053 11396 13057 11452
rect 13057 11396 13113 11452
rect 13113 11396 13117 11452
rect 13053 11392 13117 11396
rect 3917 10908 3981 10912
rect 3917 10852 3921 10908
rect 3921 10852 3977 10908
rect 3977 10852 3981 10908
rect 3917 10848 3981 10852
rect 3997 10908 4061 10912
rect 3997 10852 4001 10908
rect 4001 10852 4057 10908
rect 4057 10852 4061 10908
rect 3997 10848 4061 10852
rect 4077 10908 4141 10912
rect 4077 10852 4081 10908
rect 4081 10852 4137 10908
rect 4137 10852 4141 10908
rect 4077 10848 4141 10852
rect 4157 10908 4221 10912
rect 4157 10852 4161 10908
rect 4161 10852 4217 10908
rect 4217 10852 4221 10908
rect 4157 10848 4221 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 15778 10908 15842 10912
rect 15778 10852 15782 10908
rect 15782 10852 15838 10908
rect 15838 10852 15842 10908
rect 15778 10848 15842 10852
rect 15858 10908 15922 10912
rect 15858 10852 15862 10908
rect 15862 10852 15918 10908
rect 15918 10852 15922 10908
rect 15858 10848 15922 10852
rect 15938 10908 16002 10912
rect 15938 10852 15942 10908
rect 15942 10852 15998 10908
rect 15998 10852 16002 10908
rect 15938 10848 16002 10852
rect 16018 10908 16082 10912
rect 16018 10852 16022 10908
rect 16022 10852 16078 10908
rect 16078 10852 16082 10908
rect 16018 10848 16082 10852
rect 6882 10364 6946 10368
rect 6882 10308 6886 10364
rect 6886 10308 6942 10364
rect 6942 10308 6946 10364
rect 6882 10304 6946 10308
rect 6962 10364 7026 10368
rect 6962 10308 6966 10364
rect 6966 10308 7022 10364
rect 7022 10308 7026 10364
rect 6962 10304 7026 10308
rect 7042 10364 7106 10368
rect 7042 10308 7046 10364
rect 7046 10308 7102 10364
rect 7102 10308 7106 10364
rect 7042 10304 7106 10308
rect 7122 10364 7186 10368
rect 7122 10308 7126 10364
rect 7126 10308 7182 10364
rect 7182 10308 7186 10364
rect 7122 10304 7186 10308
rect 12813 10364 12877 10368
rect 12813 10308 12817 10364
rect 12817 10308 12873 10364
rect 12873 10308 12877 10364
rect 12813 10304 12877 10308
rect 12893 10364 12957 10368
rect 12893 10308 12897 10364
rect 12897 10308 12953 10364
rect 12953 10308 12957 10364
rect 12893 10304 12957 10308
rect 12973 10364 13037 10368
rect 12973 10308 12977 10364
rect 12977 10308 13033 10364
rect 13033 10308 13037 10364
rect 12973 10304 13037 10308
rect 13053 10364 13117 10368
rect 13053 10308 13057 10364
rect 13057 10308 13113 10364
rect 13113 10308 13117 10364
rect 13053 10304 13117 10308
rect 12388 9828 12452 9892
rect 3917 9820 3981 9824
rect 3917 9764 3921 9820
rect 3921 9764 3977 9820
rect 3977 9764 3981 9820
rect 3917 9760 3981 9764
rect 3997 9820 4061 9824
rect 3997 9764 4001 9820
rect 4001 9764 4057 9820
rect 4057 9764 4061 9820
rect 3997 9760 4061 9764
rect 4077 9820 4141 9824
rect 4077 9764 4081 9820
rect 4081 9764 4137 9820
rect 4137 9764 4141 9820
rect 4077 9760 4141 9764
rect 4157 9820 4221 9824
rect 4157 9764 4161 9820
rect 4161 9764 4217 9820
rect 4217 9764 4221 9820
rect 4157 9760 4221 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 15778 9820 15842 9824
rect 15778 9764 15782 9820
rect 15782 9764 15838 9820
rect 15838 9764 15842 9820
rect 15778 9760 15842 9764
rect 15858 9820 15922 9824
rect 15858 9764 15862 9820
rect 15862 9764 15918 9820
rect 15918 9764 15922 9820
rect 15858 9760 15922 9764
rect 15938 9820 16002 9824
rect 15938 9764 15942 9820
rect 15942 9764 15998 9820
rect 15998 9764 16002 9820
rect 15938 9760 16002 9764
rect 16018 9820 16082 9824
rect 16018 9764 16022 9820
rect 16022 9764 16078 9820
rect 16078 9764 16082 9820
rect 16018 9760 16082 9764
rect 6882 9276 6946 9280
rect 6882 9220 6886 9276
rect 6886 9220 6942 9276
rect 6942 9220 6946 9276
rect 6882 9216 6946 9220
rect 6962 9276 7026 9280
rect 6962 9220 6966 9276
rect 6966 9220 7022 9276
rect 7022 9220 7026 9276
rect 6962 9216 7026 9220
rect 7042 9276 7106 9280
rect 7042 9220 7046 9276
rect 7046 9220 7102 9276
rect 7102 9220 7106 9276
rect 7042 9216 7106 9220
rect 7122 9276 7186 9280
rect 7122 9220 7126 9276
rect 7126 9220 7182 9276
rect 7182 9220 7186 9276
rect 7122 9216 7186 9220
rect 12813 9276 12877 9280
rect 12813 9220 12817 9276
rect 12817 9220 12873 9276
rect 12873 9220 12877 9276
rect 12813 9216 12877 9220
rect 12893 9276 12957 9280
rect 12893 9220 12897 9276
rect 12897 9220 12953 9276
rect 12953 9220 12957 9276
rect 12893 9216 12957 9220
rect 12973 9276 13037 9280
rect 12973 9220 12977 9276
rect 12977 9220 13033 9276
rect 13033 9220 13037 9276
rect 12973 9216 13037 9220
rect 13053 9276 13117 9280
rect 13053 9220 13057 9276
rect 13057 9220 13113 9276
rect 13113 9220 13117 9276
rect 13053 9216 13117 9220
rect 12388 9012 12452 9076
rect 13492 9012 13556 9076
rect 3917 8732 3981 8736
rect 3917 8676 3921 8732
rect 3921 8676 3977 8732
rect 3977 8676 3981 8732
rect 3917 8672 3981 8676
rect 3997 8732 4061 8736
rect 3997 8676 4001 8732
rect 4001 8676 4057 8732
rect 4057 8676 4061 8732
rect 3997 8672 4061 8676
rect 4077 8732 4141 8736
rect 4077 8676 4081 8732
rect 4081 8676 4137 8732
rect 4137 8676 4141 8732
rect 4077 8672 4141 8676
rect 4157 8732 4221 8736
rect 4157 8676 4161 8732
rect 4161 8676 4217 8732
rect 4217 8676 4221 8732
rect 4157 8672 4221 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 15778 8732 15842 8736
rect 15778 8676 15782 8732
rect 15782 8676 15838 8732
rect 15838 8676 15842 8732
rect 15778 8672 15842 8676
rect 15858 8732 15922 8736
rect 15858 8676 15862 8732
rect 15862 8676 15918 8732
rect 15918 8676 15922 8732
rect 15858 8672 15922 8676
rect 15938 8732 16002 8736
rect 15938 8676 15942 8732
rect 15942 8676 15998 8732
rect 15998 8676 16002 8732
rect 15938 8672 16002 8676
rect 16018 8732 16082 8736
rect 16018 8676 16022 8732
rect 16022 8676 16078 8732
rect 16078 8676 16082 8732
rect 16018 8672 16082 8676
rect 13308 8468 13372 8532
rect 6882 8188 6946 8192
rect 6882 8132 6886 8188
rect 6886 8132 6942 8188
rect 6942 8132 6946 8188
rect 6882 8128 6946 8132
rect 6962 8188 7026 8192
rect 6962 8132 6966 8188
rect 6966 8132 7022 8188
rect 7022 8132 7026 8188
rect 6962 8128 7026 8132
rect 7042 8188 7106 8192
rect 7042 8132 7046 8188
rect 7046 8132 7102 8188
rect 7102 8132 7106 8188
rect 7042 8128 7106 8132
rect 7122 8188 7186 8192
rect 7122 8132 7126 8188
rect 7126 8132 7182 8188
rect 7182 8132 7186 8188
rect 7122 8128 7186 8132
rect 12813 8188 12877 8192
rect 12813 8132 12817 8188
rect 12817 8132 12873 8188
rect 12873 8132 12877 8188
rect 12813 8128 12877 8132
rect 12893 8188 12957 8192
rect 12893 8132 12897 8188
rect 12897 8132 12953 8188
rect 12953 8132 12957 8188
rect 12893 8128 12957 8132
rect 12973 8188 13037 8192
rect 12973 8132 12977 8188
rect 12977 8132 13033 8188
rect 13033 8132 13037 8188
rect 12973 8128 13037 8132
rect 13053 8188 13117 8192
rect 13053 8132 13057 8188
rect 13057 8132 13113 8188
rect 13113 8132 13117 8188
rect 13053 8128 13117 8132
rect 3372 7924 3436 7988
rect 3917 7644 3981 7648
rect 3917 7588 3921 7644
rect 3921 7588 3977 7644
rect 3977 7588 3981 7644
rect 3917 7584 3981 7588
rect 3997 7644 4061 7648
rect 3997 7588 4001 7644
rect 4001 7588 4057 7644
rect 4057 7588 4061 7644
rect 3997 7584 4061 7588
rect 4077 7644 4141 7648
rect 4077 7588 4081 7644
rect 4081 7588 4137 7644
rect 4137 7588 4141 7644
rect 4077 7584 4141 7588
rect 4157 7644 4221 7648
rect 4157 7588 4161 7644
rect 4161 7588 4217 7644
rect 4217 7588 4221 7644
rect 4157 7584 4221 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 15778 7644 15842 7648
rect 15778 7588 15782 7644
rect 15782 7588 15838 7644
rect 15838 7588 15842 7644
rect 15778 7584 15842 7588
rect 15858 7644 15922 7648
rect 15858 7588 15862 7644
rect 15862 7588 15918 7644
rect 15918 7588 15922 7644
rect 15858 7584 15922 7588
rect 15938 7644 16002 7648
rect 15938 7588 15942 7644
rect 15942 7588 15998 7644
rect 15998 7588 16002 7644
rect 15938 7584 16002 7588
rect 16018 7644 16082 7648
rect 16018 7588 16022 7644
rect 16022 7588 16078 7644
rect 16078 7588 16082 7644
rect 16018 7584 16082 7588
rect 11468 7244 11532 7308
rect 12572 7108 12636 7172
rect 6882 7100 6946 7104
rect 6882 7044 6886 7100
rect 6886 7044 6942 7100
rect 6942 7044 6946 7100
rect 6882 7040 6946 7044
rect 6962 7100 7026 7104
rect 6962 7044 6966 7100
rect 6966 7044 7022 7100
rect 7022 7044 7026 7100
rect 6962 7040 7026 7044
rect 7042 7100 7106 7104
rect 7042 7044 7046 7100
rect 7046 7044 7102 7100
rect 7102 7044 7106 7100
rect 7042 7040 7106 7044
rect 7122 7100 7186 7104
rect 7122 7044 7126 7100
rect 7126 7044 7182 7100
rect 7182 7044 7186 7100
rect 7122 7040 7186 7044
rect 12813 7100 12877 7104
rect 12813 7044 12817 7100
rect 12817 7044 12873 7100
rect 12873 7044 12877 7100
rect 12813 7040 12877 7044
rect 12893 7100 12957 7104
rect 12893 7044 12897 7100
rect 12897 7044 12953 7100
rect 12953 7044 12957 7100
rect 12893 7040 12957 7044
rect 12973 7100 13037 7104
rect 12973 7044 12977 7100
rect 12977 7044 13033 7100
rect 13033 7044 13037 7100
rect 12973 7040 13037 7044
rect 13053 7100 13117 7104
rect 13053 7044 13057 7100
rect 13057 7044 13113 7100
rect 13113 7044 13117 7100
rect 13053 7040 13117 7044
rect 3917 6556 3981 6560
rect 3917 6500 3921 6556
rect 3921 6500 3977 6556
rect 3977 6500 3981 6556
rect 3917 6496 3981 6500
rect 3997 6556 4061 6560
rect 3997 6500 4001 6556
rect 4001 6500 4057 6556
rect 4057 6500 4061 6556
rect 3997 6496 4061 6500
rect 4077 6556 4141 6560
rect 4077 6500 4081 6556
rect 4081 6500 4137 6556
rect 4137 6500 4141 6556
rect 4077 6496 4141 6500
rect 4157 6556 4221 6560
rect 4157 6500 4161 6556
rect 4161 6500 4217 6556
rect 4217 6500 4221 6556
rect 4157 6496 4221 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 15778 6556 15842 6560
rect 15778 6500 15782 6556
rect 15782 6500 15838 6556
rect 15838 6500 15842 6556
rect 15778 6496 15842 6500
rect 15858 6556 15922 6560
rect 15858 6500 15862 6556
rect 15862 6500 15918 6556
rect 15918 6500 15922 6556
rect 15858 6496 15922 6500
rect 15938 6556 16002 6560
rect 15938 6500 15942 6556
rect 15942 6500 15998 6556
rect 15998 6500 16002 6556
rect 15938 6496 16002 6500
rect 16018 6556 16082 6560
rect 16018 6500 16022 6556
rect 16022 6500 16078 6556
rect 16078 6500 16082 6556
rect 16018 6496 16082 6500
rect 3372 6156 3436 6220
rect 6882 6012 6946 6016
rect 6882 5956 6886 6012
rect 6886 5956 6942 6012
rect 6942 5956 6946 6012
rect 6882 5952 6946 5956
rect 6962 6012 7026 6016
rect 6962 5956 6966 6012
rect 6966 5956 7022 6012
rect 7022 5956 7026 6012
rect 6962 5952 7026 5956
rect 7042 6012 7106 6016
rect 7042 5956 7046 6012
rect 7046 5956 7102 6012
rect 7102 5956 7106 6012
rect 7042 5952 7106 5956
rect 7122 6012 7186 6016
rect 7122 5956 7126 6012
rect 7126 5956 7182 6012
rect 7182 5956 7186 6012
rect 7122 5952 7186 5956
rect 12813 6012 12877 6016
rect 12813 5956 12817 6012
rect 12817 5956 12873 6012
rect 12873 5956 12877 6012
rect 12813 5952 12877 5956
rect 12893 6012 12957 6016
rect 12893 5956 12897 6012
rect 12897 5956 12953 6012
rect 12953 5956 12957 6012
rect 12893 5952 12957 5956
rect 12973 6012 13037 6016
rect 12973 5956 12977 6012
rect 12977 5956 13033 6012
rect 13033 5956 13037 6012
rect 12973 5952 13037 5956
rect 13053 6012 13117 6016
rect 13053 5956 13057 6012
rect 13057 5956 13113 6012
rect 13113 5956 13117 6012
rect 13053 5952 13117 5956
rect 13492 5944 13556 5948
rect 13492 5888 13542 5944
rect 13542 5888 13556 5944
rect 13492 5884 13556 5888
rect 3372 5748 3436 5812
rect 3917 5468 3981 5472
rect 3917 5412 3921 5468
rect 3921 5412 3977 5468
rect 3977 5412 3981 5468
rect 3917 5408 3981 5412
rect 3997 5468 4061 5472
rect 3997 5412 4001 5468
rect 4001 5412 4057 5468
rect 4057 5412 4061 5468
rect 3997 5408 4061 5412
rect 4077 5468 4141 5472
rect 4077 5412 4081 5468
rect 4081 5412 4137 5468
rect 4137 5412 4141 5468
rect 4077 5408 4141 5412
rect 4157 5468 4221 5472
rect 4157 5412 4161 5468
rect 4161 5412 4217 5468
rect 4217 5412 4221 5468
rect 4157 5408 4221 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 15778 5468 15842 5472
rect 15778 5412 15782 5468
rect 15782 5412 15838 5468
rect 15838 5412 15842 5468
rect 15778 5408 15842 5412
rect 15858 5468 15922 5472
rect 15858 5412 15862 5468
rect 15862 5412 15918 5468
rect 15918 5412 15922 5468
rect 15858 5408 15922 5412
rect 15938 5468 16002 5472
rect 15938 5412 15942 5468
rect 15942 5412 15998 5468
rect 15998 5412 16002 5468
rect 15938 5408 16002 5412
rect 16018 5468 16082 5472
rect 16018 5412 16022 5468
rect 16022 5412 16078 5468
rect 16078 5412 16082 5468
rect 16018 5408 16082 5412
rect 12572 5204 12636 5268
rect 6882 4924 6946 4928
rect 6882 4868 6886 4924
rect 6886 4868 6942 4924
rect 6942 4868 6946 4924
rect 6882 4864 6946 4868
rect 6962 4924 7026 4928
rect 6962 4868 6966 4924
rect 6966 4868 7022 4924
rect 7022 4868 7026 4924
rect 6962 4864 7026 4868
rect 7042 4924 7106 4928
rect 7042 4868 7046 4924
rect 7046 4868 7102 4924
rect 7102 4868 7106 4924
rect 7042 4864 7106 4868
rect 7122 4924 7186 4928
rect 7122 4868 7126 4924
rect 7126 4868 7182 4924
rect 7182 4868 7186 4924
rect 7122 4864 7186 4868
rect 12813 4924 12877 4928
rect 12813 4868 12817 4924
rect 12817 4868 12873 4924
rect 12873 4868 12877 4924
rect 12813 4864 12877 4868
rect 12893 4924 12957 4928
rect 12893 4868 12897 4924
rect 12897 4868 12953 4924
rect 12953 4868 12957 4924
rect 12893 4864 12957 4868
rect 12973 4924 13037 4928
rect 12973 4868 12977 4924
rect 12977 4868 13033 4924
rect 13033 4868 13037 4924
rect 12973 4864 13037 4868
rect 13053 4924 13117 4928
rect 13053 4868 13057 4924
rect 13057 4868 13113 4924
rect 13113 4868 13117 4924
rect 13053 4864 13117 4868
rect 13308 4388 13372 4452
rect 3917 4380 3981 4384
rect 3917 4324 3921 4380
rect 3921 4324 3977 4380
rect 3977 4324 3981 4380
rect 3917 4320 3981 4324
rect 3997 4380 4061 4384
rect 3997 4324 4001 4380
rect 4001 4324 4057 4380
rect 4057 4324 4061 4380
rect 3997 4320 4061 4324
rect 4077 4380 4141 4384
rect 4077 4324 4081 4380
rect 4081 4324 4137 4380
rect 4137 4324 4141 4380
rect 4077 4320 4141 4324
rect 4157 4380 4221 4384
rect 4157 4324 4161 4380
rect 4161 4324 4217 4380
rect 4217 4324 4221 4380
rect 4157 4320 4221 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 15778 4380 15842 4384
rect 15778 4324 15782 4380
rect 15782 4324 15838 4380
rect 15838 4324 15842 4380
rect 15778 4320 15842 4324
rect 15858 4380 15922 4384
rect 15858 4324 15862 4380
rect 15862 4324 15918 4380
rect 15918 4324 15922 4380
rect 15858 4320 15922 4324
rect 15938 4380 16002 4384
rect 15938 4324 15942 4380
rect 15942 4324 15998 4380
rect 15998 4324 16002 4380
rect 15938 4320 16002 4324
rect 16018 4380 16082 4384
rect 16018 4324 16022 4380
rect 16022 4324 16078 4380
rect 16078 4324 16082 4380
rect 16018 4320 16082 4324
rect 11468 3844 11532 3908
rect 6882 3836 6946 3840
rect 6882 3780 6886 3836
rect 6886 3780 6942 3836
rect 6942 3780 6946 3836
rect 6882 3776 6946 3780
rect 6962 3836 7026 3840
rect 6962 3780 6966 3836
rect 6966 3780 7022 3836
rect 7022 3780 7026 3836
rect 6962 3776 7026 3780
rect 7042 3836 7106 3840
rect 7042 3780 7046 3836
rect 7046 3780 7102 3836
rect 7102 3780 7106 3836
rect 7042 3776 7106 3780
rect 7122 3836 7186 3840
rect 7122 3780 7126 3836
rect 7126 3780 7182 3836
rect 7182 3780 7186 3836
rect 7122 3776 7186 3780
rect 12813 3836 12877 3840
rect 12813 3780 12817 3836
rect 12817 3780 12873 3836
rect 12873 3780 12877 3836
rect 12813 3776 12877 3780
rect 12893 3836 12957 3840
rect 12893 3780 12897 3836
rect 12897 3780 12953 3836
rect 12953 3780 12957 3836
rect 12893 3776 12957 3780
rect 12973 3836 13037 3840
rect 12973 3780 12977 3836
rect 12977 3780 13033 3836
rect 13033 3780 13037 3836
rect 12973 3776 13037 3780
rect 13053 3836 13117 3840
rect 13053 3780 13057 3836
rect 13057 3780 13113 3836
rect 13113 3780 13117 3836
rect 13053 3776 13117 3780
rect 3917 3292 3981 3296
rect 3917 3236 3921 3292
rect 3921 3236 3977 3292
rect 3977 3236 3981 3292
rect 3917 3232 3981 3236
rect 3997 3292 4061 3296
rect 3997 3236 4001 3292
rect 4001 3236 4057 3292
rect 4057 3236 4061 3292
rect 3997 3232 4061 3236
rect 4077 3292 4141 3296
rect 4077 3236 4081 3292
rect 4081 3236 4137 3292
rect 4137 3236 4141 3292
rect 4077 3232 4141 3236
rect 4157 3292 4221 3296
rect 4157 3236 4161 3292
rect 4161 3236 4217 3292
rect 4217 3236 4221 3292
rect 4157 3232 4221 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 15778 3292 15842 3296
rect 15778 3236 15782 3292
rect 15782 3236 15838 3292
rect 15838 3236 15842 3292
rect 15778 3232 15842 3236
rect 15858 3292 15922 3296
rect 15858 3236 15862 3292
rect 15862 3236 15918 3292
rect 15918 3236 15922 3292
rect 15858 3232 15922 3236
rect 15938 3292 16002 3296
rect 15938 3236 15942 3292
rect 15942 3236 15998 3292
rect 15998 3236 16002 3292
rect 15938 3232 16002 3236
rect 16018 3292 16082 3296
rect 16018 3236 16022 3292
rect 16022 3236 16078 3292
rect 16078 3236 16082 3292
rect 16018 3232 16082 3236
rect 6882 2748 6946 2752
rect 6882 2692 6886 2748
rect 6886 2692 6942 2748
rect 6942 2692 6946 2748
rect 6882 2688 6946 2692
rect 6962 2748 7026 2752
rect 6962 2692 6966 2748
rect 6966 2692 7022 2748
rect 7022 2692 7026 2748
rect 6962 2688 7026 2692
rect 7042 2748 7106 2752
rect 7042 2692 7046 2748
rect 7046 2692 7102 2748
rect 7102 2692 7106 2748
rect 7042 2688 7106 2692
rect 7122 2748 7186 2752
rect 7122 2692 7126 2748
rect 7126 2692 7182 2748
rect 7182 2692 7186 2748
rect 7122 2688 7186 2692
rect 12813 2748 12877 2752
rect 12813 2692 12817 2748
rect 12817 2692 12873 2748
rect 12873 2692 12877 2748
rect 12813 2688 12877 2692
rect 12893 2748 12957 2752
rect 12893 2692 12897 2748
rect 12897 2692 12953 2748
rect 12953 2692 12957 2748
rect 12893 2688 12957 2692
rect 12973 2748 13037 2752
rect 12973 2692 12977 2748
rect 12977 2692 13033 2748
rect 13033 2692 13037 2748
rect 12973 2688 13037 2692
rect 13053 2748 13117 2752
rect 13053 2692 13057 2748
rect 13057 2692 13113 2748
rect 13113 2692 13117 2748
rect 13053 2688 13117 2692
rect 3917 2204 3981 2208
rect 3917 2148 3921 2204
rect 3921 2148 3977 2204
rect 3977 2148 3981 2204
rect 3917 2144 3981 2148
rect 3997 2204 4061 2208
rect 3997 2148 4001 2204
rect 4001 2148 4057 2204
rect 4057 2148 4061 2204
rect 3997 2144 4061 2148
rect 4077 2204 4141 2208
rect 4077 2148 4081 2204
rect 4081 2148 4137 2204
rect 4137 2148 4141 2204
rect 4077 2144 4141 2148
rect 4157 2204 4221 2208
rect 4157 2148 4161 2204
rect 4161 2148 4217 2204
rect 4217 2148 4221 2204
rect 4157 2144 4221 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 15778 2204 15842 2208
rect 15778 2148 15782 2204
rect 15782 2148 15838 2204
rect 15838 2148 15842 2204
rect 15778 2144 15842 2148
rect 15858 2204 15922 2208
rect 15858 2148 15862 2204
rect 15862 2148 15918 2204
rect 15918 2148 15922 2204
rect 15858 2144 15922 2148
rect 15938 2204 16002 2208
rect 15938 2148 15942 2204
rect 15942 2148 15998 2204
rect 15998 2148 16002 2204
rect 15938 2144 16002 2148
rect 16018 2204 16082 2208
rect 16018 2148 16022 2204
rect 16022 2148 16078 2204
rect 16078 2148 16082 2204
rect 16018 2144 16082 2148
<< metal4 >>
rect 3909 14176 4229 14736
rect 3909 14112 3917 14176
rect 3981 14112 3997 14176
rect 4061 14112 4077 14176
rect 4141 14112 4157 14176
rect 4221 14112 4229 14176
rect 3909 13088 4229 14112
rect 3909 13024 3917 13088
rect 3981 13024 3997 13088
rect 4061 13024 4077 13088
rect 4141 13024 4157 13088
rect 4221 13024 4229 13088
rect 3909 12000 4229 13024
rect 3909 11936 3917 12000
rect 3981 11936 3997 12000
rect 4061 11936 4077 12000
rect 4141 11936 4157 12000
rect 4221 11936 4229 12000
rect 3909 10912 4229 11936
rect 3909 10848 3917 10912
rect 3981 10848 3997 10912
rect 4061 10848 4077 10912
rect 4141 10848 4157 10912
rect 4221 10848 4229 10912
rect 3909 9824 4229 10848
rect 3909 9760 3917 9824
rect 3981 9760 3997 9824
rect 4061 9760 4077 9824
rect 4141 9760 4157 9824
rect 4221 9760 4229 9824
rect 3909 8736 4229 9760
rect 3909 8672 3917 8736
rect 3981 8672 3997 8736
rect 4061 8672 4077 8736
rect 4141 8672 4157 8736
rect 4221 8672 4229 8736
rect 3371 7988 3437 7989
rect 3371 7924 3372 7988
rect 3436 7924 3437 7988
rect 3371 7923 3437 7924
rect 3374 6221 3434 7923
rect 3909 7648 4229 8672
rect 3909 7584 3917 7648
rect 3981 7584 3997 7648
rect 4061 7584 4077 7648
rect 4141 7584 4157 7648
rect 4221 7584 4229 7648
rect 3909 6560 4229 7584
rect 3909 6496 3917 6560
rect 3981 6496 3997 6560
rect 4061 6496 4077 6560
rect 4141 6496 4157 6560
rect 4221 6496 4229 6560
rect 3371 6220 3437 6221
rect 3371 6156 3372 6220
rect 3436 6156 3437 6220
rect 3371 6155 3437 6156
rect 3374 5813 3434 6155
rect 3371 5812 3437 5813
rect 3371 5748 3372 5812
rect 3436 5748 3437 5812
rect 3371 5747 3437 5748
rect 3909 5472 4229 6496
rect 3909 5408 3917 5472
rect 3981 5408 3997 5472
rect 4061 5408 4077 5472
rect 4141 5408 4157 5472
rect 4221 5408 4229 5472
rect 3909 4384 4229 5408
rect 3909 4320 3917 4384
rect 3981 4320 3997 4384
rect 4061 4320 4077 4384
rect 4141 4320 4157 4384
rect 4221 4320 4229 4384
rect 3909 3296 4229 4320
rect 3909 3232 3917 3296
rect 3981 3232 3997 3296
rect 4061 3232 4077 3296
rect 4141 3232 4157 3296
rect 4221 3232 4229 3296
rect 3909 2208 4229 3232
rect 3909 2144 3917 2208
rect 3981 2144 3997 2208
rect 4061 2144 4077 2208
rect 4141 2144 4157 2208
rect 4221 2144 4229 2208
rect 3909 2128 4229 2144
rect 6874 14720 7195 14736
rect 6874 14656 6882 14720
rect 6946 14656 6962 14720
rect 7026 14656 7042 14720
rect 7106 14656 7122 14720
rect 7186 14656 7195 14720
rect 6874 13632 7195 14656
rect 6874 13568 6882 13632
rect 6946 13568 6962 13632
rect 7026 13568 7042 13632
rect 7106 13568 7122 13632
rect 7186 13568 7195 13632
rect 6874 12544 7195 13568
rect 6874 12480 6882 12544
rect 6946 12480 6962 12544
rect 7026 12480 7042 12544
rect 7106 12480 7122 12544
rect 7186 12480 7195 12544
rect 6874 11456 7195 12480
rect 6874 11392 6882 11456
rect 6946 11392 6962 11456
rect 7026 11392 7042 11456
rect 7106 11392 7122 11456
rect 7186 11392 7195 11456
rect 6874 10368 7195 11392
rect 6874 10304 6882 10368
rect 6946 10304 6962 10368
rect 7026 10304 7042 10368
rect 7106 10304 7122 10368
rect 7186 10304 7195 10368
rect 6874 9280 7195 10304
rect 6874 9216 6882 9280
rect 6946 9216 6962 9280
rect 7026 9216 7042 9280
rect 7106 9216 7122 9280
rect 7186 9216 7195 9280
rect 6874 8192 7195 9216
rect 6874 8128 6882 8192
rect 6946 8128 6962 8192
rect 7026 8128 7042 8192
rect 7106 8128 7122 8192
rect 7186 8128 7195 8192
rect 6874 7104 7195 8128
rect 6874 7040 6882 7104
rect 6946 7040 6962 7104
rect 7026 7040 7042 7104
rect 7106 7040 7122 7104
rect 7186 7040 7195 7104
rect 6874 6016 7195 7040
rect 6874 5952 6882 6016
rect 6946 5952 6962 6016
rect 7026 5952 7042 6016
rect 7106 5952 7122 6016
rect 7186 5952 7195 6016
rect 6874 4928 7195 5952
rect 6874 4864 6882 4928
rect 6946 4864 6962 4928
rect 7026 4864 7042 4928
rect 7106 4864 7122 4928
rect 7186 4864 7195 4928
rect 6874 3840 7195 4864
rect 6874 3776 6882 3840
rect 6946 3776 6962 3840
rect 7026 3776 7042 3840
rect 7106 3776 7122 3840
rect 7186 3776 7195 3840
rect 6874 2752 7195 3776
rect 6874 2688 6882 2752
rect 6946 2688 6962 2752
rect 7026 2688 7042 2752
rect 7106 2688 7122 2752
rect 7186 2688 7195 2752
rect 6874 2128 7195 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 12805 14720 13125 14736
rect 12805 14656 12813 14720
rect 12877 14656 12893 14720
rect 12957 14656 12973 14720
rect 13037 14656 13053 14720
rect 13117 14656 13125 14720
rect 12805 13632 13125 14656
rect 12805 13568 12813 13632
rect 12877 13568 12893 13632
rect 12957 13568 12973 13632
rect 13037 13568 13053 13632
rect 13117 13568 13125 13632
rect 12805 12544 13125 13568
rect 12805 12480 12813 12544
rect 12877 12480 12893 12544
rect 12957 12480 12973 12544
rect 13037 12480 13053 12544
rect 13117 12480 13125 12544
rect 12805 11456 13125 12480
rect 12805 11392 12813 11456
rect 12877 11392 12893 11456
rect 12957 11392 12973 11456
rect 13037 11392 13053 11456
rect 13117 11392 13125 11456
rect 12805 10368 13125 11392
rect 12805 10304 12813 10368
rect 12877 10304 12893 10368
rect 12957 10304 12973 10368
rect 13037 10304 13053 10368
rect 13117 10304 13125 10368
rect 12387 9892 12453 9893
rect 12387 9828 12388 9892
rect 12452 9828 12453 9892
rect 12387 9827 12453 9828
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 12390 9077 12450 9827
rect 12805 9280 13125 10304
rect 12805 9216 12813 9280
rect 12877 9216 12893 9280
rect 12957 9216 12973 9280
rect 13037 9216 13053 9280
rect 13117 9216 13125 9280
rect 12387 9076 12453 9077
rect 12387 9012 12388 9076
rect 12452 9012 12453 9076
rect 12387 9011 12453 9012
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 12805 8192 13125 9216
rect 15770 14176 16091 14736
rect 15770 14112 15778 14176
rect 15842 14112 15858 14176
rect 15922 14112 15938 14176
rect 16002 14112 16018 14176
rect 16082 14112 16091 14176
rect 15770 13088 16091 14112
rect 15770 13024 15778 13088
rect 15842 13024 15858 13088
rect 15922 13024 15938 13088
rect 16002 13024 16018 13088
rect 16082 13024 16091 13088
rect 15770 12000 16091 13024
rect 15770 11936 15778 12000
rect 15842 11936 15858 12000
rect 15922 11936 15938 12000
rect 16002 11936 16018 12000
rect 16082 11936 16091 12000
rect 15770 10912 16091 11936
rect 15770 10848 15778 10912
rect 15842 10848 15858 10912
rect 15922 10848 15938 10912
rect 16002 10848 16018 10912
rect 16082 10848 16091 10912
rect 15770 9824 16091 10848
rect 15770 9760 15778 9824
rect 15842 9760 15858 9824
rect 15922 9760 15938 9824
rect 16002 9760 16018 9824
rect 16082 9760 16091 9824
rect 13491 9076 13557 9077
rect 13491 9012 13492 9076
rect 13556 9012 13557 9076
rect 13491 9011 13557 9012
rect 13307 8532 13373 8533
rect 13307 8468 13308 8532
rect 13372 8468 13373 8532
rect 13307 8467 13373 8468
rect 12805 8128 12813 8192
rect 12877 8128 12893 8192
rect 12957 8128 12973 8192
rect 13037 8128 13053 8192
rect 13117 8128 13125 8192
rect 11467 7308 11533 7309
rect 11467 7244 11468 7308
rect 11532 7244 11533 7308
rect 11467 7243 11533 7244
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 11470 3909 11530 7243
rect 12571 7172 12637 7173
rect 12571 7108 12572 7172
rect 12636 7108 12637 7172
rect 12571 7107 12637 7108
rect 12574 5269 12634 7107
rect 12805 7104 13125 8128
rect 12805 7040 12813 7104
rect 12877 7040 12893 7104
rect 12957 7040 12973 7104
rect 13037 7040 13053 7104
rect 13117 7040 13125 7104
rect 12805 6016 13125 7040
rect 12805 5952 12813 6016
rect 12877 5952 12893 6016
rect 12957 5952 12973 6016
rect 13037 5952 13053 6016
rect 13117 5952 13125 6016
rect 12571 5268 12637 5269
rect 12571 5204 12572 5268
rect 12636 5204 12637 5268
rect 12571 5203 12637 5204
rect 12805 4928 13125 5952
rect 12805 4864 12813 4928
rect 12877 4864 12893 4928
rect 12957 4864 12973 4928
rect 13037 4864 13053 4928
rect 13117 4864 13125 4928
rect 11467 3908 11533 3909
rect 11467 3844 11468 3908
rect 11532 3844 11533 3908
rect 11467 3843 11533 3844
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12805 3840 13125 4864
rect 13310 4453 13370 8467
rect 13494 5949 13554 9011
rect 15770 8736 16091 9760
rect 15770 8672 15778 8736
rect 15842 8672 15858 8736
rect 15922 8672 15938 8736
rect 16002 8672 16018 8736
rect 16082 8672 16091 8736
rect 15770 7648 16091 8672
rect 15770 7584 15778 7648
rect 15842 7584 15858 7648
rect 15922 7584 15938 7648
rect 16002 7584 16018 7648
rect 16082 7584 16091 7648
rect 15770 6560 16091 7584
rect 15770 6496 15778 6560
rect 15842 6496 15858 6560
rect 15922 6496 15938 6560
rect 16002 6496 16018 6560
rect 16082 6496 16091 6560
rect 13491 5948 13557 5949
rect 13491 5884 13492 5948
rect 13556 5884 13557 5948
rect 13491 5883 13557 5884
rect 15770 5472 16091 6496
rect 15770 5408 15778 5472
rect 15842 5408 15858 5472
rect 15922 5408 15938 5472
rect 16002 5408 16018 5472
rect 16082 5408 16091 5472
rect 13307 4452 13373 4453
rect 13307 4388 13308 4452
rect 13372 4388 13373 4452
rect 13307 4387 13373 4388
rect 12805 3776 12813 3840
rect 12877 3776 12893 3840
rect 12957 3776 12973 3840
rect 13037 3776 13053 3840
rect 13117 3776 13125 3840
rect 12805 2752 13125 3776
rect 12805 2688 12813 2752
rect 12877 2688 12893 2752
rect 12957 2688 12973 2752
rect 13037 2688 13053 2752
rect 13117 2688 13125 2752
rect 12805 2128 13125 2688
rect 15770 4384 16091 5408
rect 15770 4320 15778 4384
rect 15842 4320 15858 4384
rect 15922 4320 15938 4384
rect 16002 4320 16018 4384
rect 16082 4320 16091 4384
rect 15770 3296 16091 4320
rect 15770 3232 15778 3296
rect 15842 3232 15858 3296
rect 15922 3232 15938 3296
rect 16002 3232 16018 3296
rect 16082 3232 16091 3296
rect 15770 2208 16091 3232
rect 15770 2144 15778 2208
rect 15842 2144 15858 2208
rect 15922 2144 15938 2208
rect 16002 2144 16018 2208
rect 16082 2144 16091 2208
rect 15770 2128 16091 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_2 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1608910539
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _42_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1608910539
transform 1 0 1564 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1932 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1608910539
transform 1 0 2116 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1608910539
transform 1 0 1748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2852 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_E_FTB01
timestamp 1608910539
transform 1 0 2944 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1608910539
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1608910539
transform 1 0 2484 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1608910539
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32
timestamp 1608910539
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1608910539
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4692 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 4140 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 3404 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4232 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1608910539
transform 1 0 3864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1608910539
transform 1 0 3496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 5796 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 5244 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1608910539
transform 1 0 5060 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1608910539
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1608910539
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1608910539
transform 1 0 6348 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1608910539
transform 1 0 6164 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 5980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1608910539
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1608910539
transform 1 0 5888 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 6808 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1608910539
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_68
timestamp 1608910539
transform 1 0 7360 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 7176 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 6992 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 7452 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1608910539
transform 1 0 8188 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1608910539
transform 1 0 8004 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 7452 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 6900 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1608910539
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8832 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1608910539
transform 1 0 9016 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94
timestamp 1608910539
transform 1 0 9752 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 10212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 9844 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1608910539
transform 1 0 9844 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10672 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_1_125
timestamp 1608910539
transform 1 0 12604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 1608910539
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1608910539
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1608910539
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11500 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11408 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14076 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13524 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13984 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 13432 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12696 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_154
timestamp 1608910539
transform 1 0 15272 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_E_FTB01_A
timestamp 1608910539
transform 1 0 15088 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 15180 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1608910539
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1608910539
transform 1 0 15364 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14536 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_162 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 16008 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1608910539
transform 1 0 16192 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 15456 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_170 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 16744 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_N_FTB01_A
timestamp 1608910539
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l4_in_0__S
timestamp 1608910539
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_1_S_FTB01_A
timestamp 1608910539
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1608910539
transform 1 0 17112 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_N_FTB01
timestamp 1608910539
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1608910539
transform 1 0 17296 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1608910539
transform 1 0 18308 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1608910539
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1608910539
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_1_S_FTB01
timestamp 1608910539
transform 1 0 18032 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 18400 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1608910539
transform -1 0 18860 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1608910539
transform -1 0 18860 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1608910539
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1608910539
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_21
timestamp 1608910539
transform 1 0 3036 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1608910539
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 4048 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5520 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1608910539
transform 1 0 8096 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1608910539
transform 1 0 6992 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 8188 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8740 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1608910539
transform 1 0 7268 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1608910539
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 9660 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 11408 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _19_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 11132 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 12880 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_2_156
timestamp 1608910539
transform 1 0 15456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_146
timestamp 1608910539
transform 1 0 14536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 15272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1608910539
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1608910539
transform 1 0 14628 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1608910539
transform 1 0 16376 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1608910539
transform 1 0 15548 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_2_175
timestamp 1608910539
transform 1 0 17204 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1608910539
transform 1 0 17296 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1608910539
transform 1 0 17480 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1608910539
transform 1 0 17664 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1608910539
transform 1 0 18216 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1608910539
transform 1 0 17848 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1608910539
transform -1 0 18860 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1608910539
transform 1 0 1380 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1608910539
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1608910539
transform 1 0 2576 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1608910539
transform 1 0 1472 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1608910539
transform 1 0 2208 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1608910539
transform 1 0 1840 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_29
timestamp 1608910539
transform 1 0 3772 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3588 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 3404 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3864 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1608910539
transform 1 0 4692 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1608910539
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58
timestamp 1608910539
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 6808 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1608910539
transform 1 0 6348 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 8280 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1608910539
transform 1 0 9752 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1608910539
transform 1 0 10120 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_125
timestamp 1608910539
transform 1 0 12604 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1608910539
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10948 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1608910539
transform 1 0 13708 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1608910539
transform 1 0 12880 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_153
timestamp 1608910539
transform 1 0 15180 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14996 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15272 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1608910539
transform 1 0 14536 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_60
timestamp 1608910539
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16744 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1608910539
transform 1 0 17572 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1608910539
transform 1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1608910539
transform 1 0 18400 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1608910539
transform -1 0 18860 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_14
timestamp 1608910539
transform 1 0 2392 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1608910539
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 1472 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1608910539
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 2484 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1608910539
transform 1 0 2024 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1608910539
transform 1 0 1656 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_39
timestamp 1608910539
transform 1 0 4692 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 4324 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 4508 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4784 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_61
timestamp 1608910539
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1608910539
transform 1 0 6532 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1608910539
transform 1 0 6348 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1608910539
transform 1 0 6164 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1608910539
transform 1 0 5980 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4968 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_82
timestamp 1608910539
transform 1 0 8648 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_63
timestamp 1608910539
transform 1 0 6900 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8740 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 7176 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9844 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9660 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 10212 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_62
timestamp 1608910539
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1608910539
transform 1 0 10396 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11224 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1608910539
transform 1 0 12052 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1608910539
transform 1 0 12880 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 13708 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_63
timestamp 1608910539
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 15272 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1608910539
transform 1 0 16744 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1608910539
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16928 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1608910539
transform 1 0 17112 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1608910539
transform 1 0 17940 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp 1608910539
transform 1 0 18492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1608910539
transform -1 0 18860 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1608910539
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1608910539
transform 1 0 1748 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1608910539
transform 1 0 2576 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1608910539
transform 1 0 1380 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_38
timestamp 1608910539
transform 1 0 4600 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1608910539
transform 1 0 3404 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 4692 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1608910539
transform 1 0 4232 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1608910539
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 6164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_64
timestamp 1608910539
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1608910539
transform 1 0 7728 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6900 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1608910539
transform 1 0 8556 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_84
timestamp 1608910539
transform 1 0 8832 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10672 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 10396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8924 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_65
timestamp 1608910539
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 10856 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13892 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1608910539
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1608910539
transform 1 0 15456 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16284 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66
timestamp 1608910539
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1608910539
transform 1 0 17112 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1608910539
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 18400 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1608910539
transform -1 0 18860 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_10
timestamp 1608910539
transform 1 0 2024 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1608910539
transform 1 0 1380 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1608910539
transform 1 0 1380 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 1472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1608910539
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1608910539
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1608910539
transform 1 0 1472 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1608910539
transform 1 0 1656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1608910539
transform 1 0 2116 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1608910539
transform 1 0 2300 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 2944 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1608910539
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1608910539
transform 1 0 3128 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1608910539
transform 1 0 4416 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1608910539
transform 1 0 4784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1608910539
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1608910539
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5520 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1608910539
transform 1 0 6348 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 5060 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 6808 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_78
timestamp 1608910539
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 7176 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8188 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1608910539
transform 1 0 7360 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8372 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1608910539
transform 1 0 9660 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1608910539
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1608910539
transform 1 0 10672 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 9752 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 12052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 12236 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1608910539
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1608910539
transform 1 0 11224 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11500 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1608910539
transform 1 0 12512 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1608910539
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_126
timestamp 1608910539
transform 1 0 12696 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 13340 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 12788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13524 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12972 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13708 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13800 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_7_154
timestamp 1608910539
transform 1 0 15272 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_146
timestamp 1608910539
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1608910539
transform 1 0 15364 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1608910539
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1608910539
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15732 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1608910539
transform 1 0 16100 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16376 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1608910539
transform 1 0 17388 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1608910539
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1608910539
transform 1 0 16560 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1608910539
transform 1 0 17572 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1608910539
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1608910539
transform 1 0 18216 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1608910539
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1608910539
transform 1 0 18400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1608910539
transform -1 0 18860 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1608910539
transform -1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1608910539
transform 1 0 1380 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1608910539
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 1564 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_21
timestamp 1608910539
transform 1 0 3036 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1608910539
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1608910539
transform 1 0 3128 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4876 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6624 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 6348 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1608910539
transform 1 0 6808 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_71
timestamp 1608910539
transform 1 0 7636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 7728 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_8_93
timestamp 1608910539
transform 1 0 9660 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9200 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1608910539
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10028 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1608910539
transform 1 0 9752 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12328 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10856 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12880 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13708 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_8_146
timestamp 1608910539
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1608910539
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15456 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1608910539
transform 1 0 17756 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1608910539
transform 1 0 16928 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1608910539
transform -1 0 18860 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 2576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1608910539
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1608910539
transform 1 0 1748 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1608910539
transform 1 0 2760 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1608910539
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3588 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1608910539
transform 1 0 4600 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1608910539
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1608910539
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1608910539
transform 1 0 5428 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1608910539
transform 1 0 6256 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1608910539
transform 1 0 8096 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _16_
timestamp 1608910539
transform 1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1608910539
transform 1 0 10580 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9752 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1608910539
transform 1 0 8924 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_9_112
timestamp 1608910539
transform 1 0 11408 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1608910539
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 14076 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 13892 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 14260 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_9_159
timestamp 1608910539
transform 1 0 15732 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16100 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1608910539
transform 1 0 15824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1608910539
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1608910539
transform 1 0 18032 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1608910539
transform 1 0 18400 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1608910539
transform -1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1608910539
transform 1 0 1380 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 1472 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 1656 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1608910539
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1608910539
transform 1 0 2668 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1608910539
transform 1 0 1840 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_28
timestamp 1608910539
transform 1 0 3680 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3496 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1608910539
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1608910539
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1608910539
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5888 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_10_73
timestamp 1608910539
transform 1 0 7820 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp 1608910539
transform 1 0 7544 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1608910539
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 7636 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1608910539
transform 1 0 8096 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_87
timestamp 1608910539
transform 1 0 9108 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8924 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 9660 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1608910539
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_122
timestamp 1608910539
transform 1 0 12328 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1608910539
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 12420 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1608910539
transform 1 0 13892 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_164
timestamp 1608910539
transform 1 0 16192 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1608910539
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_148
timestamp 1608910539
transform 1 0 14720 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1608910539
transform 1 0 14812 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1608910539
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1608910539
transform 1 0 15364 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1608910539
transform 1 0 17296 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1608910539
transform 1 0 16468 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1608910539
transform 1 0 18124 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1608910539
transform 1 0 18492 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1608910539
transform -1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1608910539
transform 1 0 1380 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1608910539
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 1564 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 4508 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 3036 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1608910539
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_53
timestamp 1608910539
transform 1 0 5980 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1608910539
transform 1 0 6256 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 6072 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1608910539
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8280 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 10488 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_125
timestamp 1608910539
transform 1 0 12604 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1608910539
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1608910539
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 14168 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 12696 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1608910539
transform 1 0 13156 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 14352 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_11_160
timestamp 1608910539
transform 1 0 15824 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 16284 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1608910539
transform 1 0 15916 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1608910539
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1608910539
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1608910539
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1608910539
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1608910539
transform -1 0 18860 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1608910539
transform 1 0 1380 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1608910539
transform 1 0 1472 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1608910539
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 1656 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1608910539
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1608910539
transform 1 0 3128 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 3680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 3496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 3312 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1608910539
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_39
timestamp 1608910539
transform 1 0 4692 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_32
timestamp 1608910539
transform 1 0 4048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 4508 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 4140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 4784 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1608910539
transform 1 0 6256 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_79
timestamp 1608910539
transform 1 0 8372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_65
timestamp 1608910539
transform 1 0 7084 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1608910539
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1608910539
transform 1 0 8464 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1608910539
transform 1 0 9292 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1608910539
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1608910539
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1608910539
transform 1 0 11132 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1608910539
transform 1 0 11960 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1608910539
transform 1 0 12788 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 13616 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_154
timestamp 1608910539
transform 1 0 15272 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1608910539
transform 1 0 15088 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1608910539
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 15364 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_12_181
timestamp 1608910539
transform 1 0 17756 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_171
timestamp 1608910539
transform 1 0 16836 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1608910539
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1608910539
transform 1 0 18216 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1608910539
transform 1 0 17848 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1608910539
transform -1 0 18860 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1608910539
transform 1 0 1380 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1608910539
transform 1 0 1472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1608910539
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1608910539
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1608910539
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1608910539
transform 1 0 1656 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_12
timestamp 1608910539
transform 1 0 2208 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1608910539
transform 1 0 2300 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1608910539
transform 1 0 2852 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 1380 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp 1608910539
transform 1 0 4048 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_25
timestamp 1608910539
transform 1 0 3404 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 4140 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 3128 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1608910539
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1608910539
transform 1 0 3128 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1608910539
transform 1 0 3496 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1608910539
transform 1 0 4324 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1608910539
transform 1 0 4324 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5152 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1608910539
transform 1 0 5152 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1608910539
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 6440 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6256 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 5980 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1608910539
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1608910539
transform 1 0 6164 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 6808 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 1608910539
transform 1 0 7176 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 7268 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 8280 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 9200 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1608910539
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_94
timestamp 1608910539
transform 1 0 9752 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1608910539
transform 1 0 9844 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1608910539
transform 1 0 9844 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1608910539
transform 1 0 10672 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1608910539
transform 1 0 10672 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_14_116
timestamp 1608910539
transform 1 0 11776 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1608910539
transform 1 0 12420 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 11500 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1608910539
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11500 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 11868 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1608910539
transform 1 0 12512 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_136
timestamp 1608910539
transform 1 0 13616 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1608910539
transform 1 0 14168 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1608910539
transform 1 0 13340 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1608910539
transform 1 0 13708 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12788 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1608910539
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1608910539
transform 1 0 15364 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_top_ipin_0.prog_clk
timestamp 1608910539
transform 1 0 16376 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1608910539
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1608910539
transform 1 0 15548 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1608910539
transform 1 0 14536 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1608910539
transform 1 0 16652 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1608910539
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1608910539
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1608910539
transform 1 0 16744 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1608910539
transform 1 0 16744 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1608910539
transform 1 0 17572 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1608910539
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1608910539
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1608910539
transform 1 0 18400 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1608910539
transform -1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1608910539
transform -1 0 18860 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1608910539
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1608910539
transform 1 0 1380 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1608910539
transform 1 0 2208 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_21
timestamp 1608910539
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1608910539
transform 1 0 3128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 3956 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_49
timestamp 1608910539
transform 1 0 5612 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 5428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1608910539
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_15_80
timestamp 1608910539
transform 1 0 8464 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 8740 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_15_99
timestamp 1608910539
transform 1 0 10212 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1608910539
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1608910539
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1608910539
transform 1 0 11132 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1608910539
transform 1 0 13892 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1608910539
transform 1 0 15364 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 16192 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1608910539
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1608910539
transform 1 0 18032 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1608910539
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1608910539
transform -1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1608910539
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1608910539
transform 1 0 1656 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 1840 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1608910539
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 2208 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_16_35
timestamp 1608910539
transform 1 0 4324 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1608910539
transform 1 0 4048 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1608910539
transform 1 0 3864 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 3680 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1608910539
transform 1 0 4140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1608910539
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp 1608910539
transform 1 0 5060 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1608910539
transform 1 0 6716 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 5244 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1608910539
transform 1 0 8372 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1608910539
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_16_93
timestamp 1608910539
transform 1 0 9660 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1608910539
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 9200 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1608910539
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1608910539
transform 1 0 10212 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1608910539
transform 1 0 9936 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1608910539
transform 1 0 12512 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1608910539
transform 1 0 11684 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_138
timestamp 1608910539
transform 1 0 13800 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_133
timestamp 1608910539
transform 1 0 13340 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1608910539
transform 1 0 13616 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_150
timestamp 1608910539
transform 1 0 14904 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1608910539
transform 1 0 14720 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 14536 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1608910539
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1608910539
transform 1 0 15272 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1608910539
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1608910539
transform 1 0 17296 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1608910539
transform 1 0 16744 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1608910539
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1608910539
transform 1 0 17480 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1608910539
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1608910539
transform -1 0 18860 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_18 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 2760 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 1380 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1608910539
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1608910539
transform 1 0 1932 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_30
timestamp 1608910539
transform 1 0 3864 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1608910539
transform 1 0 5704 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_42
timestamp 1608910539
transform 1 0 4968 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1608910539
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1608910539
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1608910539
transform 1 0 5888 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_17_64
timestamp 1608910539
transform 1 0 6992 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1608910539
transform 1 0 7084 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1608910539
transform 1 0 8372 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1608910539
transform 1 0 7912 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_95
timestamp 1608910539
transform 1 0 9844 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1608910539
transform 1 0 10120 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1608910539
transform 1 0 10304 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1608910539
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1608910539
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1608910539
transform 1 0 11132 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_17_135
timestamp 1608910539
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1608910539
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 14444 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_157
timestamp 1608910539
transform 1 0 15548 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1608910539
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1608910539
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_169
timestamp 1608910539
transform 1 0 16652 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1608910539
transform 1 0 18124 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1608910539
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 18308 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1608910539
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1608910539
transform 1 0 18492 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1608910539
transform -1 0 18860 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1608910539
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1608910539
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1608910539
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1608910539
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1608910539
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1608910539
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1608910539
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1608910539
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_76
timestamp 1608910539
transform 1 0 8096 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1608910539
transform 1 0 7360 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1608910539
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_104
timestamp 1608910539
transform 1 0 10672 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1608910539
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1608910539
transform 1 0 9200 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1608910539
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1608910539
transform 1 0 9844 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_18_116
timestamp 1608910539
transform 1 0 11776 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_140
timestamp 1608910539
transform 1 0 13984 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_128
timestamp 1608910539
transform 1 0 12880 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1608910539
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1608910539
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_152
timestamp 1608910539
transform 1 0 15088 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1608910539
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1608910539
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1608910539
transform -1 0 18860 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1608910539
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1608910539
transform 1 0 1472 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1608910539
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1608910539
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01
timestamp 1608910539
transform 1 0 2024 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _32_
timestamp 1608910539
transform 1 0 1656 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_E_FTB01_A
timestamp 1608910539
transform 1 0 2576 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_18
timestamp 1608910539
transform 1 0 2760 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1608910539
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1608910539
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1608910539
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_30
timestamp 1608910539
transform 1 0 3864 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1608910539
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1608910539
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1608910539
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1608910539
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1608910539
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1608910539
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1608910539
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1608910539
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1608910539
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1608910539
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1608910539
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1608910539
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1608910539
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1608910539
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1608910539
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1608910539
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1608910539
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1608910539
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1608910539
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1608910539
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1608910539
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1608910539
transform 1 0 14076 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1608910539
transform 1 0 12972 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1608910539
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_166
timestamp 1608910539
transform 1 0 16376 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1608910539
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_159
timestamp 1608910539
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_147
timestamp 1608910539
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1608910539
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_185
timestamp 1608910539
transform 1 0 18124 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1608910539
transform 1 0 17112 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1608910539
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_171
timestamp 1608910539
transform 1 0 16836 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_E_FTB01_A
timestamp 1608910539
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_S_FTB01_A
timestamp 1608910539
transform 1 0 17388 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1608910539
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  clk_3_E_FTB01
timestamp 1608910539
transform 1 0 18032 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_1_S_FTB01
timestamp 1608910539
transform 1 0 17572 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1608910539
transform 1 0 18492 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1608910539
transform -1 0 18860 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1608910539
transform -1 0 18860 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_19
timestamp 1608910539
transform 1 0 2852 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_W_FTB01_A
timestamp 1608910539
transform 1 0 2668 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_W_FTB01_A
timestamp 1608910539
transform 1 0 1380 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1608910539
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  clk_3_W_FTB01
timestamp 1608910539
transform 1 0 2116 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_W_FTB01
timestamp 1608910539
transform 1 0 1564 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_31
timestamp 1608910539
transform 1 0 3956 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1608910539
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_43
timestamp 1608910539
transform 1 0 5060 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1608910539
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1608910539
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1608910539
transform 1 0 6164 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1608910539
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1608910539
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_86
timestamp 1608910539
transform 1 0 9016 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_1_N_FTB01_A
timestamp 1608910539
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  clk_1_N_FTB01
timestamp 1608910539
transform 1 0 9568 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1608910539
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1608910539
transform 1 0 11224 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1608910539
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1608910539
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_159
timestamp 1608910539
transform 1 0 15732 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_147
timestamp 1608910539
transform 1 0 14628 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_167
timestamp 1608910539
transform 1 0 16468 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_W_FTB01_A
timestamp 1608910539
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1608910539
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1608910539
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1608910539
transform 1 0 16836 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_E_FTB01
timestamp 1608910539
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1608910539
transform 1 0 17388 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1608910539
transform -1 0 18860 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_19
timestamp 1608910539
transform 1 0 2852 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_W_FTB01_A
timestamp 1608910539
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_W_FTB01_A
timestamp 1608910539
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1608910539
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_W_FTB01
timestamp 1608910539
transform 1 0 2116 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1608910539
transform 1 0 1564 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1608910539
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1608910539
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_56
timestamp 1608910539
transform 1 0 6256 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1608910539
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1608910539
transform 1 0 6808 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_75
timestamp 1608910539
transform 1 0 8004 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_63
timestamp 1608910539
transform 1 0 6900 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_94
timestamp 1608910539
transform 1 0 9752 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_87
timestamp 1608910539
transform 1 0 9108 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1608910539
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_125
timestamp 1608910539
transform 1 0 12604 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_118
timestamp 1608910539
transform 1 0 11960 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_106
timestamp 1608910539
transform 1 0 10856 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1608910539
transform 1 0 12512 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1608910539
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_156
timestamp 1608910539
transform 1 0 15456 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_149
timestamp 1608910539
transform 1 0 14812 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1608910539
transform 1 0 15364 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_187
timestamp 1608910539
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1608910539
transform 1 0 18032 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_180
timestamp 1608910539
transform 1 0 17664 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_168
timestamp 1608910539
transform 1 0 16560 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_E_FTB01_A
timestamp 1608910539
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1608910539
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1608910539
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 13608 800 13728 6 REGIN_FEEDTHROUGH
port 0 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 REGOUT_FEEDTHROUGH
port 1 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 SC_IN_BOT
port 2 nsew signal input
rlabel metal2 s 1950 16400 2006 17200 6 SC_IN_TOP
port 3 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_OUT_BOT
port 4 nsew signal tristate
rlabel metal2 s 5906 16400 5962 17200 6 SC_OUT_TOP
port 5 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_0_
port 6 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_10_
port 7 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_11_
port 8 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_12_
port 9 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_13_
port 10 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_14_
port 11 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_grid_pin_15_
port 12 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_1_
port 13 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_2_
port 14 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_3_
port 15 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_4_
port 16 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_5_
port 17 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_6_
port 18 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_7_
port 19 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_8_
port 20 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_9_
port 21 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 ccff_head
port 22 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 ccff_tail
port 23 nsew signal tristate
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[0]
port 24 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[10]
port 25 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[11]
port 26 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[12]
port 27 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[13]
port 28 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[14]
port 29 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[15]
port 30 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[16]
port 31 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 32 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 33 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[19]
port 34 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[1]
port 35 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[2]
port 36 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[3]
port 37 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[4]
port 38 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[5]
port 39 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[6]
port 40 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[7]
port 41 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[8]
port 42 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[9]
port 43 nsew signal input
rlabel metal3 s 0 144 800 264 6 chanx_left_out[0]
port 44 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[10]
port 45 nsew signal tristate
rlabel metal3 s 0 3680 800 3800 6 chanx_left_out[11]
port 46 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 chanx_left_out[12]
port 47 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_out[13]
port 48 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[14]
port 49 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[15]
port 50 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 chanx_left_out[16]
port 51 nsew signal tristate
rlabel metal3 s 0 5720 800 5840 6 chanx_left_out[17]
port 52 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[18]
port 53 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[19]
port 54 nsew signal tristate
rlabel metal3 s 0 416 800 536 6 chanx_left_out[1]
port 55 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 chanx_left_out[2]
port 56 nsew signal tristate
rlabel metal3 s 0 1096 800 1216 6 chanx_left_out[3]
port 57 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[4]
port 58 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[5]
port 59 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 chanx_left_out[6]
port 60 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 chanx_left_out[7]
port 61 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 chanx_left_out[8]
port 62 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[9]
port 63 nsew signal tristate
rlabel metal3 s 19200 9664 20000 9784 6 chanx_right_in[0]
port 64 nsew signal input
rlabel metal3 s 19200 13472 20000 13592 6 chanx_right_in[10]
port 65 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[11]
port 66 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[12]
port 67 nsew signal input
rlabel metal3 s 19200 14560 20000 14680 6 chanx_right_in[13]
port 68 nsew signal input
rlabel metal3 s 19200 14968 20000 15088 6 chanx_right_in[14]
port 69 nsew signal input
rlabel metal3 s 19200 15376 20000 15496 6 chanx_right_in[15]
port 70 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 chanx_right_in[16]
port 71 nsew signal input
rlabel metal3 s 19200 16056 20000 16176 6 chanx_right_in[17]
port 72 nsew signal input
rlabel metal3 s 19200 16464 20000 16584 6 chanx_right_in[18]
port 73 nsew signal input
rlabel metal3 s 19200 16872 20000 16992 6 chanx_right_in[19]
port 74 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[1]
port 75 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[2]
port 76 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[3]
port 77 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[4]
port 78 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 chanx_right_in[5]
port 79 nsew signal input
rlabel metal3 s 19200 11840 20000 11960 6 chanx_right_in[6]
port 80 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 chanx_right_in[7]
port 81 nsew signal input
rlabel metal3 s 19200 12656 20000 12776 6 chanx_right_in[8]
port 82 nsew signal input
rlabel metal3 s 19200 13064 20000 13184 6 chanx_right_in[9]
port 83 nsew signal input
rlabel metal3 s 19200 2048 20000 2168 6 chanx_right_out[0]
port 84 nsew signal tristate
rlabel metal3 s 19200 5856 20000 5976 6 chanx_right_out[10]
port 85 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[11]
port 86 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[12]
port 87 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[13]
port 88 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[14]
port 89 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[15]
port 90 nsew signal tristate
rlabel metal3 s 19200 8032 20000 8152 6 chanx_right_out[16]
port 91 nsew signal tristate
rlabel metal3 s 19200 8440 20000 8560 6 chanx_right_out[17]
port 92 nsew signal tristate
rlabel metal3 s 19200 8848 20000 8968 6 chanx_right_out[18]
port 93 nsew signal tristate
rlabel metal3 s 19200 9256 20000 9376 6 chanx_right_out[19]
port 94 nsew signal tristate
rlabel metal3 s 19200 2320 20000 2440 6 chanx_right_out[1]
port 95 nsew signal tristate
rlabel metal3 s 19200 2728 20000 2848 6 chanx_right_out[2]
port 96 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[3]
port 97 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[4]
port 98 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[5]
port 99 nsew signal tristate
rlabel metal3 s 19200 4224 20000 4344 6 chanx_right_out[6]
port 100 nsew signal tristate
rlabel metal3 s 19200 4632 20000 4752 6 chanx_right_out[7]
port 101 nsew signal tristate
rlabel metal3 s 19200 5040 20000 5160 6 chanx_right_out[8]
port 102 nsew signal tristate
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[9]
port 103 nsew signal tristate
rlabel metal2 s 9862 16400 9918 17200 6 clk_1_N_out
port 104 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 clk_1_S_out
port 105 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 clk_1_W_in
port 106 nsew signal input
rlabel metal3 s 19200 1640 20000 1760 6 clk_2_E_out
port 107 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 clk_2_W_in
port 108 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 clk_2_W_out
port 109 nsew signal tristate
rlabel metal3 s 19200 1232 20000 1352 6 clk_3_E_out
port 110 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 clk_3_W_in
port 111 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 clk_3_W_out
port 112 nsew signal tristate
rlabel metal2 s 13910 16400 13966 17200 6 prog_clk_0_N_in
port 113 nsew signal input
rlabel metal2 s 17866 16400 17922 17200 6 prog_clk_0_W_out
port 114 nsew signal tristate
rlabel metal3 s 19200 824 20000 944 6 prog_clk_1_N_out
port 115 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_1_S_out
port 116 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 prog_clk_1_W_in
port 117 nsew signal input
rlabel metal3 s 19200 416 20000 536 6 prog_clk_2_E_out
port 118 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 prog_clk_2_W_in
port 119 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 prog_clk_2_W_out
port 120 nsew signal tristate
rlabel metal3 s 19200 144 20000 264 6 prog_clk_3_E_out
port 121 nsew signal tristate
rlabel metal3 s 0 15240 800 15360 6 prog_clk_3_W_in
port 122 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 prog_clk_3_W_out
port 123 nsew signal tristate
rlabel metal4 s 15771 2128 16091 14736 6 VPWR
port 124 nsew power bidirectional
rlabel metal4 s 9840 2128 10160 14736 6 VPWR
port 125 nsew power bidirectional
rlabel metal4 s 3909 2128 4229 14736 6 VPWR
port 126 nsew power bidirectional
rlabel metal4 s 12805 2128 13125 14736 6 VGND
port 127 nsew ground bidirectional
rlabel metal4 s 6875 2128 7195 14736 6 VGND
port 128 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
