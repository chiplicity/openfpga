magic
tech sky130A
magscale 1 2
timestamp 1606931033
<< locali >>
rect 2329 13855 2363 14025
rect 20453 13855 20487 13957
rect 6653 12699 6687 12869
rect 2789 11747 2823 11781
rect 2731 11713 2823 11747
rect 15393 11611 15427 11781
rect 7481 11135 7515 11305
rect 12173 10591 12207 10761
rect 10425 9435 10459 9537
rect 15025 9027 15059 9129
rect 12173 8347 12207 8449
rect 15209 7395 15243 7497
rect 13001 6715 13035 6817
rect 12633 5559 12667 5729
rect 17233 4607 17267 4709
rect 11713 3927 11747 4029
rect 3341 2839 3375 3145
<< viali >>
rect 1961 19465 1995 19499
rect 6009 19465 6043 19499
rect 19165 19465 19199 19499
rect 20729 19465 20763 19499
rect 1777 19261 1811 19295
rect 2329 19261 2363 19295
rect 5825 19261 5859 19295
rect 18981 19261 19015 19295
rect 20545 19261 20579 19295
rect 2513 19125 2547 19159
rect 1961 18921 1995 18955
rect 6377 18853 6411 18887
rect 18429 18853 18463 18887
rect 1777 18785 1811 18819
rect 6101 18785 6135 18819
rect 18153 18785 18187 18819
rect 1961 18377 1995 18411
rect 20729 18377 20763 18411
rect 1777 18173 1811 18207
rect 20545 18173 20579 18207
rect 1869 17833 1903 17867
rect 2513 17765 2547 17799
rect 19993 17765 20027 17799
rect 1685 17697 1719 17731
rect 2237 17697 2271 17731
rect 19717 17697 19751 17731
rect 1961 17289 1995 17323
rect 20729 17289 20763 17323
rect 1777 17085 1811 17119
rect 20545 17085 20579 17119
rect 1961 16745 1995 16779
rect 20453 16745 20487 16779
rect 1777 16609 1811 16643
rect 20269 16609 20303 16643
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 3433 16201 3467 16235
rect 13553 16201 13587 16235
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 1777 15997 1811 16031
rect 2329 15997 2363 16031
rect 3249 15997 3283 16031
rect 13369 15997 13403 16031
rect 19993 15997 20027 16031
rect 20545 15997 20579 16031
rect 1961 15657 1995 15691
rect 2513 15657 2547 15691
rect 20453 15657 20487 15691
rect 4353 15589 4387 15623
rect 12817 15589 12851 15623
rect 1777 15521 1811 15555
rect 2329 15521 2363 15555
rect 4077 15521 4111 15555
rect 12541 15521 12575 15555
rect 20269 15521 20303 15555
rect 2513 15113 2547 15147
rect 20177 15113 20211 15147
rect 20729 15113 20763 15147
rect 1961 15045 1995 15079
rect 13737 15045 13771 15079
rect 19625 15045 19659 15079
rect 14381 14977 14415 15011
rect 1777 14909 1811 14943
rect 2329 14909 2363 14943
rect 2973 14909 3007 14943
rect 19441 14909 19475 14943
rect 19993 14909 20027 14943
rect 20545 14909 20579 14943
rect 3240 14841 3274 14875
rect 14105 14841 14139 14875
rect 4353 14773 4387 14807
rect 14197 14773 14231 14807
rect 1685 14569 1719 14603
rect 4261 14569 4295 14603
rect 13461 14569 13495 14603
rect 2329 14501 2363 14535
rect 12050 14501 12084 14535
rect 13829 14501 13863 14535
rect 16221 14501 16255 14535
rect 17018 14501 17052 14535
rect 19993 14501 20027 14535
rect 1501 14433 1535 14467
rect 2053 14433 2087 14467
rect 3157 14433 3191 14467
rect 4077 14433 4111 14467
rect 9945 14433 9979 14467
rect 13921 14433 13955 14467
rect 16129 14433 16163 14467
rect 19165 14433 19199 14467
rect 19717 14433 19751 14467
rect 3249 14365 3283 14399
rect 3433 14365 3467 14399
rect 9689 14365 9723 14399
rect 11805 14365 11839 14399
rect 14105 14365 14139 14399
rect 16313 14365 16347 14399
rect 16773 14365 16807 14399
rect 2789 14297 2823 14331
rect 11069 14229 11103 14263
rect 13185 14229 13219 14263
rect 15761 14229 15795 14263
rect 18153 14229 18187 14263
rect 19349 14229 19383 14263
rect 2329 14025 2363 14059
rect 14565 14025 14599 14059
rect 18981 14025 19015 14059
rect 19533 14025 19567 14059
rect 1961 13889 1995 13923
rect 5457 13957 5491 13991
rect 12081 13957 12115 13991
rect 16497 13957 16531 13991
rect 20453 13957 20487 13991
rect 4077 13889 4111 13923
rect 7481 13889 7515 13923
rect 8401 13889 8435 13923
rect 10701 13889 10735 13923
rect 13185 13889 13219 13923
rect 17049 13889 17083 13923
rect 20821 13889 20855 13923
rect 1685 13821 1719 13855
rect 2329 13821 2363 13855
rect 2421 13821 2455 13855
rect 4333 13821 4367 13855
rect 7297 13821 7331 13855
rect 10968 13821 11002 13855
rect 13452 13821 13486 13855
rect 14841 13821 14875 13855
rect 15097 13821 15131 13855
rect 18061 13821 18095 13855
rect 18797 13821 18831 13855
rect 19349 13821 19383 13855
rect 19901 13821 19935 13855
rect 20177 13821 20211 13855
rect 20453 13821 20487 13855
rect 20637 13821 20671 13855
rect 2688 13753 2722 13787
rect 7205 13753 7239 13787
rect 7849 13753 7883 13787
rect 8646 13753 8680 13787
rect 16865 13753 16899 13787
rect 17509 13753 17543 13787
rect 18337 13753 18371 13787
rect 3801 13685 3835 13719
rect 6837 13685 6871 13719
rect 9781 13685 9815 13719
rect 16221 13685 16255 13719
rect 16957 13685 16991 13719
rect 1593 13481 1627 13515
rect 1961 13481 1995 13515
rect 2973 13481 3007 13515
rect 4261 13481 4295 13515
rect 5089 13481 5123 13515
rect 5181 13481 5215 13515
rect 6285 13481 6319 13515
rect 6653 13481 6687 13515
rect 8677 13481 8711 13515
rect 10149 13481 10183 13515
rect 16957 13481 16991 13515
rect 9689 13413 9723 13447
rect 11529 13413 11563 13447
rect 11621 13413 11655 13447
rect 15844 13413 15878 13447
rect 1409 13345 1443 13379
rect 2329 13345 2363 13379
rect 3341 13345 3375 13379
rect 4077 13345 4111 13379
rect 6745 13345 6779 13379
rect 7564 13345 7598 13379
rect 10517 13345 10551 13379
rect 10609 13345 10643 13379
rect 13093 13345 13127 13379
rect 13360 13345 13394 13379
rect 15577 13345 15611 13379
rect 17785 13345 17819 13379
rect 18052 13345 18086 13379
rect 19809 13345 19843 13379
rect 19901 13345 19935 13379
rect 2421 13277 2455 13311
rect 2605 13277 2639 13311
rect 3433 13277 3467 13311
rect 3525 13277 3559 13311
rect 5365 13277 5399 13311
rect 6837 13277 6871 13311
rect 7297 13277 7331 13311
rect 10793 13277 10827 13311
rect 11805 13277 11839 13311
rect 12541 13277 12575 13311
rect 14749 13277 14783 13311
rect 19993 13277 20027 13311
rect 4721 13141 4755 13175
rect 11161 13141 11195 13175
rect 14473 13141 14507 13175
rect 19165 13141 19199 13175
rect 19441 13141 19475 13175
rect 2513 12937 2547 12971
rect 3801 12937 3835 12971
rect 6837 12937 6871 12971
rect 9045 12937 9079 12971
rect 11069 12937 11103 12971
rect 13829 12937 13863 12971
rect 16589 12937 16623 12971
rect 20913 12937 20947 12971
rect 6193 12869 6227 12903
rect 6653 12869 6687 12903
rect 7849 12869 7883 12903
rect 15577 12869 15611 12903
rect 1961 12801 1995 12835
rect 2973 12801 3007 12835
rect 3157 12801 3191 12835
rect 4353 12801 4387 12835
rect 4813 12801 4847 12835
rect 1777 12733 1811 12767
rect 4261 12733 4295 12767
rect 7389 12801 7423 12835
rect 8309 12801 8343 12835
rect 8493 12801 8527 12835
rect 9505 12801 9539 12835
rect 9597 12801 9631 12835
rect 10609 12801 10643 12835
rect 11621 12801 11655 12835
rect 13001 12801 13035 12835
rect 14289 12801 14323 12835
rect 14473 12801 14507 12835
rect 16129 12801 16163 12835
rect 17141 12801 17175 12835
rect 18245 12801 18279 12835
rect 20177 12801 20211 12835
rect 12817 12733 12851 12767
rect 14197 12733 14231 12767
rect 18512 12733 18546 12767
rect 19993 12733 20027 12767
rect 20729 12733 20763 12767
rect 5080 12665 5114 12699
rect 6653 12665 6687 12699
rect 7297 12665 7331 12699
rect 8217 12665 8251 12699
rect 9413 12665 9447 12699
rect 10517 12665 10551 12699
rect 11437 12665 11471 12699
rect 11529 12665 11563 12699
rect 16037 12665 16071 12699
rect 2881 12597 2915 12631
rect 4169 12597 4203 12631
rect 7205 12597 7239 12631
rect 10057 12597 10091 12631
rect 10425 12597 10459 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 15945 12597 15979 12631
rect 16957 12597 16991 12631
rect 17049 12597 17083 12631
rect 19625 12597 19659 12631
rect 2421 12393 2455 12427
rect 3617 12393 3651 12427
rect 5457 12393 5491 12427
rect 7941 12393 7975 12427
rect 12909 12393 12943 12427
rect 14105 12393 14139 12427
rect 15945 12393 15979 12427
rect 16405 12393 16439 12427
rect 17325 12393 17359 12427
rect 18337 12393 18371 12427
rect 19165 12393 19199 12427
rect 1869 12325 1903 12359
rect 6552 12325 6586 12359
rect 19533 12325 19567 12359
rect 20913 12325 20947 12359
rect 1777 12257 1811 12291
rect 2789 12257 2823 12291
rect 3433 12257 3467 12291
rect 4333 12257 4367 12291
rect 8309 12257 8343 12291
rect 10149 12257 10183 12291
rect 10793 12257 10827 12291
rect 11060 12257 11094 12291
rect 12817 12257 12851 12291
rect 13461 12257 13495 12291
rect 14473 12257 14507 12291
rect 16313 12257 16347 12291
rect 18981 12257 19015 12291
rect 19625 12257 19659 12291
rect 20269 12257 20303 12291
rect 2053 12189 2087 12223
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 4077 12189 4111 12223
rect 6285 12189 6319 12223
rect 8401 12189 8435 12223
rect 8493 12189 8527 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 13001 12189 13035 12223
rect 14565 12189 14599 12223
rect 14749 12189 14783 12223
rect 16497 12189 16531 12223
rect 17417 12189 17451 12223
rect 17509 12189 17543 12223
rect 18429 12189 18463 12223
rect 18613 12189 18647 12223
rect 19717 12189 19751 12223
rect 7665 12121 7699 12155
rect 12173 12121 12207 12155
rect 16957 12121 16991 12155
rect 20453 12121 20487 12155
rect 1409 12053 1443 12087
rect 9781 12053 9815 12087
rect 12449 12053 12483 12087
rect 17969 12053 18003 12087
rect 11805 11849 11839 11883
rect 13461 11849 13495 11883
rect 16957 11849 16991 11883
rect 18061 11849 18095 11883
rect 20913 11849 20947 11883
rect 2789 11781 2823 11815
rect 4997 11781 5031 11815
rect 7481 11781 7515 11815
rect 8493 11781 8527 11815
rect 15301 11781 15335 11815
rect 15393 11781 15427 11815
rect 2513 11713 2547 11747
rect 2697 11713 2731 11747
rect 4261 11713 4295 11747
rect 5549 11713 5583 11747
rect 8033 11713 8067 11747
rect 8769 11713 8803 11747
rect 13001 11713 13035 11747
rect 2881 11645 2915 11679
rect 3157 11645 3191 11679
rect 5365 11645 5399 11679
rect 5457 11645 5491 11679
rect 6193 11645 6227 11679
rect 7849 11645 7883 11679
rect 8677 11645 8711 11679
rect 10425 11645 10459 11679
rect 12817 11645 12851 11679
rect 13645 11645 13679 11679
rect 13921 11645 13955 11679
rect 14188 11645 14222 11679
rect 15577 11713 15611 11747
rect 18521 11713 18555 11747
rect 18705 11713 18739 11747
rect 17233 11645 17267 11679
rect 19073 11645 19107 11679
rect 19340 11645 19374 11679
rect 20729 11645 20763 11679
rect 9036 11577 9070 11611
rect 10670 11577 10704 11611
rect 12909 11577 12943 11611
rect 15393 11577 15427 11611
rect 15844 11577 15878 11611
rect 17509 11577 17543 11611
rect 1869 11509 1903 11543
rect 2237 11509 2271 11543
rect 2329 11509 2363 11543
rect 3617 11509 3651 11543
rect 3985 11509 4019 11543
rect 4077 11509 4111 11543
rect 6009 11509 6043 11543
rect 7941 11509 7975 11543
rect 10149 11509 10183 11543
rect 12449 11509 12483 11543
rect 18429 11509 18463 11543
rect 20453 11509 20487 11543
rect 3525 11305 3559 11339
rect 7297 11305 7331 11339
rect 7481 11305 7515 11339
rect 8033 11305 8067 11339
rect 8585 11305 8619 11339
rect 12909 11305 12943 11339
rect 15301 11305 15335 11339
rect 16313 11305 16347 11339
rect 18797 11305 18831 11339
rect 20269 11305 20303 11339
rect 1869 11169 1903 11203
rect 2136 11169 2170 11203
rect 4261 11169 4295 11203
rect 4528 11169 4562 11203
rect 6173 11169 6207 11203
rect 9045 11237 9079 11271
rect 10977 11237 11011 11271
rect 11796 11237 11830 11271
rect 15669 11237 15703 11271
rect 17132 11237 17166 11271
rect 7941 11169 7975 11203
rect 8953 11169 8987 11203
rect 10057 11169 10091 11203
rect 10701 11169 10735 11203
rect 13369 11169 13403 11203
rect 13636 11169 13670 11203
rect 19165 11169 19199 11203
rect 20177 11169 20211 11203
rect 5917 11101 5951 11135
rect 7481 11101 7515 11135
rect 8125 11101 8159 11135
rect 9229 11101 9263 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11529 11101 11563 11135
rect 15761 11101 15795 11135
rect 15945 11101 15979 11135
rect 16865 11101 16899 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 20361 11101 20395 11135
rect 3249 11033 3283 11067
rect 5641 11033 5675 11067
rect 7573 11033 7607 11067
rect 9689 11033 9723 11067
rect 14749 11033 14783 11067
rect 18245 11033 18279 11067
rect 19809 11033 19843 11067
rect 2053 10761 2087 10795
rect 3065 10761 3099 10795
rect 5457 10761 5491 10795
rect 8217 10761 8251 10795
rect 9045 10761 9079 10795
rect 10057 10761 10091 10795
rect 11345 10761 11379 10795
rect 12173 10761 12207 10795
rect 14289 10761 14323 10795
rect 16497 10761 16531 10795
rect 19441 10761 19475 10795
rect 2513 10625 2547 10659
rect 2697 10625 2731 10659
rect 3617 10625 3651 10659
rect 6193 10625 6227 10659
rect 6285 10625 6319 10659
rect 6837 10625 6871 10659
rect 9597 10625 9631 10659
rect 10609 10625 10643 10659
rect 11897 10625 11931 10659
rect 17509 10693 17543 10727
rect 12449 10625 12483 10659
rect 14841 10625 14875 10659
rect 16037 10625 16071 10659
rect 17141 10625 17175 10659
rect 18061 10625 18095 10659
rect 3433 10557 3467 10591
rect 4077 10557 4111 10591
rect 9505 10557 9539 10591
rect 11805 10557 11839 10591
rect 12173 10557 12207 10591
rect 12716 10557 12750 10591
rect 17693 10557 17727 10591
rect 19717 10557 19751 10591
rect 19973 10557 20007 10591
rect 4344 10489 4378 10523
rect 6101 10489 6135 10523
rect 7104 10489 7138 10523
rect 8585 10489 8619 10523
rect 9413 10489 9447 10523
rect 14749 10489 14783 10523
rect 15853 10489 15887 10523
rect 18328 10489 18362 10523
rect 2421 10421 2455 10455
rect 3525 10421 3559 10455
rect 5733 10421 5767 10455
rect 10425 10421 10459 10455
rect 10517 10421 10551 10455
rect 11713 10421 11747 10455
rect 13829 10421 13863 10455
rect 14657 10421 14691 10455
rect 15485 10421 15519 10455
rect 15945 10421 15979 10455
rect 16865 10421 16899 10455
rect 16957 10421 16991 10455
rect 21097 10421 21131 10455
rect 4261 10217 4295 10251
rect 4629 10217 4663 10251
rect 5273 10217 5307 10251
rect 8125 10217 8159 10251
rect 8585 10217 8619 10251
rect 11069 10217 11103 10251
rect 11621 10217 11655 10251
rect 11989 10217 12023 10251
rect 12633 10217 12667 10251
rect 13093 10217 13127 10251
rect 14841 10217 14875 10251
rect 15853 10217 15887 10251
rect 16497 10217 16531 10251
rect 16865 10217 16899 10251
rect 17509 10217 17543 10251
rect 20361 10217 20395 10251
rect 4721 10149 4755 10183
rect 8493 10149 8527 10183
rect 13001 10149 13035 10183
rect 15945 10149 15979 10183
rect 16957 10149 16991 10183
rect 17969 10149 18003 10183
rect 1777 10081 1811 10115
rect 2044 10081 2078 10115
rect 5641 10081 5675 10115
rect 6736 10081 6770 10115
rect 9689 10081 9723 10115
rect 9956 10081 9990 10115
rect 13645 10081 13679 10115
rect 14565 10081 14599 10115
rect 15025 10081 15059 10115
rect 17877 10081 17911 10115
rect 18705 10081 18739 10115
rect 18972 10081 19006 10115
rect 4905 10013 4939 10047
rect 5733 10013 5767 10047
rect 5825 10013 5859 10047
rect 6469 10013 6503 10047
rect 8677 10013 8711 10047
rect 12081 10013 12115 10047
rect 12173 10013 12207 10047
rect 13185 10013 13219 10047
rect 13829 10013 13863 10047
rect 16037 10013 16071 10047
rect 17049 10013 17083 10047
rect 18153 10013 18187 10047
rect 7849 9945 7883 9979
rect 14381 9945 14415 9979
rect 15485 9945 15519 9979
rect 3157 9877 3191 9911
rect 20085 9877 20119 9911
rect 1869 9673 1903 9707
rect 10241 9673 10275 9707
rect 10517 9673 10551 9707
rect 14197 9673 14231 9707
rect 2881 9605 2915 9639
rect 5549 9605 5583 9639
rect 6837 9605 6871 9639
rect 16957 9605 16991 9639
rect 2329 9537 2363 9571
rect 2513 9537 2547 9571
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 4537 9537 4571 9571
rect 6193 9537 6227 9571
rect 7481 9537 7515 9571
rect 8309 9537 8343 9571
rect 8401 9537 8435 9571
rect 8861 9537 8895 9571
rect 10425 9537 10459 9571
rect 11069 9537 11103 9571
rect 11805 9537 11839 9571
rect 11989 9537 12023 9571
rect 14841 9537 14875 9571
rect 15761 9537 15795 9571
rect 17509 9537 17543 9571
rect 19717 9537 19751 9571
rect 2237 9469 2271 9503
rect 4353 9469 4387 9503
rect 5917 9469 5951 9503
rect 10977 9469 11011 9503
rect 12449 9469 12483 9503
rect 19984 9469 20018 9503
rect 8217 9401 8251 9435
rect 9128 9401 9162 9435
rect 10425 9401 10459 9435
rect 12716 9401 12750 9435
rect 14657 9401 14691 9435
rect 15577 9401 15611 9435
rect 16221 9401 16255 9435
rect 3249 9333 3283 9367
rect 3985 9333 4019 9367
rect 4445 9333 4479 9367
rect 6009 9333 6043 9367
rect 7205 9333 7239 9367
rect 7297 9333 7331 9367
rect 7849 9333 7883 9367
rect 10885 9333 10919 9367
rect 11345 9333 11379 9367
rect 11713 9333 11747 9367
rect 13829 9333 13863 9367
rect 14565 9333 14599 9367
rect 15209 9333 15243 9367
rect 15669 9333 15703 9367
rect 17325 9333 17359 9367
rect 17417 9333 17451 9367
rect 21097 9333 21131 9367
rect 2053 9129 2087 9163
rect 2421 9129 2455 9163
rect 3065 9129 3099 9163
rect 4445 9129 4479 9163
rect 13921 9129 13955 9163
rect 14197 9129 14231 9163
rect 15025 9129 15059 9163
rect 16681 9129 16715 9163
rect 19809 9129 19843 9163
rect 20453 9129 20487 9163
rect 9045 9061 9079 9095
rect 12449 9061 12483 9095
rect 17325 9061 17359 9095
rect 4813 8993 4847 9027
rect 5457 8993 5491 9027
rect 6193 8993 6227 9027
rect 6460 8993 6494 9027
rect 8033 8993 8067 9027
rect 8493 8993 8527 9027
rect 8953 8993 8987 9027
rect 10057 8993 10091 9027
rect 10701 8993 10735 9027
rect 12541 8993 12575 9027
rect 12808 8993 12842 9027
rect 14565 8993 14599 9027
rect 15025 8993 15059 9027
rect 15557 8993 15591 9027
rect 18696 8993 18730 9027
rect 20269 8993 20303 9027
rect 2513 8925 2547 8959
rect 2697 8925 2731 8959
rect 4905 8925 4939 8959
rect 5089 8925 5123 8959
rect 9137 8925 9171 8959
rect 10149 8925 10183 8959
rect 10241 8925 10275 8959
rect 14657 8925 14691 8959
rect 14841 8925 14875 8959
rect 15301 8925 15335 8959
rect 17417 8925 17451 8959
rect 17509 8925 17543 8959
rect 18429 8925 18463 8959
rect 7573 8857 7607 8891
rect 7849 8857 7883 8891
rect 8309 8789 8343 8823
rect 8585 8789 8619 8823
rect 9689 8789 9723 8823
rect 16957 8789 16991 8823
rect 4169 8585 4203 8619
rect 6837 8585 6871 8619
rect 9873 8585 9907 8619
rect 12081 8585 12115 8619
rect 18981 8585 19015 8619
rect 14841 8517 14875 8551
rect 15209 8517 15243 8551
rect 4721 8449 4755 8483
rect 5825 8449 5859 8483
rect 7297 8449 7331 8483
rect 7481 8449 7515 8483
rect 8033 8449 8067 8483
rect 12173 8449 12207 8483
rect 13001 8449 13035 8483
rect 15669 8449 15703 8483
rect 15761 8449 15795 8483
rect 17417 8449 17451 8483
rect 19625 8449 19659 8483
rect 20545 8449 20579 8483
rect 1869 8381 1903 8415
rect 4537 8381 4571 8415
rect 8493 8381 8527 8415
rect 10701 8381 10735 8415
rect 13461 8381 13495 8415
rect 17141 8381 17175 8415
rect 2136 8313 2170 8347
rect 5641 8313 5675 8347
rect 7205 8313 7239 8347
rect 8760 8313 8794 8347
rect 10968 8313 11002 8347
rect 12173 8313 12207 8347
rect 12909 8313 12943 8347
rect 13728 8313 13762 8347
rect 15577 8313 15611 8347
rect 17233 8313 17267 8347
rect 19349 8313 19383 8347
rect 20361 8313 20395 8347
rect 3249 8245 3283 8279
rect 4629 8245 4663 8279
rect 5181 8245 5215 8279
rect 5549 8245 5583 8279
rect 6285 8245 6319 8279
rect 12449 8245 12483 8279
rect 12817 8245 12851 8279
rect 16773 8245 16807 8279
rect 19441 8245 19475 8279
rect 19993 8245 20027 8279
rect 20453 8245 20487 8279
rect 1961 8041 1995 8075
rect 2973 8041 3007 8075
rect 4537 8041 4571 8075
rect 5273 8041 5307 8075
rect 5641 8041 5675 8075
rect 6745 8041 6779 8075
rect 7389 8041 7423 8075
rect 8953 8041 8987 8075
rect 9045 8041 9079 8075
rect 10149 8041 10183 8075
rect 10609 8041 10643 8075
rect 13369 8041 13403 8075
rect 14197 8041 14231 8075
rect 14565 8041 14599 8075
rect 19073 8041 19107 8075
rect 19717 8041 19751 8075
rect 20913 8041 20947 8075
rect 2329 7973 2363 8007
rect 3433 7973 3467 8007
rect 7757 7973 7791 8007
rect 11989 7973 12023 8007
rect 13737 7973 13771 8007
rect 16028 7973 16062 8007
rect 17960 7973 17994 8007
rect 3341 7905 3375 7939
rect 4445 7905 4479 7939
rect 7849 7905 7883 7939
rect 10517 7905 10551 7939
rect 11897 7905 11931 7939
rect 12909 7905 12943 7939
rect 15669 7905 15703 7939
rect 20085 7905 20119 7939
rect 2421 7837 2455 7871
rect 2605 7837 2639 7871
rect 3617 7837 3651 7871
rect 4629 7837 4663 7871
rect 5733 7837 5767 7871
rect 5917 7837 5951 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 7941 7837 7975 7871
rect 9137 7837 9171 7871
rect 10701 7837 10735 7871
rect 12081 7837 12115 7871
rect 13001 7837 13035 7871
rect 13093 7837 13127 7871
rect 13829 7837 13863 7871
rect 14013 7837 14047 7871
rect 14657 7837 14691 7871
rect 14749 7837 14783 7871
rect 15761 7837 15795 7871
rect 17693 7837 17727 7871
rect 20177 7837 20211 7871
rect 20361 7837 20395 7871
rect 6377 7769 6411 7803
rect 8585 7769 8619 7803
rect 12541 7769 12575 7803
rect 4077 7701 4111 7735
rect 11529 7701 11563 7735
rect 15485 7701 15519 7735
rect 17141 7701 17175 7735
rect 2145 7497 2179 7531
rect 4905 7497 4939 7531
rect 9873 7497 9907 7531
rect 10149 7497 10183 7531
rect 15025 7497 15059 7531
rect 15209 7497 15243 7531
rect 17693 7497 17727 7531
rect 18705 7497 18739 7531
rect 7941 7429 7975 7463
rect 2789 7361 2823 7395
rect 3709 7361 3743 7395
rect 5457 7361 5491 7395
rect 7481 7361 7515 7395
rect 10701 7361 10735 7395
rect 11713 7361 11747 7395
rect 13001 7361 13035 7395
rect 15209 7361 15243 7395
rect 15853 7361 15887 7395
rect 19257 7361 19291 7395
rect 20361 7361 20395 7395
rect 3525 7293 3559 7327
rect 8125 7293 8159 7327
rect 8493 7293 8527 7327
rect 8760 7293 8794 7327
rect 12817 7293 12851 7327
rect 13645 7293 13679 7327
rect 16313 7293 16347 7327
rect 18153 7293 18187 7327
rect 20729 7293 20763 7327
rect 2513 7225 2547 7259
rect 7389 7225 7423 7259
rect 11621 7225 11655 7259
rect 13912 7225 13946 7259
rect 15761 7225 15795 7259
rect 16580 7225 16614 7259
rect 19073 7225 19107 7259
rect 2605 7157 2639 7191
rect 3157 7157 3191 7191
rect 3617 7157 3651 7191
rect 5273 7157 5307 7191
rect 5365 7157 5399 7191
rect 6929 7157 6963 7191
rect 7297 7157 7331 7191
rect 10517 7157 10551 7191
rect 10609 7157 10643 7191
rect 11161 7157 11195 7191
rect 11529 7157 11563 7191
rect 12449 7157 12483 7191
rect 12909 7157 12943 7191
rect 15301 7157 15335 7191
rect 15669 7157 15703 7191
rect 19165 7157 19199 7191
rect 19717 7157 19751 7191
rect 20085 7157 20119 7191
rect 20177 7157 20211 7191
rect 20913 7157 20947 7191
rect 3065 6953 3099 6987
rect 7573 6953 7607 6987
rect 9873 6953 9907 6987
rect 16589 6953 16623 6987
rect 19901 6953 19935 6987
rect 8585 6885 8619 6919
rect 10241 6885 10275 6919
rect 13553 6885 13587 6919
rect 14565 6885 14599 6919
rect 17509 6885 17543 6919
rect 18889 6885 18923 6919
rect 1685 6817 1719 6851
rect 1952 6817 1986 6851
rect 4988 6817 5022 6851
rect 8677 6817 8711 6851
rect 11336 6817 11370 6851
rect 12909 6817 12943 6851
rect 13001 6817 13035 6851
rect 14657 6817 14691 6851
rect 15301 6817 15335 6851
rect 16037 6817 16071 6851
rect 16497 6817 16531 6851
rect 18981 6817 19015 6851
rect 4721 6749 4755 6783
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 8861 6749 8895 6783
rect 10333 6749 10367 6783
rect 10425 6749 10459 6783
rect 11069 6749 11103 6783
rect 13645 6749 13679 6783
rect 13829 6749 13863 6783
rect 14749 6749 14783 6783
rect 16681 6749 16715 6783
rect 17601 6749 17635 6783
rect 17785 6749 17819 6783
rect 19073 6749 19107 6783
rect 19993 6749 20027 6783
rect 20177 6749 20211 6783
rect 13001 6681 13035 6715
rect 13185 6681 13219 6715
rect 14197 6681 14231 6715
rect 15853 6681 15887 6715
rect 16129 6681 16163 6715
rect 17141 6681 17175 6715
rect 18521 6681 18555 6715
rect 19533 6681 19567 6715
rect 6101 6613 6135 6647
rect 7205 6613 7239 6647
rect 8217 6613 8251 6647
rect 12449 6613 12483 6647
rect 12725 6613 12759 6647
rect 3525 6409 3559 6443
rect 4905 6409 4939 6443
rect 6837 6409 6871 6443
rect 17601 6409 17635 6443
rect 20269 6409 20303 6443
rect 5917 6341 5951 6375
rect 11161 6341 11195 6375
rect 2145 6273 2179 6307
rect 4353 6273 4387 6307
rect 5365 6273 5399 6307
rect 5457 6273 5491 6307
rect 6285 6273 6319 6307
rect 7481 6273 7515 6307
rect 11897 6273 11931 6307
rect 16681 6273 16715 6307
rect 18705 6273 18739 6307
rect 19625 6273 19659 6307
rect 20821 6273 20855 6307
rect 6101 6205 6135 6239
rect 8125 6205 8159 6239
rect 9781 6205 9815 6239
rect 12449 6205 12483 6239
rect 12716 6205 12750 6239
rect 14381 6205 14415 6239
rect 16497 6205 16531 6239
rect 17417 6205 17451 6239
rect 19441 6205 19475 6239
rect 20729 6205 20763 6239
rect 2412 6137 2446 6171
rect 4169 6137 4203 6171
rect 8370 6137 8404 6171
rect 10026 6137 10060 6171
rect 14648 6137 14682 6171
rect 18429 6137 18463 6171
rect 1685 6069 1719 6103
rect 3801 6069 3835 6103
rect 4261 6069 4295 6103
rect 5273 6069 5307 6103
rect 7205 6069 7239 6103
rect 7297 6069 7331 6103
rect 9505 6069 9539 6103
rect 13829 6069 13863 6103
rect 15761 6069 15795 6103
rect 16037 6069 16071 6103
rect 16405 6069 16439 6103
rect 18061 6069 18095 6103
rect 18521 6069 18555 6103
rect 19073 6069 19107 6103
rect 19533 6069 19567 6103
rect 20637 6069 20671 6103
rect 1961 5865 1995 5899
rect 2329 5865 2363 5899
rect 5825 5865 5859 5899
rect 6193 5865 6227 5899
rect 6285 5865 6319 5899
rect 8953 5865 8987 5899
rect 10701 5865 10735 5899
rect 12081 5865 12115 5899
rect 17325 5865 17359 5899
rect 19257 5865 19291 5899
rect 4322 5797 4356 5831
rect 7104 5797 7138 5831
rect 11069 5797 11103 5831
rect 16190 5797 16224 5831
rect 17868 5797 17902 5831
rect 10057 5729 10091 5763
rect 12633 5729 12667 5763
rect 12725 5729 12759 5763
rect 12992 5729 13026 5763
rect 14381 5729 14415 5763
rect 19625 5729 19659 5763
rect 20269 5729 20303 5763
rect 2421 5661 2455 5695
rect 2605 5661 2639 5695
rect 4084 5661 4118 5695
rect 6377 5661 6411 5695
rect 6837 5661 6871 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 11161 5661 11195 5695
rect 11345 5661 11379 5695
rect 12173 5661 12207 5695
rect 12357 5661 12391 5695
rect 15945 5661 15979 5695
rect 17601 5661 17635 5695
rect 19717 5661 19751 5695
rect 19809 5661 19843 5695
rect 5457 5525 5491 5559
rect 8217 5525 8251 5559
rect 8585 5525 8619 5559
rect 9689 5525 9723 5559
rect 11713 5525 11747 5559
rect 12633 5525 12667 5559
rect 14105 5525 14139 5559
rect 18981 5525 19015 5559
rect 20453 5525 20487 5559
rect 2053 5321 2087 5355
rect 7297 5321 7331 5355
rect 8585 5321 8619 5355
rect 10149 5321 10183 5355
rect 13093 5321 13127 5355
rect 17141 5321 17175 5355
rect 18061 5321 18095 5355
rect 21005 5321 21039 5355
rect 17601 5253 17635 5287
rect 2605 5185 2639 5219
rect 5365 5185 5399 5219
rect 5549 5185 5583 5219
rect 7849 5185 7883 5219
rect 9137 5185 9171 5219
rect 10793 5185 10827 5219
rect 11713 5185 11747 5219
rect 13645 5185 13679 5219
rect 14565 5185 14599 5219
rect 18613 5185 18647 5219
rect 5273 5117 5307 5151
rect 7757 5117 7791 5151
rect 8493 5117 8527 5151
rect 9045 5117 9079 5151
rect 12449 5117 12483 5151
rect 13461 5117 13495 5151
rect 14381 5117 14415 5151
rect 15209 5117 15243 5151
rect 15761 5117 15795 5151
rect 16028 5117 16062 5151
rect 17417 5117 17451 5151
rect 18521 5117 18555 5151
rect 19073 5117 19107 5151
rect 19625 5117 19659 5151
rect 11529 5049 11563 5083
rect 15025 5049 15059 5083
rect 18429 5049 18463 5083
rect 19870 5049 19904 5083
rect 2421 4981 2455 5015
rect 2513 4981 2547 5015
rect 4905 4981 4939 5015
rect 7665 4981 7699 5015
rect 8309 4981 8343 5015
rect 8953 4981 8987 5015
rect 10517 4981 10551 5015
rect 10609 4981 10643 5015
rect 11161 4981 11195 5015
rect 11621 4981 11655 5015
rect 12633 4981 12667 5015
rect 13553 4981 13587 5015
rect 14013 4981 14047 5015
rect 14473 4981 14507 5015
rect 15393 4981 15427 5015
rect 19257 4981 19291 5015
rect 3709 4777 3743 4811
rect 7205 4777 7239 4811
rect 7573 4777 7607 4811
rect 9689 4777 9723 4811
rect 11161 4777 11195 4811
rect 12081 4777 12115 4811
rect 12173 4777 12207 4811
rect 17785 4777 17819 4811
rect 19809 4777 19843 4811
rect 4620 4709 4654 4743
rect 11069 4709 11103 4743
rect 13636 4709 13670 4743
rect 17233 4709 17267 4743
rect 18674 4709 18708 4743
rect 20361 4709 20395 4743
rect 2329 4641 2363 4675
rect 2596 4641 2630 4675
rect 4353 4641 4387 4675
rect 6377 4641 6411 4675
rect 8585 4641 8619 4675
rect 10057 4641 10091 4675
rect 12817 4641 12851 4675
rect 15669 4641 15703 4675
rect 16773 4641 16807 4675
rect 20085 4641 20119 4675
rect 6469 4573 6503 4607
rect 6561 4573 6595 4607
rect 7665 4573 7699 4607
rect 7757 4573 7791 4607
rect 8677 4573 8711 4607
rect 8769 4573 8803 4607
rect 10149 4573 10183 4607
rect 10241 4573 10275 4607
rect 11345 4573 11379 4607
rect 12357 4573 12391 4607
rect 13369 4573 13403 4607
rect 16865 4573 16899 4607
rect 17049 4573 17083 4607
rect 17233 4573 17267 4607
rect 17877 4573 17911 4607
rect 17969 4573 18003 4607
rect 18429 4573 18463 4607
rect 6009 4505 6043 4539
rect 16405 4505 16439 4539
rect 5733 4437 5767 4471
rect 8217 4437 8251 4471
rect 10701 4437 10735 4471
rect 11713 4437 11747 4471
rect 13001 4437 13035 4471
rect 14749 4437 14783 4471
rect 15853 4437 15887 4471
rect 17417 4437 17451 4471
rect 3249 4233 3283 4267
rect 9045 4233 9079 4267
rect 16865 4233 16899 4267
rect 1869 4097 1903 4131
rect 4077 4097 4111 4131
rect 4997 4097 5031 4131
rect 5181 4097 5215 4131
rect 6101 4097 6135 4131
rect 7665 4097 7699 4131
rect 9689 4097 9723 4131
rect 11897 4097 11931 4131
rect 12909 4097 12943 4131
rect 13001 4097 13035 4131
rect 16497 4097 16531 4131
rect 17509 4097 17543 4131
rect 18705 4097 18739 4131
rect 19717 4097 19751 4131
rect 20637 4097 20671 4131
rect 2136 4029 2170 4063
rect 7932 4029 7966 4063
rect 9413 4029 9447 4063
rect 10241 4029 10275 4063
rect 10508 4029 10542 4063
rect 11713 4029 11747 4063
rect 13737 4029 13771 4063
rect 16221 4029 16255 4063
rect 17233 4029 17267 4063
rect 19441 4029 19475 4063
rect 20453 4029 20487 4063
rect 3893 3961 3927 3995
rect 12817 3961 12851 3995
rect 14004 3961 14038 3995
rect 16313 3961 16347 3995
rect 18429 3961 18463 3995
rect 3525 3893 3559 3927
rect 3985 3893 4019 3927
rect 4537 3893 4571 3927
rect 4905 3893 4939 3927
rect 5549 3893 5583 3927
rect 5917 3893 5951 3927
rect 6009 3893 6043 3927
rect 11621 3893 11655 3927
rect 11713 3893 11747 3927
rect 12449 3893 12483 3927
rect 15117 3893 15151 3927
rect 15393 3893 15427 3927
rect 15853 3893 15887 3927
rect 17325 3893 17359 3927
rect 18061 3893 18095 3927
rect 18521 3893 18555 3927
rect 19073 3893 19107 3927
rect 19533 3893 19567 3927
rect 20085 3893 20119 3927
rect 20545 3893 20579 3927
rect 3065 3689 3099 3723
rect 10977 3689 11011 3723
rect 11529 3689 11563 3723
rect 11897 3689 11931 3723
rect 13001 3689 13035 3723
rect 14565 3689 14599 3723
rect 15301 3689 15335 3723
rect 15669 3689 15703 3723
rect 15761 3689 15795 3723
rect 17785 3689 17819 3723
rect 18521 3689 18555 3723
rect 18981 3689 19015 3723
rect 19809 3689 19843 3723
rect 9965 3621 9999 3655
rect 10885 3621 10919 3655
rect 11989 3621 12023 3655
rect 14657 3621 14691 3655
rect 16672 3621 16706 3655
rect 18889 3621 18923 3655
rect 2973 3553 3007 3587
rect 4445 3553 4479 3587
rect 5825 3553 5859 3587
rect 6092 3553 6126 3587
rect 8585 3553 8619 3587
rect 8677 3553 8711 3587
rect 9689 3553 9723 3587
rect 12909 3553 12943 3587
rect 13645 3553 13679 3587
rect 16405 3553 16439 3587
rect 20177 3553 20211 3587
rect 3249 3485 3283 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 7481 3485 7515 3519
rect 8769 3485 8803 3519
rect 11161 3485 11195 3519
rect 12173 3485 12207 3519
rect 13093 3485 13127 3519
rect 14841 3485 14875 3519
rect 15853 3485 15887 3519
rect 18061 3485 18095 3519
rect 19073 3485 19107 3519
rect 20269 3485 20303 3519
rect 20453 3485 20487 3519
rect 2605 3417 2639 3451
rect 8217 3417 8251 3451
rect 10517 3417 10551 3451
rect 13829 3417 13863 3451
rect 4077 3349 4111 3383
rect 7205 3349 7239 3383
rect 12541 3349 12575 3383
rect 14197 3349 14231 3383
rect 2421 3145 2455 3179
rect 3341 3145 3375 3179
rect 4813 3145 4847 3179
rect 5733 3145 5767 3179
rect 8217 3145 8251 3179
rect 8677 3145 8711 3179
rect 16589 3145 16623 3179
rect 3065 3009 3099 3043
rect 2789 2941 2823 2975
rect 5089 3009 5123 3043
rect 6377 3009 6411 3043
rect 13645 3009 13679 3043
rect 17417 3009 17451 3043
rect 17601 3009 17635 3043
rect 18061 3009 18095 3043
rect 20453 3009 20487 3043
rect 3433 2941 3467 2975
rect 6837 2941 6871 2975
rect 8493 2941 8527 2975
rect 9045 2941 9079 2975
rect 10701 2941 10735 2975
rect 12633 2941 12667 2975
rect 13369 2941 13403 2975
rect 14105 2941 14139 2975
rect 14841 2941 14875 2975
rect 15577 2941 15611 2975
rect 16405 2941 16439 2975
rect 17325 2941 17359 2975
rect 20269 2941 20303 2975
rect 3678 2873 3712 2907
rect 7082 2873 7116 2907
rect 9312 2873 9346 2907
rect 10968 2873 11002 2907
rect 12909 2873 12943 2907
rect 14381 2873 14415 2907
rect 15117 2873 15151 2907
rect 15853 2873 15887 2907
rect 18328 2873 18362 2907
rect 2881 2805 2915 2839
rect 3341 2805 3375 2839
rect 6101 2805 6135 2839
rect 6193 2805 6227 2839
rect 10425 2805 10459 2839
rect 12081 2805 12115 2839
rect 16957 2805 16991 2839
rect 19441 2805 19475 2839
rect 4077 2601 4111 2635
rect 6285 2601 6319 2635
rect 7297 2601 7331 2635
rect 8217 2601 8251 2635
rect 8585 2601 8619 2635
rect 9781 2601 9815 2635
rect 10241 2601 10275 2635
rect 12817 2601 12851 2635
rect 14473 2601 14507 2635
rect 16221 2601 16255 2635
rect 17325 2601 17359 2635
rect 17877 2601 17911 2635
rect 18613 2601 18647 2635
rect 18981 2601 19015 2635
rect 19625 2601 19659 2635
rect 19993 2601 20027 2635
rect 6193 2533 6227 2567
rect 11069 2533 11103 2567
rect 4445 2465 4479 2499
rect 8677 2465 8711 2499
rect 10149 2465 10183 2499
rect 10793 2465 10827 2499
rect 11529 2465 11563 2499
rect 12633 2465 12667 2499
rect 13185 2465 13219 2499
rect 13737 2465 13771 2499
rect 14289 2465 14323 2499
rect 14841 2465 14875 2499
rect 15485 2465 15519 2499
rect 16037 2465 16071 2499
rect 16589 2465 16623 2499
rect 17141 2465 17175 2499
rect 17693 2465 17727 2499
rect 19073 2465 19107 2499
rect 20085 2465 20119 2499
rect 4537 2397 4571 2431
rect 4721 2397 4755 2431
rect 6469 2397 6503 2431
rect 7389 2397 7423 2431
rect 7573 2397 7607 2431
rect 8861 2397 8895 2431
rect 10333 2397 10367 2431
rect 11713 2397 11747 2431
rect 19165 2397 19199 2431
rect 20177 2397 20211 2431
rect 6929 2329 6963 2363
rect 13369 2329 13403 2363
rect 15025 2329 15059 2363
rect 5825 2261 5859 2295
rect 13921 2261 13955 2295
rect 15669 2261 15703 2295
rect 16773 2261 16807 2295
<< metal1 >>
rect 1104 20154 21620 20176
rect 1104 20102 7846 20154
rect 7898 20102 7910 20154
rect 7962 20102 7974 20154
rect 8026 20102 8038 20154
rect 8090 20102 14710 20154
rect 14762 20102 14774 20154
rect 14826 20102 14838 20154
rect 14890 20102 14902 20154
rect 14954 20102 21620 20154
rect 1104 20080 21620 20102
rect 1104 19610 21620 19632
rect 1104 19558 4414 19610
rect 4466 19558 4478 19610
rect 4530 19558 4542 19610
rect 4594 19558 4606 19610
rect 4658 19558 11278 19610
rect 11330 19558 11342 19610
rect 11394 19558 11406 19610
rect 11458 19558 11470 19610
rect 11522 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 18270 19610
rect 18322 19558 18334 19610
rect 18386 19558 21620 19610
rect 1104 19536 21620 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 5997 19499 6055 19505
rect 5997 19496 6009 19499
rect 3752 19468 6009 19496
rect 3752 19456 3758 19468
rect 5997 19465 6009 19468
rect 6043 19465 6055 19499
rect 19150 19496 19156 19508
rect 19111 19468 19156 19496
rect 5997 19459 6055 19465
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 20714 19496 20720 19508
rect 20675 19468 20720 19496
rect 20714 19456 20720 19468
rect 20772 19456 20778 19508
rect 1765 19295 1823 19301
rect 1765 19261 1777 19295
rect 1811 19261 1823 19295
rect 1765 19255 1823 19261
rect 2317 19295 2375 19301
rect 2317 19261 2329 19295
rect 2363 19292 2375 19295
rect 4798 19292 4804 19304
rect 2363 19264 4804 19292
rect 2363 19261 2375 19264
rect 2317 19255 2375 19261
rect 1780 19224 1808 19255
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 5810 19292 5816 19304
rect 5771 19264 5816 19292
rect 5810 19252 5816 19264
rect 5868 19252 5874 19304
rect 18414 19252 18420 19304
rect 18472 19292 18478 19304
rect 18969 19295 19027 19301
rect 18969 19292 18981 19295
rect 18472 19264 18981 19292
rect 18472 19252 18478 19264
rect 18969 19261 18981 19264
rect 19015 19261 19027 19295
rect 20530 19292 20536 19304
rect 20491 19264 20536 19292
rect 18969 19255 19027 19261
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 4890 19224 4896 19236
rect 1780 19196 4896 19224
rect 4890 19184 4896 19196
rect 4948 19184 4954 19236
rect 2501 19159 2559 19165
rect 2501 19125 2513 19159
rect 2547 19156 2559 19159
rect 2774 19156 2780 19168
rect 2547 19128 2780 19156
rect 2547 19125 2559 19128
rect 2501 19119 2559 19125
rect 2774 19116 2780 19128
rect 2832 19116 2838 19168
rect 1104 19066 21620 19088
rect 1104 19014 7846 19066
rect 7898 19014 7910 19066
rect 7962 19014 7974 19066
rect 8026 19014 8038 19066
rect 8090 19014 14710 19066
rect 14762 19014 14774 19066
rect 14826 19014 14838 19066
rect 14890 19014 14902 19066
rect 14954 19014 21620 19066
rect 1104 18992 21620 19014
rect 1946 18952 1952 18964
rect 1907 18924 1952 18952
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6365 18887 6423 18893
rect 6365 18884 6377 18887
rect 5868 18856 6377 18884
rect 5868 18844 5874 18856
rect 6365 18853 6377 18856
rect 6411 18853 6423 18887
rect 18414 18884 18420 18896
rect 18375 18856 18420 18884
rect 6365 18847 6423 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 1765 18819 1823 18825
rect 1765 18785 1777 18819
rect 1811 18816 1823 18819
rect 6086 18816 6092 18828
rect 1811 18788 5856 18816
rect 6047 18788 6092 18816
rect 1811 18785 1823 18788
rect 1765 18779 1823 18785
rect 5828 18760 5856 18788
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18012 18788 18153 18816
rect 18012 18776 18018 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 5810 18708 5816 18760
rect 5868 18708 5874 18760
rect 1104 18522 21620 18544
rect 1104 18470 4414 18522
rect 4466 18470 4478 18522
rect 4530 18470 4542 18522
rect 4594 18470 4606 18522
rect 4658 18470 11278 18522
rect 11330 18470 11342 18522
rect 11394 18470 11406 18522
rect 11458 18470 11470 18522
rect 11522 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 18270 18522
rect 18322 18470 18334 18522
rect 18386 18470 21620 18522
rect 1104 18448 21620 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 20714 18408 20720 18420
rect 20675 18380 20720 18408
rect 20714 18368 20720 18380
rect 20772 18368 20778 18420
rect 1762 18204 1768 18216
rect 1723 18176 1768 18204
rect 1762 18164 1768 18176
rect 1820 18164 1826 18216
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 8202 18204 8208 18216
rect 5776 18176 8208 18204
rect 5776 18164 5782 18176
rect 8202 18164 8208 18176
rect 8260 18164 8266 18216
rect 20530 18204 20536 18216
rect 20491 18176 20536 18204
rect 20530 18164 20536 18176
rect 20588 18164 20594 18216
rect 1104 17978 21620 18000
rect 1104 17926 7846 17978
rect 7898 17926 7910 17978
rect 7962 17926 7974 17978
rect 8026 17926 8038 17978
rect 8090 17926 14710 17978
rect 14762 17926 14774 17978
rect 14826 17926 14838 17978
rect 14890 17926 14902 17978
rect 14954 17926 21620 17978
rect 1104 17904 21620 17926
rect 1854 17864 1860 17876
rect 1815 17836 1860 17864
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 1762 17756 1768 17808
rect 1820 17796 1826 17808
rect 2501 17799 2559 17805
rect 2501 17796 2513 17799
rect 1820 17768 2513 17796
rect 1820 17756 1826 17768
rect 2501 17765 2513 17768
rect 2547 17765 2559 17799
rect 2501 17759 2559 17765
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 20530 17796 20536 17808
rect 20027 17768 20536 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 20530 17756 20536 17768
rect 20588 17756 20594 17808
rect 1673 17731 1731 17737
rect 1673 17697 1685 17731
rect 1719 17697 1731 17731
rect 1673 17691 1731 17697
rect 2225 17731 2283 17737
rect 2225 17697 2237 17731
rect 2271 17728 2283 17731
rect 6638 17728 6644 17740
rect 2271 17700 6644 17728
rect 2271 17697 2283 17700
rect 2225 17691 2283 17697
rect 1688 17660 1716 17691
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 19702 17728 19708 17740
rect 19663 17700 19708 17728
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 7466 17660 7472 17672
rect 1688 17632 7472 17660
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 1104 17434 21620 17456
rect 1104 17382 4414 17434
rect 4466 17382 4478 17434
rect 4530 17382 4542 17434
rect 4594 17382 4606 17434
rect 4658 17382 11278 17434
rect 11330 17382 11342 17434
rect 11394 17382 11406 17434
rect 11458 17382 11470 17434
rect 11522 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 18270 17434
rect 18322 17382 18334 17434
rect 18386 17382 21620 17434
rect 1104 17360 21620 17382
rect 1670 17280 1676 17332
rect 1728 17320 1734 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1728 17292 1961 17320
rect 1728 17280 1734 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 20714 17320 20720 17332
rect 20675 17292 20720 17320
rect 1949 17283 2007 17289
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 1765 17119 1823 17125
rect 1765 17085 1777 17119
rect 1811 17116 1823 17119
rect 6454 17116 6460 17128
rect 1811 17088 6460 17116
rect 1811 17085 1823 17088
rect 1765 17079 1823 17085
rect 6454 17076 6460 17088
rect 6512 17076 6518 17128
rect 19978 17076 19984 17128
rect 20036 17116 20042 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20036 17088 20545 17116
rect 20036 17076 20042 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 1104 16890 21620 16912
rect 1104 16838 7846 16890
rect 7898 16838 7910 16890
rect 7962 16838 7974 16890
rect 8026 16838 8038 16890
rect 8090 16838 14710 16890
rect 14762 16838 14774 16890
rect 14826 16838 14838 16890
rect 14890 16838 14902 16890
rect 14954 16838 21620 16890
rect 1104 16816 21620 16838
rect 1946 16776 1952 16788
rect 1907 16748 1952 16776
rect 1946 16736 1952 16748
rect 2004 16736 2010 16788
rect 20438 16776 20444 16788
rect 20399 16748 20444 16776
rect 20438 16736 20444 16748
rect 20496 16736 20502 16788
rect 1765 16643 1823 16649
rect 1765 16609 1777 16643
rect 1811 16640 1823 16643
rect 5350 16640 5356 16652
rect 1811 16612 5356 16640
rect 1811 16609 1823 16612
rect 1765 16603 1823 16609
rect 5350 16600 5356 16612
rect 5408 16600 5414 16652
rect 20257 16643 20315 16649
rect 20257 16609 20269 16643
rect 20303 16640 20315 16643
rect 20530 16640 20536 16652
rect 20303 16612 20536 16640
rect 20303 16609 20315 16612
rect 20257 16603 20315 16609
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 1104 16346 21620 16368
rect 1104 16294 4414 16346
rect 4466 16294 4478 16346
rect 4530 16294 4542 16346
rect 4594 16294 4606 16346
rect 4658 16294 11278 16346
rect 11330 16294 11342 16346
rect 11394 16294 11406 16346
rect 11458 16294 11470 16346
rect 11522 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 18270 16346
rect 18322 16294 18334 16346
rect 18386 16294 21620 16346
rect 1104 16272 21620 16294
rect 1946 16232 1952 16244
rect 1907 16204 1952 16232
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 2314 16192 2320 16244
rect 2372 16232 2378 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 2372 16204 2513 16232
rect 2372 16192 2378 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 3418 16232 3424 16244
rect 3379 16204 3424 16232
rect 2501 16195 2559 16201
rect 3418 16192 3424 16204
rect 3476 16192 3482 16244
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 17862 16232 17868 16244
rect 13587 16204 17868 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 17862 16192 17868 16204
rect 17920 16192 17926 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20806 16232 20812 16244
rect 20763 16204 20812 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 7282 16096 7288 16108
rect 2332 16068 7288 16096
rect 2332 16037 2360 16068
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 1765 16031 1823 16037
rect 1765 15997 1777 16031
rect 1811 15997 1823 16031
rect 1765 15991 1823 15997
rect 2317 16031 2375 16037
rect 2317 15997 2329 16031
rect 2363 15997 2375 16031
rect 3234 16028 3240 16040
rect 3195 16000 3240 16028
rect 2317 15991 2375 15997
rect 1780 15960 1808 15991
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 12802 15988 12808 16040
rect 12860 16028 12866 16040
rect 13357 16031 13415 16037
rect 13357 16028 13369 16031
rect 12860 16000 13369 16028
rect 12860 15988 12866 16000
rect 13357 15997 13369 16000
rect 13403 15997 13415 16031
rect 13357 15991 13415 15997
rect 19886 15988 19892 16040
rect 19944 16028 19950 16040
rect 19981 16031 20039 16037
rect 19981 16028 19993 16031
rect 19944 16000 19993 16028
rect 19944 15988 19950 16000
rect 19981 15997 19993 16000
rect 20027 15997 20039 16031
rect 19981 15991 20039 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 5442 15960 5448 15972
rect 1780 15932 5448 15960
rect 5442 15920 5448 15932
rect 5500 15920 5506 15972
rect 19794 15920 19800 15972
rect 19852 15960 19858 15972
rect 20548 15960 20576 15991
rect 19852 15932 20576 15960
rect 19852 15920 19858 15932
rect 1104 15802 21620 15824
rect 1104 15750 7846 15802
rect 7898 15750 7910 15802
rect 7962 15750 7974 15802
rect 8026 15750 8038 15802
rect 8090 15750 14710 15802
rect 14762 15750 14774 15802
rect 14826 15750 14838 15802
rect 14890 15750 14902 15802
rect 14954 15750 21620 15802
rect 1104 15728 21620 15750
rect 1946 15688 1952 15700
rect 1907 15660 1952 15688
rect 1946 15648 1952 15660
rect 2004 15648 2010 15700
rect 2498 15688 2504 15700
rect 2459 15660 2504 15688
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 20438 15688 20444 15700
rect 20399 15660 20444 15688
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 3234 15580 3240 15632
rect 3292 15620 3298 15632
rect 4341 15623 4399 15629
rect 4341 15620 4353 15623
rect 3292 15592 4353 15620
rect 3292 15580 3298 15592
rect 4341 15589 4353 15592
rect 4387 15589 4399 15623
rect 12802 15620 12808 15632
rect 12763 15592 12808 15620
rect 4341 15583 4399 15589
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 1765 15555 1823 15561
rect 1765 15521 1777 15555
rect 1811 15521 1823 15555
rect 1765 15515 1823 15521
rect 2317 15555 2375 15561
rect 2317 15521 2329 15555
rect 2363 15521 2375 15555
rect 2317 15515 2375 15521
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4246 15552 4252 15564
rect 4111 15524 4252 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 1780 15416 1808 15515
rect 2332 15484 2360 15515
rect 4246 15512 4252 15524
rect 4304 15512 4310 15564
rect 12526 15552 12532 15564
rect 12487 15524 12532 15552
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 20070 15512 20076 15564
rect 20128 15552 20134 15564
rect 20257 15555 20315 15561
rect 20257 15552 20269 15555
rect 20128 15524 20269 15552
rect 20128 15512 20134 15524
rect 20257 15521 20269 15524
rect 20303 15521 20315 15555
rect 20257 15515 20315 15521
rect 5074 15484 5080 15496
rect 2332 15456 5080 15484
rect 5074 15444 5080 15456
rect 5132 15444 5138 15496
rect 4154 15416 4160 15428
rect 1780 15388 4160 15416
rect 4154 15376 4160 15388
rect 4212 15376 4218 15428
rect 1104 15258 21620 15280
rect 1104 15206 4414 15258
rect 4466 15206 4478 15258
rect 4530 15206 4542 15258
rect 4594 15206 4606 15258
rect 4658 15206 11278 15258
rect 11330 15206 11342 15258
rect 11394 15206 11406 15258
rect 11458 15206 11470 15258
rect 11522 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 18270 15258
rect 18322 15206 18334 15258
rect 18386 15206 21620 15258
rect 1104 15184 21620 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15144 2559 15147
rect 2774 15144 2780 15156
rect 2547 15116 2780 15144
rect 2547 15113 2559 15116
rect 2501 15107 2559 15113
rect 2774 15104 2780 15116
rect 2832 15104 2838 15156
rect 20165 15147 20223 15153
rect 20165 15113 20177 15147
rect 20211 15144 20223 15147
rect 20254 15144 20260 15156
rect 20211 15116 20260 15144
rect 20211 15113 20223 15116
rect 20165 15107 20223 15113
rect 20254 15104 20260 15116
rect 20312 15104 20318 15156
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 20717 15147 20775 15153
rect 20717 15144 20729 15147
rect 20680 15116 20729 15144
rect 20680 15104 20686 15116
rect 20717 15113 20729 15116
rect 20763 15113 20775 15147
rect 20717 15107 20775 15113
rect 1946 15076 1952 15088
rect 1907 15048 1952 15076
rect 1946 15036 1952 15048
rect 2004 15036 2010 15088
rect 13725 15079 13783 15085
rect 13725 15045 13737 15079
rect 13771 15076 13783 15079
rect 15378 15076 15384 15088
rect 13771 15048 15384 15076
rect 13771 15045 13783 15048
rect 13725 15039 13783 15045
rect 15378 15036 15384 15048
rect 15436 15036 15442 15088
rect 19610 15076 19616 15088
rect 19571 15048 19616 15076
rect 19610 15036 19616 15048
rect 19668 15036 19674 15088
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 15008 14427 15011
rect 14550 15008 14556 15020
rect 14415 14980 14556 15008
rect 14415 14977 14427 14980
rect 14369 14971 14427 14977
rect 14550 14968 14556 14980
rect 14608 14968 14614 15020
rect 20346 14968 20352 15020
rect 20404 15008 20410 15020
rect 20622 15008 20628 15020
rect 20404 14980 20628 15008
rect 20404 14968 20410 14980
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 1762 14940 1768 14952
rect 1723 14912 1768 14940
rect 1762 14900 1768 14912
rect 1820 14900 1826 14952
rect 2317 14943 2375 14949
rect 2317 14909 2329 14943
rect 2363 14940 2375 14943
rect 2590 14940 2596 14952
rect 2363 14912 2596 14940
rect 2363 14909 2375 14912
rect 2317 14903 2375 14909
rect 2590 14900 2596 14912
rect 2648 14900 2654 14952
rect 2774 14900 2780 14952
rect 2832 14940 2838 14952
rect 2961 14943 3019 14949
rect 2961 14940 2973 14943
rect 2832 14912 2973 14940
rect 2832 14900 2838 14912
rect 2961 14909 2973 14912
rect 3007 14909 3019 14943
rect 19426 14940 19432 14952
rect 19387 14912 19432 14940
rect 2961 14903 3019 14909
rect 19426 14900 19432 14912
rect 19484 14900 19490 14952
rect 19981 14943 20039 14949
rect 19981 14909 19993 14943
rect 20027 14909 20039 14943
rect 19981 14903 20039 14909
rect 20533 14943 20591 14949
rect 20533 14909 20545 14943
rect 20579 14909 20591 14943
rect 20533 14903 20591 14909
rect 3228 14875 3286 14881
rect 3228 14841 3240 14875
rect 3274 14872 3286 14875
rect 3786 14872 3792 14884
rect 3274 14844 3792 14872
rect 3274 14841 3286 14844
rect 3228 14835 3286 14841
rect 3786 14832 3792 14844
rect 3844 14832 3850 14884
rect 14090 14872 14096 14884
rect 14051 14844 14096 14872
rect 14090 14832 14096 14844
rect 14148 14832 14154 14884
rect 14274 14832 14280 14884
rect 14332 14872 14338 14884
rect 19996 14872 20024 14903
rect 14332 14844 20024 14872
rect 14332 14832 14338 14844
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 4341 14807 4399 14813
rect 4341 14804 4353 14807
rect 4212 14776 4353 14804
rect 4212 14764 4218 14776
rect 4341 14773 4353 14776
rect 4387 14773 4399 14807
rect 14182 14804 14188 14816
rect 14143 14776 14188 14804
rect 4341 14767 4399 14773
rect 14182 14764 14188 14776
rect 14240 14764 14246 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 20548 14804 20576 14903
rect 16264 14776 20576 14804
rect 16264 14764 16270 14776
rect 1104 14714 21620 14736
rect 1104 14662 7846 14714
rect 7898 14662 7910 14714
rect 7962 14662 7974 14714
rect 8026 14662 8038 14714
rect 8090 14662 14710 14714
rect 14762 14662 14774 14714
rect 14826 14662 14838 14714
rect 14890 14662 14902 14714
rect 14954 14662 21620 14714
rect 1104 14640 21620 14662
rect 1670 14600 1676 14612
rect 1631 14572 1676 14600
rect 1670 14560 1676 14572
rect 1728 14560 1734 14612
rect 3142 14560 3148 14612
rect 3200 14600 3206 14612
rect 4249 14603 4307 14609
rect 4249 14600 4261 14603
rect 3200 14572 4261 14600
rect 3200 14560 3206 14572
rect 4249 14569 4261 14572
rect 4295 14569 4307 14603
rect 4249 14563 4307 14569
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 13449 14603 13507 14609
rect 5132 14572 12204 14600
rect 5132 14560 5138 14572
rect 1762 14492 1768 14544
rect 1820 14532 1826 14544
rect 2317 14535 2375 14541
rect 2317 14532 2329 14535
rect 1820 14504 2329 14532
rect 1820 14492 1826 14504
rect 2317 14501 2329 14504
rect 2363 14501 2375 14535
rect 2317 14495 2375 14501
rect 8202 14492 8208 14544
rect 8260 14532 8266 14544
rect 12038 14535 12096 14541
rect 12038 14532 12050 14535
rect 8260 14504 12050 14532
rect 8260 14492 8266 14504
rect 12038 14501 12050 14504
rect 12084 14501 12096 14535
rect 12176 14532 12204 14572
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 14182 14600 14188 14612
rect 13495 14572 14188 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14182 14560 14188 14572
rect 14240 14560 14246 14612
rect 18874 14600 18880 14612
rect 15028 14572 18880 14600
rect 13817 14535 13875 14541
rect 12176 14504 13308 14532
rect 12038 14495 12096 14501
rect 1486 14464 1492 14476
rect 1447 14436 1492 14464
rect 1486 14424 1492 14436
rect 1544 14424 1550 14476
rect 2041 14467 2099 14473
rect 2041 14433 2053 14467
rect 2087 14464 2099 14467
rect 2087 14436 2820 14464
rect 2087 14433 2099 14436
rect 2041 14427 2099 14433
rect 2792 14337 2820 14436
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 2924 14436 3157 14464
rect 2924 14424 2930 14436
rect 3145 14433 3157 14436
rect 3191 14433 3203 14467
rect 3145 14427 3203 14433
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 5258 14464 5264 14476
rect 4111 14436 5264 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 9766 14424 9772 14476
rect 9824 14464 9830 14476
rect 9933 14467 9991 14473
rect 9933 14464 9945 14467
rect 9824 14436 9945 14464
rect 9824 14424 9830 14436
rect 9933 14433 9945 14436
rect 9979 14433 9991 14467
rect 13280 14464 13308 14504
rect 13817 14501 13829 14535
rect 13863 14532 13875 14535
rect 13998 14532 14004 14544
rect 13863 14504 14004 14532
rect 13863 14501 13875 14504
rect 13817 14495 13875 14501
rect 13998 14492 14004 14504
rect 14056 14492 14062 14544
rect 13909 14467 13967 14473
rect 13909 14464 13921 14467
rect 13280 14436 13921 14464
rect 9933 14427 9991 14433
rect 13909 14433 13921 14436
rect 13955 14464 13967 14467
rect 15028 14464 15056 14572
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 16206 14532 16212 14544
rect 13955 14436 15056 14464
rect 15120 14504 16212 14532
rect 13955 14433 13967 14436
rect 13909 14427 13967 14433
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 4154 14396 4160 14408
rect 3467 14368 4160 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 8444 14368 9689 14396
rect 8444 14356 8450 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 11790 14396 11796 14408
rect 10744 14368 11796 14396
rect 10744 14356 10750 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14458 14396 14464 14408
rect 14139 14368 14464 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14297 2835 14331
rect 15120 14328 15148 14504
rect 16206 14492 16212 14504
rect 16264 14492 16270 14544
rect 16942 14492 16948 14544
rect 17000 14541 17006 14544
rect 17000 14535 17064 14541
rect 17000 14501 17018 14535
rect 17052 14501 17064 14535
rect 17000 14495 17064 14501
rect 17000 14492 17006 14495
rect 19426 14492 19432 14544
rect 19484 14532 19490 14544
rect 19981 14535 20039 14541
rect 19981 14532 19993 14535
rect 19484 14504 19993 14532
rect 19484 14492 19490 14504
rect 19981 14501 19993 14504
rect 20027 14501 20039 14535
rect 19981 14495 20039 14501
rect 16117 14467 16175 14473
rect 16117 14433 16129 14467
rect 16163 14464 16175 14467
rect 17494 14464 17500 14476
rect 16163 14436 17500 14464
rect 16163 14433 16175 14436
rect 16117 14427 16175 14433
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 19153 14467 19211 14473
rect 19153 14433 19165 14467
rect 19199 14464 19211 14467
rect 19610 14464 19616 14476
rect 19199 14436 19616 14464
rect 19199 14433 19211 14436
rect 19153 14427 19211 14433
rect 19610 14424 19616 14436
rect 19668 14424 19674 14476
rect 19705 14467 19763 14473
rect 19705 14433 19717 14467
rect 19751 14433 19763 14467
rect 19705 14427 19763 14433
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16761 14399 16819 14405
rect 16356 14368 16401 14396
rect 16356 14356 16362 14368
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 2777 14291 2835 14297
rect 12728 14300 15148 14328
rect 12728 14272 12756 14300
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 16776 14328 16804 14359
rect 19518 14356 19524 14408
rect 19576 14396 19582 14408
rect 19720 14396 19748 14427
rect 19576 14368 19748 14396
rect 19576 14356 19582 14368
rect 15620 14300 16804 14328
rect 15620 14288 15626 14300
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11057 14263 11115 14269
rect 11057 14260 11069 14263
rect 11020 14232 11069 14260
rect 11020 14220 11026 14232
rect 11057 14229 11069 14232
rect 11103 14229 11115 14263
rect 11057 14223 11115 14229
rect 12710 14220 12716 14272
rect 12768 14220 12774 14272
rect 13173 14263 13231 14269
rect 13173 14229 13185 14263
rect 13219 14260 13231 14263
rect 13630 14260 13636 14272
rect 13219 14232 13636 14260
rect 13219 14229 13231 14232
rect 13173 14223 13231 14229
rect 13630 14220 13636 14232
rect 13688 14220 13694 14272
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14260 15807 14263
rect 16758 14260 16764 14272
rect 15795 14232 16764 14260
rect 15795 14229 15807 14232
rect 15749 14223 15807 14229
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 18141 14263 18199 14269
rect 18141 14229 18153 14263
rect 18187 14260 18199 14263
rect 18506 14260 18512 14272
rect 18187 14232 18512 14260
rect 18187 14229 18199 14232
rect 18141 14223 18199 14229
rect 18506 14220 18512 14232
rect 18564 14220 18570 14272
rect 19334 14260 19340 14272
rect 19295 14232 19340 14260
rect 19334 14220 19340 14232
rect 19392 14220 19398 14272
rect 1104 14170 21620 14192
rect 1104 14118 4414 14170
rect 4466 14118 4478 14170
rect 4530 14118 4542 14170
rect 4594 14118 4606 14170
rect 4658 14118 11278 14170
rect 11330 14118 11342 14170
rect 11394 14118 11406 14170
rect 11458 14118 11470 14170
rect 11522 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 18270 14170
rect 18322 14118 18334 14170
rect 18386 14118 21620 14170
rect 1104 14096 21620 14118
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14056 2375 14059
rect 2774 14056 2780 14068
rect 2363 14028 2780 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 2774 14016 2780 14028
rect 2832 14056 2838 14068
rect 3510 14056 3516 14068
rect 2832 14028 3516 14056
rect 2832 14016 2838 14028
rect 3510 14016 3516 14028
rect 3568 14056 3574 14068
rect 14550 14056 14556 14068
rect 3568 14028 4108 14056
rect 14511 14028 14556 14056
rect 3568 14016 3574 14028
rect 4080 13929 4108 14028
rect 14550 14016 14556 14028
rect 14608 14016 14614 14068
rect 18966 14056 18972 14068
rect 18927 14028 18972 14056
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19242 14016 19248 14068
rect 19300 14056 19306 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 19300 14028 19533 14056
rect 19300 14016 19306 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 5445 13991 5503 13997
rect 5445 13988 5457 13991
rect 5224 13960 5457 13988
rect 5224 13948 5230 13960
rect 5445 13957 5457 13960
rect 5491 13957 5503 13991
rect 5445 13951 5503 13957
rect 12069 13991 12127 13997
rect 12069 13957 12081 13991
rect 12115 13988 12127 13991
rect 12986 13988 12992 14000
rect 12115 13960 12992 13988
rect 12115 13957 12127 13960
rect 12069 13951 12127 13957
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 4065 13923 4123 13929
rect 1995 13892 2544 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2130 13852 2136 13864
rect 1719 13824 2136 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13852 2375 13855
rect 2409 13855 2467 13861
rect 2409 13852 2421 13855
rect 2363 13824 2421 13852
rect 2363 13821 2375 13824
rect 2317 13815 2375 13821
rect 2409 13821 2421 13824
rect 2455 13821 2467 13855
rect 2516 13852 2544 13892
rect 4065 13889 4077 13923
rect 4111 13889 4123 13923
rect 4065 13883 4123 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 8386 13920 8392 13932
rect 8347 13892 8392 13920
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 10686 13920 10692 13932
rect 10647 13892 10692 13920
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 13078 13920 13084 13932
rect 11848 13892 13084 13920
rect 11848 13880 11854 13892
rect 13078 13880 13084 13892
rect 13136 13920 13142 13932
rect 13173 13923 13231 13929
rect 13173 13920 13185 13923
rect 13136 13892 13185 13920
rect 13136 13880 13142 13892
rect 13173 13889 13185 13892
rect 13219 13889 13231 13923
rect 14568 13920 14596 14016
rect 16485 13991 16543 13997
rect 16485 13957 16497 13991
rect 16531 13957 16543 13991
rect 16485 13951 16543 13957
rect 14568 13892 14964 13920
rect 13173 13883 13231 13889
rect 3142 13852 3148 13864
rect 2516 13824 3148 13852
rect 2409 13815 2467 13821
rect 3142 13812 3148 13824
rect 3200 13812 3206 13864
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4321 13855 4379 13861
rect 4321 13852 4333 13855
rect 4212 13824 4333 13852
rect 4212 13812 4218 13824
rect 4321 13821 4333 13824
rect 4367 13821 4379 13855
rect 4321 13815 4379 13821
rect 5626 13812 5632 13864
rect 5684 13852 5690 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 5684 13824 7297 13852
rect 5684 13812 5690 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 10962 13861 10968 13864
rect 10956 13852 10968 13861
rect 10836 13824 10968 13852
rect 10836 13812 10842 13824
rect 10956 13815 10968 13824
rect 10962 13812 10968 13815
rect 11020 13812 11026 13864
rect 13440 13855 13498 13861
rect 13440 13821 13452 13855
rect 13486 13852 13498 13855
rect 14458 13852 14464 13864
rect 13486 13824 14464 13852
rect 13486 13821 13498 13824
rect 13440 13815 13498 13821
rect 14458 13812 14464 13824
rect 14516 13812 14522 13864
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13821 14887 13855
rect 14936 13852 14964 13892
rect 15085 13855 15143 13861
rect 15085 13852 15097 13855
rect 14936 13824 15097 13852
rect 14829 13815 14887 13821
rect 15085 13821 15097 13824
rect 15131 13821 15143 13855
rect 16500 13852 16528 13951
rect 19150 13948 19156 14000
rect 19208 13988 19214 14000
rect 20441 13991 20499 13997
rect 20441 13988 20453 13991
rect 19208 13960 20453 13988
rect 19208 13948 19214 13960
rect 20441 13957 20453 13960
rect 20487 13957 20499 13991
rect 20441 13951 20499 13957
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 17000 13892 17049 13920
rect 17000 13880 17006 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 20809 13923 20867 13929
rect 20809 13920 20821 13923
rect 17037 13883 17095 13889
rect 18800 13892 20821 13920
rect 18800 13861 18828 13892
rect 20809 13889 20821 13892
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 16500 13824 18061 13852
rect 15085 13815 15143 13821
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19426 13852 19432 13864
rect 19383 13824 19432 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 2676 13787 2734 13793
rect 2676 13753 2688 13787
rect 2722 13784 2734 13787
rect 3050 13784 3056 13796
rect 2722 13756 3056 13784
rect 2722 13753 2734 13756
rect 2676 13747 2734 13753
rect 3050 13744 3056 13756
rect 3108 13744 3114 13796
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 7193 13787 7251 13793
rect 5500 13756 6960 13784
rect 5500 13744 5506 13756
rect 3786 13716 3792 13728
rect 3747 13688 3792 13716
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 6822 13716 6828 13728
rect 6783 13688 6828 13716
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 6932 13716 6960 13756
rect 7193 13753 7205 13787
rect 7239 13784 7251 13787
rect 7837 13787 7895 13793
rect 7837 13784 7849 13787
rect 7239 13756 7849 13784
rect 7239 13753 7251 13756
rect 7193 13747 7251 13753
rect 7837 13753 7849 13756
rect 7883 13753 7895 13787
rect 7837 13747 7895 13753
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 8634 13787 8692 13793
rect 8634 13784 8646 13787
rect 8536 13756 8646 13784
rect 8536 13744 8542 13756
rect 8634 13753 8646 13756
rect 8680 13753 8692 13787
rect 8634 13747 8692 13753
rect 8754 13744 8760 13796
rect 8812 13784 8818 13796
rect 14550 13784 14556 13796
rect 8812 13756 14556 13784
rect 8812 13744 8818 13756
rect 14550 13744 14556 13756
rect 14608 13744 14614 13796
rect 14844 13784 14872 13815
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13852 19947 13855
rect 20162 13852 20168 13864
rect 19935 13824 20024 13852
rect 20123 13824 20168 13852
rect 19935 13821 19947 13824
rect 19889 13815 19947 13821
rect 15562 13784 15568 13796
rect 14844 13756 15568 13784
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 16758 13744 16764 13796
rect 16816 13784 16822 13796
rect 16853 13787 16911 13793
rect 16853 13784 16865 13787
rect 16816 13756 16865 13784
rect 16816 13744 16822 13756
rect 16853 13753 16865 13756
rect 16899 13753 16911 13787
rect 17494 13784 17500 13796
rect 17455 13756 17500 13784
rect 16853 13747 16911 13753
rect 17494 13744 17500 13756
rect 17552 13744 17558 13796
rect 17586 13744 17592 13796
rect 17644 13784 17650 13796
rect 18325 13787 18383 13793
rect 18325 13784 18337 13787
rect 17644 13756 18337 13784
rect 17644 13744 17650 13756
rect 18325 13753 18337 13756
rect 18371 13753 18383 13787
rect 19996 13784 20024 13824
rect 20162 13812 20168 13824
rect 20220 13812 20226 13864
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 20625 13855 20683 13861
rect 20625 13852 20637 13855
rect 20487 13824 20637 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 20625 13821 20637 13824
rect 20671 13821 20683 13855
rect 20625 13815 20683 13821
rect 20254 13784 20260 13796
rect 19996 13756 20260 13784
rect 18325 13747 18383 13753
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 9582 13716 9588 13728
rect 6932 13688 9588 13716
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 9766 13716 9772 13728
rect 9727 13688 9772 13716
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 10410 13676 10416 13728
rect 10468 13716 10474 13728
rect 15930 13716 15936 13728
rect 10468 13688 15936 13716
rect 10468 13676 10474 13688
rect 15930 13676 15936 13688
rect 15988 13676 15994 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 16632 13688 16957 13716
rect 16632 13676 16638 13688
rect 16945 13685 16957 13688
rect 16991 13685 17003 13719
rect 16945 13679 17003 13685
rect 1104 13626 21620 13648
rect 1104 13574 7846 13626
rect 7898 13574 7910 13626
rect 7962 13574 7974 13626
rect 8026 13574 8038 13626
rect 8090 13574 14710 13626
rect 14762 13574 14774 13626
rect 14826 13574 14838 13626
rect 14890 13574 14902 13626
rect 14954 13574 21620 13626
rect 1104 13552 21620 13574
rect 1578 13512 1584 13524
rect 1539 13484 1584 13512
rect 1578 13472 1584 13484
rect 1636 13472 1642 13524
rect 1949 13515 2007 13521
rect 1949 13481 1961 13515
rect 1995 13512 2007 13515
rect 2866 13512 2872 13524
rect 1995 13484 2872 13512
rect 1995 13481 2007 13484
rect 1949 13475 2007 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 2961 13515 3019 13521
rect 2961 13481 2973 13515
rect 3007 13512 3019 13515
rect 3234 13512 3240 13524
rect 3007 13484 3240 13512
rect 3007 13481 3019 13484
rect 2961 13475 3019 13481
rect 3234 13472 3240 13484
rect 3292 13472 3298 13524
rect 3326 13472 3332 13524
rect 3384 13512 3390 13524
rect 4249 13515 4307 13521
rect 4249 13512 4261 13515
rect 3384 13484 4261 13512
rect 3384 13472 3390 13484
rect 4249 13481 4261 13484
rect 4295 13481 4307 13515
rect 5074 13512 5080 13524
rect 5035 13484 5080 13512
rect 4249 13475 4307 13481
rect 5074 13472 5080 13484
rect 5132 13472 5138 13524
rect 5169 13515 5227 13521
rect 5169 13481 5181 13515
rect 5215 13512 5227 13515
rect 5442 13512 5448 13524
rect 5215 13484 5448 13512
rect 5215 13481 5227 13484
rect 5169 13475 5227 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6086 13472 6092 13524
rect 6144 13512 6150 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 6144 13484 6285 13512
rect 6144 13472 6150 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6273 13475 6331 13481
rect 6641 13515 6699 13521
rect 6641 13481 6653 13515
rect 6687 13512 6699 13515
rect 6822 13512 6828 13524
rect 6687 13484 6828 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 6822 13472 6828 13484
rect 6880 13472 6886 13524
rect 8665 13515 8723 13521
rect 8665 13481 8677 13515
rect 8711 13512 8723 13515
rect 8754 13512 8760 13524
rect 8711 13484 8760 13512
rect 8711 13481 8723 13484
rect 8665 13475 8723 13481
rect 8680 13444 8708 13475
rect 8754 13472 8760 13484
rect 8812 13472 8818 13524
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10183 13484 14504 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 6656 13416 8708 13444
rect 9677 13447 9735 13453
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1946 13376 1952 13388
rect 1443 13348 1952 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1946 13336 1952 13348
rect 2004 13336 2010 13388
rect 2314 13376 2320 13388
rect 2275 13348 2320 13376
rect 2314 13336 2320 13348
rect 2372 13336 2378 13388
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 3878 13376 3884 13388
rect 3375 13348 3884 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4062 13376 4068 13388
rect 4023 13348 4068 13376
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 2406 13308 2412 13320
rect 2367 13280 2412 13308
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13277 2651 13311
rect 3418 13308 3424 13320
rect 3379 13280 3424 13308
rect 2593 13271 2651 13277
rect 2608 13240 2636 13271
rect 3418 13268 3424 13280
rect 3476 13268 3482 13320
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 3786 13308 3792 13320
rect 3559 13280 3792 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 3528 13240 3556 13271
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 6656 13308 6684 13416
rect 9677 13413 9689 13447
rect 9723 13444 9735 13447
rect 11517 13447 11575 13453
rect 11517 13444 11529 13447
rect 9723 13416 11529 13444
rect 9723 13413 9735 13416
rect 9677 13407 9735 13413
rect 11517 13413 11529 13416
rect 11563 13413 11575 13447
rect 11517 13407 11575 13413
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 14274 13444 14280 13456
rect 11664 13416 14280 13444
rect 11664 13404 11670 13416
rect 14274 13404 14280 13416
rect 14332 13404 14338 13456
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 7374 13376 7380 13388
rect 6779 13348 7380 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7558 13385 7564 13388
rect 7552 13376 7564 13385
rect 7519 13348 7564 13376
rect 7552 13339 7564 13348
rect 7558 13336 7564 13339
rect 7616 13336 7622 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 9088 13348 10517 13376
rect 9088 13336 9094 13348
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13376 10655 13379
rect 10962 13376 10968 13388
rect 10643 13348 10968 13376
rect 10643 13345 10655 13348
rect 10597 13339 10655 13345
rect 10962 13336 10968 13348
rect 11020 13336 11026 13388
rect 13078 13376 13084 13388
rect 13039 13348 13084 13376
rect 13078 13336 13084 13348
rect 13136 13336 13142 13388
rect 13354 13385 13360 13388
rect 13348 13339 13360 13385
rect 13412 13376 13418 13388
rect 14476 13376 14504 13484
rect 14550 13472 14556 13524
rect 14608 13512 14614 13524
rect 16942 13512 16948 13524
rect 14608 13484 16344 13512
rect 16903 13484 16948 13512
rect 14608 13472 14614 13484
rect 15832 13447 15890 13453
rect 15832 13413 15844 13447
rect 15878 13444 15890 13447
rect 16206 13444 16212 13456
rect 15878 13416 16212 13444
rect 15878 13413 15890 13416
rect 15832 13407 15890 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 16316 13444 16344 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17126 13444 17132 13456
rect 16316 13416 17132 13444
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 19518 13444 19524 13456
rect 17880 13416 19524 13444
rect 15562 13376 15568 13388
rect 13412 13348 13448 13376
rect 14476 13348 15424 13376
rect 15523 13348 15568 13376
rect 13354 13336 13360 13339
rect 13412 13336 13418 13348
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6656 13280 6837 13308
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 7285 13311 7343 13317
rect 7285 13277 7297 13311
rect 7331 13277 7343 13311
rect 10778 13308 10784 13320
rect 10739 13280 10784 13308
rect 7285 13271 7343 13277
rect 2608 13212 3556 13240
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 6178 13240 6184 13252
rect 4028 13212 6184 13240
rect 4028 13200 4034 13212
rect 6178 13200 6184 13212
rect 6236 13200 6242 13252
rect 4706 13172 4712 13184
rect 4667 13144 4712 13172
rect 4706 13132 4712 13144
rect 4764 13132 4770 13184
rect 6822 13132 6828 13184
rect 6880 13172 6886 13184
rect 7300 13172 7328 13271
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 11790 13308 11796 13320
rect 11751 13280 11796 13308
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 12802 13308 12808 13320
rect 12575 13280 12808 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 12802 13268 12808 13280
rect 12860 13268 12866 13320
rect 14182 13268 14188 13320
rect 14240 13308 14246 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 14240 13280 14749 13308
rect 14240 13268 14246 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 8386 13200 8392 13252
rect 8444 13200 8450 13252
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 10594 13240 10600 13252
rect 8536 13212 10600 13240
rect 8536 13200 8542 13212
rect 10594 13200 10600 13212
rect 10652 13240 10658 13252
rect 11808 13240 11836 13268
rect 10652 13212 11836 13240
rect 10652 13200 10658 13212
rect 8404 13172 8432 13200
rect 6880 13144 8432 13172
rect 6880 13132 6886 13144
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 11149 13175 11207 13181
rect 11149 13172 11161 13175
rect 9456 13144 11161 13172
rect 9456 13132 9462 13144
rect 11149 13141 11161 13144
rect 11195 13141 11207 13175
rect 14458 13172 14464 13184
rect 14419 13144 14464 13172
rect 11149 13135 11207 13141
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 15396 13172 15424 13348
rect 15562 13336 15568 13348
rect 15620 13376 15626 13388
rect 17770 13376 17776 13388
rect 15620 13348 17776 13376
rect 15620 13336 15626 13348
rect 17770 13336 17776 13348
rect 17828 13336 17834 13388
rect 17880 13308 17908 13416
rect 19518 13404 19524 13416
rect 19576 13404 19582 13456
rect 18040 13379 18098 13385
rect 18040 13345 18052 13379
rect 18086 13376 18098 13379
rect 18506 13376 18512 13388
rect 18086 13348 18512 13376
rect 18086 13345 18098 13348
rect 18040 13339 18098 13345
rect 18506 13336 18512 13348
rect 18564 13376 18570 13388
rect 18564 13348 18828 13376
rect 18564 13336 18570 13348
rect 17788 13280 17908 13308
rect 18800 13308 18828 13348
rect 19242 13336 19248 13388
rect 19300 13376 19306 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 19300 13348 19809 13376
rect 19300 13336 19306 13348
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 19889 13379 19947 13385
rect 19889 13345 19901 13379
rect 19935 13376 19947 13379
rect 20346 13376 20352 13388
rect 19935 13348 20352 13376
rect 19935 13345 19947 13348
rect 19889 13339 19947 13345
rect 20346 13336 20352 13348
rect 20404 13336 20410 13388
rect 19981 13311 20039 13317
rect 19981 13308 19993 13311
rect 18800 13280 19993 13308
rect 17788 13172 17816 13280
rect 19981 13277 19993 13280
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 15396 13144 17816 13172
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 19153 13175 19211 13181
rect 19153 13172 19165 13175
rect 18564 13144 19165 13172
rect 18564 13132 18570 13144
rect 19153 13141 19165 13144
rect 19199 13141 19211 13175
rect 19153 13135 19211 13141
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 19429 13175 19487 13181
rect 19429 13172 19441 13175
rect 19392 13144 19441 13172
rect 19392 13132 19398 13144
rect 19429 13141 19441 13144
rect 19475 13141 19487 13175
rect 19429 13135 19487 13141
rect 1104 13082 21620 13104
rect 1104 13030 4414 13082
rect 4466 13030 4478 13082
rect 4530 13030 4542 13082
rect 4594 13030 4606 13082
rect 4658 13030 11278 13082
rect 11330 13030 11342 13082
rect 11394 13030 11406 13082
rect 11458 13030 11470 13082
rect 11522 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 18270 13082
rect 18322 13030 18334 13082
rect 18386 13030 21620 13082
rect 1104 13008 21620 13030
rect 2406 12928 2412 12980
rect 2464 12968 2470 12980
rect 2501 12971 2559 12977
rect 2501 12968 2513 12971
rect 2464 12940 2513 12968
rect 2464 12928 2470 12940
rect 2501 12937 2513 12940
rect 2547 12937 2559 12971
rect 2501 12931 2559 12937
rect 3418 12928 3424 12980
rect 3476 12968 3482 12980
rect 3789 12971 3847 12977
rect 3789 12968 3801 12971
rect 3476 12940 3801 12968
rect 3476 12928 3482 12940
rect 3789 12937 3801 12940
rect 3835 12937 3847 12971
rect 3789 12931 3847 12937
rect 3878 12928 3884 12980
rect 3936 12968 3942 12980
rect 6825 12971 6883 12977
rect 6825 12968 6837 12971
rect 3936 12940 6837 12968
rect 3936 12928 3942 12940
rect 6825 12937 6837 12940
rect 6871 12937 6883 12971
rect 9030 12968 9036 12980
rect 8991 12940 9036 12968
rect 6825 12931 6883 12937
rect 9030 12928 9036 12940
rect 9088 12928 9094 12980
rect 9766 12928 9772 12980
rect 9824 12968 9830 12980
rect 9824 12940 10824 12968
rect 9824 12928 9830 12940
rect 3510 12860 3516 12912
rect 3568 12900 3574 12912
rect 6178 12900 6184 12912
rect 3568 12872 4844 12900
rect 6091 12872 6184 12900
rect 3568 12860 3574 12872
rect 1946 12832 1952 12844
rect 1907 12804 1952 12832
rect 1946 12792 1952 12804
rect 2004 12792 2010 12844
rect 2958 12832 2964 12844
rect 2919 12804 2964 12832
rect 2958 12792 2964 12804
rect 3016 12792 3022 12844
rect 3050 12792 3056 12844
rect 3108 12832 3114 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 3108 12804 3157 12832
rect 3108 12792 3114 12804
rect 3145 12801 3157 12804
rect 3191 12832 3203 12835
rect 3970 12832 3976 12844
rect 3191 12804 3976 12832
rect 3191 12801 3203 12804
rect 3145 12795 3203 12801
rect 3970 12792 3976 12804
rect 4028 12832 4034 12844
rect 4816 12841 4844 12872
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 6641 12903 6699 12909
rect 6641 12869 6653 12903
rect 6687 12900 6699 12903
rect 7837 12903 7895 12909
rect 6687 12872 7512 12900
rect 6687 12869 6699 12872
rect 6641 12863 6699 12869
rect 4341 12835 4399 12841
rect 4341 12832 4353 12835
rect 4028 12804 4353 12832
rect 4028 12792 4034 12804
rect 4341 12801 4353 12804
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 6196 12832 6224 12860
rect 7377 12835 7435 12841
rect 7377 12832 7389 12835
rect 6196 12804 7389 12832
rect 4801 12795 4859 12801
rect 7377 12801 7389 12804
rect 7423 12801 7435 12835
rect 7484 12832 7512 12872
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 10502 12900 10508 12912
rect 7883 12872 10508 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 8297 12835 8355 12841
rect 8297 12832 8309 12835
rect 7484 12804 8309 12832
rect 7377 12795 7435 12801
rect 8297 12801 8309 12804
rect 8343 12801 8355 12835
rect 8478 12832 8484 12844
rect 8439 12804 8484 12832
rect 8297 12795 8355 12801
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 9490 12832 9496 12844
rect 9451 12804 9496 12832
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9585 12835 9643 12841
rect 9585 12801 9597 12835
rect 9631 12832 9643 12835
rect 9766 12832 9772 12844
rect 9631 12804 9772 12832
rect 9631 12801 9643 12804
rect 9585 12795 9643 12801
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 10594 12832 10600 12844
rect 10555 12804 10600 12832
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 10796 12832 10824 12940
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 11020 12940 11069 12968
rect 11020 12928 11026 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 11057 12931 11115 12937
rect 13817 12971 13875 12977
rect 13817 12937 13829 12971
rect 13863 12968 13875 12971
rect 14090 12968 14096 12980
rect 13863 12940 14096 12968
rect 13863 12937 13875 12940
rect 13817 12931 13875 12937
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 16574 12968 16580 12980
rect 16535 12940 16580 12968
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 20898 12968 20904 12980
rect 20859 12940 20904 12968
rect 20898 12928 20904 12940
rect 20956 12928 20962 12980
rect 15565 12903 15623 12909
rect 15565 12869 15577 12903
rect 15611 12900 15623 12903
rect 17310 12900 17316 12912
rect 15611 12872 17316 12900
rect 15611 12869 15623 12872
rect 15565 12863 15623 12869
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 10796 12804 11621 12832
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 12986 12832 12992 12844
rect 12947 12804 12992 12832
rect 11609 12795 11667 12801
rect 12986 12792 12992 12804
rect 13044 12792 13050 12844
rect 14274 12832 14280 12844
rect 14235 12804 14280 12832
rect 14274 12792 14280 12804
rect 14332 12792 14338 12844
rect 14458 12832 14464 12844
rect 14419 12804 14464 12832
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 15838 12792 15844 12844
rect 15896 12832 15902 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15896 12804 16129 12832
rect 15896 12792 15902 12804
rect 16117 12801 16129 12804
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 17129 12835 17187 12841
rect 17129 12832 17141 12835
rect 16264 12804 17141 12832
rect 16264 12792 16270 12804
rect 17129 12801 17141 12804
rect 17175 12801 17187 12835
rect 17129 12795 17187 12801
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17828 12804 18245 12832
rect 17828 12792 17834 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 19610 12792 19616 12844
rect 19668 12832 19674 12844
rect 20165 12835 20223 12841
rect 20165 12832 20177 12835
rect 19668 12804 20177 12832
rect 19668 12792 19674 12804
rect 20165 12801 20177 12804
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 1762 12764 1768 12776
rect 1723 12736 1768 12764
rect 1762 12724 1768 12736
rect 1820 12724 1826 12776
rect 2976 12764 3004 12792
rect 3878 12764 3884 12776
rect 2976 12736 3884 12764
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 4249 12767 4307 12773
rect 4249 12733 4261 12767
rect 4295 12764 4307 12767
rect 4706 12764 4712 12776
rect 4295 12736 4712 12764
rect 4295 12733 4307 12736
rect 4249 12727 4307 12733
rect 4706 12724 4712 12736
rect 4764 12724 4770 12776
rect 12434 12764 12440 12776
rect 4908 12736 12440 12764
rect 3510 12656 3516 12708
rect 3568 12696 3574 12708
rect 3694 12696 3700 12708
rect 3568 12668 3700 12696
rect 3568 12656 3574 12668
rect 3694 12656 3700 12668
rect 3752 12656 3758 12708
rect 3970 12656 3976 12708
rect 4028 12696 4034 12708
rect 4908 12696 4936 12736
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 14182 12764 14188 12776
rect 14143 12736 14188 12764
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 15930 12724 15936 12776
rect 15988 12764 15994 12776
rect 18506 12773 18512 12776
rect 18500 12764 18512 12773
rect 15988 12736 16160 12764
rect 18467 12736 18512 12764
rect 15988 12724 15994 12736
rect 4028 12668 4936 12696
rect 5068 12699 5126 12705
rect 4028 12656 4034 12668
rect 5068 12665 5080 12699
rect 5114 12696 5126 12699
rect 5442 12696 5448 12708
rect 5114 12668 5448 12696
rect 5114 12665 5126 12668
rect 5068 12659 5126 12665
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 5552 12668 6653 12696
rect 2498 12588 2504 12640
rect 2556 12628 2562 12640
rect 2869 12631 2927 12637
rect 2869 12628 2881 12631
rect 2556 12600 2881 12628
rect 2556 12588 2562 12600
rect 2869 12597 2881 12600
rect 2915 12597 2927 12631
rect 2869 12591 2927 12597
rect 4157 12631 4215 12637
rect 4157 12597 4169 12631
rect 4203 12628 4215 12631
rect 4706 12628 4712 12640
rect 4203 12600 4712 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4706 12588 4712 12600
rect 4764 12628 4770 12640
rect 5552 12628 5580 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 7285 12699 7343 12705
rect 7285 12665 7297 12699
rect 7331 12696 7343 12699
rect 7650 12696 7656 12708
rect 7331 12668 7656 12696
rect 7331 12665 7343 12668
rect 7285 12659 7343 12665
rect 7650 12656 7656 12668
rect 7708 12696 7714 12708
rect 8205 12699 8263 12705
rect 8205 12696 8217 12699
rect 7708 12668 8217 12696
rect 7708 12656 7714 12668
rect 8205 12665 8217 12668
rect 8251 12665 8263 12699
rect 9398 12696 9404 12708
rect 9359 12668 9404 12696
rect 8205 12659 8263 12665
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 10318 12696 10324 12708
rect 9508 12668 10324 12696
rect 4764 12600 5580 12628
rect 7193 12631 7251 12637
rect 4764 12588 4770 12600
rect 7193 12597 7205 12631
rect 7239 12628 7251 12631
rect 9508 12628 9536 12668
rect 10318 12656 10324 12668
rect 10376 12696 10382 12708
rect 10505 12699 10563 12705
rect 10505 12696 10517 12699
rect 10376 12668 10517 12696
rect 10376 12656 10382 12668
rect 10505 12665 10517 12668
rect 10551 12665 10563 12699
rect 10505 12659 10563 12665
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 11425 12699 11483 12705
rect 11425 12696 11437 12699
rect 10652 12668 11437 12696
rect 10652 12656 10658 12668
rect 11425 12665 11437 12668
rect 11471 12665 11483 12699
rect 11425 12659 11483 12665
rect 11517 12699 11575 12705
rect 11517 12665 11529 12699
rect 11563 12696 11575 12699
rect 15102 12696 15108 12708
rect 11563 12668 15108 12696
rect 11563 12665 11575 12668
rect 11517 12659 11575 12665
rect 15102 12656 15108 12668
rect 15160 12656 15166 12708
rect 15194 12656 15200 12708
rect 15252 12696 15258 12708
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 15252 12668 16037 12696
rect 15252 12656 15258 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 16132 12696 16160 12736
rect 18500 12727 18512 12736
rect 18506 12724 18512 12727
rect 18564 12724 18570 12776
rect 18782 12724 18788 12776
rect 18840 12764 18846 12776
rect 19981 12767 20039 12773
rect 19981 12764 19993 12767
rect 18840 12736 19993 12764
rect 18840 12724 18846 12736
rect 19981 12733 19993 12736
rect 20027 12733 20039 12767
rect 19981 12727 20039 12733
rect 20622 12724 20628 12776
rect 20680 12764 20686 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20680 12736 20729 12764
rect 20680 12724 20686 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 19886 12696 19892 12708
rect 16132 12668 19892 12696
rect 16025 12659 16083 12665
rect 19886 12656 19892 12668
rect 19944 12656 19950 12708
rect 7239 12600 9536 12628
rect 7239 12597 7251 12600
rect 7193 12591 7251 12597
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 10045 12631 10103 12637
rect 10045 12628 10057 12631
rect 9640 12600 10057 12628
rect 9640 12588 9646 12600
rect 10045 12597 10057 12600
rect 10091 12597 10103 12631
rect 10410 12628 10416 12640
rect 10371 12600 10416 12628
rect 10045 12591 10103 12597
rect 10410 12588 10416 12600
rect 10468 12588 10474 12640
rect 11974 12588 11980 12640
rect 12032 12628 12038 12640
rect 12437 12631 12495 12637
rect 12437 12628 12449 12631
rect 12032 12600 12449 12628
rect 12032 12588 12038 12600
rect 12437 12597 12449 12600
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 12710 12588 12716 12640
rect 12768 12628 12774 12640
rect 12897 12631 12955 12637
rect 12897 12628 12909 12631
rect 12768 12600 12909 12628
rect 12768 12588 12774 12600
rect 12897 12597 12909 12600
rect 12943 12597 12955 12631
rect 15930 12628 15936 12640
rect 15891 12600 15936 12628
rect 12897 12591 12955 12597
rect 15930 12588 15936 12600
rect 15988 12588 15994 12640
rect 16666 12588 16672 12640
rect 16724 12628 16730 12640
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 16724 12600 16957 12628
rect 16724 12588 16730 12600
rect 16945 12597 16957 12600
rect 16991 12597 17003 12631
rect 16945 12591 17003 12597
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 19610 12628 19616 12640
rect 17092 12600 17137 12628
rect 19571 12600 19616 12628
rect 17092 12588 17098 12600
rect 19610 12588 19616 12600
rect 19668 12588 19674 12640
rect 1104 12538 21620 12560
rect 1104 12486 7846 12538
rect 7898 12486 7910 12538
rect 7962 12486 7974 12538
rect 8026 12486 8038 12538
rect 8090 12486 14710 12538
rect 14762 12486 14774 12538
rect 14826 12486 14838 12538
rect 14890 12486 14902 12538
rect 14954 12486 21620 12538
rect 1104 12464 21620 12486
rect 2314 12384 2320 12436
rect 2372 12424 2378 12436
rect 2409 12427 2467 12433
rect 2409 12424 2421 12427
rect 2372 12396 2421 12424
rect 2372 12384 2378 12396
rect 2409 12393 2421 12396
rect 2455 12393 2467 12427
rect 3602 12424 3608 12436
rect 3563 12396 3608 12424
rect 2409 12387 2467 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 5442 12424 5448 12436
rect 5403 12396 5448 12424
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 7374 12384 7380 12436
rect 7432 12424 7438 12436
rect 7929 12427 7987 12433
rect 7929 12424 7941 12427
rect 7432 12396 7941 12424
rect 7432 12384 7438 12396
rect 7929 12393 7941 12396
rect 7975 12393 7987 12427
rect 7929 12387 7987 12393
rect 8036 12396 12388 12424
rect 1857 12359 1915 12365
rect 1857 12325 1869 12359
rect 1903 12356 1915 12359
rect 2958 12356 2964 12368
rect 1903 12328 2964 12356
rect 1903 12325 1915 12328
rect 1857 12319 1915 12325
rect 2958 12316 2964 12328
rect 3016 12316 3022 12368
rect 4154 12316 4160 12368
rect 4212 12356 4218 12368
rect 5074 12356 5080 12368
rect 4212 12328 5080 12356
rect 4212 12316 4218 12328
rect 5074 12316 5080 12328
rect 5132 12316 5138 12368
rect 6540 12359 6598 12365
rect 6540 12325 6552 12359
rect 6586 12356 6598 12359
rect 7006 12356 7012 12368
rect 6586 12328 7012 12356
rect 6586 12325 6598 12328
rect 6540 12319 6598 12325
rect 7006 12316 7012 12328
rect 7064 12316 7070 12368
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 7834 12356 7840 12368
rect 7524 12328 7840 12356
rect 7524 12316 7530 12328
rect 7834 12316 7840 12328
rect 7892 12316 7898 12368
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12257 1823 12291
rect 1765 12251 1823 12257
rect 1394 12084 1400 12096
rect 1355 12056 1400 12084
rect 1394 12044 1400 12056
rect 1452 12044 1458 12096
rect 1780 12084 1808 12251
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 3142 12248 3148 12300
rect 3200 12288 3206 12300
rect 3421 12291 3479 12297
rect 3421 12288 3433 12291
rect 3200 12260 3433 12288
rect 3200 12248 3206 12260
rect 3421 12257 3433 12260
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 3510 12248 3516 12300
rect 3568 12288 3574 12300
rect 4321 12291 4379 12297
rect 4321 12288 4333 12291
rect 3568 12260 4333 12288
rect 3568 12248 3574 12260
rect 4321 12257 4333 12260
rect 4367 12257 4379 12291
rect 4321 12251 4379 12257
rect 5258 12248 5264 12300
rect 5316 12288 5322 12300
rect 8036 12288 8064 12396
rect 8202 12316 8208 12368
rect 8260 12356 8266 12368
rect 12360 12356 12388 12396
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12897 12427 12955 12433
rect 12897 12424 12909 12427
rect 12492 12396 12909 12424
rect 12492 12384 12498 12396
rect 12897 12393 12909 12396
rect 12943 12393 12955 12427
rect 12897 12387 12955 12393
rect 14093 12427 14151 12433
rect 14093 12393 14105 12427
rect 14139 12424 14151 12427
rect 15194 12424 15200 12436
rect 14139 12396 15200 12424
rect 14139 12393 14151 12396
rect 14093 12387 14151 12393
rect 15194 12384 15200 12396
rect 15252 12384 15258 12436
rect 15930 12424 15936 12436
rect 15891 12396 15936 12424
rect 15930 12384 15936 12396
rect 15988 12384 15994 12436
rect 16022 12384 16028 12436
rect 16080 12424 16086 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16080 12396 16405 12424
rect 16080 12384 16086 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 17034 12424 17040 12436
rect 16393 12387 16451 12393
rect 16500 12396 17040 12424
rect 16500 12356 16528 12396
rect 17034 12384 17040 12396
rect 17092 12384 17098 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 18325 12427 18383 12433
rect 18325 12393 18337 12427
rect 18371 12424 18383 12427
rect 19153 12427 19211 12433
rect 19153 12424 19165 12427
rect 18371 12396 19165 12424
rect 18371 12393 18383 12396
rect 18325 12387 18383 12393
rect 19153 12393 19165 12396
rect 19199 12393 19211 12427
rect 20346 12424 20352 12436
rect 19153 12387 19211 12393
rect 19444 12396 20352 12424
rect 8260 12328 10272 12356
rect 12360 12328 16528 12356
rect 8260 12316 8266 12328
rect 5316 12260 8064 12288
rect 8297 12291 8355 12297
rect 5316 12248 5322 12260
rect 8297 12257 8309 12291
rect 8343 12288 8355 12291
rect 8570 12288 8576 12300
rect 8343 12260 8576 12288
rect 8343 12257 8355 12260
rect 8297 12251 8355 12257
rect 8570 12248 8576 12260
rect 8628 12248 8634 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10244 12232 10272 12328
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 19444 12356 19472 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 16632 12328 19472 12356
rect 19521 12359 19579 12365
rect 16632 12316 16638 12328
rect 19521 12325 19533 12359
rect 19567 12356 19579 12359
rect 20901 12359 20959 12365
rect 20901 12356 20913 12359
rect 19567 12328 20913 12356
rect 19567 12325 19579 12328
rect 19521 12319 19579 12325
rect 20901 12325 20913 12328
rect 20947 12325 20959 12359
rect 20901 12319 20959 12325
rect 10686 12248 10692 12300
rect 10744 12288 10750 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10744 12260 10793 12288
rect 10744 12248 10750 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 11048 12291 11106 12297
rect 11048 12288 11060 12291
rect 10781 12251 10839 12257
rect 10888 12260 11060 12288
rect 2038 12220 2044 12232
rect 1999 12192 2044 12220
rect 2038 12180 2044 12192
rect 2096 12180 2102 12232
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 3050 12220 3056 12232
rect 3011 12192 3056 12220
rect 2869 12183 2927 12189
rect 2884 12152 2912 12183
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 3694 12180 3700 12232
rect 3752 12220 3758 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3752 12192 4077 12220
rect 3752 12180 3758 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5960 12192 6285 12220
rect 5960 12180 5966 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7524 12192 8401 12220
rect 7524 12180 7530 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 10226 12220 10232 12232
rect 10187 12192 10232 12220
rect 8481 12183 8539 12189
rect 3142 12152 3148 12164
rect 2884 12124 3148 12152
rect 3142 12112 3148 12124
rect 3200 12112 3206 12164
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 7653 12155 7711 12161
rect 7653 12152 7665 12155
rect 7616 12124 7665 12152
rect 7616 12112 7622 12124
rect 7653 12121 7665 12124
rect 7699 12152 7711 12155
rect 8496 12152 8524 12183
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12220 10471 12223
rect 10888 12220 10916 12260
rect 11048 12257 11060 12260
rect 11094 12288 11106 12291
rect 11790 12288 11796 12300
rect 11094 12260 11796 12288
rect 11094 12257 11106 12260
rect 11048 12251 11106 12257
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 12805 12291 12863 12297
rect 12805 12257 12817 12291
rect 12851 12288 12863 12291
rect 13449 12291 13507 12297
rect 13449 12288 13461 12291
rect 12851 12260 13461 12288
rect 12851 12257 12863 12260
rect 12805 12251 12863 12257
rect 13449 12257 13461 12260
rect 13495 12257 13507 12291
rect 14458 12288 14464 12300
rect 14419 12260 14464 12288
rect 13449 12251 13507 12257
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 16301 12291 16359 12297
rect 16301 12288 16313 12291
rect 16172 12260 16313 12288
rect 16172 12248 16178 12260
rect 16301 12257 16313 12260
rect 16347 12257 16359 12291
rect 16301 12251 16359 12257
rect 17770 12248 17776 12300
rect 17828 12288 17834 12300
rect 18969 12291 19027 12297
rect 18969 12288 18981 12291
rect 17828 12260 18981 12288
rect 17828 12248 17834 12260
rect 18969 12257 18981 12260
rect 19015 12288 19027 12291
rect 19613 12291 19671 12297
rect 19613 12288 19625 12291
rect 19015 12260 19625 12288
rect 19015 12257 19027 12260
rect 18969 12251 19027 12257
rect 19613 12257 19625 12260
rect 19659 12288 19671 12291
rect 19659 12260 20116 12288
rect 19659 12257 19671 12260
rect 19613 12251 19671 12257
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 10459 12192 10916 12220
rect 12176 12192 13001 12220
rect 10459 12189 10471 12192
rect 10413 12183 10471 12189
rect 10502 12152 10508 12164
rect 7699 12124 8524 12152
rect 8588 12124 10508 12152
rect 7699 12121 7711 12124
rect 7653 12115 7711 12121
rect 3050 12084 3056 12096
rect 1780 12056 3056 12084
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3878 12044 3884 12096
rect 3936 12084 3942 12096
rect 8588 12084 8616 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12176 12161 12204 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 13170 12180 13176 12232
rect 13228 12220 13234 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 13228 12192 14565 12220
rect 13228 12180 13234 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14734 12220 14740 12232
rect 14647 12192 14740 12220
rect 14553 12183 14611 12189
rect 14734 12180 14740 12192
rect 14792 12220 14798 12232
rect 16482 12220 16488 12232
rect 14792 12192 16488 12220
rect 14792 12180 14798 12192
rect 16482 12180 16488 12192
rect 16540 12180 16546 12232
rect 17402 12220 17408 12232
rect 17363 12192 17408 12220
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17494 12180 17500 12232
rect 17552 12220 17558 12232
rect 17552 12192 17597 12220
rect 17552 12180 17558 12192
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18012 12192 18429 12220
rect 18012 12180 18018 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12220 18659 12223
rect 19518 12220 19524 12232
rect 18647 12192 19524 12220
rect 18647 12189 18659 12192
rect 18601 12183 18659 12189
rect 19518 12180 19524 12192
rect 19576 12180 19582 12232
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12189 19763 12223
rect 20088 12220 20116 12260
rect 20162 12248 20168 12300
rect 20220 12288 20226 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 20220 12260 20269 12288
rect 20220 12248 20226 12260
rect 20257 12257 20269 12260
rect 20303 12257 20315 12291
rect 20257 12251 20315 12257
rect 20622 12220 20628 12232
rect 20088 12192 20628 12220
rect 19705 12183 19763 12189
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 11940 12124 12173 12152
rect 11940 12112 11946 12124
rect 12161 12121 12173 12124
rect 12207 12121 12219 12155
rect 12161 12115 12219 12121
rect 16945 12155 17003 12161
rect 16945 12121 16957 12155
rect 16991 12152 17003 12155
rect 18782 12152 18788 12164
rect 16991 12124 18788 12152
rect 16991 12121 17003 12124
rect 16945 12115 17003 12121
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 18874 12112 18880 12164
rect 18932 12152 18938 12164
rect 19720 12152 19748 12183
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20438 12152 20444 12164
rect 18932 12124 19748 12152
rect 20399 12124 20444 12152
rect 18932 12112 18938 12124
rect 20438 12112 20444 12124
rect 20496 12112 20502 12164
rect 3936 12056 8616 12084
rect 9769 12087 9827 12093
rect 3936 12044 3942 12056
rect 9769 12053 9781 12087
rect 9815 12084 9827 12087
rect 11698 12084 11704 12096
rect 9815 12056 11704 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 12437 12087 12495 12093
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12802 12084 12808 12096
rect 12483 12056 12808 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17957 12087 18015 12093
rect 17957 12084 17969 12087
rect 17276 12056 17969 12084
rect 17276 12044 17282 12056
rect 17957 12053 17969 12056
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 18892 12084 18920 12112
rect 18564 12056 18920 12084
rect 18564 12044 18570 12056
rect 1104 11994 21620 12016
rect 1104 11942 4414 11994
rect 4466 11942 4478 11994
rect 4530 11942 4542 11994
rect 4594 11942 4606 11994
rect 4658 11942 11278 11994
rect 11330 11942 11342 11994
rect 11394 11942 11406 11994
rect 11458 11942 11470 11994
rect 11522 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 18270 11994
rect 18322 11942 18334 11994
rect 18386 11942 21620 11994
rect 1104 11920 21620 11942
rect 4062 11840 4068 11892
rect 4120 11880 4126 11892
rect 11790 11880 11796 11892
rect 4120 11852 11376 11880
rect 11751 11852 11796 11880
rect 4120 11840 4126 11852
rect 2777 11815 2835 11821
rect 2777 11781 2789 11815
rect 2823 11812 2835 11815
rect 4985 11815 5043 11821
rect 2823 11784 4292 11812
rect 2823 11781 2835 11784
rect 2777 11775 2835 11781
rect 2038 11704 2044 11756
rect 2096 11744 2102 11756
rect 4264 11753 4292 11784
rect 4985 11781 4997 11815
rect 5031 11812 5043 11815
rect 6178 11812 6184 11824
rect 5031 11784 6184 11812
rect 5031 11781 5043 11784
rect 4985 11775 5043 11781
rect 6178 11772 6184 11784
rect 6236 11772 6242 11824
rect 7466 11812 7472 11824
rect 7427 11784 7472 11812
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 7668 11784 8156 11812
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 2096 11716 2513 11744
rect 2096 11704 2102 11716
rect 2501 11713 2513 11716
rect 2547 11744 2559 11747
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2547 11716 2697 11744
rect 2547 11713 2559 11716
rect 2501 11707 2559 11713
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5224 11716 5549 11744
rect 5224 11704 5230 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 7098 11744 7104 11756
rect 5537 11707 5595 11713
rect 6104 11716 7104 11744
rect 2869 11679 2927 11685
rect 2869 11645 2881 11679
rect 2915 11676 2927 11679
rect 3145 11679 3203 11685
rect 2915 11648 3096 11676
rect 2915 11645 2927 11648
rect 2869 11639 2927 11645
rect 3068 11608 3096 11648
rect 3145 11645 3157 11679
rect 3191 11676 3203 11679
rect 3970 11676 3976 11688
rect 3191 11648 3976 11676
rect 3191 11645 3203 11648
rect 3145 11639 3203 11645
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 5258 11636 5264 11688
rect 5316 11676 5322 11688
rect 5353 11679 5411 11685
rect 5353 11676 5365 11679
rect 5316 11648 5365 11676
rect 5316 11636 5322 11648
rect 5353 11645 5365 11648
rect 5399 11645 5411 11679
rect 5353 11639 5411 11645
rect 5442 11636 5448 11688
rect 5500 11676 5506 11688
rect 6104 11676 6132 11716
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 5500 11648 6132 11676
rect 6181 11679 6239 11685
rect 5500 11636 5506 11648
rect 6181 11645 6193 11679
rect 6227 11676 6239 11679
rect 7668 11676 7696 11784
rect 8018 11744 8024 11756
rect 7979 11716 8024 11744
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 7837 11679 7895 11685
rect 7837 11676 7849 11679
rect 6227 11648 7696 11676
rect 7760 11648 7849 11676
rect 6227 11645 6239 11648
rect 6181 11639 6239 11645
rect 3326 11608 3332 11620
rect 3068 11580 3332 11608
rect 3326 11568 3332 11580
rect 3384 11568 3390 11620
rect 6914 11608 6920 11620
rect 3620 11580 6920 11608
rect 1854 11540 1860 11552
rect 1815 11512 1860 11540
rect 1854 11500 1860 11512
rect 1912 11500 1918 11552
rect 2222 11540 2228 11552
rect 2183 11512 2228 11540
rect 2222 11500 2228 11512
rect 2280 11500 2286 11552
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 3620 11549 3648 11580
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7006 11568 7012 11620
rect 7064 11608 7070 11620
rect 7760 11608 7788 11648
rect 7837 11645 7849 11648
rect 7883 11645 7895 11679
rect 8128 11676 8156 11784
rect 8386 11772 8392 11824
rect 8444 11812 8450 11824
rect 8481 11815 8539 11821
rect 8481 11812 8493 11815
rect 8444 11784 8493 11812
rect 8444 11772 8450 11784
rect 8481 11781 8493 11784
rect 8527 11812 8539 11815
rect 11348 11812 11376 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 13078 11840 13084 11892
rect 13136 11880 13142 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13136 11852 13461 11880
rect 13136 11840 13142 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 15010 11840 15016 11892
rect 15068 11880 15074 11892
rect 16850 11880 16856 11892
rect 15068 11852 16856 11880
rect 15068 11840 15074 11852
rect 16850 11840 16856 11852
rect 16908 11840 16914 11892
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 17494 11880 17500 11892
rect 16991 11852 17500 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17954 11840 17960 11892
rect 18012 11880 18018 11892
rect 18049 11883 18107 11889
rect 18049 11880 18061 11883
rect 18012 11852 18061 11880
rect 18012 11840 18018 11852
rect 18049 11849 18061 11852
rect 18095 11849 18107 11883
rect 19334 11880 19340 11892
rect 18049 11843 18107 11849
rect 18524 11852 19340 11880
rect 12710 11812 12716 11824
rect 8527 11784 8800 11812
rect 11348 11784 12716 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 8772 11753 8800 11784
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 15289 11815 15347 11821
rect 15289 11781 15301 11815
rect 15335 11812 15347 11815
rect 15381 11815 15439 11821
rect 15381 11812 15393 11815
rect 15335 11784 15393 11812
rect 15335 11781 15347 11784
rect 15289 11775 15347 11781
rect 15381 11781 15393 11784
rect 15427 11781 15439 11815
rect 15381 11775 15439 11781
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 8478 11676 8484 11688
rect 8128 11648 8484 11676
rect 7837 11639 7895 11645
rect 8478 11636 8484 11648
rect 8536 11676 8542 11688
rect 8665 11679 8723 11685
rect 8665 11676 8677 11679
rect 8536 11648 8677 11676
rect 8536 11636 8542 11648
rect 8665 11645 8677 11648
rect 8711 11645 8723 11679
rect 8772 11676 8800 11707
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 12986 11744 12992 11756
rect 10100 11716 10548 11744
rect 12947 11716 12992 11744
rect 10100 11704 10106 11716
rect 9490 11676 9496 11688
rect 8772 11648 9496 11676
rect 8665 11639 8723 11645
rect 9490 11636 9496 11648
rect 9548 11676 9554 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 9548 11648 10425 11676
rect 9548 11636 9554 11648
rect 10413 11645 10425 11648
rect 10459 11645 10471 11679
rect 10520 11676 10548 11716
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 15562 11744 15568 11756
rect 15523 11716 15568 11744
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 18524 11753 18552 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20901 11883 20959 11889
rect 20901 11849 20913 11883
rect 20947 11880 20959 11883
rect 20990 11880 20996 11892
rect 20947 11852 20996 11880
rect 20947 11849 20959 11852
rect 20901 11843 20959 11849
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 18509 11747 18567 11753
rect 16868 11716 18000 11744
rect 11606 11676 11612 11688
rect 10520 11648 11612 11676
rect 10413 11639 10471 11645
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 13633 11679 13691 11685
rect 13633 11645 13645 11679
rect 13679 11676 13691 11679
rect 13814 11676 13820 11688
rect 13679 11648 13820 11676
rect 13679 11645 13691 11648
rect 13633 11639 13691 11645
rect 13814 11636 13820 11648
rect 13872 11636 13878 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14176 11679 14234 11685
rect 14176 11645 14188 11679
rect 14222 11676 14234 11679
rect 14734 11676 14740 11688
rect 14222 11648 14740 11676
rect 14222 11645 14234 11648
rect 14176 11639 14234 11645
rect 7064 11580 7788 11608
rect 9024 11611 9082 11617
rect 7064 11568 7070 11580
rect 9024 11577 9036 11611
rect 9070 11608 9082 11611
rect 9582 11608 9588 11620
rect 9070 11580 9588 11608
rect 9070 11577 9082 11580
rect 9024 11571 9082 11577
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 10658 11611 10716 11617
rect 10658 11608 10670 11611
rect 10244 11580 10670 11608
rect 10244 11552 10272 11580
rect 10658 11577 10670 11580
rect 10704 11577 10716 11611
rect 10658 11571 10716 11577
rect 12342 11568 12348 11620
rect 12400 11608 12406 11620
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12400 11580 12909 11608
rect 12400 11568 12406 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 13924 11608 13952 11639
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15580 11676 15608 11704
rect 16868 11688 16896 11716
rect 16850 11676 16856 11688
rect 14844 11648 16856 11676
rect 14844 11608 14872 11648
rect 16850 11636 16856 11648
rect 16908 11636 16914 11688
rect 17218 11676 17224 11688
rect 17179 11648 17224 11676
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 17972 11676 18000 11716
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18509 11707 18567 11713
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11744 18751 11747
rect 18874 11744 18880 11756
rect 18739 11716 18880 11744
rect 18739 11713 18751 11716
rect 18693 11707 18751 11713
rect 18874 11704 18880 11716
rect 18932 11704 18938 11756
rect 19061 11679 19119 11685
rect 19061 11676 19073 11679
rect 17972 11648 19073 11676
rect 19061 11645 19073 11648
rect 19107 11645 19119 11679
rect 19061 11639 19119 11645
rect 19328 11679 19386 11685
rect 19328 11645 19340 11679
rect 19374 11676 19386 11679
rect 19610 11676 19616 11688
rect 19374 11648 19616 11676
rect 19374 11645 19386 11648
rect 19328 11639 19386 11645
rect 19610 11636 19616 11648
rect 19668 11636 19674 11688
rect 20070 11636 20076 11688
rect 20128 11676 20134 11688
rect 20438 11676 20444 11688
rect 20128 11648 20444 11676
rect 20128 11636 20134 11648
rect 20438 11636 20444 11648
rect 20496 11636 20502 11688
rect 20714 11676 20720 11688
rect 20675 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11636 20778 11688
rect 15838 11617 15844 11620
rect 13924 11580 14872 11608
rect 15381 11611 15439 11617
rect 12897 11571 12955 11577
rect 15381 11577 15393 11611
rect 15427 11608 15439 11611
rect 15832 11608 15844 11617
rect 15427 11580 15844 11608
rect 15427 11577 15439 11580
rect 15381 11571 15439 11577
rect 15832 11571 15844 11580
rect 15838 11568 15844 11571
rect 15896 11568 15902 11620
rect 16574 11568 16580 11620
rect 16632 11608 16638 11620
rect 17497 11611 17555 11617
rect 17497 11608 17509 11611
rect 16632 11580 17509 11608
rect 16632 11568 16638 11580
rect 17497 11577 17509 11580
rect 17543 11577 17555 11611
rect 17497 11571 17555 11577
rect 3605 11543 3663 11549
rect 2372 11512 2417 11540
rect 2372 11500 2378 11512
rect 3605 11509 3617 11543
rect 3651 11509 3663 11543
rect 3970 11540 3976 11552
rect 3931 11512 3976 11540
rect 3605 11503 3663 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4065 11543 4123 11549
rect 4065 11509 4077 11543
rect 4111 11540 4123 11543
rect 4154 11540 4160 11552
rect 4111 11512 4160 11540
rect 4111 11509 4123 11512
rect 4065 11503 4123 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 5997 11543 6055 11549
rect 5997 11540 6009 11543
rect 5960 11512 6009 11540
rect 5960 11500 5966 11512
rect 5997 11509 6009 11512
rect 6043 11509 6055 11543
rect 5997 11503 6055 11509
rect 6454 11500 6460 11552
rect 6512 11540 6518 11552
rect 7742 11540 7748 11552
rect 6512 11512 7748 11540
rect 6512 11500 6518 11512
rect 7742 11500 7748 11512
rect 7800 11500 7806 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8202 11540 8208 11552
rect 7975 11512 8208 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 10042 11540 10048 11552
rect 8444 11512 10048 11540
rect 8444 11500 8450 11512
rect 10042 11500 10048 11512
rect 10100 11500 10106 11552
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10226 11540 10232 11552
rect 10183 11512 10232 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 12437 11543 12495 11549
rect 12437 11509 12449 11543
rect 12483 11540 12495 11543
rect 13354 11540 13360 11552
rect 12483 11512 13360 11540
rect 12483 11509 12495 11512
rect 12437 11503 12495 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 17586 11540 17592 11552
rect 16264 11512 17592 11540
rect 16264 11500 16270 11512
rect 17586 11500 17592 11512
rect 17644 11500 17650 11552
rect 18417 11543 18475 11549
rect 18417 11509 18429 11543
rect 18463 11540 18475 11543
rect 18506 11540 18512 11552
rect 18463 11512 18512 11540
rect 18463 11509 18475 11512
rect 18417 11503 18475 11509
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 19426 11500 19432 11552
rect 19484 11540 19490 11552
rect 20441 11543 20499 11549
rect 20441 11540 20453 11543
rect 19484 11512 20453 11540
rect 19484 11500 19490 11512
rect 20441 11509 20453 11512
rect 20487 11509 20499 11543
rect 20441 11503 20499 11509
rect 1104 11450 21620 11472
rect 1104 11398 7846 11450
rect 7898 11398 7910 11450
rect 7962 11398 7974 11450
rect 8026 11398 8038 11450
rect 8090 11398 14710 11450
rect 14762 11398 14774 11450
rect 14826 11398 14838 11450
rect 14890 11398 14902 11450
rect 14954 11398 21620 11450
rect 1104 11376 21620 11398
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3513 11339 3571 11345
rect 3513 11336 3525 11339
rect 2832 11308 3525 11336
rect 2832 11296 2838 11308
rect 3513 11305 3525 11308
rect 3559 11305 3571 11339
rect 3513 11299 3571 11305
rect 6730 11296 6736 11348
rect 6788 11336 6794 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 6788 11308 7297 11336
rect 6788 11296 6794 11308
rect 7285 11305 7297 11308
rect 7331 11336 7343 11339
rect 7469 11339 7527 11345
rect 7469 11336 7481 11339
rect 7331 11308 7481 11336
rect 7331 11305 7343 11308
rect 7285 11299 7343 11305
rect 7469 11305 7481 11308
rect 7515 11305 7527 11339
rect 7469 11299 7527 11305
rect 7742 11296 7748 11348
rect 7800 11336 7806 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7800 11308 8033 11336
rect 7800 11296 7806 11308
rect 8021 11305 8033 11308
rect 8067 11336 8079 11339
rect 8294 11336 8300 11348
rect 8067 11308 8300 11336
rect 8067 11305 8079 11308
rect 8021 11299 8079 11305
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 10870 11336 10876 11348
rect 8720 11308 10876 11336
rect 8720 11296 8726 11308
rect 10870 11296 10876 11308
rect 10928 11296 10934 11348
rect 12802 11336 12808 11348
rect 10980 11308 12808 11336
rect 3234 11268 3240 11280
rect 1872 11240 3240 11268
rect 1872 11209 1900 11240
rect 3234 11228 3240 11240
rect 3292 11268 3298 11280
rect 5902 11268 5908 11280
rect 3292 11240 3740 11268
rect 3292 11228 3298 11240
rect 3712 11212 3740 11240
rect 4264 11240 5908 11268
rect 1857 11203 1915 11209
rect 1857 11169 1869 11203
rect 1903 11169 1915 11203
rect 1857 11163 1915 11169
rect 2124 11203 2182 11209
rect 2124 11169 2136 11203
rect 2170 11200 2182 11203
rect 2682 11200 2688 11212
rect 2170 11172 2688 11200
rect 2170 11169 2182 11172
rect 2124 11163 2182 11169
rect 2682 11160 2688 11172
rect 2740 11160 2746 11212
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 4062 11200 4068 11212
rect 3752 11172 4068 11200
rect 3752 11160 3758 11172
rect 4062 11160 4068 11172
rect 4120 11200 4126 11212
rect 4264 11209 4292 11240
rect 5902 11228 5908 11240
rect 5960 11228 5966 11280
rect 5994 11228 6000 11280
rect 6052 11268 6058 11280
rect 8386 11268 8392 11280
rect 6052 11240 8392 11268
rect 6052 11228 6058 11240
rect 8386 11228 8392 11240
rect 8444 11228 8450 11280
rect 9030 11268 9036 11280
rect 8991 11240 9036 11268
rect 9030 11228 9036 11240
rect 9088 11228 9094 11280
rect 10778 11268 10784 11280
rect 9416 11240 10784 11268
rect 4249 11203 4307 11209
rect 4249 11200 4261 11203
rect 4120 11172 4261 11200
rect 4120 11160 4126 11172
rect 4249 11169 4261 11172
rect 4295 11169 4307 11203
rect 4249 11163 4307 11169
rect 4516 11203 4574 11209
rect 4516 11169 4528 11203
rect 4562 11200 4574 11203
rect 5442 11200 5448 11212
rect 4562 11172 5448 11200
rect 4562 11169 4574 11172
rect 4516 11163 4574 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 6161 11203 6219 11209
rect 6161 11200 6173 11203
rect 5644 11172 6173 11200
rect 3237 11067 3295 11073
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 3510 11064 3516 11076
rect 3283 11036 3516 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 3510 11024 3516 11036
rect 3568 11024 3574 11076
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5644 11073 5672 11172
rect 6161 11169 6173 11172
rect 6207 11169 6219 11203
rect 6161 11163 6219 11169
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7929 11203 7987 11209
rect 7929 11200 7941 11203
rect 7340 11172 7941 11200
rect 7340 11160 7346 11172
rect 7929 11169 7941 11172
rect 7975 11200 7987 11203
rect 7975 11172 8892 11200
rect 7975 11169 7987 11172
rect 7929 11163 7987 11169
rect 5902 11132 5908 11144
rect 5863 11104 5908 11132
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 7515 11104 8125 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 5629 11067 5687 11073
rect 5629 11064 5641 11067
rect 5592 11036 5641 11064
rect 5592 11024 5598 11036
rect 5629 11033 5641 11036
rect 5675 11033 5687 11067
rect 7561 11067 7619 11073
rect 5629 11027 5687 11033
rect 7208 11036 7420 11064
rect 3694 10956 3700 11008
rect 3752 10996 3758 11008
rect 7208 10996 7236 11036
rect 3752 10968 7236 10996
rect 7392 10996 7420 11036
rect 7561 11033 7573 11067
rect 7607 11064 7619 11067
rect 8202 11064 8208 11076
rect 7607 11036 8208 11064
rect 7607 11033 7619 11036
rect 7561 11027 7619 11033
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 8864 11064 8892 11172
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 8996 11172 9041 11200
rect 8996 11160 9002 11172
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11132 9275 11135
rect 9306 11132 9312 11144
rect 9263 11104 9312 11132
rect 9263 11101 9275 11104
rect 9217 11095 9275 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9416 11064 9444 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 10980 11277 11008 11308
rect 12802 11296 12808 11308
rect 12860 11296 12866 11348
rect 12897 11339 12955 11345
rect 12897 11305 12909 11339
rect 12943 11336 12955 11339
rect 12986 11336 12992 11348
rect 12943 11308 12992 11336
rect 12943 11305 12955 11308
rect 12897 11299 12955 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 15286 11336 15292 11348
rect 15247 11308 15292 11336
rect 15286 11296 15292 11308
rect 15344 11296 15350 11348
rect 16114 11296 16120 11348
rect 16172 11336 16178 11348
rect 16301 11339 16359 11345
rect 16301 11336 16313 11339
rect 16172 11308 16313 11336
rect 16172 11296 16178 11308
rect 16301 11305 16313 11308
rect 16347 11305 16359 11339
rect 18785 11339 18843 11345
rect 16301 11299 16359 11305
rect 17052 11308 18736 11336
rect 10965 11271 11023 11277
rect 10965 11237 10977 11271
rect 11011 11237 11023 11271
rect 10965 11231 11023 11237
rect 11784 11271 11842 11277
rect 11784 11237 11796 11271
rect 11830 11268 11842 11271
rect 11882 11268 11888 11280
rect 11830 11240 11888 11268
rect 11830 11237 11842 11240
rect 11784 11231 11842 11237
rect 11882 11228 11888 11240
rect 11940 11228 11946 11280
rect 12434 11228 12440 11280
rect 12492 11268 12498 11280
rect 15657 11271 15715 11277
rect 15657 11268 15669 11271
rect 12492 11240 15669 11268
rect 12492 11228 12498 11240
rect 15657 11237 15669 11240
rect 15703 11237 15715 11271
rect 15657 11231 15715 11237
rect 15930 11228 15936 11280
rect 15988 11268 15994 11280
rect 17052 11268 17080 11308
rect 15988 11240 17080 11268
rect 17120 11271 17178 11277
rect 15988 11228 15994 11240
rect 17120 11237 17132 11271
rect 17166 11268 17178 11271
rect 17494 11268 17500 11280
rect 17166 11240 17500 11268
rect 17166 11237 17178 11240
rect 17120 11231 17178 11237
rect 17494 11228 17500 11240
rect 17552 11228 17558 11280
rect 18708 11268 18736 11308
rect 18785 11305 18797 11339
rect 18831 11336 18843 11339
rect 20257 11339 20315 11345
rect 20257 11336 20269 11339
rect 18831 11308 20269 11336
rect 18831 11305 18843 11308
rect 18785 11299 18843 11305
rect 20257 11305 20269 11308
rect 20303 11305 20315 11339
rect 20257 11299 20315 11305
rect 20530 11268 20536 11280
rect 18708 11240 20536 11268
rect 20530 11228 20536 11240
rect 20588 11228 20594 11280
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9732 11172 10057 11200
rect 9732 11160 9738 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 10045 11163 10103 11169
rect 10428 11172 10701 11200
rect 10134 11132 10140 11144
rect 10095 11104 10140 11132
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10226 11092 10232 11144
rect 10284 11132 10290 11144
rect 10284 11104 10329 11132
rect 10284 11092 10290 11104
rect 8864 11036 9444 11064
rect 9677 11067 9735 11073
rect 9677 11033 9689 11067
rect 9723 11064 9735 11067
rect 10428 11064 10456 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 13078 11200 13084 11212
rect 10689 11163 10747 11169
rect 12544 11172 13084 11200
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 10652 11104 11529 11132
rect 10652 11092 10658 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 9723 11036 10456 11064
rect 9723 11033 9735 11036
rect 9677 11027 9735 11033
rect 12250 10996 12256 11008
rect 7392 10968 12256 10996
rect 3752 10956 3758 10968
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12544 10996 12572 11172
rect 13078 11160 13084 11172
rect 13136 11200 13142 11212
rect 13630 11209 13636 11212
rect 13357 11203 13415 11209
rect 13357 11200 13369 11203
rect 13136 11172 13369 11200
rect 13136 11160 13142 11172
rect 13357 11169 13369 11172
rect 13403 11169 13415 11203
rect 13624 11200 13636 11209
rect 13591 11172 13636 11200
rect 13357 11163 13415 11169
rect 13624 11163 13636 11172
rect 13630 11160 13636 11163
rect 13688 11160 13694 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 19153 11203 19211 11209
rect 19153 11200 19165 11203
rect 13964 11172 19165 11200
rect 13964 11160 13970 11172
rect 19153 11169 19165 11172
rect 19199 11169 19211 11203
rect 19153 11163 19211 11169
rect 19794 11160 19800 11212
rect 19852 11160 19858 11212
rect 20162 11200 20168 11212
rect 20123 11172 20168 11200
rect 20162 11160 20168 11172
rect 20220 11160 20226 11212
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13262 11132 13268 11144
rect 12860 11104 13268 11132
rect 12860 11092 12866 11104
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 15010 11132 15016 11144
rect 14516 11104 15016 11132
rect 14516 11092 14522 11104
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15746 11132 15752 11144
rect 15707 11104 15752 11132
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16022 11132 16028 11144
rect 15979 11104 16028 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 14737 11067 14795 11073
rect 14737 11033 14749 11067
rect 14783 11064 14795 11067
rect 15948 11064 15976 11095
rect 16022 11092 16028 11104
rect 16080 11132 16086 11144
rect 16482 11132 16488 11144
rect 16080 11104 16488 11132
rect 16080 11092 16086 11104
rect 16482 11092 16488 11104
rect 16540 11092 16546 11144
rect 16850 11132 16856 11144
rect 16811 11104 16856 11132
rect 16850 11092 16856 11104
rect 16908 11092 16914 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19426 11132 19432 11144
rect 19387 11104 19432 11132
rect 19426 11092 19432 11104
rect 19484 11092 19490 11144
rect 19812 11132 19840 11160
rect 20346 11132 20352 11144
rect 19720 11104 19840 11132
rect 20307 11104 20352 11132
rect 14783 11036 15976 11064
rect 18233 11067 18291 11073
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 18233 11033 18245 11067
rect 18279 11064 18291 11067
rect 18874 11064 18880 11076
rect 18279 11036 18880 11064
rect 18279 11033 18291 11036
rect 18233 11027 18291 11033
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 12492 10968 12572 10996
rect 12492 10956 12498 10968
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 13538 10996 13544 11008
rect 12860 10968 13544 10996
rect 12860 10956 12866 10968
rect 13538 10956 13544 10968
rect 13596 10996 13602 11008
rect 19720 10996 19748 11104
rect 20346 11092 20352 11104
rect 20404 11092 20410 11144
rect 19797 11067 19855 11073
rect 19797 11033 19809 11067
rect 19843 11064 19855 11067
rect 19886 11064 19892 11076
rect 19843 11036 19892 11064
rect 19843 11033 19855 11036
rect 19797 11027 19855 11033
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 13596 10968 19748 10996
rect 13596 10956 13602 10968
rect 1104 10906 21620 10928
rect 1104 10854 4414 10906
rect 4466 10854 4478 10906
rect 4530 10854 4542 10906
rect 4594 10854 4606 10906
rect 4658 10854 11278 10906
rect 11330 10854 11342 10906
rect 11394 10854 11406 10906
rect 11458 10854 11470 10906
rect 11522 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 18270 10906
rect 18322 10854 18334 10906
rect 18386 10854 21620 10906
rect 1104 10832 21620 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 2041 10795 2099 10801
rect 2041 10792 2053 10795
rect 1820 10764 2053 10792
rect 1820 10752 1826 10764
rect 2041 10761 2053 10764
rect 2087 10761 2099 10795
rect 2041 10755 2099 10761
rect 2958 10752 2964 10804
rect 3016 10792 3022 10804
rect 3053 10795 3111 10801
rect 3053 10792 3065 10795
rect 3016 10764 3065 10792
rect 3016 10752 3022 10764
rect 3053 10761 3065 10764
rect 3099 10761 3111 10795
rect 5442 10792 5448 10804
rect 3053 10755 3111 10761
rect 4080 10764 5304 10792
rect 5403 10764 5448 10792
rect 4080 10724 4108 10764
rect 2516 10696 4108 10724
rect 5276 10724 5304 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7616 10764 8217 10792
rect 7616 10752 7622 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9674 10792 9680 10804
rect 9079 10764 9680 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 5350 10724 5356 10736
rect 5276 10696 5356 10724
rect 2516 10665 2544 10696
rect 5350 10684 5356 10696
rect 5408 10684 5414 10736
rect 5460 10724 5488 10752
rect 8220 10724 8248 10755
rect 9674 10752 9680 10764
rect 9732 10752 9738 10804
rect 10045 10795 10103 10801
rect 10045 10761 10057 10795
rect 10091 10792 10103 10795
rect 10134 10792 10140 10804
rect 10091 10764 10140 10792
rect 10091 10761 10103 10764
rect 10045 10755 10103 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 11333 10795 11391 10801
rect 11333 10761 11345 10795
rect 11379 10792 11391 10795
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11379 10764 12173 10792
rect 11379 10761 11391 10764
rect 11333 10755 11391 10761
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 14277 10795 14335 10801
rect 14277 10761 14289 10795
rect 14323 10792 14335 10795
rect 15746 10792 15752 10804
rect 14323 10764 15752 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16485 10795 16543 10801
rect 16485 10792 16497 10795
rect 15847 10764 16497 10792
rect 9306 10724 9312 10736
rect 5460 10696 6316 10724
rect 8220 10696 9312 10724
rect 2501 10659 2559 10665
rect 2501 10625 2513 10659
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3510 10656 3516 10668
rect 2731 10628 3516 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3602 10616 3608 10668
rect 3660 10656 3666 10668
rect 3660 10628 3705 10656
rect 3660 10616 3666 10628
rect 3878 10616 3884 10668
rect 3936 10656 3942 10668
rect 6178 10656 6184 10668
rect 3936 10628 4200 10656
rect 6139 10628 6184 10656
rect 3936 10616 3942 10628
rect 2222 10548 2228 10600
rect 2280 10588 2286 10600
rect 2866 10588 2872 10600
rect 2280 10560 2872 10588
rect 2280 10548 2286 10560
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3142 10548 3148 10600
rect 3200 10588 3206 10600
rect 3421 10591 3479 10597
rect 3421 10588 3433 10591
rect 3200 10560 3433 10588
rect 3200 10548 3206 10560
rect 3421 10557 3433 10560
rect 3467 10588 3479 10591
rect 4062 10588 4068 10600
rect 3467 10560 3924 10588
rect 4023 10560 4068 10588
rect 3467 10557 3479 10560
rect 3421 10551 3479 10557
rect 3896 10532 3924 10560
rect 4062 10548 4068 10560
rect 4120 10548 4126 10600
rect 4172 10588 4200 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6288 10665 6316 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 15102 10684 15108 10736
rect 15160 10724 15166 10736
rect 15847 10724 15875 10764
rect 16485 10761 16497 10764
rect 16531 10761 16543 10795
rect 17126 10792 17132 10804
rect 17039 10764 17132 10792
rect 16485 10755 16543 10761
rect 17126 10752 17132 10764
rect 17184 10792 17190 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 17184 10764 19441 10792
rect 17184 10752 17190 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 15160 10696 15875 10724
rect 15160 10684 15166 10696
rect 6273 10659 6331 10665
rect 6273 10625 6285 10659
rect 6319 10625 6331 10659
rect 6822 10656 6828 10668
rect 6783 10628 6828 10656
rect 6273 10619 6331 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 9582 10656 9588 10668
rect 9543 10628 9588 10656
rect 9582 10616 9588 10628
rect 9640 10656 9646 10668
rect 10597 10659 10655 10665
rect 10597 10656 10609 10659
rect 9640 10628 10609 10656
rect 9640 10616 9646 10628
rect 10597 10625 10609 10628
rect 10643 10625 10655 10659
rect 11882 10656 11888 10668
rect 11843 10628 11888 10656
rect 10597 10619 10655 10625
rect 11882 10616 11888 10628
rect 11940 10616 11946 10668
rect 12434 10656 12440 10668
rect 12395 10628 12440 10656
rect 12434 10616 12440 10628
rect 12492 10616 12498 10668
rect 13630 10616 13636 10668
rect 13688 10656 13694 10668
rect 14829 10659 14887 10665
rect 14829 10656 14841 10659
rect 13688 10628 14841 10656
rect 13688 10616 13694 10628
rect 14829 10625 14841 10628
rect 14875 10656 14887 10659
rect 15654 10656 15660 10668
rect 14875 10628 15660 10656
rect 14875 10625 14887 10628
rect 14829 10619 14887 10625
rect 15654 10616 15660 10628
rect 15712 10616 15718 10668
rect 16022 10656 16028 10668
rect 15983 10628 16028 10656
rect 16022 10616 16028 10628
rect 16080 10616 16086 10668
rect 17144 10665 17172 10752
rect 17218 10684 17224 10736
rect 17276 10724 17282 10736
rect 17497 10727 17555 10733
rect 17497 10724 17509 10727
rect 17276 10696 17509 10724
rect 17276 10684 17282 10696
rect 17497 10693 17509 10696
rect 17543 10693 17555 10727
rect 17497 10687 17555 10693
rect 17129 10659 17187 10665
rect 17129 10625 17141 10659
rect 17175 10625 17187 10659
rect 17512 10656 17540 10687
rect 18049 10659 18107 10665
rect 18049 10656 18061 10659
rect 17512 10628 18061 10656
rect 17129 10619 17187 10625
rect 18049 10625 18061 10628
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 4172 10560 9505 10588
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 11793 10591 11851 10597
rect 11793 10588 11805 10591
rect 11756 10560 11805 10588
rect 11756 10548 11762 10560
rect 11793 10557 11805 10560
rect 11839 10557 11851 10591
rect 11793 10551 11851 10557
rect 12161 10591 12219 10597
rect 12161 10557 12173 10591
rect 12207 10588 12219 10591
rect 12342 10588 12348 10600
rect 12207 10560 12348 10588
rect 12207 10557 12219 10560
rect 12161 10551 12219 10557
rect 12342 10548 12348 10560
rect 12400 10548 12406 10600
rect 12704 10591 12762 10597
rect 12704 10557 12716 10591
rect 12750 10588 12762 10591
rect 12986 10588 12992 10600
rect 12750 10560 12992 10588
rect 12750 10557 12762 10560
rect 12704 10551 12762 10557
rect 12986 10548 12992 10560
rect 13044 10548 13050 10600
rect 15102 10548 15108 10600
rect 15160 10588 15166 10600
rect 17681 10591 17739 10597
rect 17681 10588 17693 10591
rect 15160 10560 17693 10588
rect 15160 10548 15166 10560
rect 17681 10557 17693 10560
rect 17727 10557 17739 10591
rect 18064 10588 18092 10619
rect 19426 10616 19432 10668
rect 19484 10656 19490 10668
rect 19484 10628 19840 10656
rect 19484 10616 19490 10628
rect 18598 10588 18604 10600
rect 18064 10560 18604 10588
rect 17681 10551 17739 10557
rect 18598 10548 18604 10560
rect 18656 10588 18662 10600
rect 19702 10588 19708 10600
rect 18656 10560 19708 10588
rect 18656 10548 18662 10560
rect 19702 10548 19708 10560
rect 19760 10548 19766 10600
rect 19812 10588 19840 10628
rect 19961 10591 20019 10597
rect 19961 10588 19973 10591
rect 19812 10560 19973 10588
rect 19961 10557 19973 10560
rect 20007 10557 20019 10591
rect 19961 10551 20019 10557
rect 3878 10480 3884 10532
rect 3936 10480 3942 10532
rect 4332 10523 4390 10529
rect 4332 10489 4344 10523
rect 4378 10520 4390 10523
rect 5166 10520 5172 10532
rect 4378 10492 5172 10520
rect 4378 10489 4390 10492
rect 4332 10483 4390 10489
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 5258 10480 5264 10532
rect 5316 10520 5322 10532
rect 6089 10523 6147 10529
rect 6089 10520 6101 10523
rect 5316 10492 6101 10520
rect 5316 10480 5322 10492
rect 6089 10489 6101 10492
rect 6135 10489 6147 10523
rect 7092 10523 7150 10529
rect 7092 10520 7104 10523
rect 6089 10483 6147 10489
rect 6932 10492 7104 10520
rect 6932 10464 6960 10492
rect 7092 10489 7104 10492
rect 7138 10489 7150 10523
rect 8573 10523 8631 10529
rect 7092 10483 7150 10489
rect 7484 10492 8340 10520
rect 2406 10452 2412 10464
rect 2367 10424 2412 10452
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6914 10412 6920 10464
rect 6972 10412 6978 10464
rect 7006 10412 7012 10464
rect 7064 10452 7070 10464
rect 7484 10452 7512 10492
rect 7064 10424 7512 10452
rect 8312 10452 8340 10492
rect 8573 10489 8585 10523
rect 8619 10520 8631 10523
rect 9401 10523 9459 10529
rect 9401 10520 9413 10523
rect 8619 10492 9413 10520
rect 8619 10489 8631 10492
rect 8573 10483 8631 10489
rect 9401 10489 9413 10492
rect 9447 10489 9459 10523
rect 12618 10520 12624 10532
rect 9401 10483 9459 10489
rect 10428 10492 12624 10520
rect 9858 10452 9864 10464
rect 8312 10424 9864 10452
rect 7064 10412 7070 10424
rect 9858 10412 9864 10424
rect 9916 10412 9922 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10428 10461 10456 10492
rect 12618 10480 12624 10492
rect 12676 10480 12682 10532
rect 14737 10523 14795 10529
rect 14737 10489 14749 10523
rect 14783 10520 14795 10523
rect 15746 10520 15752 10532
rect 14783 10492 15752 10520
rect 14783 10489 14795 10492
rect 14737 10483 14795 10489
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 15841 10523 15899 10529
rect 15841 10489 15853 10523
rect 15887 10520 15899 10523
rect 16758 10520 16764 10532
rect 15887 10492 16764 10520
rect 15887 10489 15899 10492
rect 15841 10483 15899 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 18322 10529 18328 10532
rect 18316 10520 18328 10529
rect 18283 10492 18328 10520
rect 18316 10483 18328 10492
rect 18322 10480 18328 10483
rect 18380 10480 18386 10532
rect 10413 10455 10471 10461
rect 10413 10452 10425 10455
rect 10008 10424 10425 10452
rect 10008 10412 10014 10424
rect 10413 10421 10425 10424
rect 10459 10421 10471 10455
rect 10413 10415 10471 10421
rect 10502 10412 10508 10464
rect 10560 10452 10566 10464
rect 11698 10452 11704 10464
rect 10560 10424 10605 10452
rect 11659 10424 11704 10452
rect 10560 10412 10566 10424
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11790 10412 11796 10464
rect 11848 10452 11854 10464
rect 13817 10455 13875 10461
rect 13817 10452 13829 10455
rect 11848 10424 13829 10452
rect 11848 10412 11854 10424
rect 13817 10421 13829 10424
rect 13863 10421 13875 10455
rect 13817 10415 13875 10421
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14645 10455 14703 10461
rect 14645 10452 14657 10455
rect 13964 10424 14657 10452
rect 13964 10412 13970 10424
rect 14645 10421 14657 10424
rect 14691 10421 14703 10455
rect 15470 10452 15476 10464
rect 15431 10424 15476 10452
rect 14645 10415 14703 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 15933 10455 15991 10461
rect 15933 10421 15945 10455
rect 15979 10452 15991 10455
rect 16390 10452 16396 10464
rect 15979 10424 16396 10452
rect 15979 10421 15991 10424
rect 15933 10415 15991 10421
rect 16390 10412 16396 10424
rect 16448 10412 16454 10464
rect 16850 10452 16856 10464
rect 16811 10424 16856 10452
rect 16850 10412 16856 10424
rect 16908 10412 16914 10464
rect 16945 10455 17003 10461
rect 16945 10421 16957 10455
rect 16991 10452 17003 10455
rect 17494 10452 17500 10464
rect 16991 10424 17500 10452
rect 16991 10421 17003 10424
rect 16945 10415 17003 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 20346 10412 20352 10464
rect 20404 10452 20410 10464
rect 21085 10455 21143 10461
rect 21085 10452 21097 10455
rect 20404 10424 21097 10452
rect 20404 10412 20410 10424
rect 21085 10421 21097 10424
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 1104 10362 21620 10384
rect 1104 10310 7846 10362
rect 7898 10310 7910 10362
rect 7962 10310 7974 10362
rect 8026 10310 8038 10362
rect 8090 10310 14710 10362
rect 14762 10310 14774 10362
rect 14826 10310 14838 10362
rect 14890 10310 14902 10362
rect 14954 10310 21620 10362
rect 1104 10288 21620 10310
rect 4246 10248 4252 10260
rect 4207 10220 4252 10248
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 5261 10251 5319 10257
rect 5261 10248 5273 10251
rect 4663 10220 5273 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 5261 10217 5273 10220
rect 5307 10217 5319 10251
rect 5261 10211 5319 10217
rect 5350 10208 5356 10260
rect 5408 10248 5414 10260
rect 8113 10251 8171 10257
rect 8113 10248 8125 10251
rect 5408 10220 8125 10248
rect 5408 10208 5414 10220
rect 8113 10217 8125 10220
rect 8159 10217 8171 10251
rect 8113 10211 8171 10217
rect 8294 10208 8300 10260
rect 8352 10248 8358 10260
rect 8573 10251 8631 10257
rect 8573 10248 8585 10251
rect 8352 10220 8585 10248
rect 8352 10208 8358 10220
rect 8573 10217 8585 10220
rect 8619 10217 8631 10251
rect 8573 10211 8631 10217
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 11057 10251 11115 10257
rect 11057 10248 11069 10251
rect 9640 10220 11069 10248
rect 9640 10208 9646 10220
rect 11057 10217 11069 10220
rect 11103 10217 11115 10251
rect 11057 10211 11115 10217
rect 11609 10251 11667 10257
rect 11609 10217 11621 10251
rect 11655 10217 11667 10251
rect 11974 10248 11980 10260
rect 11935 10220 11980 10248
rect 11609 10211 11667 10217
rect 3234 10180 3240 10192
rect 1780 10152 3240 10180
rect 1780 10121 1808 10152
rect 3234 10140 3240 10152
rect 3292 10140 3298 10192
rect 4709 10183 4767 10189
rect 4709 10149 4721 10183
rect 4755 10180 4767 10183
rect 5718 10180 5724 10192
rect 4755 10152 5724 10180
rect 4755 10149 4767 10152
rect 4709 10143 4767 10149
rect 5718 10140 5724 10152
rect 5776 10140 5782 10192
rect 7374 10140 7380 10192
rect 7432 10180 7438 10192
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 7432 10152 8493 10180
rect 7432 10140 7438 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 10778 10180 10784 10192
rect 8481 10143 8539 10149
rect 10244 10152 10784 10180
rect 10244 10124 10272 10152
rect 10778 10140 10784 10152
rect 10836 10140 10842 10192
rect 11624 10180 11652 10211
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 12621 10251 12679 10257
rect 12621 10248 12633 10251
rect 12584 10220 12633 10248
rect 12584 10208 12590 10220
rect 12621 10217 12633 10220
rect 12667 10217 12679 10251
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 12621 10211 12679 10217
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14829 10251 14887 10257
rect 14829 10248 14841 10251
rect 13872 10220 14841 10248
rect 13872 10208 13878 10220
rect 14829 10217 14841 10220
rect 14875 10248 14887 10251
rect 15102 10248 15108 10260
rect 14875 10220 15108 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15286 10208 15292 10260
rect 15344 10248 15350 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15344 10220 15853 10248
rect 15344 10208 15350 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16485 10251 16543 10257
rect 16485 10248 16497 10251
rect 16448 10220 16497 10248
rect 16448 10208 16454 10220
rect 16485 10217 16497 10220
rect 16531 10217 16543 10251
rect 16485 10211 16543 10217
rect 16853 10251 16911 10257
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17218 10248 17224 10260
rect 16899 10220 17224 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17218 10208 17224 10220
rect 17276 10208 17282 10260
rect 17494 10248 17500 10260
rect 17455 10220 17500 10248
rect 17494 10208 17500 10220
rect 17552 10208 17558 10260
rect 20162 10208 20168 10260
rect 20220 10248 20226 10260
rect 20349 10251 20407 10257
rect 20349 10248 20361 10251
rect 20220 10220 20361 10248
rect 20220 10208 20226 10220
rect 20349 10217 20361 10220
rect 20395 10217 20407 10251
rect 20349 10211 20407 10217
rect 12989 10183 13047 10189
rect 12989 10180 13001 10183
rect 11624 10152 13001 10180
rect 12989 10149 13001 10152
rect 13035 10149 13047 10183
rect 14458 10180 14464 10192
rect 12989 10143 13047 10149
rect 13096 10152 14464 10180
rect 2038 10121 2044 10124
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10081 1823 10115
rect 2032 10112 2044 10121
rect 1999 10084 2044 10112
rect 1765 10075 1823 10081
rect 2032 10075 2044 10084
rect 2038 10072 2044 10075
rect 2096 10072 2102 10124
rect 3510 10072 3516 10124
rect 3568 10112 3574 10124
rect 4246 10112 4252 10124
rect 3568 10084 4252 10112
rect 3568 10072 3574 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 5629 10115 5687 10121
rect 5629 10112 5641 10115
rect 4856 10084 5641 10112
rect 4856 10072 4862 10084
rect 5629 10081 5641 10084
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 6724 10115 6782 10121
rect 6724 10081 6736 10115
rect 6770 10112 6782 10115
rect 7558 10112 7564 10124
rect 6770 10084 7564 10112
rect 6770 10081 6782 10084
rect 6724 10075 6782 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7668 10084 7972 10112
rect 4893 10047 4951 10053
rect 4893 10013 4905 10047
rect 4939 10044 4951 10047
rect 5534 10044 5540 10056
rect 4939 10016 5540 10044
rect 4939 10013 4951 10016
rect 4893 10007 4951 10013
rect 5534 10004 5540 10016
rect 5592 10004 5598 10056
rect 5718 10044 5724 10056
rect 5679 10016 5724 10044
rect 5718 10004 5724 10016
rect 5776 10004 5782 10056
rect 5813 10047 5871 10053
rect 5813 10013 5825 10047
rect 5859 10013 5871 10047
rect 5813 10007 5871 10013
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 5350 9976 5356 9988
rect 4672 9948 5356 9976
rect 4672 9936 4678 9948
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 5442 9936 5448 9988
rect 5500 9976 5506 9988
rect 5828 9976 5856 10007
rect 5902 10004 5908 10056
rect 5960 10044 5966 10056
rect 6178 10044 6184 10056
rect 5960 10016 6184 10044
rect 5960 10004 5966 10016
rect 6178 10004 6184 10016
rect 6236 10044 6242 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6236 10016 6469 10044
rect 6236 10004 6242 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 7668 9976 7696 10084
rect 7944 10044 7972 10084
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 9490 10112 9496 10124
rect 8444 10084 9496 10112
rect 8444 10072 8450 10084
rect 9490 10072 9496 10084
rect 9548 10112 9554 10124
rect 9677 10115 9735 10121
rect 9677 10112 9689 10115
rect 9548 10084 9689 10112
rect 9548 10072 9554 10084
rect 9677 10081 9689 10084
rect 9723 10081 9735 10115
rect 9677 10075 9735 10081
rect 9944 10115 10002 10121
rect 9944 10081 9956 10115
rect 9990 10112 10002 10115
rect 10226 10112 10232 10124
rect 9990 10084 10232 10112
rect 9990 10081 10002 10084
rect 9944 10075 10002 10081
rect 10226 10072 10232 10084
rect 10284 10072 10290 10124
rect 11054 10072 11060 10124
rect 11112 10112 11118 10124
rect 11698 10112 11704 10124
rect 11112 10084 11704 10112
rect 11112 10072 11118 10084
rect 11698 10072 11704 10084
rect 11756 10112 11762 10124
rect 13096 10112 13124 10152
rect 14458 10140 14464 10152
rect 14516 10140 14522 10192
rect 15470 10140 15476 10192
rect 15528 10180 15534 10192
rect 15933 10183 15991 10189
rect 15933 10180 15945 10183
rect 15528 10152 15945 10180
rect 15528 10140 15534 10152
rect 15933 10149 15945 10152
rect 15979 10149 15991 10183
rect 15933 10143 15991 10149
rect 16945 10183 17003 10189
rect 16945 10149 16957 10183
rect 16991 10180 17003 10183
rect 17957 10183 18015 10189
rect 17957 10180 17969 10183
rect 16991 10152 17969 10180
rect 16991 10149 17003 10152
rect 16945 10143 17003 10149
rect 17957 10149 17969 10152
rect 18003 10180 18015 10183
rect 19058 10180 19064 10192
rect 18003 10152 19064 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 19058 10140 19064 10152
rect 19116 10180 19122 10192
rect 20622 10180 20628 10192
rect 19116 10152 20628 10180
rect 19116 10140 19122 10152
rect 20622 10140 20628 10152
rect 20680 10140 20686 10192
rect 11756 10084 13124 10112
rect 11756 10072 11762 10084
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13412 10084 13645 10112
rect 13412 10072 13418 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 13633 10075 13691 10081
rect 13998 10072 14004 10124
rect 14056 10112 14062 10124
rect 14553 10115 14611 10121
rect 14553 10112 14565 10115
rect 14056 10084 14565 10112
rect 14056 10072 14062 10084
rect 14553 10081 14565 10084
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 15194 10112 15200 10124
rect 15059 10084 15200 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 7944 10016 8677 10044
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 5500 9948 5856 9976
rect 7392 9948 7696 9976
rect 5500 9936 5506 9948
rect 3142 9908 3148 9920
rect 3055 9880 3148 9908
rect 3142 9868 3148 9880
rect 3200 9908 3206 9920
rect 7392 9908 7420 9948
rect 7742 9936 7748 9988
rect 7800 9976 7806 9988
rect 7837 9979 7895 9985
rect 7837 9976 7849 9979
rect 7800 9948 7849 9976
rect 7800 9936 7806 9948
rect 7837 9945 7849 9948
rect 7883 9945 7895 9979
rect 7837 9939 7895 9945
rect 7926 9936 7932 9988
rect 7984 9976 7990 9988
rect 8478 9976 8484 9988
rect 7984 9948 8484 9976
rect 7984 9936 7990 9948
rect 8478 9936 8484 9948
rect 8536 9936 8542 9988
rect 12084 9976 12112 10007
rect 12158 10004 12164 10056
rect 12216 10044 12222 10056
rect 12216 10016 12261 10044
rect 12216 10004 12222 10016
rect 12710 10004 12716 10056
rect 12768 10044 12774 10056
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12768 10016 13185 10044
rect 12768 10004 12774 10016
rect 13173 10013 13185 10016
rect 13219 10013 13231 10047
rect 13173 10007 13231 10013
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 13817 10047 13875 10053
rect 13817 10044 13829 10047
rect 13780 10016 13829 10044
rect 13780 10004 13786 10016
rect 13817 10013 13829 10016
rect 13863 10013 13875 10047
rect 13817 10007 13875 10013
rect 12250 9976 12256 9988
rect 12084 9948 12256 9976
rect 12250 9936 12256 9948
rect 12308 9936 12314 9988
rect 12342 9936 12348 9988
rect 12400 9976 12406 9988
rect 14369 9979 14427 9985
rect 12400 9948 12664 9976
rect 12400 9936 12406 9948
rect 3200 9880 7420 9908
rect 3200 9868 3206 9880
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 10962 9908 10968 9920
rect 7524 9880 10968 9908
rect 7524 9868 7530 9880
rect 10962 9868 10968 9880
rect 11020 9868 11026 9920
rect 12636 9908 12664 9948
rect 14369 9945 14381 9979
rect 14415 9976 14427 9979
rect 15028 9976 15056 10075
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 15712 10084 17080 10112
rect 15712 10072 15718 10084
rect 17052 10056 17080 10084
rect 17494 10072 17500 10124
rect 17552 10112 17558 10124
rect 17865 10115 17923 10121
rect 17865 10112 17877 10115
rect 17552 10084 17877 10112
rect 17552 10072 17558 10084
rect 17865 10081 17877 10084
rect 17911 10081 17923 10115
rect 17865 10075 17923 10081
rect 18598 10072 18604 10124
rect 18656 10112 18662 10124
rect 18693 10115 18751 10121
rect 18693 10112 18705 10115
rect 18656 10084 18705 10112
rect 18656 10072 18662 10084
rect 18693 10081 18705 10084
rect 18739 10081 18751 10115
rect 18693 10075 18751 10081
rect 18960 10115 19018 10121
rect 18960 10081 18972 10115
rect 19006 10112 19018 10115
rect 19794 10112 19800 10124
rect 19006 10084 19800 10112
rect 19006 10081 19018 10084
rect 18960 10075 19018 10081
rect 19794 10072 19800 10084
rect 19852 10072 19858 10124
rect 15838 10004 15844 10056
rect 15896 10044 15902 10056
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15896 10016 16037 10044
rect 15896 10004 15902 10016
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 17034 10044 17040 10056
rect 16947 10016 17040 10044
rect 16025 10007 16083 10013
rect 17034 10004 17040 10016
rect 17092 10004 17098 10056
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10044 18199 10047
rect 18322 10044 18328 10056
rect 18187 10016 18328 10044
rect 18187 10013 18199 10016
rect 18141 10007 18199 10013
rect 18322 10004 18328 10016
rect 18380 10044 18386 10056
rect 18380 10016 18644 10044
rect 18380 10004 18386 10016
rect 14415 9948 15056 9976
rect 15473 9979 15531 9985
rect 14415 9945 14427 9948
rect 14369 9939 14427 9945
rect 15473 9945 15485 9979
rect 15519 9976 15531 9979
rect 17402 9976 17408 9988
rect 15519 9948 17408 9976
rect 15519 9945 15531 9948
rect 15473 9939 15531 9945
rect 17402 9936 17408 9948
rect 17460 9936 17466 9988
rect 18046 9936 18052 9988
rect 18104 9936 18110 9988
rect 13630 9908 13636 9920
rect 12636 9880 13636 9908
rect 13630 9868 13636 9880
rect 13688 9908 13694 9920
rect 18064 9908 18092 9936
rect 13688 9880 18092 9908
rect 18616 9908 18644 10016
rect 20073 9911 20131 9917
rect 20073 9908 20085 9911
rect 18616 9880 20085 9908
rect 13688 9868 13694 9880
rect 20073 9877 20085 9880
rect 20119 9877 20131 9911
rect 20073 9871 20131 9877
rect 1104 9818 21620 9840
rect 1104 9766 4414 9818
rect 4466 9766 4478 9818
rect 4530 9766 4542 9818
rect 4594 9766 4606 9818
rect 4658 9766 11278 9818
rect 11330 9766 11342 9818
rect 11394 9766 11406 9818
rect 11458 9766 11470 9818
rect 11522 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 18270 9818
rect 18322 9766 18334 9818
rect 18386 9766 21620 9818
rect 1104 9744 21620 9766
rect 1857 9707 1915 9713
rect 1857 9673 1869 9707
rect 1903 9704 1915 9707
rect 2406 9704 2412 9716
rect 1903 9676 2412 9704
rect 1903 9673 1915 9676
rect 1857 9667 1915 9673
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2682 9704 2688 9716
rect 2595 9676 2688 9704
rect 2682 9664 2688 9676
rect 2740 9704 2746 9716
rect 3142 9704 3148 9716
rect 2740 9676 3148 9704
rect 2740 9664 2746 9676
rect 3142 9664 3148 9676
rect 3200 9664 3206 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 7466 9704 7472 9716
rect 4120 9676 7472 9704
rect 4120 9664 4126 9676
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 7834 9664 7840 9716
rect 7892 9704 7898 9716
rect 10226 9704 10232 9716
rect 7892 9676 10088 9704
rect 10187 9676 10232 9704
rect 7892 9664 7898 9676
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 2317 9571 2375 9577
rect 2317 9568 2329 9571
rect 1912 9540 2329 9568
rect 1912 9528 1918 9540
rect 2317 9537 2329 9540
rect 2363 9537 2375 9571
rect 2317 9531 2375 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2700 9568 2728 9664
rect 2866 9636 2872 9648
rect 2827 9608 2872 9636
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 4890 9636 4896 9648
rect 3344 9608 4896 9636
rect 3344 9577 3372 9608
rect 4890 9596 4896 9608
rect 4948 9596 4954 9648
rect 4982 9596 4988 9648
rect 5040 9636 5046 9648
rect 5442 9636 5448 9648
rect 5040 9608 5448 9636
rect 5040 9596 5046 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5537 9639 5595 9645
rect 5537 9605 5549 9639
rect 5583 9636 5595 9639
rect 5626 9636 5632 9648
rect 5583 9608 5632 9636
rect 5583 9605 5595 9608
rect 5537 9599 5595 9605
rect 5626 9596 5632 9608
rect 5684 9596 5690 9648
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 6696 9608 6837 9636
rect 6696 9596 6702 9608
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 6972 9608 7512 9636
rect 6972 9596 6978 9608
rect 2547 9540 2728 9568
rect 3329 9571 3387 9577
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9568 3479 9571
rect 3602 9568 3608 9580
rect 3467 9540 3608 9568
rect 3467 9537 3479 9540
rect 3421 9531 3479 9537
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 2225 9503 2283 9509
rect 2225 9500 2237 9503
rect 1452 9472 2237 9500
rect 1452 9460 1458 9472
rect 2225 9469 2237 9472
rect 2271 9469 2283 9503
rect 2225 9463 2283 9469
rect 2682 9460 2688 9512
rect 2740 9500 2746 9512
rect 3436 9500 3464 9531
rect 3602 9528 3608 9540
rect 3660 9568 3666 9580
rect 4525 9571 4583 9577
rect 4525 9568 4537 9571
rect 3660 9540 4537 9568
rect 3660 9528 3666 9540
rect 4525 9537 4537 9540
rect 4571 9537 4583 9571
rect 4525 9531 4583 9537
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 7282 9568 7288 9580
rect 6227 9540 7288 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7484 9577 7512 9608
rect 7558 9596 7564 9648
rect 7616 9636 7622 9648
rect 10060 9636 10088 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 10502 9704 10508 9716
rect 10463 9676 10508 9704
rect 10502 9664 10508 9676
rect 10560 9664 10566 9716
rect 12342 9704 12348 9716
rect 10612 9676 12348 9704
rect 10612 9636 10640 9676
rect 12342 9664 12348 9676
rect 12400 9664 12406 9716
rect 12618 9704 12624 9716
rect 12452 9676 12624 9704
rect 12452 9636 12480 9676
rect 12618 9664 12624 9676
rect 12676 9704 12682 9716
rect 12802 9704 12808 9716
rect 12676 9676 12808 9704
rect 12676 9664 12682 9676
rect 12802 9664 12808 9676
rect 12860 9664 12866 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14231 9676 17080 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 7616 9608 8432 9636
rect 10060 9608 10640 9636
rect 10704 9608 11836 9636
rect 7616 9596 7622 9608
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 7742 9568 7748 9580
rect 7515 9540 7748 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 7742 9528 7748 9540
rect 7800 9528 7806 9580
rect 8202 9528 8208 9580
rect 8260 9568 8266 9580
rect 8404 9577 8432 9608
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 8260 9540 8309 9568
rect 8260 9528 8266 9540
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 8389 9571 8447 9577
rect 8389 9537 8401 9571
rect 8435 9537 8447 9571
rect 8389 9531 8447 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8536 9540 8861 9568
rect 8536 9528 8542 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 8849 9531 8907 9537
rect 10060 9540 10425 9568
rect 2740 9472 3464 9500
rect 2740 9460 2746 9472
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 4246 9500 4252 9512
rect 3752 9472 4252 9500
rect 3752 9460 3758 9472
rect 4246 9460 4252 9472
rect 4304 9500 4310 9512
rect 4341 9503 4399 9509
rect 4341 9500 4353 9503
rect 4304 9472 4353 9500
rect 4304 9460 4310 9472
rect 4341 9469 4353 9472
rect 4387 9469 4399 9503
rect 4341 9463 4399 9469
rect 4430 9460 4436 9512
rect 4488 9500 4494 9512
rect 5905 9503 5963 9509
rect 5905 9500 5917 9503
rect 4488 9472 5917 9500
rect 4488 9460 4494 9472
rect 5905 9469 5917 9472
rect 5951 9469 5963 9503
rect 5905 9463 5963 9469
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 10060 9500 10088 9540
rect 10413 9537 10425 9540
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10704 9500 10732 9608
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11808 9577 11836 9608
rect 11992 9608 12480 9636
rect 11992 9577 12020 9608
rect 16758 9596 16764 9648
rect 16816 9636 16822 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16816 9608 16957 9636
rect 16816 9596 16822 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 17052 9636 17080 9676
rect 17126 9664 17132 9716
rect 17184 9704 17190 9716
rect 20070 9704 20076 9716
rect 17184 9676 20076 9704
rect 17184 9664 17190 9676
rect 20070 9664 20076 9676
rect 20128 9664 20134 9716
rect 19610 9636 19616 9648
rect 17052 9608 19616 9636
rect 16945 9599 17003 9605
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 11057 9571 11115 9577
rect 11057 9568 11069 9571
rect 10836 9540 11069 9568
rect 10836 9528 10842 9540
rect 11057 9537 11069 9540
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9537 12035 9571
rect 14829 9571 14887 9577
rect 11977 9531 12035 9537
rect 12268 9540 12572 9568
rect 6052 9472 10088 9500
rect 10152 9472 10732 9500
rect 6052 9460 6058 9472
rect 7098 9432 7104 9444
rect 3988 9404 7104 9432
rect 2958 9324 2964 9376
rect 3016 9364 3022 9376
rect 3988 9373 4016 9404
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 7466 9392 7472 9444
rect 7524 9432 7530 9444
rect 8205 9435 8263 9441
rect 8205 9432 8217 9435
rect 7524 9404 8217 9432
rect 7524 9392 7530 9404
rect 8205 9401 8217 9404
rect 8251 9401 8263 9435
rect 8205 9395 8263 9401
rect 9116 9435 9174 9441
rect 9116 9401 9128 9435
rect 9162 9432 9174 9435
rect 9858 9432 9864 9444
rect 9162 9404 9864 9432
rect 9162 9401 9174 9404
rect 9116 9395 9174 9401
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 3237 9367 3295 9373
rect 3237 9364 3249 9367
rect 3016 9336 3249 9364
rect 3016 9324 3022 9336
rect 3237 9333 3249 9336
rect 3283 9333 3295 9367
rect 3237 9327 3295 9333
rect 3973 9367 4031 9373
rect 3973 9333 3985 9367
rect 4019 9333 4031 9367
rect 4430 9364 4436 9376
rect 4391 9336 4436 9364
rect 3973 9327 4031 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5997 9367 6055 9373
rect 5997 9364 6009 9367
rect 4672 9336 6009 9364
rect 4672 9324 4678 9336
rect 5997 9333 6009 9336
rect 6043 9333 6055 9367
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 5997 9327 6055 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7331 9336 7849 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 10152 9364 10180 9472
rect 10870 9460 10876 9512
rect 10928 9500 10934 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 10928 9472 10977 9500
rect 10928 9460 10934 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 12268 9500 12296 9540
rect 10965 9463 11023 9469
rect 11072 9472 12296 9500
rect 10413 9435 10471 9441
rect 10413 9401 10425 9435
rect 10459 9432 10471 9435
rect 11072 9432 11100 9472
rect 12342 9460 12348 9512
rect 12400 9500 12406 9512
rect 12437 9503 12495 9509
rect 12437 9500 12449 9503
rect 12400 9472 12449 9500
rect 12400 9460 12406 9472
rect 12437 9469 12449 9472
rect 12483 9469 12495 9503
rect 12544 9500 12572 9540
rect 14829 9537 14841 9571
rect 14875 9568 14887 9571
rect 15654 9568 15660 9580
rect 14875 9540 15660 9568
rect 14875 9537 14887 9540
rect 14829 9531 14887 9537
rect 15654 9528 15660 9540
rect 15712 9528 15718 9580
rect 15746 9528 15752 9580
rect 15804 9568 15810 9580
rect 15804 9540 15849 9568
rect 15804 9528 15810 9540
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 17092 9540 17509 9568
rect 17092 9528 17098 9540
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 19702 9568 19708 9580
rect 19663 9540 19708 9568
rect 17497 9531 17555 9537
rect 19702 9528 19708 9540
rect 19760 9528 19766 9580
rect 19972 9503 20030 9509
rect 12544 9472 16344 9500
rect 12437 9463 12495 9469
rect 12526 9432 12532 9444
rect 10459 9404 11100 9432
rect 11348 9404 12532 9432
rect 10459 9401 10471 9404
rect 10413 9395 10471 9401
rect 8352 9336 10180 9364
rect 8352 9324 8358 9336
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10284 9336 10885 9364
rect 10284 9324 10290 9336
rect 10873 9333 10885 9336
rect 10919 9364 10931 9367
rect 10962 9364 10968 9376
rect 10919 9336 10968 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11348 9373 11376 9404
rect 12526 9392 12532 9404
rect 12584 9392 12590 9444
rect 12710 9441 12716 9444
rect 12704 9432 12716 9441
rect 12671 9404 12716 9432
rect 12704 9395 12716 9404
rect 12710 9392 12716 9395
rect 12768 9392 12774 9444
rect 13446 9392 13452 9444
rect 13504 9432 13510 9444
rect 14182 9432 14188 9444
rect 13504 9404 14188 9432
rect 13504 9392 13510 9404
rect 14182 9392 14188 9404
rect 14240 9392 14246 9444
rect 14645 9435 14703 9441
rect 14645 9401 14657 9435
rect 14691 9432 14703 9435
rect 15102 9432 15108 9444
rect 14691 9404 15108 9432
rect 14691 9401 14703 9404
rect 14645 9395 14703 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 16209 9435 16267 9441
rect 16209 9432 16221 9435
rect 15611 9404 16221 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16209 9401 16221 9404
rect 16255 9401 16267 9435
rect 16316 9432 16344 9472
rect 19972 9469 19984 9503
rect 20018 9500 20030 9503
rect 20346 9500 20352 9512
rect 20018 9472 20352 9500
rect 20018 9469 20030 9472
rect 19972 9463 20030 9469
rect 20346 9460 20352 9472
rect 20404 9460 20410 9512
rect 16316 9404 21128 9432
rect 16209 9395 16267 9401
rect 11333 9367 11391 9373
rect 11333 9333 11345 9367
rect 11379 9333 11391 9367
rect 11698 9364 11704 9376
rect 11659 9336 11704 9364
rect 11333 9327 11391 9333
rect 11698 9324 11704 9336
rect 11756 9324 11762 9376
rect 13814 9364 13820 9376
rect 13775 9336 13820 9364
rect 13814 9324 13820 9336
rect 13872 9324 13878 9376
rect 14550 9364 14556 9376
rect 14511 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15286 9364 15292 9376
rect 15243 9336 15292 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15528 9336 15669 9364
rect 15528 9324 15534 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 17310 9364 17316 9376
rect 17271 9336 17316 9364
rect 15657 9327 15715 9333
rect 17310 9324 17316 9336
rect 17368 9324 17374 9376
rect 17405 9367 17463 9373
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17494 9364 17500 9376
rect 17451 9336 17500 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 21100 9373 21128 9404
rect 21085 9367 21143 9373
rect 21085 9333 21097 9367
rect 21131 9333 21143 9367
rect 21085 9327 21143 9333
rect 1104 9274 21620 9296
rect 1104 9222 7846 9274
rect 7898 9222 7910 9274
rect 7962 9222 7974 9274
rect 8026 9222 8038 9274
rect 8090 9222 14710 9274
rect 14762 9222 14774 9274
rect 14826 9222 14838 9274
rect 14890 9222 14902 9274
rect 14954 9222 21620 9274
rect 1104 9200 21620 9222
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2314 9160 2320 9172
rect 2087 9132 2320 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 2314 9120 2320 9132
rect 2372 9120 2378 9172
rect 2409 9163 2467 9169
rect 2409 9129 2421 9163
rect 2455 9160 2467 9163
rect 2498 9160 2504 9172
rect 2455 9132 2504 9160
rect 2455 9129 2467 9132
rect 2409 9123 2467 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 3050 9160 3056 9172
rect 3011 9132 3056 9160
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 4433 9163 4491 9169
rect 4433 9129 4445 9163
rect 4479 9160 4491 9163
rect 4798 9160 4804 9172
rect 4479 9132 4804 9160
rect 4479 9129 4491 9132
rect 4433 9123 4491 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 8404 9132 12480 9160
rect 3418 9052 3424 9104
rect 3476 9092 3482 9104
rect 8294 9092 8300 9104
rect 3476 9064 8300 9092
rect 3476 9052 3482 9064
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 4614 9024 4620 9036
rect 2608 8996 4620 9024
rect 2608 8968 2636 8996
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4801 9027 4859 9033
rect 4801 8993 4813 9027
rect 4847 9024 4859 9027
rect 5445 9027 5503 9033
rect 5445 9024 5457 9027
rect 4847 8996 5457 9024
rect 4847 8993 4859 8996
rect 4801 8987 4859 8993
rect 5445 8993 5457 8996
rect 5491 8993 5503 9027
rect 6178 9024 6184 9036
rect 6139 8996 6184 9024
rect 5445 8987 5503 8993
rect 6178 8984 6184 8996
rect 6236 8984 6242 9036
rect 6448 9027 6506 9033
rect 6448 8993 6460 9027
rect 6494 9024 6506 9027
rect 6730 9024 6736 9036
rect 6494 8996 6736 9024
rect 6494 8993 6506 8996
rect 6448 8987 6506 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8202 9024 8208 9036
rect 8067 8996 8208 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8404 9024 8432 9132
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8628 9064 9045 9092
rect 8628 9052 8634 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 11606 9092 11612 9104
rect 9033 9055 9091 9061
rect 9784 9064 11612 9092
rect 8481 9027 8539 9033
rect 8481 9024 8493 9027
rect 8404 8996 8493 9024
rect 8481 8993 8493 8996
rect 8527 8993 8539 9027
rect 8481 8987 8539 8993
rect 8941 9027 8999 9033
rect 8941 8993 8953 9027
rect 8987 8993 8999 9027
rect 8941 8987 8999 8993
rect 2501 8959 2559 8965
rect 2501 8925 2513 8959
rect 2547 8956 2559 8959
rect 2590 8956 2596 8968
rect 2547 8928 2596 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 2590 8916 2596 8928
rect 2648 8916 2654 8968
rect 2682 8916 2688 8968
rect 2740 8956 2746 8968
rect 4890 8956 4896 8968
rect 2740 8928 2785 8956
rect 4851 8928 4896 8956
rect 2740 8916 2746 8928
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 5077 8959 5135 8965
rect 5077 8925 5089 8959
rect 5123 8956 5135 8959
rect 5166 8956 5172 8968
rect 5123 8928 5172 8956
rect 5123 8925 5135 8928
rect 5077 8919 5135 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8956 8956 8984 8987
rect 8168 8928 8984 8956
rect 8168 8916 8174 8928
rect 9030 8916 9036 8968
rect 9088 8956 9094 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 9088 8928 9137 8956
rect 9088 8916 9094 8928
rect 9125 8925 9137 8928
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 6178 8888 6184 8900
rect 4488 8860 6184 8888
rect 4488 8848 4494 8860
rect 6178 8848 6184 8860
rect 6236 8848 6242 8900
rect 7558 8888 7564 8900
rect 7519 8860 7564 8888
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 7837 8891 7895 8897
rect 7837 8888 7849 8891
rect 7800 8860 7849 8888
rect 7800 8848 7806 8860
rect 7837 8857 7849 8860
rect 7883 8857 7895 8891
rect 9784 8888 9812 9064
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 12452 9101 12480 9132
rect 12710 9120 12716 9172
rect 12768 9160 12774 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 12768 9132 13921 9160
rect 12768 9120 12774 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 14185 9163 14243 9169
rect 14185 9129 14197 9163
rect 14231 9160 14243 9163
rect 14550 9160 14556 9172
rect 14231 9132 14556 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 15013 9163 15071 9169
rect 15013 9129 15025 9163
rect 15059 9160 15071 9163
rect 15286 9160 15292 9172
rect 15059 9132 15292 9160
rect 15059 9129 15071 9132
rect 15013 9123 15071 9129
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 15654 9120 15660 9172
rect 15712 9160 15718 9172
rect 16022 9160 16028 9172
rect 15712 9132 16028 9160
rect 15712 9120 15718 9132
rect 16022 9120 16028 9132
rect 16080 9160 16086 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16080 9132 16681 9160
rect 16080 9120 16086 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 19794 9160 19800 9172
rect 19755 9132 19800 9160
rect 16669 9123 16727 9129
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20036 9132 20453 9160
rect 20036 9120 20042 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 12437 9095 12495 9101
rect 12437 9061 12449 9095
rect 12483 9092 12495 9095
rect 13998 9092 14004 9104
rect 12483 9064 14004 9092
rect 12483 9061 12495 9064
rect 12437 9055 12495 9061
rect 13998 9052 14004 9064
rect 14056 9052 14062 9104
rect 15746 9092 15752 9104
rect 14476 9064 15752 9092
rect 10042 9024 10048 9036
rect 10003 8996 10048 9024
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 10689 9027 10747 9033
rect 10689 8993 10701 9027
rect 10735 9024 10747 9027
rect 10962 9024 10968 9036
rect 10735 8996 10968 9024
rect 10735 8993 10747 8996
rect 10689 8987 10747 8993
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 12529 9027 12587 9033
rect 12529 8993 12541 9027
rect 12575 9024 12587 9027
rect 12618 9024 12624 9036
rect 12575 8996 12624 9024
rect 12575 8993 12587 8996
rect 12529 8987 12587 8993
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12796 9027 12854 9033
rect 12796 8993 12808 9027
rect 12842 9024 12854 9027
rect 13170 9024 13176 9036
rect 12842 8996 13176 9024
rect 12842 8993 12854 8996
rect 12796 8987 12854 8993
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 14476 9024 14504 9064
rect 15746 9052 15752 9064
rect 15804 9052 15810 9104
rect 17310 9092 17316 9104
rect 17223 9064 17316 9092
rect 17310 9052 17316 9064
rect 17368 9092 17374 9104
rect 18598 9092 18604 9104
rect 17368 9064 18604 9092
rect 17368 9052 17374 9064
rect 18598 9052 18604 9064
rect 18656 9052 18662 9104
rect 13872 8996 14504 9024
rect 14553 9027 14611 9033
rect 13872 8984 13878 8996
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 15013 9027 15071 9033
rect 15013 9024 15025 9027
rect 14599 8996 15025 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 15013 8993 15025 8996
rect 15059 8993 15071 9027
rect 15545 9027 15603 9033
rect 15545 9024 15557 9027
rect 15013 8987 15071 8993
rect 15212 8996 15557 9024
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10229 8959 10287 8965
rect 10229 8925 10241 8959
rect 10275 8925 10287 8959
rect 10229 8919 10287 8925
rect 7837 8851 7895 8857
rect 7935 8860 9812 8888
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 7935 8820 7963 8860
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10244 8888 10272 8919
rect 13906 8916 13912 8968
rect 13964 8956 13970 8968
rect 14645 8959 14703 8965
rect 14645 8956 14657 8959
rect 13964 8928 14657 8956
rect 13964 8916 13970 8928
rect 14645 8925 14657 8928
rect 14691 8925 14703 8959
rect 14826 8956 14832 8968
rect 14787 8928 14832 8956
rect 14645 8919 14703 8925
rect 14826 8916 14832 8928
rect 14884 8956 14890 8968
rect 15212 8956 15240 8996
rect 15545 8993 15557 8996
rect 15591 8993 15603 9027
rect 15764 9024 15792 9052
rect 18684 9027 18742 9033
rect 15764 8996 17540 9024
rect 15545 8987 15603 8993
rect 14884 8928 15240 8956
rect 14884 8916 14890 8928
rect 15286 8916 15292 8968
rect 15344 8956 15350 8968
rect 15344 8928 15389 8956
rect 15344 8916 15350 8928
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17512 8965 17540 8996
rect 18684 8993 18696 9027
rect 18730 9024 18742 9027
rect 19058 9024 19064 9036
rect 18730 8996 19064 9024
rect 18730 8993 18742 8996
rect 18684 8987 18742 8993
rect 19058 8984 19064 8996
rect 19116 8984 19122 9036
rect 19610 8984 19616 9036
rect 19668 9024 19674 9036
rect 20257 9027 20315 9033
rect 20257 9024 20269 9027
rect 19668 8996 20269 9024
rect 19668 8984 19674 8996
rect 20257 8993 20269 8996
rect 20303 8993 20315 9027
rect 20257 8987 20315 8993
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17368 8928 17417 8956
rect 17368 8916 17374 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 17497 8959 17555 8965
rect 17497 8925 17509 8959
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 17644 8928 18429 8956
rect 17644 8916 17650 8928
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 9916 8860 10272 8888
rect 9916 8848 9922 8860
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 11698 8888 11704 8900
rect 10560 8860 11704 8888
rect 10560 8848 10566 8860
rect 11698 8848 11704 8860
rect 11756 8848 11762 8900
rect 12066 8848 12072 8900
rect 12124 8888 12130 8900
rect 12342 8888 12348 8900
rect 12124 8860 12348 8888
rect 12124 8848 12130 8860
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 16224 8860 17356 8888
rect 4120 8792 7963 8820
rect 4120 8780 4126 8792
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8297 8823 8355 8829
rect 8297 8820 8309 8823
rect 8260 8792 8309 8820
rect 8260 8780 8266 8792
rect 8297 8789 8309 8792
rect 8343 8789 8355 8823
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8297 8783 8355 8789
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 9677 8823 9735 8829
rect 9677 8789 9689 8823
rect 9723 8820 9735 8823
rect 10778 8820 10784 8832
rect 9723 8792 10784 8820
rect 9723 8789 9735 8792
rect 9677 8783 9735 8789
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 16224 8820 16252 8860
rect 16942 8820 16948 8832
rect 10928 8792 16252 8820
rect 16903 8792 16948 8820
rect 10928 8780 10934 8792
rect 16942 8780 16948 8792
rect 17000 8780 17006 8832
rect 17328 8820 17356 8860
rect 18782 8820 18788 8832
rect 17328 8792 18788 8820
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 1104 8730 21620 8752
rect 1104 8678 4414 8730
rect 4466 8678 4478 8730
rect 4530 8678 4542 8730
rect 4594 8678 4606 8730
rect 4658 8678 11278 8730
rect 11330 8678 11342 8730
rect 11394 8678 11406 8730
rect 11458 8678 11470 8730
rect 11522 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 18270 8730
rect 18322 8678 18334 8730
rect 18386 8678 21620 8730
rect 1104 8656 21620 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 3234 8616 3240 8628
rect 2096 8588 3240 8616
rect 2096 8576 2102 8588
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 4154 8616 4160 8628
rect 4115 8588 4160 8616
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 5074 8576 5080 8628
rect 5132 8616 5138 8628
rect 6638 8616 6644 8628
rect 5132 8588 6644 8616
rect 5132 8576 5138 8588
rect 6638 8576 6644 8588
rect 6696 8576 6702 8628
rect 6825 8619 6883 8625
rect 6825 8585 6837 8619
rect 6871 8616 6883 8619
rect 7190 8616 7196 8628
rect 6871 8588 7196 8616
rect 6871 8585 6883 8588
rect 6825 8579 6883 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 9674 8616 9680 8628
rect 8496 8588 9680 8616
rect 4062 8508 4068 8560
rect 4120 8548 4126 8560
rect 8496 8548 8524 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 9858 8616 9864 8628
rect 9819 8588 9864 8616
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 12069 8619 12127 8625
rect 12069 8585 12081 8619
rect 12115 8616 12127 8619
rect 12158 8616 12164 8628
rect 12115 8588 12164 8616
rect 12115 8585 12127 8588
rect 12069 8579 12127 8585
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 17954 8616 17960 8628
rect 12492 8588 17960 8616
rect 12492 8576 12498 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18969 8619 19027 8625
rect 18969 8585 18981 8619
rect 19015 8616 19027 8619
rect 19150 8616 19156 8628
rect 19015 8588 19156 8616
rect 19015 8585 19027 8588
rect 18969 8579 19027 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 4120 8520 8524 8548
rect 12176 8548 12204 8576
rect 14826 8548 14832 8560
rect 12176 8520 13124 8548
rect 14739 8520 14832 8548
rect 4120 8508 4126 8520
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 3752 8452 4721 8480
rect 3752 8440 3758 8452
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 5994 8480 6000 8492
rect 5859 8452 6000 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 5994 8440 6000 8452
rect 6052 8440 6058 8492
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7285 8483 7343 8489
rect 7285 8480 7297 8483
rect 6880 8452 7297 8480
rect 6880 8440 6886 8452
rect 7285 8449 7297 8452
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 7558 8480 7564 8492
rect 7515 8452 7564 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 8110 8480 8116 8492
rect 8067 8452 8116 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8480 12219 8483
rect 12802 8480 12808 8492
rect 12207 8452 12808 8480
rect 12207 8449 12219 8452
rect 12161 8443 12219 8449
rect 12802 8440 12808 8452
rect 12860 8480 12866 8492
rect 12986 8480 12992 8492
rect 12860 8452 12992 8480
rect 12860 8440 12866 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13096 8480 13124 8520
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 15102 8508 15108 8560
rect 15160 8548 15166 8560
rect 15197 8551 15255 8557
rect 15197 8548 15209 8551
rect 15160 8520 15209 8548
rect 15160 8508 15166 8520
rect 15197 8517 15209 8520
rect 15243 8517 15255 8551
rect 16942 8548 16948 8560
rect 15197 8511 15255 8517
rect 15304 8520 15516 8548
rect 13170 8480 13176 8492
rect 13083 8452 13176 8480
rect 13170 8440 13176 8452
rect 13228 8480 13234 8492
rect 14844 8480 14872 8508
rect 15304 8480 15332 8520
rect 13228 8452 13584 8480
rect 14844 8452 15332 8480
rect 13228 8440 13234 8452
rect 1670 8372 1676 8424
rect 1728 8412 1734 8424
rect 1857 8415 1915 8421
rect 1857 8412 1869 8415
rect 1728 8384 1869 8412
rect 1728 8372 1734 8384
rect 1857 8381 1869 8384
rect 1903 8381 1915 8415
rect 1857 8375 1915 8381
rect 4525 8415 4583 8421
rect 4525 8381 4537 8415
rect 4571 8412 4583 8415
rect 5442 8412 5448 8424
rect 4571 8384 5448 8412
rect 4571 8381 4583 8384
rect 4525 8375 4583 8381
rect 5442 8372 5448 8384
rect 5500 8372 5506 8424
rect 6362 8372 6368 8424
rect 6420 8412 6426 8424
rect 8478 8412 8484 8424
rect 6420 8384 7144 8412
rect 8439 8384 8484 8412
rect 6420 8372 6426 8384
rect 2124 8347 2182 8353
rect 2124 8313 2136 8347
rect 2170 8344 2182 8347
rect 2682 8344 2688 8356
rect 2170 8316 2688 8344
rect 2170 8313 2182 8316
rect 2124 8307 2182 8313
rect 2682 8304 2688 8316
rect 2740 8304 2746 8356
rect 5074 8304 5080 8356
rect 5132 8304 5138 8356
rect 5629 8347 5687 8353
rect 5629 8313 5641 8347
rect 5675 8344 5687 8347
rect 6086 8344 6092 8356
rect 5675 8316 5764 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 3234 8276 3240 8288
rect 3195 8248 3240 8276
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 4617 8279 4675 8285
rect 4617 8245 4629 8279
rect 4663 8276 4675 8279
rect 5083 8276 5111 8304
rect 4663 8248 5111 8276
rect 5169 8279 5227 8285
rect 4663 8245 4675 8248
rect 4617 8239 4675 8245
rect 5169 8245 5181 8279
rect 5215 8276 5227 8279
rect 5442 8276 5448 8288
rect 5215 8248 5448 8276
rect 5215 8245 5227 8248
rect 5169 8239 5227 8245
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 5736 8276 5764 8316
rect 5920 8316 6092 8344
rect 5920 8276 5948 8316
rect 6086 8304 6092 8316
rect 6144 8344 6150 8356
rect 6546 8344 6552 8356
rect 6144 8316 6552 8344
rect 6144 8304 6150 8316
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7116 8344 7144 8384
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 10594 8412 10600 8424
rect 8588 8384 10600 8412
rect 7193 8347 7251 8353
rect 7193 8344 7205 8347
rect 7116 8316 7205 8344
rect 7193 8313 7205 8316
rect 7239 8313 7251 8347
rect 7193 8307 7251 8313
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 8588 8344 8616 8384
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 12618 8412 12624 8424
rect 10735 8384 12624 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 12618 8372 12624 8384
rect 12676 8412 12682 8424
rect 13449 8415 13507 8421
rect 12676 8384 13216 8412
rect 12676 8372 12682 8384
rect 13188 8356 13216 8384
rect 13449 8381 13461 8415
rect 13495 8381 13507 8415
rect 13556 8412 13584 8452
rect 13998 8412 14004 8424
rect 13556 8384 14004 8412
rect 13449 8375 13507 8381
rect 7616 8316 8616 8344
rect 8748 8347 8806 8353
rect 7616 8304 7622 8316
rect 8748 8313 8760 8347
rect 8794 8344 8806 8347
rect 9122 8344 9128 8356
rect 8794 8316 9128 8344
rect 8794 8313 8806 8316
rect 8748 8307 8806 8313
rect 9122 8304 9128 8316
rect 9180 8304 9186 8356
rect 9306 8304 9312 8356
rect 9364 8344 9370 8356
rect 10502 8344 10508 8356
rect 9364 8316 10508 8344
rect 9364 8304 9370 8316
rect 10502 8304 10508 8316
rect 10560 8304 10566 8356
rect 10956 8347 11014 8353
rect 10956 8313 10968 8347
rect 11002 8344 11014 8347
rect 12161 8347 12219 8353
rect 12161 8344 12173 8347
rect 11002 8316 12173 8344
rect 11002 8313 11014 8316
rect 10956 8307 11014 8313
rect 12161 8313 12173 8316
rect 12207 8313 12219 8347
rect 12161 8307 12219 8313
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12768 8316 12909 8344
rect 12768 8304 12774 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 12897 8307 12955 8313
rect 13170 8304 13176 8356
rect 13228 8344 13234 8356
rect 13464 8344 13492 8375
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 15488 8412 15516 8520
rect 15672 8520 16948 8548
rect 15672 8489 15700 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17034 8508 17040 8560
rect 17092 8548 17098 8560
rect 18506 8548 18512 8560
rect 17092 8520 18512 8548
rect 17092 8508 17098 8520
rect 18506 8508 18512 8520
rect 18564 8508 18570 8560
rect 15657 8483 15715 8489
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17678 8480 17684 8492
rect 17451 8452 17684 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 15764 8412 15792 8443
rect 17678 8440 17684 8452
rect 17736 8440 17742 8492
rect 19613 8483 19671 8489
rect 19613 8449 19625 8483
rect 19659 8480 19671 8483
rect 19794 8480 19800 8492
rect 19659 8452 19800 8480
rect 19659 8449 19671 8452
rect 19613 8443 19671 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 20530 8480 20536 8492
rect 20491 8452 20536 8480
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 15488 8384 15792 8412
rect 16114 8372 16120 8424
rect 16172 8412 16178 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 16172 8384 17141 8412
rect 16172 8372 16178 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17129 8375 17187 8381
rect 13228 8316 13492 8344
rect 13716 8347 13774 8353
rect 13228 8304 13234 8316
rect 13716 8313 13728 8347
rect 13762 8344 13774 8347
rect 13814 8344 13820 8356
rect 13762 8316 13820 8344
rect 13762 8313 13774 8316
rect 13716 8307 13774 8313
rect 13814 8304 13820 8316
rect 13872 8304 13878 8356
rect 15562 8344 15568 8356
rect 15523 8316 15568 8344
rect 15562 8304 15568 8316
rect 15620 8304 15626 8356
rect 17218 8344 17224 8356
rect 17179 8316 17224 8344
rect 17218 8304 17224 8316
rect 17276 8304 17282 8356
rect 18966 8344 18972 8356
rect 17328 8316 18972 8344
rect 6270 8276 6276 8288
rect 5592 8248 5637 8276
rect 5736 8248 5948 8276
rect 6231 8248 6276 8276
rect 5592 8236 5598 8248
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 6638 8236 6644 8288
rect 6696 8276 6702 8288
rect 11974 8276 11980 8288
rect 6696 8248 11980 8276
rect 6696 8236 6702 8248
rect 11974 8236 11980 8248
rect 12032 8236 12038 8288
rect 12250 8236 12256 8288
rect 12308 8276 12314 8288
rect 12437 8279 12495 8285
rect 12437 8276 12449 8279
rect 12308 8248 12449 8276
rect 12308 8236 12314 8248
rect 12437 8245 12449 8248
rect 12483 8245 12495 8279
rect 12437 8239 12495 8245
rect 12805 8279 12863 8285
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13538 8276 13544 8288
rect 12851 8248 13544 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13538 8236 13544 8248
rect 13596 8236 13602 8288
rect 16761 8279 16819 8285
rect 16761 8245 16773 8279
rect 16807 8276 16819 8279
rect 17328 8276 17356 8316
rect 18966 8304 18972 8316
rect 19024 8304 19030 8356
rect 19334 8344 19340 8356
rect 19295 8316 19340 8344
rect 19334 8304 19340 8316
rect 19392 8304 19398 8356
rect 20349 8347 20407 8353
rect 20349 8313 20361 8347
rect 20395 8344 20407 8347
rect 20898 8344 20904 8356
rect 20395 8316 20904 8344
rect 20395 8313 20407 8316
rect 20349 8307 20407 8313
rect 20898 8304 20904 8316
rect 20956 8304 20962 8356
rect 16807 8248 17356 8276
rect 16807 8245 16819 8248
rect 16761 8239 16819 8245
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 19978 8276 19984 8288
rect 19484 8248 19529 8276
rect 19939 8248 19984 8276
rect 19484 8236 19490 8248
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 20438 8276 20444 8288
rect 20399 8248 20444 8276
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 1104 8186 21620 8208
rect 1104 8134 7846 8186
rect 7898 8134 7910 8186
rect 7962 8134 7974 8186
rect 8026 8134 8038 8186
rect 8090 8134 14710 8186
rect 14762 8134 14774 8186
rect 14826 8134 14838 8186
rect 14890 8134 14902 8186
rect 14954 8134 21620 8186
rect 1104 8112 21620 8134
rect 1946 8072 1952 8084
rect 1907 8044 1952 8072
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2961 8075 3019 8081
rect 2961 8041 2973 8075
rect 3007 8072 3019 8075
rect 3970 8072 3976 8084
rect 3007 8044 3976 8072
rect 3007 8041 3019 8044
rect 2961 8035 3019 8041
rect 3970 8032 3976 8044
rect 4028 8032 4034 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4525 8075 4583 8081
rect 4525 8072 4537 8075
rect 4304 8044 4537 8072
rect 4304 8032 4310 8044
rect 4525 8041 4537 8044
rect 4571 8041 4583 8075
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 4525 8035 4583 8041
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6328 8044 6745 8072
rect 6328 8032 6334 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 7374 8072 7380 8084
rect 7335 8044 7380 8072
rect 6733 8035 6791 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8294 8072 8300 8084
rect 7616 8044 8300 8072
rect 7616 8032 7622 8044
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 8570 8032 8576 8084
rect 8628 8072 8634 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8628 8044 8953 8072
rect 8628 8032 8634 8044
rect 8941 8041 8953 8044
rect 8987 8041 8999 8075
rect 8941 8035 8999 8041
rect 9033 8075 9091 8081
rect 9033 8041 9045 8075
rect 9079 8072 9091 8075
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9079 8044 10149 8072
rect 9079 8041 9091 8044
rect 9033 8035 9091 8041
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10560 8044 10609 8072
rect 10560 8032 10566 8044
rect 10597 8041 10609 8044
rect 10643 8072 10655 8075
rect 12066 8072 12072 8084
rect 10643 8044 12072 8072
rect 10643 8041 10655 8044
rect 10597 8035 10655 8041
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13357 8075 13415 8081
rect 13357 8072 13369 8075
rect 13136 8044 13369 8072
rect 13136 8032 13142 8044
rect 13357 8041 13369 8044
rect 13403 8041 13415 8075
rect 13357 8035 13415 8041
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13504 8044 13860 8072
rect 13504 8032 13510 8044
rect 2317 8007 2375 8013
rect 2317 7973 2329 8007
rect 2363 8004 2375 8007
rect 3050 8004 3056 8016
rect 2363 7976 3056 8004
rect 2363 7973 2375 7976
rect 2317 7967 2375 7973
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 3418 8004 3424 8016
rect 3379 7976 3424 8004
rect 3418 7964 3424 7976
rect 3476 7964 3482 8016
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 7745 8007 7803 8013
rect 7745 8004 7757 8007
rect 3568 7976 7757 8004
rect 3568 7964 3574 7976
rect 7745 7973 7757 7976
rect 7791 7973 7803 8007
rect 7745 7967 7803 7973
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 10870 8004 10876 8016
rect 8904 7976 10876 8004
rect 8904 7964 8910 7976
rect 10870 7964 10876 7976
rect 10928 7964 10934 8016
rect 11977 8007 12035 8013
rect 11977 7973 11989 8007
rect 12023 8004 12035 8007
rect 12342 8004 12348 8016
rect 12023 7976 12348 8004
rect 12023 7973 12035 7976
rect 11977 7967 12035 7973
rect 12342 7964 12348 7976
rect 12400 8004 12406 8016
rect 12400 7976 12480 8004
rect 12400 7964 12406 7976
rect 3329 7939 3387 7945
rect 3329 7905 3341 7939
rect 3375 7936 3387 7939
rect 3970 7936 3976 7948
rect 3375 7908 3976 7936
rect 3375 7905 3387 7908
rect 3329 7899 3387 7905
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4433 7939 4491 7945
rect 4433 7936 4445 7939
rect 4212 7908 4445 7936
rect 4212 7896 4218 7908
rect 4433 7905 4445 7908
rect 4479 7936 4491 7939
rect 5074 7936 5080 7948
rect 4479 7908 5080 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 5074 7896 5080 7908
rect 5132 7896 5138 7948
rect 6638 7936 6644 7948
rect 5828 7908 6644 7936
rect 5828 7880 5856 7908
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 6730 7896 6736 7948
rect 6788 7936 6794 7948
rect 6788 7908 6960 7936
rect 6788 7896 6794 7908
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2682 7868 2688 7880
rect 2639 7840 2688 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2682 7828 2688 7840
rect 2740 7868 2746 7880
rect 3605 7871 3663 7877
rect 3605 7868 3617 7871
rect 2740 7840 3617 7868
rect 2740 7828 2746 7840
rect 3605 7837 3617 7840
rect 3651 7868 3663 7871
rect 3694 7868 3700 7880
rect 3651 7840 3700 7868
rect 3651 7837 3663 7840
rect 3605 7831 3663 7837
rect 3694 7828 3700 7840
rect 3752 7828 3758 7880
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4617 7871 4675 7877
rect 4617 7868 4629 7871
rect 3844 7840 4629 7868
rect 3844 7828 3850 7840
rect 4617 7837 4629 7840
rect 4663 7837 4675 7871
rect 4617 7831 4675 7837
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5534 7868 5540 7880
rect 5408 7840 5540 7868
rect 5408 7828 5414 7840
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 5810 7868 5816 7880
rect 5767 7840 5816 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7837 5963 7871
rect 5905 7831 5963 7837
rect 3234 7760 3240 7812
rect 3292 7800 3298 7812
rect 3292 7772 4200 7800
rect 3292 7760 3298 7772
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 4065 7735 4123 7741
rect 4065 7732 4077 7735
rect 3568 7704 4077 7732
rect 3568 7692 3574 7704
rect 4065 7701 4077 7704
rect 4111 7701 4123 7735
rect 4172 7732 4200 7772
rect 5166 7760 5172 7812
rect 5224 7800 5230 7812
rect 5920 7800 5948 7831
rect 6546 7828 6552 7880
rect 6604 7868 6610 7880
rect 6932 7877 6960 7908
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7837 7939 7895 7945
rect 7837 7936 7849 7939
rect 7156 7908 7849 7936
rect 7156 7896 7162 7908
rect 7837 7905 7849 7908
rect 7883 7905 7895 7939
rect 7837 7899 7895 7905
rect 9674 7896 9680 7948
rect 9732 7936 9738 7948
rect 10410 7936 10416 7948
rect 9732 7908 10416 7936
rect 9732 7896 9738 7908
rect 10410 7896 10416 7908
rect 10468 7936 10474 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10468 7908 10517 7936
rect 10468 7896 10474 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 11146 7896 11152 7948
rect 11204 7936 11210 7948
rect 11606 7936 11612 7948
rect 11204 7908 11612 7936
rect 11204 7896 11210 7908
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 11885 7939 11943 7945
rect 11885 7905 11897 7939
rect 11931 7936 11943 7939
rect 12452 7936 12480 7976
rect 12526 7964 12532 8016
rect 12584 8004 12590 8016
rect 13725 8007 13783 8013
rect 13725 8004 13737 8007
rect 12584 7976 13737 8004
rect 12584 7964 12590 7976
rect 13725 7973 13737 7976
rect 13771 7973 13783 8007
rect 13832 8004 13860 8044
rect 13906 8032 13912 8084
rect 13964 8072 13970 8084
rect 14185 8075 14243 8081
rect 14185 8072 14197 8075
rect 13964 8044 14197 8072
rect 13964 8032 13970 8044
rect 14185 8041 14197 8044
rect 14231 8041 14243 8075
rect 14550 8072 14556 8084
rect 14511 8044 14556 8072
rect 14185 8035 14243 8041
rect 14550 8032 14556 8044
rect 14608 8032 14614 8084
rect 19058 8072 19064 8084
rect 19019 8044 19064 8072
rect 19058 8032 19064 8044
rect 19116 8032 19122 8084
rect 19705 8075 19763 8081
rect 19705 8041 19717 8075
rect 19751 8072 19763 8075
rect 20438 8072 20444 8084
rect 19751 8044 20444 8072
rect 19751 8041 19763 8044
rect 19705 8035 19763 8041
rect 20438 8032 20444 8044
rect 20496 8032 20502 8084
rect 20898 8072 20904 8084
rect 20859 8044 20904 8072
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 14090 8004 14096 8016
rect 13832 7976 14096 8004
rect 13725 7967 13783 7973
rect 14090 7964 14096 7976
rect 14148 7964 14154 8016
rect 16022 8013 16028 8016
rect 16016 8004 16028 8013
rect 15983 7976 16028 8004
rect 16016 7967 16028 7976
rect 16022 7964 16028 7967
rect 16080 7964 16086 8016
rect 17678 7964 17684 8016
rect 17736 8004 17742 8016
rect 17948 8007 18006 8013
rect 17948 8004 17960 8007
rect 17736 7976 17960 8004
rect 17736 7964 17742 7976
rect 17948 7973 17960 7976
rect 17994 8004 18006 8007
rect 20530 8004 20536 8016
rect 17994 7976 20536 8004
rect 17994 7973 18006 7976
rect 17948 7967 18006 7973
rect 20530 7964 20536 7976
rect 20588 7964 20594 8016
rect 12802 7936 12808 7948
rect 11931 7908 12204 7936
rect 12452 7908 12808 7936
rect 11931 7905 11943 7908
rect 11885 7899 11943 7905
rect 12176 7880 12204 7908
rect 12802 7896 12808 7908
rect 12860 7896 12866 7948
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13538 7936 13544 7948
rect 12943 7908 13544 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 13964 7908 14780 7936
rect 13964 7896 13970 7908
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6604 7840 6837 7868
rect 6604 7828 6610 7840
rect 6825 7837 6837 7840
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 9122 7868 9128 7880
rect 9083 7840 9128 7868
rect 7929 7831 7987 7837
rect 6362 7800 6368 7812
rect 5224 7772 5948 7800
rect 6323 7772 6368 7800
rect 5224 7760 5230 7772
rect 6362 7760 6368 7772
rect 6420 7760 6426 7812
rect 7944 7732 7972 7831
rect 9122 7828 9128 7840
rect 9180 7828 9186 7880
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7837 10747 7871
rect 10689 7831 10747 7837
rect 8573 7803 8631 7809
rect 8573 7769 8585 7803
rect 8619 7800 8631 7803
rect 10042 7800 10048 7812
rect 8619 7772 10048 7800
rect 8619 7769 8631 7772
rect 8573 7763 8631 7769
rect 10042 7760 10048 7772
rect 10100 7760 10106 7812
rect 4172 7704 7972 7732
rect 4065 7695 4123 7701
rect 9030 7692 9036 7744
rect 9088 7732 9094 7744
rect 10704 7732 10732 7831
rect 11790 7828 11796 7880
rect 11848 7868 11854 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11848 7840 12081 7868
rect 11848 7828 11854 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 12158 7828 12164 7880
rect 12216 7828 12222 7880
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12768 7840 13001 7868
rect 12768 7828 12774 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 13078 7828 13084 7880
rect 13136 7868 13142 7880
rect 13817 7871 13875 7877
rect 13136 7840 13181 7868
rect 13136 7828 13142 7840
rect 13817 7837 13829 7871
rect 13863 7837 13875 7871
rect 13998 7868 14004 7880
rect 13959 7840 14004 7868
rect 13817 7831 13875 7837
rect 12529 7803 12587 7809
rect 12529 7769 12541 7803
rect 12575 7800 12587 7803
rect 13832 7800 13860 7831
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 14752 7877 14780 7908
rect 15194 7896 15200 7948
rect 15252 7936 15258 7948
rect 15657 7939 15715 7945
rect 15657 7936 15669 7939
rect 15252 7908 15669 7936
rect 15252 7896 15258 7908
rect 15657 7905 15669 7908
rect 15703 7905 15715 7939
rect 15657 7899 15715 7905
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 19610 7936 19616 7948
rect 16356 7908 19616 7936
rect 16356 7896 16362 7908
rect 19610 7896 19616 7908
rect 19668 7896 19674 7948
rect 20073 7939 20131 7945
rect 20073 7905 20085 7939
rect 20119 7936 20131 7939
rect 20714 7936 20720 7948
rect 20119 7908 20720 7936
rect 20119 7905 20131 7908
rect 20073 7899 20131 7905
rect 14645 7871 14703 7877
rect 14645 7868 14657 7871
rect 14148 7840 14657 7868
rect 14148 7828 14154 7840
rect 14645 7837 14657 7840
rect 14691 7837 14703 7871
rect 14645 7831 14703 7837
rect 14737 7871 14795 7877
rect 14737 7837 14749 7871
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 15746 7868 15752 7880
rect 15344 7840 15752 7868
rect 15344 7828 15350 7840
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 17586 7828 17592 7880
rect 17644 7868 17650 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 17644 7840 17693 7868
rect 17644 7828 17650 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 20088 7868 20116 7899
rect 20714 7896 20720 7908
rect 20772 7896 20778 7948
rect 19208 7840 20116 7868
rect 19208 7828 19214 7840
rect 20162 7828 20168 7880
rect 20220 7868 20226 7880
rect 20349 7871 20407 7877
rect 20220 7840 20265 7868
rect 20220 7828 20226 7840
rect 20349 7837 20361 7871
rect 20395 7837 20407 7871
rect 20349 7831 20407 7837
rect 12575 7772 13860 7800
rect 12575 7769 12587 7772
rect 12529 7763 12587 7769
rect 9088 7704 10732 7732
rect 11517 7735 11575 7741
rect 9088 7692 9094 7704
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 12802 7732 12808 7744
rect 11563 7704 12808 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 12802 7692 12808 7704
rect 12860 7692 12866 7744
rect 15473 7735 15531 7741
rect 15473 7701 15485 7735
rect 15519 7732 15531 7735
rect 15746 7732 15752 7744
rect 15519 7704 15752 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 15746 7692 15752 7704
rect 15804 7692 15810 7744
rect 17126 7732 17132 7744
rect 17087 7704 17132 7732
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17862 7692 17868 7744
rect 17920 7732 17926 7744
rect 20364 7732 20392 7831
rect 20438 7732 20444 7744
rect 17920 7704 20444 7732
rect 17920 7692 17926 7704
rect 20438 7692 20444 7704
rect 20496 7692 20502 7744
rect 1104 7642 21620 7664
rect 1104 7590 4414 7642
rect 4466 7590 4478 7642
rect 4530 7590 4542 7642
rect 4594 7590 4606 7642
rect 4658 7590 11278 7642
rect 11330 7590 11342 7642
rect 11394 7590 11406 7642
rect 11458 7590 11470 7642
rect 11522 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 18270 7642
rect 18322 7590 18334 7642
rect 18386 7590 21620 7642
rect 1104 7568 21620 7590
rect 2130 7528 2136 7540
rect 2091 7500 2136 7528
rect 2130 7488 2136 7500
rect 2188 7488 2194 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 4154 7528 4160 7540
rect 3108 7500 4160 7528
rect 3108 7488 3114 7500
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5718 7528 5724 7540
rect 4939 7500 5724 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 8846 7528 8852 7540
rect 6696 7500 8852 7528
rect 6696 7488 6702 7500
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9180 7500 9873 7528
rect 9180 7488 9186 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 10134 7528 10140 7540
rect 10095 7500 10140 7528
rect 9861 7491 9919 7497
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 3786 7460 3792 7472
rect 3660 7432 3792 7460
rect 3660 7420 3666 7432
rect 3786 7420 3792 7432
rect 3844 7420 3850 7472
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7429 7987 7463
rect 7929 7423 7987 7429
rect 2774 7352 2780 7404
rect 2832 7392 2838 7404
rect 2832 7364 2877 7392
rect 2832 7352 2838 7364
rect 3050 7352 3056 7404
rect 3108 7392 3114 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3108 7364 3709 7392
rect 3108 7352 3114 7364
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4028 7364 5304 7392
rect 4028 7352 4034 7364
rect 3510 7324 3516 7336
rect 3471 7296 3516 7324
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 5276 7324 5304 7364
rect 5350 7352 5356 7404
rect 5408 7392 5414 7404
rect 5445 7395 5503 7401
rect 5445 7392 5457 7395
rect 5408 7364 5457 7392
rect 5408 7352 5414 7364
rect 5445 7361 5457 7364
rect 5491 7361 5503 7395
rect 5445 7355 5503 7361
rect 5626 7352 5632 7404
rect 5684 7392 5690 7404
rect 7006 7392 7012 7404
rect 5684 7364 7012 7392
rect 5684 7352 5690 7364
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 7098 7352 7104 7404
rect 7156 7392 7162 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7156 7364 7481 7392
rect 7156 7352 7162 7364
rect 7469 7361 7481 7364
rect 7515 7361 7527 7395
rect 7944 7392 7972 7423
rect 8018 7392 8024 7404
rect 7944 7364 8024 7392
rect 7469 7355 7527 7361
rect 8018 7352 8024 7364
rect 8076 7352 8082 7404
rect 9876 7392 9904 7491
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 14274 7488 14280 7540
rect 14332 7528 14338 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14332 7500 15025 7528
rect 14332 7488 14338 7500
rect 15013 7497 15025 7500
rect 15059 7528 15071 7531
rect 15197 7531 15255 7537
rect 15197 7528 15209 7531
rect 15059 7500 15209 7528
rect 15059 7497 15071 7500
rect 15013 7491 15071 7497
rect 15197 7497 15209 7500
rect 15243 7497 15255 7531
rect 17678 7528 17684 7540
rect 17639 7500 17684 7528
rect 15197 7491 15255 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18693 7531 18751 7537
rect 18693 7497 18705 7531
rect 18739 7528 18751 7531
rect 19426 7528 19432 7540
rect 18739 7500 19432 7528
rect 18739 7497 18751 7500
rect 18693 7491 18751 7497
rect 19426 7488 19432 7500
rect 19484 7488 19490 7540
rect 19794 7488 19800 7540
rect 19852 7528 19858 7540
rect 20162 7528 20168 7540
rect 19852 7500 20168 7528
rect 19852 7488 19858 7500
rect 20162 7488 20168 7500
rect 20220 7528 20226 7540
rect 20346 7528 20352 7540
rect 20220 7500 20352 7528
rect 20220 7488 20226 7500
rect 20346 7488 20352 7500
rect 20404 7488 20410 7540
rect 14642 7420 14648 7472
rect 14700 7460 14706 7472
rect 14700 7432 16344 7460
rect 14700 7420 14706 7432
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 9876 7364 10701 7392
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11701 7395 11759 7401
rect 11701 7392 11713 7395
rect 11204 7364 11713 7392
rect 11204 7352 11210 7364
rect 11701 7361 11713 7364
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 12618 7352 12624 7404
rect 12676 7392 12682 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12676 7364 13001 7392
rect 12676 7352 12682 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 15243 7364 15853 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 16316 7392 16344 7432
rect 16316 7364 16436 7392
rect 15841 7355 15899 7361
rect 8113 7327 8171 7333
rect 5276 7296 8064 7324
rect 1946 7216 1952 7268
rect 2004 7256 2010 7268
rect 2501 7259 2559 7265
rect 2501 7256 2513 7259
rect 2004 7228 2513 7256
rect 2004 7216 2010 7228
rect 2501 7225 2513 7228
rect 2547 7225 2559 7259
rect 2501 7219 2559 7225
rect 3786 7216 3792 7268
rect 3844 7256 3850 7268
rect 7377 7259 7435 7265
rect 7377 7256 7389 7259
rect 3844 7228 7389 7256
rect 3844 7216 3850 7228
rect 7377 7225 7389 7228
rect 7423 7225 7435 7259
rect 8036 7256 8064 7296
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 8202 7324 8208 7336
rect 8159 7296 8208 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 8478 7324 8484 7336
rect 8439 7296 8484 7324
rect 8478 7284 8484 7296
rect 8536 7284 8542 7336
rect 8748 7327 8806 7333
rect 8748 7293 8760 7327
rect 8794 7324 8806 7327
rect 9030 7324 9036 7336
rect 8794 7296 9036 7324
rect 8794 7293 8806 7296
rect 8748 7287 8806 7293
rect 9030 7284 9036 7296
rect 9088 7284 9094 7336
rect 9306 7284 9312 7336
rect 9364 7324 9370 7336
rect 10226 7324 10232 7336
rect 9364 7296 10232 7324
rect 9364 7284 9370 7296
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 12434 7284 12440 7336
rect 12492 7284 12498 7336
rect 12802 7324 12808 7336
rect 12763 7296 12808 7324
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13170 7324 13176 7336
rect 12952 7296 13176 7324
rect 12952 7284 12958 7296
rect 13170 7284 13176 7296
rect 13228 7324 13234 7336
rect 13633 7327 13691 7333
rect 13633 7324 13645 7327
rect 13228 7296 13645 7324
rect 13228 7284 13234 7296
rect 13633 7293 13645 7296
rect 13679 7293 13691 7327
rect 13633 7287 13691 7293
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7293 16359 7327
rect 16408 7324 16436 7364
rect 19058 7352 19064 7404
rect 19116 7392 19122 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 19116 7364 19257 7392
rect 19116 7352 19122 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7392 20407 7395
rect 20530 7392 20536 7404
rect 20395 7364 20536 7392
rect 20395 7361 20407 7364
rect 20349 7355 20407 7361
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 18141 7327 18199 7333
rect 16408 7296 18092 7324
rect 16301 7287 16359 7293
rect 8036 7228 8248 7256
rect 7377 7219 7435 7225
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 3145 7191 3203 7197
rect 3145 7188 3157 7191
rect 2639 7160 3157 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 3145 7157 3157 7160
rect 3191 7157 3203 7191
rect 3145 7151 3203 7157
rect 3605 7191 3663 7197
rect 3605 7157 3617 7191
rect 3651 7188 3663 7191
rect 4798 7188 4804 7200
rect 3651 7160 4804 7188
rect 3651 7157 3663 7160
rect 3605 7151 3663 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5353 7191 5411 7197
rect 5353 7157 5365 7191
rect 5399 7188 5411 7191
rect 6638 7188 6644 7200
rect 5399 7160 6644 7188
rect 5399 7157 5411 7160
rect 5353 7151 5411 7157
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 6914 7188 6920 7200
rect 6875 7160 6920 7188
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7282 7188 7288 7200
rect 7243 7160 7288 7188
rect 7282 7148 7288 7160
rect 7340 7148 7346 7200
rect 8220 7188 8248 7228
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 11054 7256 11060 7268
rect 8352 7228 11060 7256
rect 8352 7216 8358 7228
rect 11054 7216 11060 7228
rect 11112 7216 11118 7268
rect 11609 7259 11667 7265
rect 11609 7225 11621 7259
rect 11655 7256 11667 7259
rect 12452 7256 12480 7284
rect 12710 7256 12716 7268
rect 11655 7228 12716 7256
rect 11655 7225 11667 7228
rect 11609 7219 11667 7225
rect 12710 7216 12716 7228
rect 12768 7216 12774 7268
rect 13906 7265 13912 7268
rect 13900 7256 13912 7265
rect 13867 7228 13912 7256
rect 13900 7219 13912 7228
rect 13906 7216 13912 7219
rect 13964 7216 13970 7268
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14826 7256 14832 7268
rect 14056 7228 14832 7256
rect 14056 7216 14062 7228
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 15194 7216 15200 7268
rect 15252 7256 15258 7268
rect 15749 7259 15807 7265
rect 15749 7256 15761 7259
rect 15252 7228 15761 7256
rect 15252 7216 15258 7228
rect 15749 7225 15761 7228
rect 15795 7225 15807 7259
rect 15749 7219 15807 7225
rect 15838 7216 15844 7268
rect 15896 7256 15902 7268
rect 16316 7256 16344 7287
rect 15896 7228 16344 7256
rect 15896 7216 15902 7228
rect 9950 7188 9956 7200
rect 8220 7160 9956 7188
rect 9950 7148 9956 7160
rect 10008 7148 10014 7200
rect 10502 7188 10508 7200
rect 10463 7160 10508 7188
rect 10502 7148 10508 7160
rect 10560 7148 10566 7200
rect 10597 7191 10655 7197
rect 10597 7157 10609 7191
rect 10643 7188 10655 7191
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 10643 7160 11161 7188
rect 10643 7157 10655 7160
rect 10597 7151 10655 7157
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11149 7151 11207 7157
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 11698 7188 11704 7200
rect 11563 7160 11704 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 11698 7148 11704 7160
rect 11756 7148 11762 7200
rect 12437 7191 12495 7197
rect 12437 7157 12449 7191
rect 12483 7188 12495 7191
rect 12526 7188 12532 7200
rect 12483 7160 12532 7188
rect 12483 7157 12495 7160
rect 12437 7151 12495 7157
rect 12526 7148 12532 7160
rect 12584 7148 12590 7200
rect 12802 7148 12808 7200
rect 12860 7188 12866 7200
rect 12897 7191 12955 7197
rect 12897 7188 12909 7191
rect 12860 7160 12909 7188
rect 12860 7148 12866 7160
rect 12897 7157 12909 7160
rect 12943 7157 12955 7191
rect 12897 7151 12955 7157
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 15160 7160 15301 7188
rect 15160 7148 15166 7160
rect 15289 7157 15301 7160
rect 15335 7157 15347 7191
rect 15654 7188 15660 7200
rect 15615 7160 15660 7188
rect 15289 7151 15347 7157
rect 15654 7148 15660 7160
rect 15712 7148 15718 7200
rect 16316 7188 16344 7228
rect 16568 7259 16626 7265
rect 16568 7225 16580 7259
rect 16614 7256 16626 7259
rect 16666 7256 16672 7268
rect 16614 7228 16672 7256
rect 16614 7225 16626 7228
rect 16568 7219 16626 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 18064 7256 18092 7296
rect 18141 7293 18153 7327
rect 18187 7324 18199 7327
rect 19426 7324 19432 7336
rect 18187 7296 19432 7324
rect 18187 7293 18199 7296
rect 18141 7287 18199 7293
rect 19426 7284 19432 7296
rect 19484 7284 19490 7336
rect 20714 7324 20720 7336
rect 20675 7296 20720 7324
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 18782 7256 18788 7268
rect 18064 7228 18788 7256
rect 18782 7216 18788 7228
rect 18840 7216 18846 7268
rect 19061 7259 19119 7265
rect 19061 7225 19073 7259
rect 19107 7256 19119 7259
rect 19518 7256 19524 7268
rect 19107 7228 19524 7256
rect 19107 7225 19119 7228
rect 19061 7219 19119 7225
rect 19518 7216 19524 7228
rect 19576 7216 19582 7268
rect 17586 7188 17592 7200
rect 16316 7160 17592 7188
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 19153 7191 19211 7197
rect 19153 7157 19165 7191
rect 19199 7188 19211 7191
rect 19705 7191 19763 7197
rect 19705 7188 19717 7191
rect 19199 7160 19717 7188
rect 19199 7157 19211 7160
rect 19153 7151 19211 7157
rect 19705 7157 19717 7160
rect 19751 7157 19763 7191
rect 20070 7188 20076 7200
rect 20031 7160 20076 7188
rect 19705 7151 19763 7157
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20162 7148 20168 7200
rect 20220 7188 20226 7200
rect 20901 7191 20959 7197
rect 20220 7160 20265 7188
rect 20220 7148 20226 7160
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 21082 7188 21088 7200
rect 20947 7160 21088 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 21082 7148 21088 7160
rect 21140 7148 21146 7200
rect 1104 7098 21620 7120
rect 1104 7046 7846 7098
rect 7898 7046 7910 7098
rect 7962 7046 7974 7098
rect 8026 7046 8038 7098
rect 8090 7046 14710 7098
rect 14762 7046 14774 7098
rect 14826 7046 14838 7098
rect 14890 7046 14902 7098
rect 14954 7046 21620 7098
rect 1104 7024 21620 7046
rect 3050 6984 3056 6996
rect 3011 6956 3056 6984
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 6972 6956 7573 6984
rect 6972 6944 6978 6956
rect 7561 6953 7573 6956
rect 7607 6953 7619 6987
rect 7561 6947 7619 6953
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 10502 6984 10508 6996
rect 9907 6956 10508 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 11256 6956 11928 6984
rect 2406 6876 2412 6928
rect 2464 6916 2470 6928
rect 5350 6916 5356 6928
rect 2464 6888 5356 6916
rect 2464 6876 2470 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 6362 6876 6368 6928
rect 6420 6916 6426 6928
rect 8573 6919 8631 6925
rect 8573 6916 8585 6919
rect 6420 6888 8585 6916
rect 6420 6876 6426 6888
rect 8573 6885 8585 6888
rect 8619 6885 8631 6919
rect 8573 6879 8631 6885
rect 9030 6876 9036 6928
rect 9088 6916 9094 6928
rect 9088 6888 10180 6916
rect 9088 6876 9094 6888
rect 1670 6848 1676 6860
rect 1631 6820 1676 6848
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 1940 6851 1998 6857
rect 1940 6817 1952 6851
rect 1986 6848 1998 6851
rect 2222 6848 2228 6860
rect 1986 6820 2228 6848
rect 1986 6817 1998 6820
rect 1940 6811 1998 6817
rect 2222 6808 2228 6820
rect 2280 6808 2286 6860
rect 4976 6851 5034 6857
rect 4976 6817 4988 6851
rect 5022 6848 5034 6851
rect 5994 6848 6000 6860
rect 5022 6820 6000 6848
rect 5022 6817 5034 6820
rect 4976 6811 5034 6817
rect 5994 6808 6000 6820
rect 6052 6808 6058 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 6328 6820 8677 6848
rect 6328 6808 6334 6820
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 10152 6848 10180 6888
rect 10226 6876 10232 6928
rect 10284 6916 10290 6928
rect 11256 6916 11284 6956
rect 10284 6888 11284 6916
rect 11900 6916 11928 6956
rect 12250 6944 12256 6996
rect 12308 6984 12314 6996
rect 16577 6987 16635 6993
rect 16577 6984 16589 6987
rect 12308 6956 16589 6984
rect 12308 6944 12314 6956
rect 16577 6953 16589 6956
rect 16623 6953 16635 6987
rect 16577 6947 16635 6953
rect 17402 6944 17408 6996
rect 17460 6984 17466 6996
rect 19889 6987 19947 6993
rect 19889 6984 19901 6987
rect 17460 6956 19901 6984
rect 17460 6944 17466 6956
rect 19889 6953 19901 6956
rect 19935 6953 19947 6987
rect 19889 6947 19947 6953
rect 13541 6919 13599 6925
rect 13541 6916 13553 6919
rect 11900 6888 13553 6916
rect 10284 6876 10290 6888
rect 13541 6885 13553 6888
rect 13587 6885 13599 6919
rect 13541 6879 13599 6885
rect 13814 6876 13820 6928
rect 13872 6876 13878 6928
rect 14553 6919 14611 6925
rect 14553 6885 14565 6919
rect 14599 6916 14611 6919
rect 14599 6888 15332 6916
rect 14599 6885 14611 6888
rect 14553 6879 14611 6885
rect 11146 6848 11152 6860
rect 10152 6820 11152 6848
rect 8665 6811 8723 6817
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4709 6783 4767 6789
rect 4709 6780 4721 6783
rect 4212 6752 4721 6780
rect 4212 6740 4218 6752
rect 4709 6749 4721 6752
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7190 6780 7196 6792
rect 6972 6752 7196 6780
rect 6972 6740 6978 6752
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 7650 6780 7656 6792
rect 7611 6752 7656 6780
rect 7650 6740 7656 6752
rect 7708 6740 7714 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8294 6780 8300 6792
rect 7883 6752 8300 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8294 6740 8300 6752
rect 8352 6740 8358 6792
rect 10428 6789 10456 6820
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11324 6851 11382 6857
rect 11324 6817 11336 6851
rect 11370 6848 11382 6851
rect 11790 6848 11796 6860
rect 11370 6820 11796 6848
rect 11370 6817 11382 6820
rect 11324 6811 11382 6817
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 12897 6851 12955 6857
rect 12897 6817 12909 6851
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 12989 6851 13047 6857
rect 12989 6817 13001 6851
rect 13035 6848 13047 6851
rect 13832 6848 13860 6876
rect 13035 6820 13860 6848
rect 13035 6817 13047 6820
rect 12989 6811 13047 6817
rect 8849 6783 8907 6789
rect 8849 6749 8861 6783
rect 8895 6780 8907 6783
rect 10321 6783 10379 6789
rect 8895 6752 10272 6780
rect 8895 6749 8907 6752
rect 8849 6743 8907 6749
rect 7006 6672 7012 6724
rect 7064 6712 7070 6724
rect 10134 6712 10140 6724
rect 7064 6684 10140 6712
rect 7064 6672 7070 6684
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 5442 6604 5448 6656
rect 5500 6644 5506 6656
rect 6089 6647 6147 6653
rect 6089 6644 6101 6647
rect 5500 6616 6101 6644
rect 5500 6604 5506 6616
rect 6089 6613 6101 6616
rect 6135 6613 6147 6647
rect 7190 6644 7196 6656
rect 7151 6616 7196 6644
rect 6089 6607 6147 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 8205 6647 8263 6653
rect 8205 6613 8217 6647
rect 8251 6644 8263 6647
rect 9766 6644 9772 6656
rect 8251 6616 9772 6644
rect 8251 6613 8263 6616
rect 8205 6607 8263 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10244 6644 10272 6752
rect 10321 6749 10333 6783
rect 10367 6749 10379 6783
rect 10321 6743 10379 6749
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 11054 6780 11060 6792
rect 11015 6752 11060 6780
rect 10413 6743 10471 6749
rect 10336 6712 10364 6743
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 12912 6780 12940 6811
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 15304 6857 15332 6888
rect 15470 6876 15476 6928
rect 15528 6916 15534 6928
rect 17497 6919 17555 6925
rect 17497 6916 17509 6919
rect 15528 6888 17509 6916
rect 15528 6876 15534 6888
rect 17497 6885 17509 6888
rect 17543 6885 17555 6919
rect 17497 6879 17555 6885
rect 18877 6919 18935 6925
rect 18877 6885 18889 6919
rect 18923 6916 18935 6919
rect 19978 6916 19984 6928
rect 18923 6888 19984 6916
rect 18923 6885 18935 6888
rect 18877 6879 18935 6885
rect 19978 6876 19984 6888
rect 20036 6876 20042 6928
rect 15289 6851 15347 6857
rect 14700 6820 14745 6848
rect 14700 6808 14706 6820
rect 15289 6817 15301 6851
rect 15335 6817 15347 6851
rect 15289 6811 15347 6817
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16025 6851 16083 6857
rect 16025 6848 16037 6851
rect 15804 6820 16037 6848
rect 15804 6808 15810 6820
rect 16025 6817 16037 6820
rect 16071 6817 16083 6851
rect 16025 6811 16083 6817
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 16485 6851 16543 6857
rect 16485 6848 16497 6851
rect 16448 6820 16497 6848
rect 16448 6808 16454 6820
rect 16485 6817 16497 6820
rect 16531 6817 16543 6851
rect 18966 6848 18972 6860
rect 18927 6820 18972 6848
rect 16485 6811 16543 6817
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 13630 6780 13636 6792
rect 12912 6752 13124 6780
rect 13591 6752 13636 6780
rect 10502 6712 10508 6724
rect 10336 6684 10508 6712
rect 10502 6672 10508 6684
rect 10560 6672 10566 6724
rect 12989 6715 13047 6721
rect 12989 6712 13001 6715
rect 11992 6684 13001 6712
rect 11992 6644 12020 6684
rect 12989 6681 13001 6684
rect 13035 6681 13047 6715
rect 12989 6675 13047 6681
rect 10244 6616 12020 6644
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12618 6644 12624 6656
rect 12483 6616 12624 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12618 6604 12624 6616
rect 12676 6604 12682 6656
rect 12713 6647 12771 6653
rect 12713 6613 12725 6647
rect 12759 6644 12771 6647
rect 12894 6644 12900 6656
rect 12759 6616 12900 6644
rect 12759 6613 12771 6616
rect 12713 6607 12771 6613
rect 12894 6604 12900 6616
rect 12952 6604 12958 6656
rect 13096 6644 13124 6752
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6780 13875 6783
rect 13906 6780 13912 6792
rect 13863 6752 13912 6780
rect 13863 6749 13875 6752
rect 13817 6743 13875 6749
rect 13906 6740 13912 6752
rect 13964 6780 13970 6792
rect 14550 6780 14556 6792
rect 13964 6752 14556 6780
rect 13964 6740 13970 6752
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14734 6780 14740 6792
rect 14695 6752 14740 6780
rect 14734 6740 14740 6752
rect 14792 6740 14798 6792
rect 16666 6780 16672 6792
rect 16579 6752 16672 6780
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16942 6740 16948 6792
rect 17000 6780 17006 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17000 6752 17601 6780
rect 17000 6740 17006 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6780 17831 6783
rect 17862 6780 17868 6792
rect 17819 6752 17868 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 13173 6715 13231 6721
rect 13173 6681 13185 6715
rect 13219 6712 13231 6715
rect 13998 6712 14004 6724
rect 13219 6684 14004 6712
rect 13219 6681 13231 6684
rect 13173 6675 13231 6681
rect 13998 6672 14004 6684
rect 14056 6672 14062 6724
rect 14185 6715 14243 6721
rect 14185 6681 14197 6715
rect 14231 6712 14243 6715
rect 15654 6712 15660 6724
rect 14231 6684 15660 6712
rect 14231 6681 14243 6684
rect 14185 6675 14243 6681
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 15838 6712 15844 6724
rect 15799 6684 15844 6712
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 16114 6712 16120 6724
rect 16075 6684 16120 6712
rect 16114 6672 16120 6684
rect 16172 6672 16178 6724
rect 15746 6644 15752 6656
rect 13096 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16684 6644 16712 6740
rect 17129 6715 17187 6721
rect 17129 6681 17141 6715
rect 17175 6712 17187 6715
rect 17218 6712 17224 6724
rect 17175 6684 17224 6712
rect 17175 6681 17187 6684
rect 17129 6675 17187 6681
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17678 6644 17684 6656
rect 16684 6616 17684 6644
rect 17678 6604 17684 6616
rect 17736 6644 17742 6656
rect 17788 6644 17816 6743
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19978 6780 19984 6792
rect 19116 6752 19161 6780
rect 19939 6752 19984 6780
rect 19116 6740 19122 6752
rect 19978 6740 19984 6752
rect 20036 6740 20042 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6780 20223 6783
rect 20530 6780 20536 6792
rect 20211 6752 20536 6780
rect 20211 6749 20223 6752
rect 20165 6743 20223 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 18509 6715 18567 6721
rect 18509 6681 18521 6715
rect 18555 6712 18567 6715
rect 19334 6712 19340 6724
rect 18555 6684 19340 6712
rect 18555 6681 18567 6684
rect 18509 6675 18567 6681
rect 19334 6672 19340 6684
rect 19392 6672 19398 6724
rect 19518 6712 19524 6724
rect 19479 6684 19524 6712
rect 19518 6672 19524 6684
rect 19576 6672 19582 6724
rect 17736 6616 17816 6644
rect 17736 6604 17742 6616
rect 1104 6554 21620 6576
rect 1104 6502 4414 6554
rect 4466 6502 4478 6554
rect 4530 6502 4542 6554
rect 4594 6502 4606 6554
rect 4658 6502 11278 6554
rect 11330 6502 11342 6554
rect 11394 6502 11406 6554
rect 11458 6502 11470 6554
rect 11522 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 18270 6554
rect 18322 6502 18334 6554
rect 18386 6502 21620 6554
rect 1104 6480 21620 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3513 6443 3571 6449
rect 3513 6440 3525 6443
rect 2832 6412 3525 6440
rect 2832 6400 2838 6412
rect 3513 6409 3525 6412
rect 3559 6440 3571 6443
rect 4062 6440 4068 6452
rect 3559 6412 4068 6440
rect 3559 6409 3571 6412
rect 3513 6403 3571 6409
rect 4062 6400 4068 6412
rect 4120 6400 4126 6452
rect 4798 6400 4804 6452
rect 4856 6440 4862 6452
rect 4893 6443 4951 6449
rect 4893 6440 4905 6443
rect 4856 6412 4905 6440
rect 4856 6400 4862 6412
rect 4893 6409 4905 6412
rect 4939 6409 4951 6443
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 4893 6403 4951 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 8846 6440 8852 6452
rect 7248 6412 8852 6440
rect 7248 6400 7254 6412
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 12342 6440 12348 6452
rect 11940 6412 12348 6440
rect 11940 6400 11946 6412
rect 12342 6400 12348 6412
rect 12400 6400 12406 6452
rect 12618 6400 12624 6452
rect 12676 6440 12682 6452
rect 16390 6440 16396 6452
rect 12676 6412 16396 6440
rect 12676 6400 12682 6412
rect 16390 6400 16396 6412
rect 16448 6400 16454 6452
rect 17589 6443 17647 6449
rect 17589 6409 17601 6443
rect 17635 6440 17647 6443
rect 18690 6440 18696 6452
rect 17635 6412 18696 6440
rect 17635 6409 17647 6412
rect 17589 6403 17647 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 20162 6400 20168 6452
rect 20220 6440 20226 6452
rect 20257 6443 20315 6449
rect 20257 6440 20269 6443
rect 20220 6412 20269 6440
rect 20220 6400 20226 6412
rect 20257 6409 20269 6412
rect 20303 6409 20315 6443
rect 20257 6403 20315 6409
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 5905 6375 5963 6381
rect 5905 6372 5917 6375
rect 4212 6344 5917 6372
rect 4212 6332 4218 6344
rect 5905 6341 5917 6344
rect 5951 6341 5963 6375
rect 5905 6335 5963 6341
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 11146 6372 11152 6384
rect 6788 6344 7512 6372
rect 11107 6344 11152 6372
rect 6788 6332 6794 6344
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 2130 6304 2136 6316
rect 1728 6276 2136 6304
rect 1728 6264 1734 6276
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 3602 6236 3608 6248
rect 2280 6208 3608 6236
rect 2280 6196 2286 6208
rect 3602 6196 3608 6208
rect 3660 6236 3666 6248
rect 4356 6236 4384 6267
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5353 6307 5411 6313
rect 5353 6304 5365 6307
rect 5224 6276 5365 6304
rect 5224 6264 5230 6276
rect 5353 6273 5365 6276
rect 5399 6273 5411 6307
rect 5353 6267 5411 6273
rect 5442 6264 5448 6316
rect 5500 6304 5506 6316
rect 6273 6307 6331 6313
rect 5500 6276 5593 6304
rect 5500 6264 5506 6276
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7282 6304 7288 6316
rect 6319 6276 7288 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7484 6313 7512 6344
rect 11146 6332 11152 6344
rect 11204 6332 11210 6384
rect 11330 6332 11336 6384
rect 11388 6372 11394 6384
rect 11974 6372 11980 6384
rect 11388 6344 11980 6372
rect 11388 6332 11394 6344
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 15654 6332 15660 6384
rect 15712 6372 15718 6384
rect 19794 6372 19800 6384
rect 15712 6344 19800 6372
rect 15712 6332 15718 6344
rect 19794 6332 19800 6344
rect 19852 6332 19858 6384
rect 7469 6307 7527 6313
rect 7469 6273 7481 6307
rect 7515 6304 7527 6307
rect 7558 6304 7564 6316
rect 7515 6276 7564 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 11885 6307 11943 6313
rect 9456 6276 9904 6304
rect 9456 6264 9462 6276
rect 5460 6236 5488 6264
rect 3660 6208 5488 6236
rect 6089 6239 6147 6245
rect 3660 6196 3666 6208
rect 6089 6205 6101 6239
rect 6135 6205 6147 6239
rect 6089 6199 6147 6205
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6236 8171 6239
rect 9769 6239 9827 6245
rect 9769 6236 9781 6239
rect 8159 6208 9781 6236
rect 8159 6205 8171 6208
rect 8113 6199 8171 6205
rect 2400 6171 2458 6177
rect 2400 6137 2412 6171
rect 2446 6168 2458 6171
rect 3050 6168 3056 6180
rect 2446 6140 3056 6168
rect 2446 6137 2458 6140
rect 2400 6131 2458 6137
rect 3050 6128 3056 6140
rect 3108 6128 3114 6180
rect 4157 6171 4215 6177
rect 4157 6168 4169 6171
rect 3344 6140 4169 6168
rect 1673 6103 1731 6109
rect 1673 6069 1685 6103
rect 1719 6100 1731 6103
rect 3344 6100 3372 6140
rect 4157 6137 4169 6140
rect 4203 6137 4215 6171
rect 4157 6131 4215 6137
rect 5074 6128 5080 6180
rect 5132 6168 5138 6180
rect 6104 6168 6132 6199
rect 8496 6180 8524 6208
rect 9769 6205 9781 6208
rect 9815 6205 9827 6239
rect 9876 6236 9904 6276
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 12066 6304 12072 6316
rect 11931 6276 12072 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16172 6276 16681 6304
rect 16172 6264 16178 6276
rect 16669 6273 16681 6276
rect 16715 6304 16727 6307
rect 17126 6304 17132 6316
rect 16715 6276 17132 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 17126 6264 17132 6276
rect 17184 6304 17190 6316
rect 17586 6304 17592 6316
rect 17184 6276 17592 6304
rect 17184 6264 17190 6276
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18693 6307 18751 6313
rect 18693 6304 18705 6307
rect 17920 6276 18705 6304
rect 17920 6264 17926 6276
rect 18693 6273 18705 6276
rect 18739 6304 18751 6307
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 18739 6276 19625 6304
rect 18739 6273 18751 6276
rect 18693 6267 18751 6273
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 20809 6307 20867 6313
rect 20809 6304 20821 6307
rect 20496 6276 20821 6304
rect 20496 6264 20502 6276
rect 20809 6273 20821 6276
rect 20855 6273 20867 6307
rect 20809 6267 20867 6273
rect 9876 6208 11008 6236
rect 9769 6199 9827 6205
rect 8202 6168 8208 6180
rect 5132 6140 5396 6168
rect 6104 6140 8208 6168
rect 5132 6128 5138 6140
rect 3786 6100 3792 6112
rect 1719 6072 3372 6100
rect 3747 6072 3792 6100
rect 1719 6069 1731 6072
rect 1673 6063 1731 6069
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 3878 6060 3884 6112
rect 3936 6100 3942 6112
rect 4249 6103 4307 6109
rect 4249 6100 4261 6103
rect 3936 6072 4261 6100
rect 3936 6060 3942 6072
rect 4249 6069 4261 6072
rect 4295 6069 4307 6103
rect 5258 6100 5264 6112
rect 5219 6072 5264 6100
rect 4249 6063 4307 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5368 6100 5396 6140
rect 8202 6128 8208 6140
rect 8260 6128 8266 6180
rect 8294 6128 8300 6180
rect 8352 6177 8358 6180
rect 8352 6171 8416 6177
rect 8352 6137 8370 6171
rect 8404 6137 8416 6171
rect 8352 6131 8416 6137
rect 8352 6128 8358 6131
rect 8478 6128 8484 6180
rect 8536 6128 8542 6180
rect 9398 6168 9404 6180
rect 8588 6140 9404 6168
rect 7193 6103 7251 6109
rect 7193 6100 7205 6103
rect 5368 6072 7205 6100
rect 7193 6069 7205 6072
rect 7239 6069 7251 6103
rect 7193 6063 7251 6069
rect 7285 6103 7343 6109
rect 7285 6069 7297 6103
rect 7331 6100 7343 6103
rect 8588 6100 8616 6140
rect 9398 6128 9404 6140
rect 9456 6128 9462 6180
rect 10014 6171 10072 6177
rect 10014 6168 10026 6171
rect 9508 6140 10026 6168
rect 7331 6072 8616 6100
rect 7331 6069 7343 6072
rect 7285 6063 7343 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9508 6109 9536 6140
rect 10014 6137 10026 6140
rect 10060 6137 10072 6171
rect 10980 6168 11008 6208
rect 11054 6196 11060 6248
rect 11112 6236 11118 6248
rect 12434 6236 12440 6248
rect 11112 6208 12440 6236
rect 11112 6196 11118 6208
rect 12434 6196 12440 6208
rect 12492 6196 12498 6248
rect 12710 6245 12716 6248
rect 12704 6236 12716 6245
rect 12671 6208 12716 6236
rect 12704 6199 12716 6208
rect 12710 6196 12716 6199
rect 12768 6196 12774 6248
rect 14274 6196 14280 6248
rect 14332 6236 14338 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14332 6208 14381 6236
rect 14332 6196 14338 6208
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 16485 6239 16543 6245
rect 16485 6236 16497 6239
rect 14369 6199 14427 6205
rect 14476 6208 16497 6236
rect 12250 6168 12256 6180
rect 10980 6140 12256 6168
rect 10014 6131 10072 6137
rect 12250 6128 12256 6140
rect 12308 6128 12314 6180
rect 14476 6168 14504 6208
rect 16485 6205 16497 6208
rect 16531 6205 16543 6239
rect 16485 6199 16543 6205
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 17276 6208 17417 6236
rect 17276 6196 17282 6208
rect 17405 6205 17417 6208
rect 17451 6205 17463 6239
rect 19426 6236 19432 6248
rect 19387 6208 19432 6236
rect 17405 6199 17463 6205
rect 19426 6196 19432 6208
rect 19484 6196 19490 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20717 6239 20775 6245
rect 20717 6236 20729 6239
rect 20680 6208 20729 6236
rect 20680 6196 20686 6208
rect 20717 6205 20729 6208
rect 20763 6205 20775 6239
rect 20717 6199 20775 6205
rect 12912 6140 14504 6168
rect 14636 6171 14694 6177
rect 9493 6103 9551 6109
rect 9493 6100 9505 6103
rect 9272 6072 9505 6100
rect 9272 6060 9278 6072
rect 9493 6069 9505 6072
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 12912 6100 12940 6140
rect 14636 6137 14648 6171
rect 14682 6168 14694 6171
rect 15102 6168 15108 6180
rect 14682 6140 15108 6168
rect 14682 6137 14694 6140
rect 14636 6131 14694 6137
rect 15102 6128 15108 6140
rect 15160 6128 15166 6180
rect 18417 6171 18475 6177
rect 18417 6168 18429 6171
rect 16040 6140 18429 6168
rect 10652 6072 12940 6100
rect 10652 6060 10658 6072
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13044 6072 13829 6100
rect 13044 6060 13050 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 16040 6109 16068 6140
rect 18417 6137 18429 6140
rect 18463 6137 18475 6171
rect 18417 6131 18475 6137
rect 18782 6128 18788 6180
rect 18840 6168 18846 6180
rect 19242 6168 19248 6180
rect 18840 6140 19248 6168
rect 18840 6128 18846 6140
rect 19242 6128 19248 6140
rect 19300 6168 19306 6180
rect 19300 6140 20668 6168
rect 19300 6128 19306 6140
rect 15749 6103 15807 6109
rect 15749 6100 15761 6103
rect 14608 6072 15761 6100
rect 14608 6060 14614 6072
rect 15749 6069 15761 6072
rect 15795 6069 15807 6103
rect 15749 6063 15807 6069
rect 16025 6103 16083 6109
rect 16025 6069 16037 6103
rect 16071 6069 16083 6103
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16025 6063 16083 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 18049 6103 18107 6109
rect 18049 6069 18061 6103
rect 18095 6100 18107 6103
rect 18322 6100 18328 6112
rect 18095 6072 18328 6100
rect 18095 6069 18107 6072
rect 18049 6063 18107 6069
rect 18322 6060 18328 6072
rect 18380 6060 18386 6112
rect 18506 6060 18512 6112
rect 18564 6100 18570 6112
rect 18564 6072 18609 6100
rect 18564 6060 18570 6072
rect 18690 6060 18696 6112
rect 18748 6100 18754 6112
rect 19061 6103 19119 6109
rect 19061 6100 19073 6103
rect 18748 6072 19073 6100
rect 18748 6060 18754 6072
rect 19061 6069 19073 6072
rect 19107 6069 19119 6103
rect 19061 6063 19119 6069
rect 19521 6103 19579 6109
rect 19521 6069 19533 6103
rect 19567 6100 19579 6103
rect 19610 6100 19616 6112
rect 19567 6072 19616 6100
rect 19567 6069 19579 6072
rect 19521 6063 19579 6069
rect 19610 6060 19616 6072
rect 19668 6060 19674 6112
rect 20640 6109 20668 6140
rect 20625 6103 20683 6109
rect 20625 6069 20637 6103
rect 20671 6069 20683 6103
rect 20625 6063 20683 6069
rect 1104 6010 21620 6032
rect 1104 5958 7846 6010
rect 7898 5958 7910 6010
rect 7962 5958 7974 6010
rect 8026 5958 8038 6010
rect 8090 5958 14710 6010
rect 14762 5958 14774 6010
rect 14826 5958 14838 6010
rect 14890 5958 14902 6010
rect 14954 5958 21620 6010
rect 1104 5936 21620 5958
rect 1946 5896 1952 5908
rect 1907 5868 1952 5896
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2317 5899 2375 5905
rect 2317 5865 2329 5899
rect 2363 5896 2375 5899
rect 3786 5896 3792 5908
rect 2363 5868 3792 5896
rect 2363 5865 2375 5868
rect 2317 5859 2375 5865
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 4028 5868 5212 5896
rect 4028 5856 4034 5868
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 4310 5831 4368 5837
rect 4310 5828 4322 5831
rect 4120 5800 4322 5828
rect 4120 5788 4126 5800
rect 4310 5797 4322 5800
rect 4356 5797 4368 5831
rect 5184 5828 5212 5868
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5316 5868 5825 5896
rect 5316 5856 5322 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 6178 5896 6184 5908
rect 6139 5868 6184 5896
rect 5813 5859 5871 5865
rect 6178 5856 6184 5868
rect 6236 5856 6242 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6454 5896 6460 5908
rect 6319 5868 6460 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 6454 5856 6460 5868
rect 6512 5896 6518 5908
rect 6512 5868 7328 5896
rect 6512 5856 6518 5868
rect 6914 5828 6920 5840
rect 5184 5800 6920 5828
rect 4310 5791 4368 5797
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 7098 5837 7104 5840
rect 7092 5828 7104 5837
rect 7059 5800 7104 5828
rect 7092 5791 7104 5800
rect 7098 5788 7104 5791
rect 7156 5788 7162 5840
rect 7300 5828 7328 5868
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8904 5868 8953 5896
rect 8904 5856 8910 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 10594 5896 10600 5908
rect 8941 5859 8999 5865
rect 9048 5868 10600 5896
rect 9048 5828 9076 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 10689 5899 10747 5905
rect 10689 5865 10701 5899
rect 10735 5896 10747 5899
rect 12069 5899 12127 5905
rect 12069 5896 12081 5899
rect 10735 5868 12081 5896
rect 10735 5865 10747 5868
rect 10689 5859 10747 5865
rect 12069 5865 12081 5868
rect 12115 5865 12127 5899
rect 12069 5859 12127 5865
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 17313 5899 17371 5905
rect 13136 5868 15700 5896
rect 13136 5856 13142 5868
rect 11057 5831 11115 5837
rect 7300 5800 9076 5828
rect 9968 5800 11008 5828
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 6730 5760 6736 5772
rect 4028 5732 6736 5760
rect 4028 5720 4034 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 6932 5760 6960 5788
rect 9968 5760 9996 5800
rect 6932 5732 9996 5760
rect 10042 5720 10048 5772
rect 10100 5760 10106 5772
rect 10980 5760 11008 5800
rect 11057 5797 11069 5831
rect 11103 5828 11115 5831
rect 12158 5828 12164 5840
rect 11103 5800 12164 5828
rect 11103 5797 11115 5800
rect 11057 5791 11115 5797
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 12894 5828 12900 5840
rect 12492 5800 12900 5828
rect 12492 5788 12498 5800
rect 12066 5760 12072 5772
rect 10100 5732 10145 5760
rect 10980 5732 12072 5760
rect 10100 5720 10106 5732
rect 12066 5720 12072 5732
rect 12124 5720 12130 5772
rect 12728 5769 12756 5800
rect 12894 5788 12900 5800
rect 12952 5828 12958 5840
rect 13446 5828 13452 5840
rect 12952 5800 13452 5828
rect 12952 5788 12958 5800
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 12986 5769 12992 5772
rect 12621 5763 12679 5769
rect 12621 5760 12633 5763
rect 12360 5732 12633 5760
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 3050 5692 3056 5704
rect 2639 5664 3056 5692
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 4062 5652 4068 5704
rect 4120 5701 4126 5704
rect 4120 5692 4130 5701
rect 4120 5664 4165 5692
rect 4120 5655 4130 5664
rect 4120 5652 4126 5655
rect 5994 5652 6000 5704
rect 6052 5692 6058 5704
rect 6365 5695 6423 5701
rect 6365 5692 6377 5695
rect 6052 5664 6377 5692
rect 6052 5652 6058 5664
rect 6365 5661 6377 5664
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6696 5664 6837 5692
rect 6696 5652 6702 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 6825 5655 6883 5661
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 9950 5584 9956 5636
rect 10008 5624 10014 5636
rect 10152 5624 10180 5655
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 11149 5695 11207 5701
rect 10284 5664 10329 5692
rect 10284 5652 10290 5664
rect 11149 5661 11161 5695
rect 11195 5692 11207 5695
rect 11238 5692 11244 5704
rect 11195 5664 11244 5692
rect 11195 5661 11207 5664
rect 11149 5655 11207 5661
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11333 5695 11391 5701
rect 11333 5661 11345 5695
rect 11379 5692 11391 5695
rect 11882 5692 11888 5704
rect 11379 5664 11888 5692
rect 11379 5661 11391 5664
rect 11333 5655 11391 5661
rect 11882 5652 11888 5664
rect 11940 5652 11946 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12360 5701 12388 5732
rect 12621 5729 12633 5732
rect 12667 5729 12679 5763
rect 12621 5723 12679 5729
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5729 12771 5763
rect 12980 5760 12992 5769
rect 12947 5732 12992 5760
rect 12713 5723 12771 5729
rect 12980 5723 12992 5732
rect 12986 5720 12992 5723
rect 13044 5720 13050 5772
rect 13998 5720 14004 5772
rect 14056 5760 14062 5772
rect 14369 5763 14427 5769
rect 14369 5760 14381 5763
rect 14056 5732 14381 5760
rect 14056 5720 14062 5732
rect 14369 5729 14381 5732
rect 14415 5729 14427 5763
rect 15672 5760 15700 5868
rect 17313 5865 17325 5899
rect 17359 5865 17371 5899
rect 17313 5859 17371 5865
rect 16114 5788 16120 5840
rect 16172 5837 16178 5840
rect 16172 5831 16236 5837
rect 16172 5797 16190 5831
rect 16224 5797 16236 5831
rect 17328 5828 17356 5859
rect 17586 5856 17592 5908
rect 17644 5896 17650 5908
rect 17644 5868 18000 5896
rect 17644 5856 17650 5868
rect 17862 5837 17868 5840
rect 17856 5828 17868 5837
rect 17328 5800 17868 5828
rect 16172 5791 16236 5797
rect 17856 5791 17868 5800
rect 16172 5788 16178 5791
rect 17862 5788 17868 5791
rect 17920 5788 17926 5840
rect 17972 5828 18000 5868
rect 18506 5856 18512 5908
rect 18564 5896 18570 5908
rect 19245 5899 19303 5905
rect 19245 5896 19257 5899
rect 18564 5868 19257 5896
rect 18564 5856 18570 5868
rect 19245 5865 19257 5868
rect 19291 5865 19303 5899
rect 19245 5859 19303 5865
rect 17972 5800 19840 5828
rect 18138 5760 18144 5772
rect 15672 5732 18144 5760
rect 14369 5723 14427 5729
rect 18138 5720 18144 5732
rect 18196 5720 18202 5772
rect 19150 5720 19156 5772
rect 19208 5760 19214 5772
rect 19613 5763 19671 5769
rect 19613 5760 19625 5763
rect 19208 5732 19625 5760
rect 19208 5720 19214 5732
rect 19613 5729 19625 5732
rect 19659 5729 19671 5763
rect 19613 5723 19671 5729
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 12032 5664 12173 5692
rect 12032 5652 12038 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12345 5695 12403 5701
rect 12345 5661 12357 5695
rect 12391 5661 12403 5695
rect 12345 5655 12403 5661
rect 13814 5652 13820 5704
rect 13872 5692 13878 5704
rect 15654 5692 15660 5704
rect 13872 5664 15660 5692
rect 13872 5652 13878 5664
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 15838 5652 15844 5704
rect 15896 5692 15902 5704
rect 15933 5695 15991 5701
rect 15933 5692 15945 5695
rect 15896 5664 15945 5692
rect 15896 5652 15902 5664
rect 15933 5661 15945 5664
rect 15979 5661 15991 5695
rect 17586 5692 17592 5704
rect 15933 5655 15991 5661
rect 16960 5664 17592 5692
rect 10870 5624 10876 5636
rect 10008 5596 10876 5624
rect 10008 5584 10014 5596
rect 10870 5584 10876 5596
rect 10928 5584 10934 5636
rect 12710 5624 12716 5636
rect 12544 5596 12716 5624
rect 5445 5559 5503 5565
rect 5445 5525 5457 5559
rect 5491 5556 5503 5559
rect 5534 5556 5540 5568
rect 5491 5528 5540 5556
rect 5491 5525 5503 5528
rect 5445 5519 5503 5525
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8294 5556 8300 5568
rect 8251 5528 8300 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 9398 5556 9404 5568
rect 8619 5528 9404 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 9674 5556 9680 5568
rect 9635 5528 9680 5556
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 11974 5556 11980 5568
rect 11747 5528 11980 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 11974 5516 11980 5528
rect 12032 5516 12038 5568
rect 12434 5516 12440 5568
rect 12492 5556 12498 5568
rect 12544 5556 12572 5596
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 14274 5584 14280 5636
rect 14332 5624 14338 5636
rect 15948 5624 15976 5655
rect 14332 5596 15976 5624
rect 14332 5584 14338 5596
rect 12492 5528 12572 5556
rect 12621 5559 12679 5565
rect 12492 5516 12498 5528
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 13630 5556 13636 5568
rect 12667 5528 13636 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 13630 5516 13636 5528
rect 13688 5556 13694 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13688 5528 14105 5556
rect 13688 5516 13694 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 15948 5556 15976 5596
rect 16960 5556 16988 5664
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 19702 5692 19708 5704
rect 19663 5664 19708 5692
rect 19702 5652 19708 5664
rect 19760 5652 19766 5704
rect 19812 5701 19840 5800
rect 20257 5763 20315 5769
rect 20257 5729 20269 5763
rect 20303 5729 20315 5763
rect 20257 5723 20315 5729
rect 19797 5695 19855 5701
rect 19797 5661 19809 5695
rect 19843 5661 19855 5695
rect 19797 5655 19855 5661
rect 19242 5584 19248 5636
rect 19300 5624 19306 5636
rect 20272 5624 20300 5723
rect 19300 5596 20300 5624
rect 19300 5584 19306 5596
rect 18966 5556 18972 5568
rect 15948 5528 16988 5556
rect 18927 5528 18972 5556
rect 14093 5519 14151 5525
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 20441 5559 20499 5565
rect 20441 5525 20453 5559
rect 20487 5556 20499 5559
rect 20990 5556 20996 5568
rect 20487 5528 20996 5556
rect 20487 5525 20499 5528
rect 20441 5519 20499 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 1104 5466 21620 5488
rect 1104 5414 4414 5466
rect 4466 5414 4478 5466
rect 4530 5414 4542 5466
rect 4594 5414 4606 5466
rect 4658 5414 11278 5466
rect 11330 5414 11342 5466
rect 11394 5414 11406 5466
rect 11458 5414 11470 5466
rect 11522 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 18270 5466
rect 18322 5414 18334 5466
rect 18386 5414 21620 5466
rect 1104 5392 21620 5414
rect 2041 5355 2099 5361
rect 2041 5321 2053 5355
rect 2087 5352 2099 5355
rect 2406 5352 2412 5364
rect 2087 5324 2412 5352
rect 2087 5321 2099 5324
rect 2041 5315 2099 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 6086 5352 6092 5364
rect 4120 5324 6092 5352
rect 4120 5312 4126 5324
rect 6086 5312 6092 5324
rect 6144 5312 6150 5364
rect 7285 5355 7343 5361
rect 7285 5321 7297 5355
rect 7331 5352 7343 5355
rect 7650 5352 7656 5364
rect 7331 5324 7656 5352
rect 7331 5321 7343 5324
rect 7285 5315 7343 5321
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8573 5355 8631 5361
rect 8573 5321 8585 5355
rect 8619 5352 8631 5355
rect 9030 5352 9036 5364
rect 8619 5324 9036 5352
rect 8619 5321 8631 5324
rect 8573 5315 8631 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 10137 5355 10195 5361
rect 10137 5321 10149 5355
rect 10183 5352 10195 5355
rect 12434 5352 12440 5364
rect 10183 5324 12440 5352
rect 10183 5321 10195 5324
rect 10137 5315 10195 5321
rect 12434 5312 12440 5324
rect 12492 5312 12498 5364
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 12636 5324 13093 5352
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 7374 5284 7380 5296
rect 6788 5256 7380 5284
rect 6788 5244 6794 5256
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 10594 5284 10600 5296
rect 7935 5256 10600 5284
rect 2222 5176 2228 5228
rect 2280 5216 2286 5228
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2280 5188 2605 5216
rect 2280 5176 2286 5188
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5040 5188 5365 5216
rect 5040 5176 5046 5188
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5534 5216 5540 5228
rect 5447 5188 5540 5216
rect 5353 5179 5411 5185
rect 5534 5176 5540 5188
rect 5592 5216 5598 5228
rect 6546 5216 6552 5228
rect 5592 5188 6552 5216
rect 5592 5176 5598 5188
rect 6546 5176 6552 5188
rect 6604 5176 6610 5228
rect 7098 5176 7104 5228
rect 7156 5216 7162 5228
rect 7650 5216 7656 5228
rect 7156 5188 7656 5216
rect 7156 5176 7162 5188
rect 7650 5176 7656 5188
rect 7708 5216 7714 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7708 5188 7849 5216
rect 7708 5176 7714 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5442 5148 5448 5160
rect 5307 5120 5448 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5718 5108 5724 5160
rect 5776 5148 5782 5160
rect 7745 5151 7803 5157
rect 7745 5148 7757 5151
rect 5776 5120 7757 5148
rect 5776 5108 5782 5120
rect 7745 5117 7757 5120
rect 7791 5148 7803 5151
rect 7935 5148 7963 5256
rect 10594 5244 10600 5256
rect 10652 5244 10658 5296
rect 11790 5284 11796 5296
rect 10796 5256 11796 5284
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 10796 5225 10824 5256
rect 11790 5244 11796 5256
rect 11848 5244 11854 5296
rect 12066 5244 12072 5296
rect 12124 5284 12130 5296
rect 12636 5284 12664 5324
rect 13081 5321 13093 5324
rect 13127 5321 13139 5355
rect 17129 5355 17187 5361
rect 17129 5352 17141 5355
rect 13081 5315 13139 5321
rect 13188 5324 17141 5352
rect 12124 5256 12664 5284
rect 12124 5244 12130 5256
rect 12710 5244 12716 5296
rect 12768 5284 12774 5296
rect 13188 5284 13216 5324
rect 17129 5321 17141 5324
rect 17175 5321 17187 5355
rect 17129 5315 17187 5321
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 17862 5352 17868 5364
rect 17736 5324 17868 5352
rect 17736 5312 17742 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 18049 5355 18107 5361
rect 18049 5352 18061 5355
rect 18012 5324 18061 5352
rect 18012 5312 18018 5324
rect 18049 5321 18061 5324
rect 18095 5321 18107 5355
rect 18049 5315 18107 5321
rect 20530 5312 20536 5364
rect 20588 5352 20594 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20588 5324 21005 5352
rect 20588 5312 20594 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 12768 5256 13216 5284
rect 12768 5244 12774 5256
rect 13814 5244 13820 5296
rect 13872 5284 13878 5296
rect 14458 5284 14464 5296
rect 13872 5256 14464 5284
rect 13872 5244 13878 5256
rect 14458 5244 14464 5256
rect 14516 5244 14522 5296
rect 17589 5287 17647 5293
rect 17589 5253 17601 5287
rect 17635 5284 17647 5287
rect 19610 5284 19616 5296
rect 17635 5256 19616 5284
rect 17635 5253 17647 5256
rect 17589 5247 17647 5253
rect 19610 5244 19616 5256
rect 19668 5244 19674 5296
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8352 5188 9137 5216
rect 8352 5176 8358 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 10781 5219 10839 5225
rect 10781 5185 10793 5219
rect 10827 5185 10839 5219
rect 10781 5179 10839 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 12728 5216 12756 5244
rect 11747 5188 12756 5216
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 12986 5176 12992 5228
rect 13044 5216 13050 5228
rect 13633 5219 13691 5225
rect 13633 5216 13645 5219
rect 13044 5188 13645 5216
rect 13044 5176 13050 5188
rect 13633 5185 13645 5188
rect 13679 5185 13691 5219
rect 14550 5216 14556 5228
rect 14511 5188 14556 5216
rect 13633 5179 13691 5185
rect 14550 5176 14556 5188
rect 14608 5176 14614 5228
rect 18601 5219 18659 5225
rect 18601 5216 18613 5219
rect 17328 5188 18613 5216
rect 7791 5120 7963 5148
rect 7791 5117 7803 5120
rect 7745 5111 7803 5117
rect 8202 5108 8208 5160
rect 8260 5148 8266 5160
rect 8481 5151 8539 5157
rect 8481 5148 8493 5151
rect 8260 5120 8493 5148
rect 8260 5108 8266 5120
rect 8481 5117 8493 5120
rect 8527 5117 8539 5151
rect 8481 5111 8539 5117
rect 9033 5151 9091 5157
rect 9033 5117 9045 5151
rect 9079 5148 9091 5151
rect 9674 5148 9680 5160
rect 9079 5120 9680 5148
rect 9079 5117 9091 5120
rect 9033 5111 9091 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 9950 5108 9956 5160
rect 10008 5148 10014 5160
rect 12437 5151 12495 5157
rect 12437 5148 12449 5151
rect 10008 5120 12449 5148
rect 10008 5108 10014 5120
rect 12437 5117 12449 5120
rect 12483 5117 12495 5151
rect 12437 5111 12495 5117
rect 13170 5108 13176 5160
rect 13228 5148 13234 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13228 5120 13461 5148
rect 13228 5108 13234 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 13538 5108 13544 5160
rect 13596 5148 13602 5160
rect 14369 5151 14427 5157
rect 14369 5148 14381 5151
rect 13596 5120 14381 5148
rect 13596 5108 13602 5120
rect 14369 5117 14381 5120
rect 14415 5117 14427 5151
rect 14369 5111 14427 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5117 15255 5151
rect 15197 5111 15255 5117
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5148 15807 5151
rect 15838 5148 15844 5160
rect 15795 5120 15844 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 2958 5080 2964 5092
rect 2424 5052 2964 5080
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2424 5021 2452 5052
rect 2958 5040 2964 5052
rect 3016 5040 3022 5092
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 11517 5083 11575 5089
rect 4028 5052 11284 5080
rect 4028 5040 4034 5052
rect 2409 5015 2467 5021
rect 2409 5012 2421 5015
rect 2372 4984 2421 5012
rect 2372 4972 2378 4984
rect 2409 4981 2421 4984
rect 2455 4981 2467 5015
rect 2409 4975 2467 4981
rect 2498 4972 2504 5024
rect 2556 5012 2562 5024
rect 4890 5012 4896 5024
rect 2556 4984 2601 5012
rect 4851 4984 4896 5012
rect 2556 4972 2562 4984
rect 4890 4972 4896 4984
rect 4948 4972 4954 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7653 5015 7711 5021
rect 7653 5012 7665 5015
rect 6972 4984 7665 5012
rect 6972 4972 6978 4984
rect 7653 4981 7665 4984
rect 7699 4981 7711 5015
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 7653 4975 7711 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8941 5015 8999 5021
rect 8941 4981 8953 5015
rect 8987 5012 8999 5015
rect 9674 5012 9680 5024
rect 8987 4984 9680 5012
rect 8987 4981 8999 4984
rect 8941 4975 8999 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 10134 4972 10140 5024
rect 10192 5012 10198 5024
rect 10505 5015 10563 5021
rect 10505 5012 10517 5015
rect 10192 4984 10517 5012
rect 10192 4972 10198 4984
rect 10505 4981 10517 4984
rect 10551 4981 10563 5015
rect 10505 4975 10563 4981
rect 10597 5015 10655 5021
rect 10597 4981 10609 5015
rect 10643 5012 10655 5015
rect 10686 5012 10692 5024
rect 10643 4984 10692 5012
rect 10643 4981 10655 4984
rect 10597 4975 10655 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11149 5015 11207 5021
rect 11149 5012 11161 5015
rect 10928 4984 11161 5012
rect 10928 4972 10934 4984
rect 11149 4981 11161 4984
rect 11195 4981 11207 5015
rect 11256 5012 11284 5052
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 11882 5080 11888 5092
rect 11563 5052 11888 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 13906 5040 13912 5092
rect 13964 5080 13970 5092
rect 15013 5083 15071 5089
rect 15013 5080 15025 5083
rect 13964 5052 15025 5080
rect 13964 5040 13970 5052
rect 15013 5049 15025 5052
rect 15059 5080 15071 5083
rect 15212 5080 15240 5111
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16016 5151 16074 5157
rect 16016 5117 16028 5151
rect 16062 5148 16074 5151
rect 17328 5148 17356 5188
rect 18601 5185 18613 5188
rect 18647 5216 18659 5219
rect 18966 5216 18972 5228
rect 18647 5188 18972 5216
rect 18647 5185 18659 5188
rect 18601 5179 18659 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 16062 5120 17356 5148
rect 17405 5151 17463 5157
rect 16062 5117 16074 5120
rect 16016 5111 16074 5117
rect 17405 5117 17417 5151
rect 17451 5148 17463 5151
rect 17954 5148 17960 5160
rect 17451 5120 17960 5148
rect 17451 5117 17463 5120
rect 17405 5111 17463 5117
rect 17954 5108 17960 5120
rect 18012 5108 18018 5160
rect 18506 5148 18512 5160
rect 18467 5120 18512 5148
rect 18506 5108 18512 5120
rect 18564 5108 18570 5160
rect 18690 5148 18696 5160
rect 18616 5120 18696 5148
rect 15059 5052 15240 5080
rect 15059 5049 15071 5052
rect 15013 5043 15071 5049
rect 17586 5040 17592 5092
rect 17644 5080 17650 5092
rect 18322 5080 18328 5092
rect 17644 5052 18328 5080
rect 17644 5040 17650 5052
rect 18322 5040 18328 5052
rect 18380 5040 18386 5092
rect 18417 5083 18475 5089
rect 18417 5049 18429 5083
rect 18463 5080 18475 5083
rect 18616 5080 18644 5120
rect 18690 5108 18696 5120
rect 18748 5108 18754 5160
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 19334 5148 19340 5160
rect 19107 5120 19340 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19334 5108 19340 5120
rect 19392 5108 19398 5160
rect 19518 5108 19524 5160
rect 19576 5148 19582 5160
rect 19613 5151 19671 5157
rect 19613 5148 19625 5151
rect 19576 5120 19625 5148
rect 19576 5108 19582 5120
rect 19613 5117 19625 5120
rect 19659 5117 19671 5151
rect 21174 5148 21180 5160
rect 19613 5111 19671 5117
rect 19720 5120 21180 5148
rect 19720 5080 19748 5120
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 18463 5052 18644 5080
rect 18708 5052 19748 5080
rect 18463 5049 18475 5052
rect 18417 5043 18475 5049
rect 11606 5012 11612 5024
rect 11256 4984 11612 5012
rect 11149 4975 11207 4981
rect 11606 4972 11612 4984
rect 11664 4972 11670 5024
rect 12621 5015 12679 5021
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12986 5012 12992 5024
rect 12667 4984 12992 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12986 4972 12992 4984
rect 13044 4972 13050 5024
rect 13354 4972 13360 5024
rect 13412 5012 13418 5024
rect 13541 5015 13599 5021
rect 13541 5012 13553 5015
rect 13412 4984 13553 5012
rect 13412 4972 13418 4984
rect 13541 4981 13553 4984
rect 13587 4981 13599 5015
rect 13998 5012 14004 5024
rect 13959 4984 14004 5012
rect 13541 4975 13599 4981
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 14274 4972 14280 5024
rect 14332 5012 14338 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 14332 4984 14473 5012
rect 14332 4972 14338 4984
rect 14461 4981 14473 4984
rect 14507 4981 14519 5015
rect 14461 4975 14519 4981
rect 15381 5015 15439 5021
rect 15381 4981 15393 5015
rect 15427 5012 15439 5015
rect 18708 5012 18736 5052
rect 19794 5040 19800 5092
rect 19852 5089 19858 5092
rect 19852 5083 19916 5089
rect 19852 5049 19870 5083
rect 19904 5049 19916 5083
rect 19852 5043 19916 5049
rect 19852 5040 19858 5043
rect 15427 4984 18736 5012
rect 15427 4981 15439 4984
rect 15381 4975 15439 4981
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19245 5015 19303 5021
rect 19245 5012 19257 5015
rect 18840 4984 19257 5012
rect 18840 4972 18846 4984
rect 19245 4981 19257 4984
rect 19291 4981 19303 5015
rect 19245 4975 19303 4981
rect 1104 4922 21620 4944
rect 1104 4870 7846 4922
rect 7898 4870 7910 4922
rect 7962 4870 7974 4922
rect 8026 4870 8038 4922
rect 8090 4870 14710 4922
rect 14762 4870 14774 4922
rect 14826 4870 14838 4922
rect 14890 4870 14902 4922
rect 14954 4870 21620 4922
rect 1104 4848 21620 4870
rect 3694 4808 3700 4820
rect 3655 4780 3700 4808
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 7193 4811 7251 4817
rect 4120 4780 6684 4808
rect 4120 4768 4126 4780
rect 3234 4740 3240 4752
rect 2332 4712 3240 4740
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2332 4681 2360 4712
rect 3234 4700 3240 4712
rect 3292 4740 3298 4752
rect 4154 4740 4160 4752
rect 3292 4712 4160 4740
rect 3292 4700 3298 4712
rect 4154 4700 4160 4712
rect 4212 4740 4218 4752
rect 4608 4743 4666 4749
rect 4212 4712 4384 4740
rect 4212 4700 4218 4712
rect 2317 4675 2375 4681
rect 2317 4672 2329 4675
rect 2188 4644 2329 4672
rect 2188 4632 2194 4644
rect 2317 4641 2329 4644
rect 2363 4641 2375 4675
rect 2317 4635 2375 4641
rect 2584 4675 2642 4681
rect 2584 4641 2596 4675
rect 2630 4672 2642 4675
rect 3142 4672 3148 4684
rect 2630 4644 3148 4672
rect 2630 4641 2642 4644
rect 2584 4635 2642 4641
rect 3142 4632 3148 4644
rect 3200 4632 3206 4684
rect 4356 4681 4384 4712
rect 4608 4709 4620 4743
rect 4654 4740 4666 4743
rect 5534 4740 5540 4752
rect 4654 4712 5540 4740
rect 4654 4709 4666 4712
rect 4608 4703 4666 4709
rect 5534 4700 5540 4712
rect 5592 4700 5598 4752
rect 6656 4740 6684 4780
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 7466 4808 7472 4820
rect 7239 4780 7472 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 7466 4768 7472 4780
rect 7524 4768 7530 4820
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 8754 4808 8760 4820
rect 7607 4780 8760 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9674 4808 9680 4820
rect 9635 4780 9680 4808
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10594 4768 10600 4820
rect 10652 4808 10658 4820
rect 11146 4808 11152 4820
rect 10652 4780 11152 4808
rect 10652 4768 10658 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 12066 4808 12072 4820
rect 12027 4780 12072 4808
rect 12066 4768 12072 4780
rect 12124 4768 12130 4820
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 15194 4808 15200 4820
rect 12207 4780 15200 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 11057 4743 11115 4749
rect 11057 4740 11069 4743
rect 6656 4712 11069 4740
rect 11057 4709 11069 4712
rect 11103 4709 11115 4743
rect 11057 4703 11115 4709
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 12176 4740 12204 4771
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 17773 4811 17831 4817
rect 17773 4777 17785 4811
rect 17819 4808 17831 4811
rect 19150 4808 19156 4820
rect 17819 4780 19156 4808
rect 17819 4777 17831 4780
rect 17773 4771 17831 4777
rect 19150 4768 19156 4780
rect 19208 4768 19214 4820
rect 19794 4808 19800 4820
rect 19755 4780 19800 4808
rect 19794 4768 19800 4780
rect 19852 4768 19858 4820
rect 13630 4749 13636 4752
rect 13624 4740 13636 4749
rect 11572 4712 12204 4740
rect 13591 4712 13636 4740
rect 11572 4700 11578 4712
rect 13624 4703 13636 4712
rect 13630 4700 13636 4703
rect 13688 4700 13694 4752
rect 17221 4743 17279 4749
rect 17221 4709 17233 4743
rect 17267 4740 17279 4743
rect 17678 4740 17684 4752
rect 17267 4712 17684 4740
rect 17267 4709 17279 4712
rect 17221 4703 17279 4709
rect 17678 4700 17684 4712
rect 17736 4740 17742 4752
rect 18662 4743 18720 4749
rect 18662 4740 18674 4743
rect 17736 4712 18674 4740
rect 17736 4700 17742 4712
rect 18662 4709 18674 4712
rect 18708 4709 18720 4743
rect 18662 4703 18720 4709
rect 19334 4700 19340 4752
rect 19392 4740 19398 4752
rect 20349 4743 20407 4749
rect 20349 4740 20361 4743
rect 19392 4712 20361 4740
rect 19392 4700 19398 4712
rect 20349 4709 20361 4712
rect 20395 4709 20407 4743
rect 20349 4703 20407 4709
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 5166 4672 5172 4684
rect 4387 4644 5172 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 8573 4675 8631 4681
rect 8573 4641 8585 4675
rect 8619 4672 8631 4675
rect 9858 4672 9864 4684
rect 8619 4644 9864 4672
rect 8619 4641 8631 4644
rect 8573 4635 8631 4641
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10042 4672 10048 4684
rect 9955 4644 10048 4672
rect 10042 4632 10048 4644
rect 10100 4672 10106 4684
rect 11790 4672 11796 4684
rect 10100 4644 11796 4672
rect 10100 4632 10106 4644
rect 11790 4632 11796 4644
rect 11848 4632 11854 4684
rect 12805 4675 12863 4681
rect 12805 4641 12817 4675
rect 12851 4641 12863 4675
rect 12805 4635 12863 4641
rect 3418 4564 3424 4616
rect 3476 4604 3482 4616
rect 4154 4604 4160 4616
rect 3476 4576 4160 4604
rect 3476 4564 3482 4576
rect 4154 4564 4160 4576
rect 4212 4564 4218 4616
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6457 4607 6515 4613
rect 6457 4604 6469 4607
rect 6328 4576 6469 4604
rect 6328 4564 6334 4576
rect 6457 4573 6469 4576
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6604 4576 6649 4604
rect 6604 4564 6610 4576
rect 7466 4564 7472 4616
rect 7524 4604 7530 4616
rect 7653 4607 7711 4613
rect 7653 4604 7665 4607
rect 7524 4576 7665 4604
rect 7524 4564 7530 4576
rect 7653 4573 7665 4576
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 8662 4604 8668 4616
rect 8623 4576 8668 4604
rect 7745 4567 7803 4573
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 5997 4539 6055 4545
rect 5997 4536 6009 4539
rect 5408 4508 6009 4536
rect 5408 4496 5414 4508
rect 5997 4505 6009 4508
rect 6043 4505 6055 4539
rect 5997 4499 6055 4505
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 6822 4536 6828 4548
rect 6420 4508 6828 4536
rect 6420 4496 6426 4508
rect 6822 4496 6828 4508
rect 6880 4496 6886 4548
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7760 4536 7788 4567
rect 8662 4564 8668 4576
rect 8720 4564 8726 4616
rect 8757 4607 8815 4613
rect 8757 4573 8769 4607
rect 8803 4573 8815 4607
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 8757 4567 8815 4573
rect 7616 4508 7788 4536
rect 7616 4496 7622 4508
rect 7926 4496 7932 4548
rect 7984 4536 7990 4548
rect 8772 4536 8800 4567
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10284 4576 10329 4604
rect 10284 4564 10290 4576
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11112 4576 11345 4604
rect 11112 4564 11118 4576
rect 11333 4573 11345 4576
rect 11379 4604 11391 4607
rect 12158 4604 12164 4616
rect 11379 4576 12164 4604
rect 11379 4573 11391 4576
rect 11333 4567 11391 4573
rect 12158 4564 12164 4576
rect 12216 4604 12222 4616
rect 12345 4607 12403 4613
rect 12345 4604 12357 4607
rect 12216 4576 12357 4604
rect 12216 4564 12222 4576
rect 12345 4573 12357 4576
rect 12391 4604 12403 4607
rect 12710 4604 12716 4616
rect 12391 4576 12716 4604
rect 12391 4573 12403 4576
rect 12345 4567 12403 4573
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 7984 4508 8800 4536
rect 7984 4496 7990 4508
rect 9766 4496 9772 4548
rect 9824 4536 9830 4548
rect 12820 4536 12848 4635
rect 15286 4632 15292 4684
rect 15344 4672 15350 4684
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15344 4644 15669 4672
rect 15344 4632 15350 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4672 16819 4675
rect 17586 4672 17592 4684
rect 16807 4644 17592 4672
rect 16807 4641 16819 4644
rect 16761 4635 16819 4641
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 18506 4672 18512 4684
rect 17880 4644 18512 4672
rect 17880 4616 17908 4644
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 18966 4632 18972 4684
rect 19024 4672 19030 4684
rect 19426 4672 19432 4684
rect 19024 4644 19432 4672
rect 19024 4632 19030 4644
rect 19426 4632 19432 4644
rect 19484 4632 19490 4684
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 20073 4675 20131 4681
rect 20073 4672 20085 4675
rect 19944 4644 20085 4672
rect 19944 4632 19950 4644
rect 20073 4641 20085 4644
rect 20119 4641 20131 4675
rect 20073 4635 20131 4641
rect 13354 4604 13360 4616
rect 13315 4576 13360 4604
rect 13354 4564 13360 4576
rect 13412 4564 13418 4616
rect 16850 4604 16856 4616
rect 16811 4576 16856 4604
rect 16850 4564 16856 4576
rect 16908 4564 16914 4616
rect 17037 4607 17095 4613
rect 17037 4573 17049 4607
rect 17083 4604 17095 4607
rect 17221 4607 17279 4613
rect 17221 4604 17233 4607
rect 17083 4576 17233 4604
rect 17083 4573 17095 4576
rect 17037 4567 17095 4573
rect 17221 4573 17233 4576
rect 17267 4573 17279 4607
rect 17862 4604 17868 4616
rect 17823 4576 17868 4604
rect 17221 4567 17279 4573
rect 17862 4564 17868 4576
rect 17920 4564 17926 4616
rect 17954 4564 17960 4616
rect 18012 4604 18018 4616
rect 18012 4576 18057 4604
rect 18012 4564 18018 4576
rect 18322 4564 18328 4616
rect 18380 4604 18386 4616
rect 18417 4607 18475 4613
rect 18417 4604 18429 4607
rect 18380 4576 18429 4604
rect 18380 4564 18386 4576
rect 18417 4573 18429 4576
rect 18463 4573 18475 4607
rect 18417 4567 18475 4573
rect 9824 4508 12848 4536
rect 16393 4539 16451 4545
rect 9824 4496 9830 4508
rect 16393 4505 16405 4539
rect 16439 4536 16451 4539
rect 16439 4508 18000 4536
rect 16439 4505 16451 4508
rect 16393 4499 16451 4505
rect 17972 4480 18000 4508
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5721 4471 5779 4477
rect 5721 4468 5733 4471
rect 5316 4440 5733 4468
rect 5316 4428 5322 4440
rect 5721 4437 5733 4440
rect 5767 4437 5779 4471
rect 5721 4431 5779 4437
rect 8205 4471 8263 4477
rect 8205 4437 8217 4471
rect 8251 4468 8263 4471
rect 9674 4468 9680 4480
rect 8251 4440 9680 4468
rect 8251 4437 8263 4440
rect 8205 4431 8263 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 10686 4468 10692 4480
rect 10647 4440 10692 4468
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 12894 4468 12900 4480
rect 11747 4440 12900 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 12894 4428 12900 4440
rect 12952 4428 12958 4480
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4468 13047 4471
rect 13630 4468 13636 4480
rect 13035 4440 13636 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14737 4471 14795 4477
rect 14737 4468 14749 4471
rect 14608 4440 14749 4468
rect 14608 4428 14614 4440
rect 14737 4437 14749 4440
rect 14783 4437 14795 4471
rect 14737 4431 14795 4437
rect 15841 4471 15899 4477
rect 15841 4437 15853 4471
rect 15887 4468 15899 4471
rect 16298 4468 16304 4480
rect 15887 4440 16304 4468
rect 15887 4437 15899 4440
rect 15841 4431 15899 4437
rect 16298 4428 16304 4440
rect 16356 4428 16362 4480
rect 17402 4468 17408 4480
rect 17363 4440 17408 4468
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 17954 4428 17960 4480
rect 18012 4428 18018 4480
rect 18432 4468 18460 4567
rect 19518 4468 19524 4480
rect 18432 4440 19524 4468
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 1104 4378 21620 4400
rect 1104 4326 4414 4378
rect 4466 4326 4478 4378
rect 4530 4326 4542 4378
rect 4594 4326 4606 4378
rect 4658 4326 11278 4378
rect 11330 4326 11342 4378
rect 11394 4326 11406 4378
rect 11458 4326 11470 4378
rect 11522 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 18270 4378
rect 18322 4326 18334 4378
rect 18386 4326 21620 4378
rect 1104 4304 21620 4326
rect 2130 4264 2136 4276
rect 1872 4236 2136 4264
rect 1872 4137 1900 4236
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 3237 4267 3295 4273
rect 3237 4264 3249 4267
rect 3200 4236 3249 4264
rect 3200 4224 3206 4236
rect 3237 4233 3249 4236
rect 3283 4264 3295 4267
rect 3602 4264 3608 4276
rect 3283 4236 3608 4264
rect 3283 4233 3295 4236
rect 3237 4227 3295 4233
rect 3602 4224 3608 4236
rect 3660 4224 3666 4276
rect 7650 4224 7656 4276
rect 7708 4264 7714 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 7708 4236 9045 4264
rect 7708 4224 7714 4236
rect 9033 4233 9045 4236
rect 9079 4264 9091 4267
rect 10226 4264 10232 4276
rect 9079 4236 10232 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 11606 4224 11612 4276
rect 11664 4264 11670 4276
rect 12526 4264 12532 4276
rect 11664 4236 12532 4264
rect 11664 4224 11670 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 16850 4264 16856 4276
rect 12636 4236 16436 4264
rect 16811 4236 16856 4264
rect 3694 4156 3700 4208
rect 3752 4196 3758 4208
rect 6270 4196 6276 4208
rect 3752 4168 6276 4196
rect 3752 4156 3758 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 10042 4196 10048 4208
rect 9600 4168 10048 4196
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4097 1915 4131
rect 4062 4128 4068 4140
rect 4023 4100 4068 4128
rect 1857 4091 1915 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4890 4088 4896 4140
rect 4948 4128 4954 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4948 4100 4997 4128
rect 4948 4088 4954 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5169 4131 5227 4137
rect 5169 4097 5181 4131
rect 5215 4128 5227 4131
rect 5258 4128 5264 4140
rect 5215 4100 5264 4128
rect 5215 4097 5227 4100
rect 5169 4091 5227 4097
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 5316 4100 6101 4128
rect 5316 4088 5322 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 6914 4128 6920 4140
rect 6696 4100 6920 4128
rect 6696 4088 6702 4100
rect 6914 4088 6920 4100
rect 6972 4128 6978 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 6972 4100 7665 4128
rect 6972 4088 6978 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 9600 4128 9628 4168
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 11716 4168 12020 4196
rect 7653 4091 7711 4097
rect 8680 4100 9628 4128
rect 9677 4131 9735 4137
rect 2124 4063 2182 4069
rect 2124 4029 2136 4063
rect 2170 4060 2182 4063
rect 3050 4060 3056 4072
rect 2170 4032 3056 4060
rect 2170 4029 2182 4032
rect 2124 4023 2182 4029
rect 3050 4020 3056 4032
rect 3108 4020 3114 4072
rect 7926 4069 7932 4072
rect 7920 4060 7932 4069
rect 3804 4032 7604 4060
rect 7887 4032 7932 4060
rect 1946 3952 1952 4004
rect 2004 3992 2010 4004
rect 3804 3992 3832 4032
rect 2004 3964 3832 3992
rect 3881 3995 3939 4001
rect 2004 3952 2010 3964
rect 3881 3961 3893 3995
rect 3927 3992 3939 3995
rect 7576 3992 7604 4032
rect 7920 4023 7932 4032
rect 7984 4060 7990 4072
rect 8202 4060 8208 4072
rect 7984 4032 8208 4060
rect 7926 4020 7932 4023
rect 7984 4020 7990 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8680 3992 8708 4100
rect 9677 4097 9689 4131
rect 9723 4128 9735 4131
rect 9766 4128 9772 4140
rect 9723 4100 9772 4128
rect 9723 4097 9735 4100
rect 9677 4091 9735 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 11716 4128 11744 4168
rect 11882 4128 11888 4140
rect 11256 4100 11744 4128
rect 11843 4100 11888 4128
rect 9398 4060 9404 4072
rect 9359 4032 9404 4060
rect 9398 4020 9404 4032
rect 9456 4020 9462 4072
rect 10226 4060 10232 4072
rect 10187 4032 10232 4060
rect 10226 4020 10232 4032
rect 10284 4020 10290 4072
rect 10496 4063 10554 4069
rect 10496 4029 10508 4063
rect 10542 4060 10554 4063
rect 11054 4060 11060 4072
rect 10542 4032 11060 4060
rect 10542 4029 10554 4032
rect 10496 4023 10554 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 3927 3964 5580 3992
rect 7576 3964 8708 3992
rect 3927 3961 3939 3964
rect 3881 3955 3939 3961
rect 3510 3924 3516 3936
rect 3471 3896 3516 3924
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 3973 3927 4031 3933
rect 3973 3893 3985 3927
rect 4019 3924 4031 3927
rect 4525 3927 4583 3933
rect 4525 3924 4537 3927
rect 4019 3896 4537 3924
rect 4019 3893 4031 3896
rect 3973 3887 4031 3893
rect 4525 3893 4537 3896
rect 4571 3893 4583 3927
rect 4525 3887 4583 3893
rect 4893 3927 4951 3933
rect 4893 3893 4905 3927
rect 4939 3924 4951 3927
rect 5350 3924 5356 3936
rect 4939 3896 5356 3924
rect 4939 3893 4951 3896
rect 4893 3887 4951 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5552 3933 5580 3964
rect 8754 3952 8760 4004
rect 8812 3992 8818 4004
rect 11256 3992 11284 4100
rect 11882 4088 11888 4100
rect 11940 4088 11946 4140
rect 11992 4128 12020 4168
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12636 4196 12664 4236
rect 12492 4168 12664 4196
rect 12728 4168 13124 4196
rect 12492 4156 12498 4168
rect 12728 4128 12756 4168
rect 12894 4128 12900 4140
rect 11992 4100 12756 4128
rect 12855 4100 12900 4128
rect 12894 4088 12900 4100
rect 12952 4088 12958 4140
rect 12989 4131 13047 4137
rect 12989 4097 13001 4131
rect 13035 4097 13047 4131
rect 13096 4128 13124 4168
rect 13096 4100 13860 4128
rect 12989 4091 13047 4097
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4060 11759 4063
rect 13004 4060 13032 4091
rect 11747 4032 13032 4060
rect 11747 4029 11759 4032
rect 11701 4023 11759 4029
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 13725 4063 13783 4069
rect 13725 4060 13737 4063
rect 13412 4032 13737 4060
rect 13412 4020 13418 4032
rect 13725 4029 13737 4032
rect 13771 4029 13783 4063
rect 13832 4060 13860 4100
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 13832 4032 16221 4060
rect 13725 4023 13783 4029
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16408 4060 16436 4236
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 17586 4224 17592 4276
rect 17644 4264 17650 4276
rect 19518 4264 19524 4276
rect 17644 4236 19524 4264
rect 17644 4224 17650 4236
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20530 4156 20536 4208
rect 20588 4196 20594 4208
rect 20588 4168 20668 4196
rect 20588 4156 20594 4168
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 16666 4128 16672 4140
rect 16531 4100 16672 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 16666 4088 16672 4100
rect 16724 4128 16730 4140
rect 17497 4131 17555 4137
rect 17497 4128 17509 4131
rect 16724 4100 17509 4128
rect 16724 4088 16730 4100
rect 17497 4097 17509 4100
rect 17543 4128 17555 4131
rect 18693 4131 18751 4137
rect 18693 4128 18705 4131
rect 17543 4100 18705 4128
rect 17543 4097 17555 4100
rect 17497 4091 17555 4097
rect 18693 4097 18705 4100
rect 18739 4128 18751 4131
rect 19334 4128 19340 4140
rect 18739 4100 19340 4128
rect 18739 4097 18751 4100
rect 18693 4091 18751 4097
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19705 4131 19763 4137
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 19794 4128 19800 4140
rect 19751 4100 19800 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 19794 4088 19800 4100
rect 19852 4088 19858 4140
rect 20640 4137 20668 4168
rect 20625 4131 20683 4137
rect 20625 4097 20637 4131
rect 20671 4097 20683 4131
rect 20625 4091 20683 4097
rect 17218 4060 17224 4072
rect 16408 4032 17224 4060
rect 16209 4023 16267 4029
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17310 4020 17316 4072
rect 17368 4060 17374 4072
rect 17586 4060 17592 4072
rect 17368 4032 17592 4060
rect 17368 4020 17374 4032
rect 17586 4020 17592 4032
rect 17644 4020 17650 4072
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 19429 4063 19487 4069
rect 19429 4060 19441 4063
rect 18012 4032 19441 4060
rect 18012 4020 18018 4032
rect 19429 4029 19441 4032
rect 19475 4029 19487 4063
rect 19429 4023 19487 4029
rect 20441 4063 20499 4069
rect 20441 4029 20453 4063
rect 20487 4060 20499 4063
rect 20530 4060 20536 4072
rect 20487 4032 20536 4060
rect 20487 4029 20499 4032
rect 20441 4023 20499 4029
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 8812 3964 11284 3992
rect 8812 3952 8818 3964
rect 11514 3952 11520 4004
rect 11572 3992 11578 4004
rect 12805 3995 12863 4001
rect 12805 3992 12817 3995
rect 11572 3964 12817 3992
rect 11572 3952 11578 3964
rect 12805 3961 12817 3964
rect 12851 3961 12863 3995
rect 12805 3955 12863 3961
rect 13992 3995 14050 4001
rect 13992 3961 14004 3995
rect 14038 3992 14050 3995
rect 14038 3964 14320 3992
rect 14038 3961 14050 3964
rect 13992 3955 14050 3961
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3893 5595 3927
rect 5537 3887 5595 3893
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5684 3896 5917 3924
rect 5684 3884 5690 3896
rect 5905 3893 5917 3896
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 10042 3924 10048 3936
rect 6043 3896 10048 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 10042 3884 10048 3896
rect 10100 3924 10106 3936
rect 11330 3924 11336 3936
rect 10100 3896 11336 3924
rect 10100 3884 10106 3896
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11606 3924 11612 3936
rect 11519 3896 11612 3924
rect 11606 3884 11612 3896
rect 11664 3924 11670 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11664 3896 11713 3924
rect 11664 3884 11670 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 14292 3924 14320 3964
rect 14366 3952 14372 4004
rect 14424 3992 14430 4004
rect 16301 3995 16359 4001
rect 16301 3992 16313 3995
rect 14424 3964 16313 3992
rect 14424 3952 14430 3964
rect 16301 3961 16313 3964
rect 16347 3961 16359 3995
rect 16301 3955 16359 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 18138 3992 18144 4004
rect 17000 3964 18144 3992
rect 17000 3952 17006 3964
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18417 3995 18475 4001
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 18598 3992 18604 4004
rect 18463 3964 18604 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 20254 3992 20260 4004
rect 19076 3964 20260 3992
rect 14550 3924 14556 3936
rect 12492 3896 12537 3924
rect 14292 3896 14556 3924
rect 12492 3884 12498 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15102 3924 15108 3936
rect 15063 3896 15108 3924
rect 15102 3884 15108 3896
rect 15160 3884 15166 3936
rect 15381 3927 15439 3933
rect 15381 3893 15393 3927
rect 15427 3924 15439 3927
rect 15654 3924 15660 3936
rect 15427 3896 15660 3924
rect 15427 3893 15439 3896
rect 15381 3887 15439 3893
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 15841 3927 15899 3933
rect 15841 3893 15853 3927
rect 15887 3924 15899 3927
rect 17126 3924 17132 3936
rect 15887 3896 17132 3924
rect 15887 3893 15899 3896
rect 15841 3887 15899 3893
rect 17126 3884 17132 3896
rect 17184 3884 17190 3936
rect 17310 3924 17316 3936
rect 17271 3896 17316 3924
rect 17310 3884 17316 3896
rect 17368 3884 17374 3936
rect 17402 3884 17408 3936
rect 17460 3924 17466 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17460 3896 18061 3924
rect 17460 3884 17466 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18506 3884 18512 3936
rect 18564 3924 18570 3936
rect 19076 3933 19104 3964
rect 20254 3952 20260 3964
rect 20312 3952 20318 4004
rect 19061 3927 19119 3933
rect 18564 3896 18609 3924
rect 18564 3884 18570 3896
rect 19061 3893 19073 3927
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 19334 3884 19340 3936
rect 19392 3924 19398 3936
rect 19521 3927 19579 3933
rect 19521 3924 19533 3927
rect 19392 3896 19533 3924
rect 19392 3884 19398 3896
rect 19521 3893 19533 3896
rect 19567 3893 19579 3927
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 19521 3887 19579 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 20533 3927 20591 3933
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 20898 3924 20904 3936
rect 20579 3896 20904 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 20898 3884 20904 3896
rect 20956 3884 20962 3936
rect 1104 3834 21620 3856
rect 1104 3782 7846 3834
rect 7898 3782 7910 3834
rect 7962 3782 7974 3834
rect 8026 3782 8038 3834
rect 8090 3782 14710 3834
rect 14762 3782 14774 3834
rect 14826 3782 14838 3834
rect 14890 3782 14902 3834
rect 14954 3782 21620 3834
rect 1104 3760 21620 3782
rect 3053 3723 3111 3729
rect 3053 3689 3065 3723
rect 3099 3720 3111 3723
rect 3510 3720 3516 3732
rect 3099 3692 3516 3720
rect 3099 3689 3111 3692
rect 3053 3683 3111 3689
rect 3510 3680 3516 3692
rect 3568 3680 3574 3732
rect 10134 3720 10140 3732
rect 4908 3692 10140 3720
rect 198 3612 204 3664
rect 256 3652 262 3664
rect 2866 3652 2872 3664
rect 256 3624 2872 3652
rect 256 3612 262 3624
rect 2866 3612 2872 3624
rect 2924 3612 2930 3664
rect 4908 3652 4936 3692
rect 10134 3680 10140 3692
rect 10192 3680 10198 3732
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10965 3723 11023 3729
rect 10965 3720 10977 3723
rect 10744 3692 10977 3720
rect 10744 3680 10750 3692
rect 10965 3689 10977 3692
rect 11011 3689 11023 3723
rect 11514 3720 11520 3732
rect 11475 3692 11520 3720
rect 10965 3683 11023 3689
rect 11514 3680 11520 3692
rect 11572 3680 11578 3732
rect 11882 3720 11888 3732
rect 11843 3692 11888 3720
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12434 3680 12440 3732
rect 12492 3720 12498 3732
rect 12989 3723 13047 3729
rect 12989 3720 13001 3723
rect 12492 3692 13001 3720
rect 12492 3680 12498 3692
rect 12989 3689 13001 3692
rect 13035 3689 13047 3723
rect 14366 3720 14372 3732
rect 12989 3683 13047 3689
rect 13096 3692 14372 3720
rect 3068 3624 4936 3652
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 2961 3587 3019 3593
rect 2961 3584 2973 3587
rect 2464 3556 2973 3584
rect 2464 3544 2470 3556
rect 2961 3553 2973 3556
rect 3007 3553 3019 3587
rect 2961 3547 3019 3553
rect 1026 3476 1032 3528
rect 1084 3516 1090 3528
rect 3068 3516 3096 3624
rect 5534 3612 5540 3664
rect 5592 3652 5598 3664
rect 7466 3652 7472 3664
rect 5592 3624 7472 3652
rect 5592 3612 5598 3624
rect 7466 3612 7472 3624
rect 7524 3652 7530 3664
rect 9950 3652 9956 3664
rect 7524 3624 9812 3652
rect 9911 3624 9956 3652
rect 7524 3612 7530 3624
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 5074 3584 5080 3596
rect 4479 3556 5080 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 5074 3544 5080 3556
rect 5132 3544 5138 3596
rect 5166 3544 5172 3596
rect 5224 3584 5230 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5224 3556 5825 3584
rect 5224 3544 5230 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 6080 3587 6138 3593
rect 6080 3553 6092 3587
rect 6126 3584 6138 3587
rect 6362 3584 6368 3596
rect 6126 3556 6368 3584
rect 6126 3553 6138 3556
rect 6080 3547 6138 3553
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 8110 3584 8116 3596
rect 7064 3556 8116 3584
rect 7064 3544 7070 3556
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8570 3584 8576 3596
rect 8531 3556 8576 3584
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 8846 3584 8852 3596
rect 8711 3556 8852 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9674 3584 9680 3596
rect 9635 3556 9680 3584
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 1084 3488 3096 3516
rect 3237 3519 3295 3525
rect 1084 3476 1090 3488
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3602 3516 3608 3528
rect 3283 3488 3608 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3602 3476 3608 3488
rect 3660 3476 3666 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 4304 3488 4537 3516
rect 4304 3476 4310 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 4890 3516 4896 3528
rect 4755 3488 4896 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 4890 3476 4896 3488
rect 4948 3516 4954 3528
rect 5258 3516 5264 3528
rect 4948 3488 5264 3516
rect 4948 3476 4954 3488
rect 5258 3476 5264 3488
rect 5316 3476 5322 3528
rect 7466 3516 7472 3528
rect 7427 3488 7472 3516
rect 7466 3476 7472 3488
rect 7524 3476 7530 3528
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 8386 3516 8392 3528
rect 7616 3488 8392 3516
rect 7616 3476 7622 3488
rect 8386 3476 8392 3488
rect 8444 3476 8450 3528
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 3326 3448 3332 3460
rect 2639 3420 3332 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 7098 3408 7104 3460
rect 7156 3448 7162 3460
rect 8205 3451 8263 3457
rect 8205 3448 8217 3451
rect 7156 3420 8217 3448
rect 7156 3408 7162 3420
rect 8205 3417 8217 3420
rect 8251 3417 8263 3451
rect 8772 3448 8800 3479
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9582 3516 9588 3528
rect 8996 3488 9588 3516
rect 8996 3476 9002 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9784 3516 9812 3624
rect 9950 3612 9956 3624
rect 10008 3612 10014 3664
rect 10152 3584 10180 3680
rect 10870 3652 10876 3664
rect 10831 3624 10876 3652
rect 10870 3612 10876 3624
rect 10928 3612 10934 3664
rect 11977 3655 12035 3661
rect 11977 3652 11989 3655
rect 10980 3624 11989 3652
rect 10980 3584 11008 3624
rect 11977 3621 11989 3624
rect 12023 3621 12035 3655
rect 13096 3652 13124 3692
rect 14366 3680 14372 3692
rect 14424 3680 14430 3732
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 15289 3723 15347 3729
rect 15289 3720 15301 3723
rect 14599 3692 15301 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 15289 3689 15301 3692
rect 15335 3689 15347 3723
rect 15654 3720 15660 3732
rect 15615 3692 15660 3720
rect 15289 3683 15347 3689
rect 15654 3680 15660 3692
rect 15712 3680 15718 3732
rect 15749 3723 15807 3729
rect 15749 3689 15761 3723
rect 15795 3720 15807 3723
rect 16482 3720 16488 3732
rect 15795 3692 16488 3720
rect 15795 3689 15807 3692
rect 15749 3683 15807 3689
rect 16482 3680 16488 3692
rect 16540 3720 16546 3732
rect 16540 3692 17632 3720
rect 16540 3680 16546 3692
rect 11977 3615 12035 3621
rect 12084 3624 13124 3652
rect 12084 3584 12112 3624
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14645 3655 14703 3661
rect 14645 3652 14657 3655
rect 14056 3624 14657 3652
rect 14056 3612 14062 3624
rect 14645 3621 14657 3624
rect 14691 3621 14703 3655
rect 14645 3615 14703 3621
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 16666 3661 16672 3664
rect 16660 3652 16672 3661
rect 15896 3624 16436 3652
rect 16627 3624 16672 3652
rect 15896 3612 15902 3624
rect 10152 3556 11008 3584
rect 11072 3556 12112 3584
rect 12897 3587 12955 3593
rect 11072 3516 11100 3556
rect 12897 3553 12909 3587
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3584 13691 3587
rect 13722 3584 13728 3596
rect 13679 3556 13728 3584
rect 13679 3553 13691 3556
rect 13633 3547 13691 3553
rect 9784 3488 11100 3516
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11606 3516 11612 3528
rect 11195 3488 11612 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12158 3516 12164 3528
rect 12119 3488 12164 3516
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 8846 3448 8852 3460
rect 8759 3420 8852 3448
rect 8205 3411 8263 3417
rect 8846 3408 8852 3420
rect 8904 3448 8910 3460
rect 10505 3451 10563 3457
rect 8904 3420 10364 3448
rect 8904 3408 8910 3420
rect 2866 3340 2872 3392
rect 2924 3380 2930 3392
rect 4065 3383 4123 3389
rect 4065 3380 4077 3383
rect 2924 3352 4077 3380
rect 2924 3340 2930 3352
rect 4065 3349 4077 3352
rect 4111 3349 4123 3383
rect 4065 3343 4123 3349
rect 7006 3340 7012 3392
rect 7064 3380 7070 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 7064 3352 7205 3380
rect 7064 3340 7070 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 9030 3340 9036 3392
rect 9088 3380 9094 3392
rect 10226 3380 10232 3392
rect 9088 3352 10232 3380
rect 9088 3340 9094 3352
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10336 3380 10364 3420
rect 10505 3417 10517 3451
rect 10551 3448 10563 3451
rect 12912 3448 12940 3547
rect 13722 3544 13728 3556
rect 13780 3544 13786 3596
rect 14550 3544 14556 3596
rect 14608 3584 14614 3596
rect 16408 3593 16436 3624
rect 16660 3615 16672 3624
rect 16666 3612 16672 3615
rect 16724 3612 16730 3664
rect 17604 3652 17632 3692
rect 17678 3680 17684 3732
rect 17736 3720 17742 3732
rect 17773 3723 17831 3729
rect 17773 3720 17785 3723
rect 17736 3692 17785 3720
rect 17736 3680 17742 3692
rect 17773 3689 17785 3692
rect 17819 3689 17831 3723
rect 18506 3720 18512 3732
rect 18467 3692 18512 3720
rect 17773 3683 17831 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 18966 3720 18972 3732
rect 18616 3692 18972 3720
rect 18230 3652 18236 3664
rect 17604 3624 18236 3652
rect 18230 3612 18236 3624
rect 18288 3612 18294 3664
rect 16393 3587 16451 3593
rect 14608 3556 15884 3584
rect 14608 3544 14614 3556
rect 13078 3516 13084 3528
rect 13039 3488 13084 3516
rect 13078 3476 13084 3488
rect 13136 3476 13142 3528
rect 14829 3519 14887 3525
rect 14829 3485 14841 3519
rect 14875 3516 14887 3519
rect 15102 3516 15108 3528
rect 14875 3488 15108 3516
rect 14875 3485 14887 3488
rect 14829 3479 14887 3485
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 15856 3525 15884 3556
rect 16393 3553 16405 3587
rect 16439 3584 16451 3587
rect 17862 3584 17868 3596
rect 16439 3556 17868 3584
rect 16439 3553 16451 3556
rect 16393 3547 16451 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18506 3544 18512 3596
rect 18564 3584 18570 3596
rect 18616 3584 18644 3692
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19242 3720 19248 3732
rect 19116 3692 19248 3720
rect 19116 3680 19122 3692
rect 19242 3680 19248 3692
rect 19300 3680 19306 3732
rect 19797 3723 19855 3729
rect 19797 3689 19809 3723
rect 19843 3720 19855 3723
rect 19978 3720 19984 3732
rect 19843 3692 19984 3720
rect 19843 3689 19855 3692
rect 19797 3683 19855 3689
rect 19978 3680 19984 3692
rect 20036 3680 20042 3732
rect 18877 3655 18935 3661
rect 18877 3621 18889 3655
rect 18923 3652 18935 3655
rect 19702 3652 19708 3664
rect 18923 3624 19708 3652
rect 18923 3621 18935 3624
rect 18877 3615 18935 3621
rect 19702 3612 19708 3624
rect 19760 3652 19766 3664
rect 20530 3652 20536 3664
rect 19760 3624 20536 3652
rect 19760 3612 19766 3624
rect 20530 3612 20536 3624
rect 20588 3612 20594 3664
rect 18564 3556 18644 3584
rect 18564 3544 18570 3556
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 20165 3587 20223 3593
rect 20165 3584 20177 3587
rect 19300 3556 20177 3584
rect 19300 3544 19306 3556
rect 20165 3553 20177 3556
rect 20211 3553 20223 3587
rect 20165 3547 20223 3553
rect 15841 3519 15899 3525
rect 15841 3485 15853 3519
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 10551 3420 12940 3448
rect 13817 3451 13875 3457
rect 10551 3417 10563 3420
rect 10505 3411 10563 3417
rect 13817 3417 13829 3451
rect 13863 3448 13875 3451
rect 15010 3448 15016 3460
rect 13863 3420 15016 3448
rect 13863 3417 13875 3420
rect 13817 3411 13875 3417
rect 15010 3408 15016 3420
rect 15068 3408 15074 3460
rect 18064 3448 18092 3479
rect 19058 3476 19064 3528
rect 19116 3516 19122 3528
rect 20257 3519 20315 3525
rect 19116 3488 19161 3516
rect 19116 3476 19122 3488
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 20257 3479 20315 3485
rect 19978 3448 19984 3460
rect 18064 3420 19984 3448
rect 19978 3408 19984 3420
rect 20036 3408 20042 3460
rect 20272 3448 20300 3479
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 20806 3448 20812 3460
rect 20272 3420 20812 3448
rect 20806 3408 20812 3420
rect 20864 3408 20870 3460
rect 10594 3380 10600 3392
rect 10336 3352 10600 3380
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 12526 3380 12532 3392
rect 12487 3352 12532 3380
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 14090 3340 14096 3392
rect 14148 3380 14154 3392
rect 14185 3383 14243 3389
rect 14185 3380 14197 3383
rect 14148 3352 14197 3380
rect 14148 3340 14154 3352
rect 14185 3349 14197 3352
rect 14231 3349 14243 3383
rect 14185 3343 14243 3349
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 20898 3380 20904 3392
rect 17644 3352 20904 3380
rect 17644 3340 17650 3352
rect 20898 3340 20904 3352
rect 20956 3340 20962 3392
rect 1104 3290 21620 3312
rect 1104 3238 4414 3290
rect 4466 3238 4478 3290
rect 4530 3238 4542 3290
rect 4594 3238 4606 3290
rect 4658 3238 11278 3290
rect 11330 3238 11342 3290
rect 11394 3238 11406 3290
rect 11458 3238 11470 3290
rect 11522 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 18270 3290
rect 18322 3238 18334 3290
rect 18386 3238 21620 3290
rect 1104 3216 21620 3238
rect 2406 3176 2412 3188
rect 2367 3148 2412 3176
rect 2406 3136 2412 3148
rect 2464 3136 2470 3188
rect 3329 3179 3387 3185
rect 3329 3176 3341 3179
rect 2516 3148 3341 3176
rect 1486 3068 1492 3120
rect 1544 3108 1550 3120
rect 2516 3108 2544 3148
rect 3329 3145 3341 3148
rect 3375 3145 3387 3179
rect 4062 3176 4068 3188
rect 3329 3139 3387 3145
rect 3436 3148 4068 3176
rect 3142 3108 3148 3120
rect 1544 3080 2544 3108
rect 2608 3080 3148 3108
rect 1544 3068 1550 3080
rect 566 3000 572 3052
rect 624 3040 630 3052
rect 2608 3040 2636 3080
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 624 3012 2636 3040
rect 624 3000 630 3012
rect 2866 3000 2872 3052
rect 2924 3000 2930 3052
rect 3050 3040 3056 3052
rect 2963 3012 3056 3040
rect 3050 3000 3056 3012
rect 3108 3040 3114 3052
rect 3436 3040 3464 3148
rect 4062 3136 4068 3148
rect 4120 3176 4126 3188
rect 4801 3179 4859 3185
rect 4801 3176 4813 3179
rect 4120 3148 4813 3176
rect 4120 3136 4126 3148
rect 4801 3145 4813 3148
rect 4847 3145 4859 3179
rect 4801 3139 4859 3145
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 8202 3176 8208 3188
rect 5767 3148 8064 3176
rect 8163 3148 8208 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 5994 3068 6000 3120
rect 6052 3108 6058 3120
rect 6730 3108 6736 3120
rect 6052 3080 6736 3108
rect 6052 3068 6058 3080
rect 6730 3068 6736 3080
rect 6788 3068 6794 3120
rect 5074 3040 5080 3052
rect 3108 3012 3464 3040
rect 5035 3012 5080 3040
rect 3108 3000 3114 3012
rect 5074 3000 5080 3012
rect 5132 3000 5138 3052
rect 6362 3040 6368 3052
rect 6275 3012 6368 3040
rect 6362 3000 6368 3012
rect 6420 3040 6426 3052
rect 8036 3040 8064 3148
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 12710 3176 12716 3188
rect 8711 3148 12716 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 16577 3179 16635 3185
rect 16577 3145 16589 3179
rect 16623 3176 16635 3179
rect 18966 3176 18972 3188
rect 16623 3148 18972 3176
rect 16623 3145 16635 3148
rect 16577 3139 16635 3145
rect 18966 3136 18972 3148
rect 19024 3136 19030 3188
rect 8478 3068 8484 3120
rect 8536 3108 8542 3120
rect 8938 3108 8944 3120
rect 8536 3080 8944 3108
rect 8536 3068 8542 3080
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 12250 3108 12256 3120
rect 11848 3080 12256 3108
rect 11848 3068 11854 3080
rect 12250 3068 12256 3080
rect 12308 3108 12314 3120
rect 17310 3108 17316 3120
rect 12308 3080 17316 3108
rect 12308 3068 12314 3080
rect 17310 3068 17316 3080
rect 17368 3068 17374 3120
rect 22094 3108 22100 3120
rect 19168 3080 22100 3108
rect 13633 3043 13691 3049
rect 6420 3012 6960 3040
rect 8036 3012 9168 3040
rect 6420 3000 6426 3012
rect 2777 2975 2835 2981
rect 2777 2941 2789 2975
rect 2823 2972 2835 2975
rect 2884 2972 2912 3000
rect 2823 2944 2912 2972
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3292 2944 3433 2972
rect 3292 2932 3298 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 6730 2972 6736 2984
rect 3421 2935 3479 2941
rect 3528 2944 6736 2972
rect 2406 2864 2412 2916
rect 2464 2904 2470 2916
rect 3528 2904 3556 2944
rect 6730 2932 6736 2944
rect 6788 2932 6794 2984
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2941 6883 2975
rect 6932 2972 6960 3012
rect 7558 2972 7564 2984
rect 6932 2944 7564 2972
rect 6825 2935 6883 2941
rect 2464 2876 3556 2904
rect 2464 2864 2470 2876
rect 3602 2864 3608 2916
rect 3660 2913 3666 2916
rect 3660 2907 3724 2913
rect 3660 2873 3678 2907
rect 3712 2873 3724 2907
rect 6638 2904 6644 2916
rect 3660 2867 3724 2873
rect 3804 2876 6644 2904
rect 3660 2864 3666 2867
rect 2869 2839 2927 2845
rect 2869 2805 2881 2839
rect 2915 2836 2927 2839
rect 3234 2836 3240 2848
rect 2915 2808 3240 2836
rect 2915 2805 2927 2808
rect 2869 2799 2927 2805
rect 3234 2796 3240 2808
rect 3292 2796 3298 2848
rect 3329 2839 3387 2845
rect 3329 2805 3341 2839
rect 3375 2836 3387 2839
rect 3804 2836 3832 2876
rect 6638 2864 6644 2876
rect 6696 2864 6702 2916
rect 6840 2904 6868 2935
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2941 8539 2975
rect 9030 2972 9036 2984
rect 8991 2944 9036 2972
rect 8481 2935 8539 2941
rect 6914 2904 6920 2916
rect 6840 2876 6920 2904
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 7006 2864 7012 2916
rect 7064 2913 7070 2916
rect 7064 2907 7128 2913
rect 7064 2873 7082 2907
rect 7116 2873 7128 2907
rect 7064 2867 7128 2873
rect 7064 2864 7070 2867
rect 3375 2808 3832 2836
rect 3375 2805 3387 2808
rect 3329 2799 3387 2805
rect 5074 2796 5080 2848
rect 5132 2836 5138 2848
rect 5810 2836 5816 2848
rect 5132 2808 5816 2836
rect 5132 2796 5138 2808
rect 5810 2796 5816 2808
rect 5868 2796 5874 2848
rect 6086 2836 6092 2848
rect 6047 2808 6092 2836
rect 6086 2796 6092 2808
rect 6144 2796 6150 2848
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 8496 2836 8524 2935
rect 9030 2932 9036 2944
rect 9088 2932 9094 2984
rect 9140 2972 9168 3012
rect 13633 3009 13645 3043
rect 13679 3040 13691 3043
rect 15470 3040 15476 3052
rect 13679 3012 15476 3040
rect 13679 3009 13691 3012
rect 13633 3003 13691 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 17402 3040 17408 3052
rect 17363 3012 17408 3040
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17589 3043 17647 3049
rect 17589 3009 17601 3043
rect 17635 3040 17647 3043
rect 17678 3040 17684 3052
rect 17635 3012 17684 3040
rect 17635 3009 17647 3012
rect 17589 3003 17647 3009
rect 17678 3000 17684 3012
rect 17736 3000 17742 3052
rect 17862 3000 17868 3052
rect 17920 3040 17926 3052
rect 18049 3043 18107 3049
rect 18049 3040 18061 3043
rect 17920 3012 18061 3040
rect 17920 3000 17926 3012
rect 18049 3009 18061 3012
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 10226 2972 10232 2984
rect 9140 2944 10232 2972
rect 10226 2932 10232 2944
rect 10284 2932 10290 2984
rect 10318 2932 10324 2984
rect 10376 2972 10382 2984
rect 10689 2975 10747 2981
rect 10689 2972 10701 2975
rect 10376 2944 10701 2972
rect 10376 2932 10382 2944
rect 10689 2941 10701 2944
rect 10735 2941 10747 2975
rect 12618 2972 12624 2984
rect 12579 2944 12624 2972
rect 10689 2935 10747 2941
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12719 2944 13369 2972
rect 9300 2907 9358 2913
rect 9300 2873 9312 2907
rect 9346 2904 9358 2907
rect 10956 2907 11014 2913
rect 9346 2876 10916 2904
rect 9346 2873 9358 2876
rect 9300 2867 9358 2873
rect 10318 2836 10324 2848
rect 6236 2808 6281 2836
rect 8496 2808 10324 2836
rect 6236 2796 6242 2808
rect 10318 2796 10324 2808
rect 10376 2796 10382 2848
rect 10413 2839 10471 2845
rect 10413 2805 10425 2839
rect 10459 2836 10471 2839
rect 10594 2836 10600 2848
rect 10459 2808 10600 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 10594 2796 10600 2808
rect 10652 2796 10658 2848
rect 10888 2836 10916 2876
rect 10956 2873 10968 2907
rect 11002 2904 11014 2907
rect 11606 2904 11612 2916
rect 11002 2876 11612 2904
rect 11002 2873 11014 2876
rect 10956 2867 11014 2873
rect 11606 2864 11612 2876
rect 11664 2864 11670 2916
rect 11974 2864 11980 2916
rect 12032 2904 12038 2916
rect 12719 2904 12747 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 14090 2972 14096 2984
rect 14051 2944 14096 2972
rect 13357 2935 13415 2941
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 14829 2975 14887 2981
rect 14829 2941 14841 2975
rect 14875 2972 14887 2975
rect 14918 2972 14924 2984
rect 14875 2944 14924 2972
rect 14875 2941 14887 2944
rect 14829 2935 14887 2941
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15436 2944 15577 2972
rect 15436 2932 15442 2944
rect 15565 2941 15577 2944
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 16393 2975 16451 2981
rect 16393 2941 16405 2975
rect 16439 2972 16451 2975
rect 17034 2972 17040 2984
rect 16439 2944 17040 2972
rect 16439 2941 16451 2944
rect 16393 2935 16451 2941
rect 17034 2932 17040 2944
rect 17092 2932 17098 2984
rect 17126 2932 17132 2984
rect 17184 2972 17190 2984
rect 17313 2975 17371 2981
rect 17313 2972 17325 2975
rect 17184 2944 17325 2972
rect 17184 2932 17190 2944
rect 17313 2941 17325 2944
rect 17359 2941 17371 2975
rect 17313 2935 17371 2941
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 18138 2972 18144 2984
rect 17552 2944 18144 2972
rect 17552 2932 17558 2944
rect 18138 2932 18144 2944
rect 18196 2932 18202 2984
rect 19168 2972 19196 3080
rect 22094 3068 22100 3080
rect 22152 3068 22158 3120
rect 20438 3040 20444 3052
rect 20399 3012 20444 3040
rect 20438 3000 20444 3012
rect 20496 3000 20502 3052
rect 18248 2944 19196 2972
rect 20257 2975 20315 2981
rect 12032 2876 12747 2904
rect 12897 2907 12955 2913
rect 12032 2864 12038 2876
rect 12897 2873 12909 2907
rect 12943 2904 12955 2907
rect 13538 2904 13544 2916
rect 12943 2876 13544 2904
rect 12943 2873 12955 2876
rect 12897 2867 12955 2873
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 14369 2907 14427 2913
rect 14369 2873 14381 2907
rect 14415 2873 14427 2907
rect 14369 2867 14427 2873
rect 12069 2839 12127 2845
rect 12069 2836 12081 2839
rect 10888 2808 12081 2836
rect 12069 2805 12081 2808
rect 12115 2836 12127 2839
rect 13078 2836 13084 2848
rect 12115 2808 13084 2836
rect 12115 2805 12127 2808
rect 12069 2799 12127 2805
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 14384 2836 14412 2867
rect 14458 2864 14464 2916
rect 14516 2904 14522 2916
rect 15105 2907 15163 2913
rect 15105 2904 15117 2907
rect 14516 2876 15117 2904
rect 14516 2864 14522 2876
rect 15105 2873 15117 2876
rect 15151 2873 15163 2907
rect 15105 2867 15163 2873
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 15252 2876 15853 2904
rect 15252 2864 15258 2876
rect 15841 2873 15853 2876
rect 15887 2873 15899 2907
rect 15841 2867 15899 2873
rect 17862 2864 17868 2916
rect 17920 2904 17926 2916
rect 18248 2904 18276 2944
rect 20257 2941 20269 2975
rect 20303 2972 20315 2975
rect 22554 2972 22560 2984
rect 20303 2944 22560 2972
rect 20303 2941 20315 2944
rect 20257 2935 20315 2941
rect 22554 2932 22560 2944
rect 22612 2932 22618 2984
rect 17920 2876 18276 2904
rect 18316 2907 18374 2913
rect 17920 2864 17926 2876
rect 18316 2873 18328 2907
rect 18362 2904 18374 2907
rect 18782 2904 18788 2916
rect 18362 2876 18788 2904
rect 18362 2873 18374 2876
rect 18316 2867 18374 2873
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 18874 2864 18880 2916
rect 18932 2904 18938 2916
rect 21634 2904 21640 2916
rect 18932 2876 21640 2904
rect 18932 2864 18938 2876
rect 21634 2864 21640 2876
rect 21692 2864 21698 2916
rect 15286 2836 15292 2848
rect 14384 2808 15292 2836
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 16945 2839 17003 2845
rect 16945 2805 16957 2839
rect 16991 2836 17003 2839
rect 19334 2836 19340 2848
rect 16991 2808 19340 2836
rect 16991 2805 17003 2808
rect 16945 2799 17003 2805
rect 19334 2796 19340 2808
rect 19392 2796 19398 2848
rect 19426 2796 19432 2848
rect 19484 2836 19490 2848
rect 20162 2836 20168 2848
rect 19484 2808 20168 2836
rect 19484 2796 19490 2808
rect 20162 2796 20168 2808
rect 20220 2796 20226 2848
rect 1104 2746 21620 2768
rect 1104 2694 7846 2746
rect 7898 2694 7910 2746
rect 7962 2694 7974 2746
rect 8026 2694 8038 2746
rect 8090 2694 14710 2746
rect 14762 2694 14774 2746
rect 14826 2694 14838 2746
rect 14890 2694 14902 2746
rect 14954 2694 21620 2746
rect 1104 2672 21620 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 4065 2635 4123 2641
rect 4065 2632 4077 2635
rect 3292 2604 4077 2632
rect 3292 2592 3298 2604
rect 4065 2601 4077 2604
rect 4111 2601 4123 2635
rect 4065 2595 4123 2601
rect 6273 2635 6331 2641
rect 6273 2601 6285 2635
rect 6319 2632 6331 2635
rect 7098 2632 7104 2644
rect 6319 2604 7104 2632
rect 6319 2601 6331 2604
rect 6273 2595 6331 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7285 2635 7343 2641
rect 7285 2601 7297 2635
rect 7331 2632 7343 2635
rect 7466 2632 7472 2644
rect 7331 2604 7472 2632
rect 7331 2601 7343 2604
rect 7285 2595 7343 2601
rect 7466 2592 7472 2604
rect 7524 2592 7530 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2601 8263 2635
rect 8570 2632 8576 2644
rect 8483 2604 8576 2632
rect 8205 2595 8263 2601
rect 3602 2524 3608 2576
rect 3660 2564 3666 2576
rect 4890 2564 4896 2576
rect 3660 2536 4896 2564
rect 3660 2524 3666 2536
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 6181 2567 6239 2573
rect 6181 2533 6193 2567
rect 6227 2564 6239 2567
rect 8220 2564 8248 2595
rect 8570 2592 8576 2604
rect 8628 2632 8634 2644
rect 9306 2632 9312 2644
rect 8628 2604 9312 2632
rect 8628 2592 8634 2604
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9769 2635 9827 2641
rect 9769 2601 9781 2635
rect 9815 2632 9827 2635
rect 9858 2632 9864 2644
rect 9815 2604 9864 2632
rect 9815 2601 9827 2604
rect 9769 2595 9827 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 10226 2632 10232 2644
rect 10187 2604 10232 2632
rect 10226 2592 10232 2604
rect 10284 2592 10290 2644
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 12805 2635 12863 2641
rect 10376 2604 10456 2632
rect 10376 2592 10382 2604
rect 6227 2536 8248 2564
rect 8312 2536 10364 2564
rect 6227 2533 6239 2536
rect 6181 2527 6239 2533
rect 3970 2456 3976 2508
rect 4028 2496 4034 2508
rect 4433 2499 4491 2505
rect 4433 2496 4445 2499
rect 4028 2468 4445 2496
rect 4028 2456 4034 2468
rect 4433 2465 4445 2468
rect 4479 2496 4491 2499
rect 4798 2496 4804 2508
rect 4479 2468 4804 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 2590 2388 2596 2440
rect 2648 2428 2654 2440
rect 4062 2428 4068 2440
rect 2648 2400 4068 2428
rect 2648 2388 2654 2400
rect 4062 2388 4068 2400
rect 4120 2428 4126 2440
rect 4525 2431 4583 2437
rect 4525 2428 4537 2431
rect 4120 2400 4537 2428
rect 4120 2388 4126 2400
rect 4525 2397 4537 2400
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 4908 2428 4936 2524
rect 7006 2496 7012 2508
rect 6472 2468 7012 2496
rect 6472 2437 6500 2468
rect 7006 2456 7012 2468
rect 7064 2496 7070 2508
rect 8312 2496 8340 2536
rect 7064 2468 8340 2496
rect 7064 2456 7070 2468
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 8665 2499 8723 2505
rect 8665 2496 8677 2499
rect 8536 2468 8677 2496
rect 8536 2456 8542 2468
rect 8665 2465 8677 2468
rect 8711 2465 8723 2499
rect 8665 2459 8723 2465
rect 10137 2499 10195 2505
rect 10137 2465 10149 2499
rect 10183 2465 10195 2499
rect 10137 2459 10195 2465
rect 4755 2400 4936 2428
rect 6457 2431 6515 2437
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 6457 2397 6469 2431
rect 6503 2397 6515 2431
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 6457 2391 6515 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7558 2428 7564 2440
rect 7471 2400 7564 2428
rect 7558 2388 7564 2400
rect 7616 2428 7622 2440
rect 8846 2428 8852 2440
rect 7616 2400 8852 2428
rect 7616 2388 7622 2400
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 2866 2320 2872 2372
rect 2924 2360 2930 2372
rect 5718 2360 5724 2372
rect 2924 2332 5724 2360
rect 2924 2320 2930 2332
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 10152 2360 10180 2459
rect 10336 2437 10364 2536
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2397 10379 2431
rect 10428 2428 10456 2604
rect 12805 2601 12817 2635
rect 12851 2632 12863 2635
rect 13998 2632 14004 2644
rect 12851 2604 14004 2632
rect 12851 2601 12863 2604
rect 12805 2595 12863 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 16209 2635 16267 2641
rect 16209 2601 16221 2635
rect 16255 2632 16267 2635
rect 17313 2635 17371 2641
rect 16255 2604 17264 2632
rect 16255 2601 16267 2604
rect 16209 2595 16267 2601
rect 11057 2567 11115 2573
rect 11057 2533 11069 2567
rect 11103 2564 11115 2567
rect 14476 2564 14504 2595
rect 16666 2564 16672 2576
rect 11103 2536 12664 2564
rect 14476 2536 16672 2564
rect 11103 2533 11115 2536
rect 11057 2527 11115 2533
rect 10778 2496 10784 2508
rect 10739 2468 10784 2496
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 12526 2496 12532 2508
rect 11563 2468 12532 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 12526 2456 12532 2468
rect 12584 2456 12590 2508
rect 12636 2505 12664 2536
rect 16666 2524 16672 2536
rect 16724 2524 16730 2576
rect 12621 2499 12679 2505
rect 12621 2465 12633 2499
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13262 2496 13268 2508
rect 13219 2468 13268 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 13538 2456 13544 2508
rect 13596 2496 13602 2508
rect 13725 2499 13783 2505
rect 13725 2496 13737 2499
rect 13596 2468 13737 2496
rect 13596 2456 13602 2468
rect 13725 2465 13737 2468
rect 13771 2465 13783 2499
rect 13725 2459 13783 2465
rect 14277 2499 14335 2505
rect 14277 2465 14289 2499
rect 14323 2496 14335 2499
rect 14458 2496 14464 2508
rect 14323 2468 14464 2496
rect 14323 2465 14335 2468
rect 14277 2459 14335 2465
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 14829 2499 14887 2505
rect 14829 2465 14841 2499
rect 14875 2496 14887 2499
rect 15194 2496 15200 2508
rect 14875 2468 15200 2496
rect 14875 2465 14887 2468
rect 14829 2459 14887 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 15470 2496 15476 2508
rect 15431 2468 15476 2496
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 16025 2499 16083 2505
rect 16025 2465 16037 2499
rect 16071 2496 16083 2499
rect 16206 2496 16212 2508
rect 16071 2468 16212 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 17129 2499 17187 2505
rect 16632 2468 16677 2496
rect 16632 2456 16638 2468
rect 17129 2465 17141 2499
rect 17175 2465 17187 2499
rect 17236 2496 17264 2604
rect 17313 2601 17325 2635
rect 17359 2601 17371 2635
rect 17862 2632 17868 2644
rect 17823 2604 17868 2632
rect 17313 2595 17371 2601
rect 17328 2564 17356 2595
rect 17862 2592 17868 2604
rect 17920 2592 17926 2644
rect 18598 2632 18604 2644
rect 18559 2604 18604 2632
rect 18598 2592 18604 2604
rect 18656 2592 18662 2644
rect 18969 2635 19027 2641
rect 18969 2601 18981 2635
rect 19015 2632 19027 2635
rect 19150 2632 19156 2644
rect 19015 2604 19156 2632
rect 19015 2601 19027 2604
rect 18969 2595 19027 2601
rect 19150 2592 19156 2604
rect 19208 2592 19214 2644
rect 19518 2592 19524 2644
rect 19576 2632 19582 2644
rect 19613 2635 19671 2641
rect 19613 2632 19625 2635
rect 19576 2604 19625 2632
rect 19576 2592 19582 2604
rect 19613 2601 19625 2604
rect 19659 2601 19671 2635
rect 19978 2632 19984 2644
rect 19939 2604 19984 2632
rect 19613 2595 19671 2601
rect 19978 2592 19984 2604
rect 20036 2592 20042 2644
rect 19426 2564 19432 2576
rect 17328 2536 19432 2564
rect 19426 2524 19432 2536
rect 19484 2524 19490 2576
rect 17586 2496 17592 2508
rect 17236 2468 17592 2496
rect 17129 2459 17187 2465
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 10428 2400 11713 2428
rect 10321 2391 10379 2397
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 17144 2428 17172 2459
rect 17586 2456 17592 2468
rect 17644 2456 17650 2508
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 18874 2496 18880 2508
rect 17727 2468 18880 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 18874 2456 18880 2468
rect 18932 2456 18938 2508
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2496 19119 2499
rect 19242 2496 19248 2508
rect 19107 2468 19248 2496
rect 19107 2465 19119 2468
rect 19061 2459 19119 2465
rect 19242 2456 19248 2468
rect 19300 2456 19306 2508
rect 20070 2496 20076 2508
rect 20031 2468 20076 2496
rect 20070 2456 20076 2468
rect 20128 2456 20134 2508
rect 17770 2428 17776 2440
rect 17144 2400 17776 2428
rect 11701 2391 11759 2397
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 19150 2428 19156 2440
rect 19111 2400 19156 2428
rect 19150 2388 19156 2400
rect 19208 2388 19214 2440
rect 20162 2428 20168 2440
rect 20123 2400 20168 2428
rect 20162 2388 20168 2400
rect 20220 2388 20226 2440
rect 6963 2332 10180 2360
rect 13357 2363 13415 2369
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 13357 2329 13369 2363
rect 13403 2360 13415 2363
rect 14366 2360 14372 2372
rect 13403 2332 14372 2360
rect 13403 2329 13415 2332
rect 13357 2323 13415 2329
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 15013 2363 15071 2369
rect 15013 2329 15025 2363
rect 15059 2360 15071 2363
rect 17126 2360 17132 2372
rect 15059 2332 17132 2360
rect 15059 2329 15071 2332
rect 15013 2323 15071 2329
rect 17126 2320 17132 2332
rect 17184 2320 17190 2372
rect 17954 2360 17960 2372
rect 17236 2332 17960 2360
rect 5813 2295 5871 2301
rect 5813 2261 5825 2295
rect 5859 2292 5871 2295
rect 8662 2292 8668 2304
rect 5859 2264 8668 2292
rect 5859 2261 5871 2264
rect 5813 2255 5871 2261
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2292 13967 2295
rect 15378 2292 15384 2304
rect 13955 2264 15384 2292
rect 13955 2261 13967 2264
rect 13909 2255 13967 2261
rect 15378 2252 15384 2264
rect 15436 2252 15442 2304
rect 15657 2295 15715 2301
rect 15657 2261 15669 2295
rect 15703 2292 15715 2295
rect 15838 2292 15844 2304
rect 15703 2264 15844 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 15838 2252 15844 2264
rect 15896 2252 15902 2304
rect 16761 2295 16819 2301
rect 16761 2261 16773 2295
rect 16807 2292 16819 2295
rect 17236 2292 17264 2332
rect 17954 2320 17960 2332
rect 18012 2320 18018 2372
rect 16807 2264 17264 2292
rect 16807 2261 16819 2264
rect 16761 2255 16819 2261
rect 1104 2202 21620 2224
rect 1104 2150 4414 2202
rect 4466 2150 4478 2202
rect 4530 2150 4542 2202
rect 4594 2150 4606 2202
rect 4658 2150 11278 2202
rect 11330 2150 11342 2202
rect 11394 2150 11406 2202
rect 11458 2150 11470 2202
rect 11522 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 18270 2202
rect 18322 2150 18334 2202
rect 18386 2150 21620 2202
rect 1104 2128 21620 2150
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 8478 2088 8484 2100
rect 6696 2060 8484 2088
rect 6696 2048 6702 2060
rect 8478 2048 8484 2060
rect 8536 2048 8542 2100
rect 6730 1980 6736 2032
rect 6788 2020 6794 2032
rect 8570 2020 8576 2032
rect 6788 1992 8576 2020
rect 6788 1980 6794 1992
rect 8570 1980 8576 1992
rect 8628 1980 8634 2032
rect 3970 1232 3976 1284
rect 4028 1272 4034 1284
rect 4982 1272 4988 1284
rect 4028 1244 4988 1272
rect 4028 1232 4034 1244
rect 4982 1232 4988 1244
rect 5040 1232 5046 1284
rect 21082 660 21088 672
rect 20272 632 21088 660
rect 20272 604 20300 632
rect 21082 620 21088 632
rect 21140 620 21146 672
rect 20254 552 20260 604
rect 20312 552 20318 604
rect 20714 552 20720 604
rect 20772 592 20778 604
rect 20990 592 20996 604
rect 20772 564 20996 592
rect 20772 552 20778 564
rect 20990 552 20996 564
rect 21048 552 21054 604
<< via1 >>
rect 7846 20102 7898 20154
rect 7910 20102 7962 20154
rect 7974 20102 8026 20154
rect 8038 20102 8090 20154
rect 14710 20102 14762 20154
rect 14774 20102 14826 20154
rect 14838 20102 14890 20154
rect 14902 20102 14954 20154
rect 4414 19558 4466 19610
rect 4478 19558 4530 19610
rect 4542 19558 4594 19610
rect 4606 19558 4658 19610
rect 11278 19558 11330 19610
rect 11342 19558 11394 19610
rect 11406 19558 11458 19610
rect 11470 19558 11522 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 18270 19558 18322 19610
rect 18334 19558 18386 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 3700 19456 3752 19508
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 20720 19499 20772 19508
rect 20720 19465 20729 19499
rect 20729 19465 20763 19499
rect 20763 19465 20772 19499
rect 20720 19456 20772 19465
rect 4804 19252 4856 19304
rect 5816 19295 5868 19304
rect 5816 19261 5825 19295
rect 5825 19261 5859 19295
rect 5859 19261 5868 19295
rect 5816 19252 5868 19261
rect 18420 19252 18472 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 4896 19184 4948 19236
rect 2780 19116 2832 19168
rect 7846 19014 7898 19066
rect 7910 19014 7962 19066
rect 7974 19014 8026 19066
rect 8038 19014 8090 19066
rect 14710 19014 14762 19066
rect 14774 19014 14826 19066
rect 14838 19014 14890 19066
rect 14902 19014 14954 19066
rect 1952 18955 2004 18964
rect 1952 18921 1961 18955
rect 1961 18921 1995 18955
rect 1995 18921 2004 18955
rect 1952 18912 2004 18921
rect 5816 18844 5868 18896
rect 18420 18887 18472 18896
rect 18420 18853 18429 18887
rect 18429 18853 18463 18887
rect 18463 18853 18472 18887
rect 18420 18844 18472 18853
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 17960 18776 18012 18828
rect 5816 18708 5868 18760
rect 4414 18470 4466 18522
rect 4478 18470 4530 18522
rect 4542 18470 4594 18522
rect 4606 18470 4658 18522
rect 11278 18470 11330 18522
rect 11342 18470 11394 18522
rect 11406 18470 11458 18522
rect 11470 18470 11522 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 18270 18470 18322 18522
rect 18334 18470 18386 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 20720 18411 20772 18420
rect 20720 18377 20729 18411
rect 20729 18377 20763 18411
rect 20763 18377 20772 18411
rect 20720 18368 20772 18377
rect 1768 18207 1820 18216
rect 1768 18173 1777 18207
rect 1777 18173 1811 18207
rect 1811 18173 1820 18207
rect 1768 18164 1820 18173
rect 5724 18164 5776 18216
rect 8208 18164 8260 18216
rect 20536 18207 20588 18216
rect 20536 18173 20545 18207
rect 20545 18173 20579 18207
rect 20579 18173 20588 18207
rect 20536 18164 20588 18173
rect 7846 17926 7898 17978
rect 7910 17926 7962 17978
rect 7974 17926 8026 17978
rect 8038 17926 8090 17978
rect 14710 17926 14762 17978
rect 14774 17926 14826 17978
rect 14838 17926 14890 17978
rect 14902 17926 14954 17978
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 1768 17756 1820 17808
rect 20536 17756 20588 17808
rect 6644 17688 6696 17740
rect 19708 17731 19760 17740
rect 19708 17697 19717 17731
rect 19717 17697 19751 17731
rect 19751 17697 19760 17731
rect 19708 17688 19760 17697
rect 7472 17620 7524 17672
rect 4414 17382 4466 17434
rect 4478 17382 4530 17434
rect 4542 17382 4594 17434
rect 4606 17382 4658 17434
rect 11278 17382 11330 17434
rect 11342 17382 11394 17434
rect 11406 17382 11458 17434
rect 11470 17382 11522 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 18270 17382 18322 17434
rect 18334 17382 18386 17434
rect 1676 17280 1728 17332
rect 20720 17323 20772 17332
rect 20720 17289 20729 17323
rect 20729 17289 20763 17323
rect 20763 17289 20772 17323
rect 20720 17280 20772 17289
rect 6460 17076 6512 17128
rect 19984 17076 20036 17128
rect 7846 16838 7898 16890
rect 7910 16838 7962 16890
rect 7974 16838 8026 16890
rect 8038 16838 8090 16890
rect 14710 16838 14762 16890
rect 14774 16838 14826 16890
rect 14838 16838 14890 16890
rect 14902 16838 14954 16890
rect 1952 16779 2004 16788
rect 1952 16745 1961 16779
rect 1961 16745 1995 16779
rect 1995 16745 2004 16779
rect 1952 16736 2004 16745
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 5356 16600 5408 16652
rect 20536 16600 20588 16652
rect 4414 16294 4466 16346
rect 4478 16294 4530 16346
rect 4542 16294 4594 16346
rect 4606 16294 4658 16346
rect 11278 16294 11330 16346
rect 11342 16294 11394 16346
rect 11406 16294 11458 16346
rect 11470 16294 11522 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 18270 16294 18322 16346
rect 18334 16294 18386 16346
rect 1952 16235 2004 16244
rect 1952 16201 1961 16235
rect 1961 16201 1995 16235
rect 1995 16201 2004 16235
rect 1952 16192 2004 16201
rect 2320 16192 2372 16244
rect 3424 16235 3476 16244
rect 3424 16201 3433 16235
rect 3433 16201 3467 16235
rect 3467 16201 3476 16235
rect 3424 16192 3476 16201
rect 17868 16192 17920 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 20812 16192 20864 16244
rect 7288 16056 7340 16108
rect 3240 16031 3292 16040
rect 3240 15997 3249 16031
rect 3249 15997 3283 16031
rect 3283 15997 3292 16031
rect 3240 15988 3292 15997
rect 12808 15988 12860 16040
rect 19892 15988 19944 16040
rect 5448 15920 5500 15972
rect 19800 15920 19852 15972
rect 7846 15750 7898 15802
rect 7910 15750 7962 15802
rect 7974 15750 8026 15802
rect 8038 15750 8090 15802
rect 14710 15750 14762 15802
rect 14774 15750 14826 15802
rect 14838 15750 14890 15802
rect 14902 15750 14954 15802
rect 1952 15691 2004 15700
rect 1952 15657 1961 15691
rect 1961 15657 1995 15691
rect 1995 15657 2004 15691
rect 1952 15648 2004 15657
rect 2504 15691 2556 15700
rect 2504 15657 2513 15691
rect 2513 15657 2547 15691
rect 2547 15657 2556 15691
rect 2504 15648 2556 15657
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 3240 15580 3292 15632
rect 12808 15623 12860 15632
rect 12808 15589 12817 15623
rect 12817 15589 12851 15623
rect 12851 15589 12860 15623
rect 12808 15580 12860 15589
rect 4252 15512 4304 15564
rect 12532 15555 12584 15564
rect 12532 15521 12541 15555
rect 12541 15521 12575 15555
rect 12575 15521 12584 15555
rect 12532 15512 12584 15521
rect 20076 15512 20128 15564
rect 5080 15444 5132 15496
rect 4160 15376 4212 15428
rect 4414 15206 4466 15258
rect 4478 15206 4530 15258
rect 4542 15206 4594 15258
rect 4606 15206 4658 15258
rect 11278 15206 11330 15258
rect 11342 15206 11394 15258
rect 11406 15206 11458 15258
rect 11470 15206 11522 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 18270 15206 18322 15258
rect 18334 15206 18386 15258
rect 2780 15104 2832 15156
rect 20260 15104 20312 15156
rect 20628 15104 20680 15156
rect 1952 15079 2004 15088
rect 1952 15045 1961 15079
rect 1961 15045 1995 15079
rect 1995 15045 2004 15079
rect 1952 15036 2004 15045
rect 15384 15036 15436 15088
rect 19616 15079 19668 15088
rect 19616 15045 19625 15079
rect 19625 15045 19659 15079
rect 19659 15045 19668 15079
rect 19616 15036 19668 15045
rect 14556 14968 14608 15020
rect 20352 14968 20404 15020
rect 20628 14968 20680 15020
rect 1768 14943 1820 14952
rect 1768 14909 1777 14943
rect 1777 14909 1811 14943
rect 1811 14909 1820 14943
rect 1768 14900 1820 14909
rect 2596 14900 2648 14952
rect 2780 14900 2832 14952
rect 19432 14943 19484 14952
rect 19432 14909 19441 14943
rect 19441 14909 19475 14943
rect 19475 14909 19484 14943
rect 19432 14900 19484 14909
rect 3792 14832 3844 14884
rect 14096 14875 14148 14884
rect 14096 14841 14105 14875
rect 14105 14841 14139 14875
rect 14139 14841 14148 14875
rect 14096 14832 14148 14841
rect 14280 14832 14332 14884
rect 4160 14764 4212 14816
rect 14188 14807 14240 14816
rect 14188 14773 14197 14807
rect 14197 14773 14231 14807
rect 14231 14773 14240 14807
rect 14188 14764 14240 14773
rect 16212 14764 16264 14816
rect 7846 14662 7898 14714
rect 7910 14662 7962 14714
rect 7974 14662 8026 14714
rect 8038 14662 8090 14714
rect 14710 14662 14762 14714
rect 14774 14662 14826 14714
rect 14838 14662 14890 14714
rect 14902 14662 14954 14714
rect 1676 14603 1728 14612
rect 1676 14569 1685 14603
rect 1685 14569 1719 14603
rect 1719 14569 1728 14603
rect 1676 14560 1728 14569
rect 3148 14560 3200 14612
rect 5080 14560 5132 14612
rect 1768 14492 1820 14544
rect 8208 14492 8260 14544
rect 14188 14560 14240 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2872 14424 2924 14476
rect 5264 14424 5316 14476
rect 9772 14424 9824 14476
rect 14004 14492 14056 14544
rect 18880 14560 18932 14612
rect 16212 14535 16264 14544
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 4160 14356 4212 14408
rect 8392 14356 8444 14408
rect 10692 14356 10744 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 14464 14356 14516 14408
rect 16212 14501 16221 14535
rect 16221 14501 16255 14535
rect 16255 14501 16264 14535
rect 16212 14492 16264 14501
rect 16948 14492 17000 14544
rect 19432 14492 19484 14544
rect 17500 14424 17552 14476
rect 19616 14424 19668 14476
rect 16304 14399 16356 14408
rect 16304 14365 16313 14399
rect 16313 14365 16347 14399
rect 16347 14365 16356 14399
rect 16304 14356 16356 14365
rect 15568 14288 15620 14340
rect 19524 14356 19576 14408
rect 10968 14220 11020 14272
rect 12716 14220 12768 14272
rect 13636 14220 13688 14272
rect 16764 14220 16816 14272
rect 18512 14220 18564 14272
rect 19340 14263 19392 14272
rect 19340 14229 19349 14263
rect 19349 14229 19383 14263
rect 19383 14229 19392 14263
rect 19340 14220 19392 14229
rect 4414 14118 4466 14170
rect 4478 14118 4530 14170
rect 4542 14118 4594 14170
rect 4606 14118 4658 14170
rect 11278 14118 11330 14170
rect 11342 14118 11394 14170
rect 11406 14118 11458 14170
rect 11470 14118 11522 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 18270 14118 18322 14170
rect 18334 14118 18386 14170
rect 2780 14016 2832 14068
rect 3516 14016 3568 14068
rect 14556 14059 14608 14068
rect 14556 14025 14565 14059
rect 14565 14025 14599 14059
rect 14599 14025 14608 14059
rect 14556 14016 14608 14025
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 19248 14016 19300 14068
rect 5172 13948 5224 14000
rect 12992 13948 13044 14000
rect 2136 13812 2188 13864
rect 7564 13880 7616 13932
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 10692 13923 10744 13932
rect 10692 13889 10701 13923
rect 10701 13889 10735 13923
rect 10735 13889 10744 13923
rect 10692 13880 10744 13889
rect 11796 13880 11848 13932
rect 13084 13880 13136 13932
rect 3148 13812 3200 13864
rect 4160 13812 4212 13864
rect 5632 13812 5684 13864
rect 10784 13812 10836 13864
rect 10968 13855 11020 13864
rect 10968 13821 11002 13855
rect 11002 13821 11020 13855
rect 10968 13812 11020 13821
rect 14464 13812 14516 13864
rect 19156 13948 19208 14000
rect 16948 13880 17000 13932
rect 3056 13744 3108 13796
rect 5448 13744 5500 13796
rect 3792 13719 3844 13728
rect 3792 13685 3801 13719
rect 3801 13685 3835 13719
rect 3835 13685 3844 13719
rect 3792 13676 3844 13685
rect 6828 13719 6880 13728
rect 6828 13685 6837 13719
rect 6837 13685 6871 13719
rect 6871 13685 6880 13719
rect 6828 13676 6880 13685
rect 8484 13744 8536 13796
rect 8760 13744 8812 13796
rect 14556 13744 14608 13796
rect 19432 13812 19484 13864
rect 20168 13855 20220 13864
rect 15568 13744 15620 13796
rect 16764 13744 16816 13796
rect 17500 13787 17552 13796
rect 17500 13753 17509 13787
rect 17509 13753 17543 13787
rect 17543 13753 17552 13787
rect 17500 13744 17552 13753
rect 17592 13744 17644 13796
rect 20168 13821 20177 13855
rect 20177 13821 20211 13855
rect 20211 13821 20220 13855
rect 20168 13812 20220 13821
rect 20260 13744 20312 13796
rect 9588 13676 9640 13728
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 10416 13676 10468 13728
rect 15936 13676 15988 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16580 13676 16632 13728
rect 7846 13574 7898 13626
rect 7910 13574 7962 13626
rect 7974 13574 8026 13626
rect 8038 13574 8090 13626
rect 14710 13574 14762 13626
rect 14774 13574 14826 13626
rect 14838 13574 14890 13626
rect 14902 13574 14954 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 2872 13472 2924 13524
rect 3240 13472 3292 13524
rect 3332 13472 3384 13524
rect 5080 13515 5132 13524
rect 5080 13481 5089 13515
rect 5089 13481 5123 13515
rect 5123 13481 5132 13515
rect 5080 13472 5132 13481
rect 5448 13472 5500 13524
rect 6092 13472 6144 13524
rect 6828 13472 6880 13524
rect 8760 13472 8812 13524
rect 1952 13336 2004 13388
rect 2320 13379 2372 13388
rect 2320 13345 2329 13379
rect 2329 13345 2363 13379
rect 2363 13345 2372 13379
rect 2320 13336 2372 13345
rect 3884 13336 3936 13388
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 2412 13311 2464 13320
rect 2412 13277 2421 13311
rect 2421 13277 2455 13311
rect 2455 13277 2464 13311
rect 2412 13268 2464 13277
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 3792 13268 3844 13320
rect 5448 13268 5500 13320
rect 11612 13447 11664 13456
rect 11612 13413 11621 13447
rect 11621 13413 11655 13447
rect 11655 13413 11664 13447
rect 11612 13404 11664 13413
rect 14280 13404 14332 13456
rect 7380 13336 7432 13388
rect 7564 13379 7616 13388
rect 7564 13345 7598 13379
rect 7598 13345 7616 13379
rect 7564 13336 7616 13345
rect 9036 13336 9088 13388
rect 10968 13336 11020 13388
rect 13084 13379 13136 13388
rect 13084 13345 13093 13379
rect 13093 13345 13127 13379
rect 13127 13345 13136 13379
rect 13084 13336 13136 13345
rect 13360 13379 13412 13388
rect 13360 13345 13394 13379
rect 13394 13345 13412 13379
rect 14556 13472 14608 13524
rect 16948 13515 17000 13524
rect 16212 13404 16264 13456
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 17132 13404 17184 13456
rect 15568 13379 15620 13388
rect 13360 13336 13412 13345
rect 10784 13311 10836 13320
rect 3976 13200 4028 13252
rect 6184 13200 6236 13252
rect 4712 13175 4764 13184
rect 4712 13141 4721 13175
rect 4721 13141 4755 13175
rect 4755 13141 4764 13175
rect 4712 13132 4764 13141
rect 6828 13132 6880 13184
rect 10784 13277 10793 13311
rect 10793 13277 10827 13311
rect 10827 13277 10836 13311
rect 10784 13268 10836 13277
rect 11796 13311 11848 13320
rect 11796 13277 11805 13311
rect 11805 13277 11839 13311
rect 11839 13277 11848 13311
rect 11796 13268 11848 13277
rect 12808 13268 12860 13320
rect 14188 13268 14240 13320
rect 8392 13200 8444 13252
rect 8484 13200 8536 13252
rect 10600 13200 10652 13252
rect 9404 13132 9456 13184
rect 14464 13175 14516 13184
rect 14464 13141 14473 13175
rect 14473 13141 14507 13175
rect 14507 13141 14516 13175
rect 14464 13132 14516 13141
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 17776 13379 17828 13388
rect 15568 13336 15620 13345
rect 17776 13345 17785 13379
rect 17785 13345 17819 13379
rect 17819 13345 17828 13379
rect 17776 13336 17828 13345
rect 19524 13404 19576 13456
rect 18512 13336 18564 13388
rect 19248 13336 19300 13388
rect 20352 13336 20404 13388
rect 18512 13132 18564 13184
rect 19340 13132 19392 13184
rect 4414 13030 4466 13082
rect 4478 13030 4530 13082
rect 4542 13030 4594 13082
rect 4606 13030 4658 13082
rect 11278 13030 11330 13082
rect 11342 13030 11394 13082
rect 11406 13030 11458 13082
rect 11470 13030 11522 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 18270 13030 18322 13082
rect 18334 13030 18386 13082
rect 2412 12928 2464 12980
rect 3424 12928 3476 12980
rect 3884 12928 3936 12980
rect 9036 12971 9088 12980
rect 9036 12937 9045 12971
rect 9045 12937 9079 12971
rect 9079 12937 9088 12971
rect 9036 12928 9088 12937
rect 9772 12928 9824 12980
rect 3516 12860 3568 12912
rect 6184 12903 6236 12912
rect 1952 12835 2004 12844
rect 1952 12801 1961 12835
rect 1961 12801 1995 12835
rect 1995 12801 2004 12835
rect 1952 12792 2004 12801
rect 2964 12835 3016 12844
rect 2964 12801 2973 12835
rect 2973 12801 3007 12835
rect 3007 12801 3016 12835
rect 2964 12792 3016 12801
rect 3056 12792 3108 12844
rect 3976 12792 4028 12844
rect 6184 12869 6193 12903
rect 6193 12869 6227 12903
rect 6227 12869 6236 12903
rect 6184 12860 6236 12869
rect 10508 12860 10560 12912
rect 8484 12835 8536 12844
rect 8484 12801 8493 12835
rect 8493 12801 8527 12835
rect 8527 12801 8536 12835
rect 8484 12792 8536 12801
rect 9496 12835 9548 12844
rect 9496 12801 9505 12835
rect 9505 12801 9539 12835
rect 9539 12801 9548 12835
rect 9496 12792 9548 12801
rect 9772 12792 9824 12844
rect 10600 12835 10652 12844
rect 10600 12801 10609 12835
rect 10609 12801 10643 12835
rect 10643 12801 10652 12835
rect 10600 12792 10652 12801
rect 10968 12928 11020 12980
rect 14096 12928 14148 12980
rect 16580 12971 16632 12980
rect 16580 12937 16589 12971
rect 16589 12937 16623 12971
rect 16623 12937 16632 12971
rect 16580 12928 16632 12937
rect 20904 12971 20956 12980
rect 20904 12937 20913 12971
rect 20913 12937 20947 12971
rect 20947 12937 20956 12971
rect 20904 12928 20956 12937
rect 17316 12860 17368 12912
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 14464 12835 14516 12844
rect 14464 12801 14473 12835
rect 14473 12801 14507 12835
rect 14507 12801 14516 12835
rect 14464 12792 14516 12801
rect 15844 12792 15896 12844
rect 16212 12792 16264 12844
rect 17776 12792 17828 12844
rect 19616 12792 19668 12844
rect 1768 12767 1820 12776
rect 1768 12733 1777 12767
rect 1777 12733 1811 12767
rect 1811 12733 1820 12767
rect 1768 12724 1820 12733
rect 3884 12724 3936 12776
rect 4712 12724 4764 12776
rect 3516 12656 3568 12708
rect 3700 12656 3752 12708
rect 3976 12656 4028 12708
rect 12440 12724 12492 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 15936 12724 15988 12776
rect 18512 12767 18564 12776
rect 5448 12656 5500 12708
rect 2504 12588 2556 12640
rect 4712 12588 4764 12640
rect 7656 12656 7708 12708
rect 9404 12699 9456 12708
rect 9404 12665 9413 12699
rect 9413 12665 9447 12699
rect 9447 12665 9456 12699
rect 9404 12656 9456 12665
rect 10324 12656 10376 12708
rect 10600 12656 10652 12708
rect 15108 12656 15160 12708
rect 15200 12656 15252 12708
rect 18512 12733 18546 12767
rect 18546 12733 18564 12767
rect 18512 12724 18564 12733
rect 18788 12724 18840 12776
rect 20628 12724 20680 12776
rect 19892 12656 19944 12708
rect 9588 12588 9640 12640
rect 10416 12631 10468 12640
rect 10416 12597 10425 12631
rect 10425 12597 10459 12631
rect 10459 12597 10468 12631
rect 10416 12588 10468 12597
rect 11980 12588 12032 12640
rect 12716 12588 12768 12640
rect 15936 12631 15988 12640
rect 15936 12597 15945 12631
rect 15945 12597 15979 12631
rect 15979 12597 15988 12631
rect 15936 12588 15988 12597
rect 16672 12588 16724 12640
rect 17040 12631 17092 12640
rect 17040 12597 17049 12631
rect 17049 12597 17083 12631
rect 17083 12597 17092 12631
rect 19616 12631 19668 12640
rect 17040 12588 17092 12597
rect 19616 12597 19625 12631
rect 19625 12597 19659 12631
rect 19659 12597 19668 12631
rect 19616 12588 19668 12597
rect 7846 12486 7898 12538
rect 7910 12486 7962 12538
rect 7974 12486 8026 12538
rect 8038 12486 8090 12538
rect 14710 12486 14762 12538
rect 14774 12486 14826 12538
rect 14838 12486 14890 12538
rect 14902 12486 14954 12538
rect 2320 12384 2372 12436
rect 3608 12427 3660 12436
rect 3608 12393 3617 12427
rect 3617 12393 3651 12427
rect 3651 12393 3660 12427
rect 3608 12384 3660 12393
rect 5448 12427 5500 12436
rect 5448 12393 5457 12427
rect 5457 12393 5491 12427
rect 5491 12393 5500 12427
rect 5448 12384 5500 12393
rect 7380 12384 7432 12436
rect 2964 12316 3016 12368
rect 4160 12316 4212 12368
rect 5080 12316 5132 12368
rect 7012 12316 7064 12368
rect 7472 12316 7524 12368
rect 7840 12316 7892 12368
rect 1400 12087 1452 12096
rect 1400 12053 1409 12087
rect 1409 12053 1443 12087
rect 1443 12053 1452 12087
rect 1400 12044 1452 12053
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 3148 12248 3200 12300
rect 3516 12248 3568 12300
rect 5264 12248 5316 12300
rect 8208 12316 8260 12368
rect 12440 12384 12492 12436
rect 15200 12384 15252 12436
rect 15936 12427 15988 12436
rect 15936 12393 15945 12427
rect 15945 12393 15979 12427
rect 15979 12393 15988 12427
rect 15936 12384 15988 12393
rect 16028 12384 16080 12436
rect 17040 12384 17092 12436
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 8576 12248 8628 12300
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 16580 12316 16632 12368
rect 20352 12384 20404 12436
rect 10692 12248 10744 12300
rect 2044 12223 2096 12232
rect 2044 12189 2053 12223
rect 2053 12189 2087 12223
rect 2087 12189 2096 12223
rect 2044 12180 2096 12189
rect 3056 12223 3108 12232
rect 3056 12189 3065 12223
rect 3065 12189 3099 12223
rect 3099 12189 3108 12223
rect 3056 12180 3108 12189
rect 3700 12180 3752 12232
rect 5908 12180 5960 12232
rect 7472 12180 7524 12232
rect 10232 12223 10284 12232
rect 3148 12112 3200 12164
rect 7564 12112 7616 12164
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 11796 12248 11848 12300
rect 14464 12291 14516 12300
rect 14464 12257 14473 12291
rect 14473 12257 14507 12291
rect 14507 12257 14516 12291
rect 14464 12248 14516 12257
rect 16120 12248 16172 12300
rect 17776 12248 17828 12300
rect 3056 12044 3108 12096
rect 3884 12044 3936 12096
rect 10508 12112 10560 12164
rect 11888 12112 11940 12164
rect 13176 12180 13228 12232
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 16488 12223 16540 12232
rect 14740 12180 14792 12189
rect 16488 12189 16497 12223
rect 16497 12189 16531 12223
rect 16531 12189 16540 12223
rect 16488 12180 16540 12189
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 17960 12180 18012 12232
rect 19524 12180 19576 12232
rect 20168 12248 20220 12300
rect 18788 12112 18840 12164
rect 18880 12112 18932 12164
rect 20628 12180 20680 12232
rect 20444 12155 20496 12164
rect 20444 12121 20453 12155
rect 20453 12121 20487 12155
rect 20487 12121 20496 12155
rect 20444 12112 20496 12121
rect 11704 12044 11756 12096
rect 12808 12044 12860 12096
rect 17224 12044 17276 12096
rect 18512 12044 18564 12096
rect 4414 11942 4466 11994
rect 4478 11942 4530 11994
rect 4542 11942 4594 11994
rect 4606 11942 4658 11994
rect 11278 11942 11330 11994
rect 11342 11942 11394 11994
rect 11406 11942 11458 11994
rect 11470 11942 11522 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 18270 11942 18322 11994
rect 18334 11942 18386 11994
rect 4068 11840 4120 11892
rect 11796 11883 11848 11892
rect 2044 11704 2096 11756
rect 6184 11772 6236 11824
rect 7472 11815 7524 11824
rect 7472 11781 7481 11815
rect 7481 11781 7515 11815
rect 7515 11781 7524 11815
rect 7472 11772 7524 11781
rect 5172 11704 5224 11756
rect 3976 11636 4028 11688
rect 5264 11636 5316 11688
rect 5448 11679 5500 11688
rect 5448 11645 5457 11679
rect 5457 11645 5491 11679
rect 5491 11645 5500 11679
rect 7104 11704 7156 11756
rect 5448 11636 5500 11645
rect 8024 11747 8076 11756
rect 8024 11713 8033 11747
rect 8033 11713 8067 11747
rect 8067 11713 8076 11747
rect 8024 11704 8076 11713
rect 3332 11568 3384 11620
rect 1860 11543 1912 11552
rect 1860 11509 1869 11543
rect 1869 11509 1903 11543
rect 1903 11509 1912 11543
rect 1860 11500 1912 11509
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 2320 11543 2372 11552
rect 2320 11509 2329 11543
rect 2329 11509 2363 11543
rect 2363 11509 2372 11543
rect 6920 11568 6972 11620
rect 7012 11568 7064 11620
rect 8392 11772 8444 11824
rect 11796 11849 11805 11883
rect 11805 11849 11839 11883
rect 11839 11849 11848 11883
rect 11796 11840 11848 11849
rect 13084 11840 13136 11892
rect 15016 11840 15068 11892
rect 16856 11840 16908 11892
rect 17500 11840 17552 11892
rect 17960 11840 18012 11892
rect 12716 11772 12768 11824
rect 8484 11636 8536 11688
rect 10048 11704 10100 11756
rect 12992 11747 13044 11756
rect 9496 11636 9548 11688
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 15568 11747 15620 11756
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 19340 11840 19392 11892
rect 20996 11840 21048 11892
rect 11612 11636 11664 11688
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13820 11636 13872 11688
rect 9588 11568 9640 11620
rect 12348 11568 12400 11620
rect 14740 11636 14792 11688
rect 16856 11636 16908 11688
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 18880 11704 18932 11756
rect 19616 11636 19668 11688
rect 20076 11636 20128 11688
rect 20444 11636 20496 11688
rect 20720 11679 20772 11688
rect 20720 11645 20729 11679
rect 20729 11645 20763 11679
rect 20763 11645 20772 11679
rect 20720 11636 20772 11645
rect 15844 11611 15896 11620
rect 15844 11577 15878 11611
rect 15878 11577 15896 11611
rect 15844 11568 15896 11577
rect 16580 11568 16632 11620
rect 2320 11500 2372 11509
rect 3976 11543 4028 11552
rect 3976 11509 3985 11543
rect 3985 11509 4019 11543
rect 4019 11509 4028 11543
rect 3976 11500 4028 11509
rect 4160 11500 4212 11552
rect 5908 11500 5960 11552
rect 6460 11500 6512 11552
rect 7748 11500 7800 11552
rect 8208 11500 8260 11552
rect 8392 11500 8444 11552
rect 10048 11500 10100 11552
rect 10232 11500 10284 11552
rect 13360 11500 13412 11552
rect 16212 11500 16264 11552
rect 17592 11500 17644 11552
rect 18512 11500 18564 11552
rect 19432 11500 19484 11552
rect 7846 11398 7898 11450
rect 7910 11398 7962 11450
rect 7974 11398 8026 11450
rect 8038 11398 8090 11450
rect 14710 11398 14762 11450
rect 14774 11398 14826 11450
rect 14838 11398 14890 11450
rect 14902 11398 14954 11450
rect 2780 11296 2832 11348
rect 6736 11296 6788 11348
rect 7748 11296 7800 11348
rect 8300 11296 8352 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 8668 11296 8720 11348
rect 10876 11296 10928 11348
rect 3240 11228 3292 11280
rect 2688 11160 2740 11212
rect 3700 11160 3752 11212
rect 4068 11160 4120 11212
rect 5908 11228 5960 11280
rect 6000 11228 6052 11280
rect 8392 11228 8444 11280
rect 9036 11271 9088 11280
rect 9036 11237 9045 11271
rect 9045 11237 9079 11271
rect 9079 11237 9088 11271
rect 9036 11228 9088 11237
rect 5448 11160 5500 11212
rect 3516 11024 3568 11076
rect 5540 11024 5592 11076
rect 7288 11160 7340 11212
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 3700 10956 3752 11008
rect 8208 11024 8260 11076
rect 8944 11203 8996 11212
rect 8944 11169 8953 11203
rect 8953 11169 8987 11203
rect 8987 11169 8996 11203
rect 8944 11160 8996 11169
rect 9312 11092 9364 11144
rect 10784 11228 10836 11280
rect 12808 11296 12860 11348
rect 12992 11296 13044 11348
rect 15292 11339 15344 11348
rect 15292 11305 15301 11339
rect 15301 11305 15335 11339
rect 15335 11305 15344 11339
rect 15292 11296 15344 11305
rect 16120 11296 16172 11348
rect 11888 11228 11940 11280
rect 12440 11228 12492 11280
rect 15936 11228 15988 11280
rect 17500 11228 17552 11280
rect 20536 11228 20588 11280
rect 9680 11160 9732 11212
rect 10140 11135 10192 11144
rect 10140 11101 10149 11135
rect 10149 11101 10183 11135
rect 10183 11101 10192 11135
rect 10140 11092 10192 11101
rect 10232 11135 10284 11144
rect 10232 11101 10241 11135
rect 10241 11101 10275 11135
rect 10275 11101 10284 11135
rect 10232 11092 10284 11101
rect 10600 11092 10652 11144
rect 12256 10956 12308 11008
rect 12440 10956 12492 11008
rect 13084 11160 13136 11212
rect 13636 11203 13688 11212
rect 13636 11169 13670 11203
rect 13670 11169 13688 11203
rect 13636 11160 13688 11169
rect 13912 11160 13964 11212
rect 19800 11160 19852 11212
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 12808 11092 12860 11144
rect 13268 11092 13320 11144
rect 14464 11092 14516 11144
rect 15016 11092 15068 11144
rect 15752 11135 15804 11144
rect 15752 11101 15761 11135
rect 15761 11101 15795 11135
rect 15795 11101 15804 11135
rect 15752 11092 15804 11101
rect 16028 11092 16080 11144
rect 16488 11092 16540 11144
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 20352 11135 20404 11144
rect 18880 11024 18932 11076
rect 12808 10956 12860 11008
rect 13544 10956 13596 11008
rect 20352 11101 20361 11135
rect 20361 11101 20395 11135
rect 20395 11101 20404 11135
rect 20352 11092 20404 11101
rect 19892 11024 19944 11076
rect 4414 10854 4466 10906
rect 4478 10854 4530 10906
rect 4542 10854 4594 10906
rect 4606 10854 4658 10906
rect 11278 10854 11330 10906
rect 11342 10854 11394 10906
rect 11406 10854 11458 10906
rect 11470 10854 11522 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 18270 10854 18322 10906
rect 18334 10854 18386 10906
rect 1768 10752 1820 10804
rect 2964 10752 3016 10804
rect 5448 10795 5500 10804
rect 5448 10761 5457 10795
rect 5457 10761 5491 10795
rect 5491 10761 5500 10795
rect 5448 10752 5500 10761
rect 7564 10752 7616 10804
rect 5356 10684 5408 10736
rect 9680 10752 9732 10804
rect 10140 10752 10192 10804
rect 15752 10752 15804 10804
rect 3516 10616 3568 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 3884 10616 3936 10668
rect 6184 10659 6236 10668
rect 2228 10548 2280 10600
rect 2872 10548 2924 10600
rect 3148 10548 3200 10600
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 9312 10684 9364 10736
rect 15108 10684 15160 10736
rect 17132 10752 17184 10804
rect 6828 10659 6880 10668
rect 6828 10625 6837 10659
rect 6837 10625 6871 10659
rect 6871 10625 6880 10659
rect 6828 10616 6880 10625
rect 9588 10659 9640 10668
rect 9588 10625 9597 10659
rect 9597 10625 9631 10659
rect 9631 10625 9640 10659
rect 9588 10616 9640 10625
rect 11888 10659 11940 10668
rect 11888 10625 11897 10659
rect 11897 10625 11931 10659
rect 11931 10625 11940 10659
rect 11888 10616 11940 10625
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 13636 10616 13688 10668
rect 15660 10616 15712 10668
rect 16028 10659 16080 10668
rect 16028 10625 16037 10659
rect 16037 10625 16071 10659
rect 16071 10625 16080 10659
rect 16028 10616 16080 10625
rect 17224 10684 17276 10736
rect 11704 10548 11756 10600
rect 12348 10548 12400 10600
rect 12992 10548 13044 10600
rect 15108 10548 15160 10600
rect 19432 10616 19484 10668
rect 18604 10548 18656 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 19708 10548 19760 10557
rect 3884 10480 3936 10532
rect 5172 10480 5224 10532
rect 5264 10480 5316 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6920 10412 6972 10464
rect 7012 10412 7064 10464
rect 9864 10412 9916 10464
rect 9956 10412 10008 10464
rect 12624 10480 12676 10532
rect 15752 10480 15804 10532
rect 16764 10480 16816 10532
rect 18328 10523 18380 10532
rect 18328 10489 18362 10523
rect 18362 10489 18380 10523
rect 18328 10480 18380 10489
rect 10508 10455 10560 10464
rect 10508 10421 10517 10455
rect 10517 10421 10551 10455
rect 10551 10421 10560 10455
rect 11704 10455 11756 10464
rect 10508 10412 10560 10421
rect 11704 10421 11713 10455
rect 11713 10421 11747 10455
rect 11747 10421 11756 10455
rect 11704 10412 11756 10421
rect 11796 10412 11848 10464
rect 13912 10412 13964 10464
rect 15476 10455 15528 10464
rect 15476 10421 15485 10455
rect 15485 10421 15519 10455
rect 15519 10421 15528 10455
rect 15476 10412 15528 10421
rect 16396 10412 16448 10464
rect 16856 10455 16908 10464
rect 16856 10421 16865 10455
rect 16865 10421 16899 10455
rect 16899 10421 16908 10455
rect 16856 10412 16908 10421
rect 17500 10412 17552 10464
rect 20352 10412 20404 10464
rect 7846 10310 7898 10362
rect 7910 10310 7962 10362
rect 7974 10310 8026 10362
rect 8038 10310 8090 10362
rect 14710 10310 14762 10362
rect 14774 10310 14826 10362
rect 14838 10310 14890 10362
rect 14902 10310 14954 10362
rect 4252 10251 4304 10260
rect 4252 10217 4261 10251
rect 4261 10217 4295 10251
rect 4295 10217 4304 10251
rect 4252 10208 4304 10217
rect 5356 10208 5408 10260
rect 8300 10208 8352 10260
rect 9588 10208 9640 10260
rect 11980 10251 12032 10260
rect 3240 10140 3292 10192
rect 5724 10140 5776 10192
rect 7380 10140 7432 10192
rect 10784 10140 10836 10192
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 12532 10208 12584 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 13820 10208 13872 10260
rect 15108 10208 15160 10260
rect 15292 10208 15344 10260
rect 16396 10208 16448 10260
rect 17224 10208 17276 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 20168 10208 20220 10260
rect 2044 10115 2096 10124
rect 2044 10081 2078 10115
rect 2078 10081 2096 10115
rect 2044 10072 2096 10081
rect 3516 10072 3568 10124
rect 4252 10072 4304 10124
rect 4804 10072 4856 10124
rect 7564 10072 7616 10124
rect 5540 10004 5592 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 4620 9936 4672 9988
rect 5356 9936 5408 9988
rect 5448 9936 5500 9988
rect 5908 10004 5960 10056
rect 6184 10004 6236 10056
rect 8392 10072 8444 10124
rect 9496 10072 9548 10124
rect 10232 10072 10284 10124
rect 11060 10072 11112 10124
rect 11704 10072 11756 10124
rect 14464 10140 14516 10192
rect 15476 10140 15528 10192
rect 19064 10140 19116 10192
rect 20628 10140 20680 10192
rect 13360 10072 13412 10124
rect 14004 10072 14056 10124
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 7748 9936 7800 9988
rect 7932 9936 7984 9988
rect 8484 9936 8536 9988
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 12716 10004 12768 10056
rect 13728 10004 13780 10056
rect 12256 9936 12308 9988
rect 12348 9936 12400 9988
rect 3148 9868 3200 9877
rect 7472 9868 7524 9920
rect 10968 9868 11020 9920
rect 15200 10072 15252 10124
rect 15660 10072 15712 10124
rect 17500 10072 17552 10124
rect 18604 10072 18656 10124
rect 19800 10072 19852 10124
rect 15844 10004 15896 10056
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 17040 10004 17092 10013
rect 18328 10004 18380 10056
rect 17408 9936 17460 9988
rect 18052 9936 18104 9988
rect 13636 9868 13688 9920
rect 4414 9766 4466 9818
rect 4478 9766 4530 9818
rect 4542 9766 4594 9818
rect 4606 9766 4658 9818
rect 11278 9766 11330 9818
rect 11342 9766 11394 9818
rect 11406 9766 11458 9818
rect 11470 9766 11522 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 18270 9766 18322 9818
rect 18334 9766 18386 9818
rect 2412 9664 2464 9716
rect 2688 9664 2740 9716
rect 3148 9664 3200 9716
rect 4068 9664 4120 9716
rect 7472 9664 7524 9716
rect 7840 9664 7892 9716
rect 10232 9707 10284 9716
rect 1860 9528 1912 9580
rect 2872 9639 2924 9648
rect 2872 9605 2881 9639
rect 2881 9605 2915 9639
rect 2915 9605 2924 9639
rect 2872 9596 2924 9605
rect 4896 9596 4948 9648
rect 4988 9596 5040 9648
rect 5448 9596 5500 9648
rect 5632 9596 5684 9648
rect 6644 9596 6696 9648
rect 6920 9596 6972 9648
rect 1400 9460 1452 9512
rect 2688 9460 2740 9512
rect 3608 9528 3660 9580
rect 7288 9528 7340 9580
rect 7564 9596 7616 9648
rect 10232 9673 10241 9707
rect 10241 9673 10275 9707
rect 10275 9673 10284 9707
rect 10232 9664 10284 9673
rect 10508 9707 10560 9716
rect 10508 9673 10517 9707
rect 10517 9673 10551 9707
rect 10551 9673 10560 9707
rect 10508 9664 10560 9673
rect 12348 9664 12400 9716
rect 12624 9664 12676 9716
rect 12808 9664 12860 9716
rect 7748 9528 7800 9580
rect 8208 9528 8260 9580
rect 8484 9528 8536 9580
rect 3700 9460 3752 9512
rect 4252 9460 4304 9512
rect 4436 9460 4488 9512
rect 6000 9460 6052 9512
rect 10784 9528 10836 9580
rect 16764 9596 16816 9648
rect 17132 9664 17184 9716
rect 20076 9664 20128 9716
rect 19616 9596 19668 9648
rect 2964 9324 3016 9376
rect 7104 9392 7156 9444
rect 7472 9392 7524 9444
rect 9864 9392 9916 9444
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 4620 9324 4672 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 8300 9324 8352 9376
rect 10876 9460 10928 9512
rect 12348 9460 12400 9512
rect 15660 9528 15712 9580
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 17040 9528 17092 9580
rect 19708 9571 19760 9580
rect 19708 9537 19717 9571
rect 19717 9537 19751 9571
rect 19751 9537 19760 9571
rect 19708 9528 19760 9537
rect 10232 9324 10284 9376
rect 10968 9324 11020 9376
rect 12532 9392 12584 9444
rect 12716 9435 12768 9444
rect 12716 9401 12750 9435
rect 12750 9401 12768 9435
rect 12716 9392 12768 9401
rect 13452 9392 13504 9444
rect 14188 9392 14240 9444
rect 15108 9392 15160 9444
rect 20352 9460 20404 9512
rect 11704 9367 11756 9376
rect 11704 9333 11713 9367
rect 11713 9333 11747 9367
rect 11747 9333 11756 9367
rect 11704 9324 11756 9333
rect 13820 9367 13872 9376
rect 13820 9333 13829 9367
rect 13829 9333 13863 9367
rect 13863 9333 13872 9367
rect 13820 9324 13872 9333
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 15292 9324 15344 9376
rect 15476 9324 15528 9376
rect 17316 9367 17368 9376
rect 17316 9333 17325 9367
rect 17325 9333 17359 9367
rect 17359 9333 17368 9367
rect 17316 9324 17368 9333
rect 17500 9324 17552 9376
rect 7846 9222 7898 9274
rect 7910 9222 7962 9274
rect 7974 9222 8026 9274
rect 8038 9222 8090 9274
rect 14710 9222 14762 9274
rect 14774 9222 14826 9274
rect 14838 9222 14890 9274
rect 14902 9222 14954 9274
rect 2320 9120 2372 9172
rect 2504 9120 2556 9172
rect 3056 9163 3108 9172
rect 3056 9129 3065 9163
rect 3065 9129 3099 9163
rect 3099 9129 3108 9163
rect 3056 9120 3108 9129
rect 4804 9120 4856 9172
rect 3424 9052 3476 9104
rect 8300 9052 8352 9104
rect 4620 8984 4672 9036
rect 6184 9027 6236 9036
rect 6184 8993 6193 9027
rect 6193 8993 6227 9027
rect 6227 8993 6236 9027
rect 6184 8984 6236 8993
rect 6736 8984 6788 9036
rect 8208 8984 8260 9036
rect 8576 9052 8628 9104
rect 2596 8916 2648 8968
rect 2688 8959 2740 8968
rect 2688 8925 2697 8959
rect 2697 8925 2731 8959
rect 2731 8925 2740 8959
rect 4896 8959 4948 8968
rect 2688 8916 2740 8925
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5172 8916 5224 8968
rect 8116 8916 8168 8968
rect 9036 8916 9088 8968
rect 4436 8848 4488 8900
rect 6184 8848 6236 8900
rect 7564 8891 7616 8900
rect 7564 8857 7573 8891
rect 7573 8857 7607 8891
rect 7607 8857 7616 8891
rect 7564 8848 7616 8857
rect 7748 8848 7800 8900
rect 11612 9052 11664 9104
rect 12716 9120 12768 9172
rect 14556 9120 14608 9172
rect 15292 9120 15344 9172
rect 15660 9120 15712 9172
rect 16028 9120 16080 9172
rect 19800 9163 19852 9172
rect 19800 9129 19809 9163
rect 19809 9129 19843 9163
rect 19843 9129 19852 9163
rect 19800 9120 19852 9129
rect 19984 9120 20036 9172
rect 14004 9052 14056 9104
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10968 8984 11020 9036
rect 12624 8984 12676 9036
rect 13176 8984 13228 9036
rect 13820 8984 13872 9036
rect 15752 9052 15804 9104
rect 17316 9095 17368 9104
rect 17316 9061 17325 9095
rect 17325 9061 17359 9095
rect 17359 9061 17368 9095
rect 17316 9052 17368 9061
rect 18604 9052 18656 9104
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 4068 8780 4120 8832
rect 9864 8848 9916 8900
rect 13912 8916 13964 8968
rect 14832 8959 14884 8968
rect 14832 8925 14841 8959
rect 14841 8925 14875 8959
rect 14875 8925 14884 8959
rect 14832 8916 14884 8925
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 17316 8916 17368 8968
rect 19064 8984 19116 9036
rect 19616 8984 19668 9036
rect 17592 8916 17644 8968
rect 10508 8848 10560 8900
rect 11704 8848 11756 8900
rect 12072 8848 12124 8900
rect 12348 8848 12400 8900
rect 8208 8780 8260 8832
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 10784 8780 10836 8832
rect 10876 8780 10928 8832
rect 16948 8823 17000 8832
rect 16948 8789 16957 8823
rect 16957 8789 16991 8823
rect 16991 8789 17000 8823
rect 16948 8780 17000 8789
rect 18788 8780 18840 8832
rect 4414 8678 4466 8730
rect 4478 8678 4530 8730
rect 4542 8678 4594 8730
rect 4606 8678 4658 8730
rect 11278 8678 11330 8730
rect 11342 8678 11394 8730
rect 11406 8678 11458 8730
rect 11470 8678 11522 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 18270 8678 18322 8730
rect 18334 8678 18386 8730
rect 2044 8576 2096 8628
rect 3240 8576 3292 8628
rect 4160 8619 4212 8628
rect 4160 8585 4169 8619
rect 4169 8585 4203 8619
rect 4203 8585 4212 8619
rect 4160 8576 4212 8585
rect 5080 8576 5132 8628
rect 6644 8576 6696 8628
rect 7196 8576 7248 8628
rect 4068 8508 4120 8560
rect 9680 8576 9732 8628
rect 9864 8619 9916 8628
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 12164 8576 12216 8628
rect 12440 8576 12492 8628
rect 17960 8576 18012 8628
rect 19156 8576 19208 8628
rect 14832 8551 14884 8560
rect 3700 8440 3752 8492
rect 6000 8440 6052 8492
rect 6828 8440 6880 8492
rect 7564 8440 7616 8492
rect 8116 8440 8168 8492
rect 12808 8440 12860 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14832 8517 14841 8551
rect 14841 8517 14875 8551
rect 14875 8517 14884 8551
rect 14832 8508 14884 8517
rect 15108 8508 15160 8560
rect 13176 8440 13228 8492
rect 1676 8372 1728 8424
rect 5448 8372 5500 8424
rect 6368 8372 6420 8424
rect 8484 8415 8536 8424
rect 2688 8304 2740 8356
rect 5080 8304 5132 8356
rect 3240 8279 3292 8288
rect 3240 8245 3249 8279
rect 3249 8245 3283 8279
rect 3283 8245 3292 8279
rect 3240 8236 3292 8245
rect 5448 8236 5500 8288
rect 5540 8279 5592 8288
rect 5540 8245 5549 8279
rect 5549 8245 5583 8279
rect 5583 8245 5592 8279
rect 6092 8304 6144 8356
rect 6552 8304 6604 8356
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 7564 8304 7616 8356
rect 10600 8372 10652 8424
rect 12624 8372 12676 8424
rect 9128 8304 9180 8356
rect 9312 8304 9364 8356
rect 10508 8304 10560 8356
rect 12716 8304 12768 8356
rect 13176 8304 13228 8356
rect 14004 8372 14056 8424
rect 16948 8508 17000 8560
rect 17040 8508 17092 8560
rect 18512 8508 18564 8560
rect 17684 8440 17736 8492
rect 19800 8440 19852 8492
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 16120 8372 16172 8424
rect 13820 8304 13872 8356
rect 15568 8347 15620 8356
rect 15568 8313 15577 8347
rect 15577 8313 15611 8347
rect 15611 8313 15620 8347
rect 15568 8304 15620 8313
rect 17224 8347 17276 8356
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 6276 8279 6328 8288
rect 5540 8236 5592 8245
rect 6276 8245 6285 8279
rect 6285 8245 6319 8279
rect 6319 8245 6328 8279
rect 6276 8236 6328 8245
rect 6644 8236 6696 8288
rect 11980 8236 12032 8288
rect 12256 8236 12308 8288
rect 13544 8236 13596 8288
rect 18972 8304 19024 8356
rect 19340 8347 19392 8356
rect 19340 8313 19349 8347
rect 19349 8313 19383 8347
rect 19383 8313 19392 8347
rect 19340 8304 19392 8313
rect 20904 8304 20956 8356
rect 19432 8279 19484 8288
rect 19432 8245 19441 8279
rect 19441 8245 19475 8279
rect 19475 8245 19484 8279
rect 19984 8279 20036 8288
rect 19432 8236 19484 8245
rect 19984 8245 19993 8279
rect 19993 8245 20027 8279
rect 20027 8245 20036 8279
rect 19984 8236 20036 8245
rect 20444 8279 20496 8288
rect 20444 8245 20453 8279
rect 20453 8245 20487 8279
rect 20487 8245 20496 8279
rect 20444 8236 20496 8245
rect 7846 8134 7898 8186
rect 7910 8134 7962 8186
rect 7974 8134 8026 8186
rect 8038 8134 8090 8186
rect 14710 8134 14762 8186
rect 14774 8134 14826 8186
rect 14838 8134 14890 8186
rect 14902 8134 14954 8186
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 3976 8032 4028 8084
rect 4252 8032 4304 8084
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 6276 8032 6328 8084
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 7564 8032 7616 8084
rect 8300 8032 8352 8084
rect 8576 8032 8628 8084
rect 10508 8032 10560 8084
rect 12072 8032 12124 8084
rect 13084 8032 13136 8084
rect 13452 8032 13504 8084
rect 3056 7964 3108 8016
rect 3424 8007 3476 8016
rect 3424 7973 3433 8007
rect 3433 7973 3467 8007
rect 3467 7973 3476 8007
rect 3424 7964 3476 7973
rect 3516 7964 3568 8016
rect 8852 7964 8904 8016
rect 10876 7964 10928 8016
rect 12348 7964 12400 8016
rect 3976 7896 4028 7948
rect 4160 7896 4212 7948
rect 5080 7896 5132 7948
rect 6644 7896 6696 7948
rect 6736 7896 6788 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2688 7828 2740 7880
rect 3700 7828 3752 7880
rect 3792 7828 3844 7880
rect 5356 7828 5408 7880
rect 5540 7828 5592 7880
rect 5816 7828 5868 7880
rect 3240 7760 3292 7812
rect 3516 7692 3568 7744
rect 5172 7760 5224 7812
rect 6552 7828 6604 7880
rect 7104 7896 7156 7948
rect 9680 7896 9732 7948
rect 10416 7896 10468 7948
rect 11152 7896 11204 7948
rect 11612 7896 11664 7948
rect 12532 7964 12584 8016
rect 13912 8032 13964 8084
rect 14556 8075 14608 8084
rect 14556 8041 14565 8075
rect 14565 8041 14599 8075
rect 14599 8041 14608 8075
rect 14556 8032 14608 8041
rect 19064 8075 19116 8084
rect 19064 8041 19073 8075
rect 19073 8041 19107 8075
rect 19107 8041 19116 8075
rect 19064 8032 19116 8041
rect 20444 8032 20496 8084
rect 20904 8075 20956 8084
rect 20904 8041 20913 8075
rect 20913 8041 20947 8075
rect 20947 8041 20956 8075
rect 20904 8032 20956 8041
rect 14096 7964 14148 8016
rect 16028 8007 16080 8016
rect 16028 7973 16062 8007
rect 16062 7973 16080 8007
rect 16028 7964 16080 7973
rect 17684 7964 17736 8016
rect 20536 7964 20588 8016
rect 12808 7896 12860 7948
rect 13544 7896 13596 7948
rect 13912 7896 13964 7948
rect 9128 7871 9180 7880
rect 6368 7803 6420 7812
rect 6368 7769 6377 7803
rect 6377 7769 6411 7803
rect 6411 7769 6420 7803
rect 6368 7760 6420 7769
rect 9128 7837 9137 7871
rect 9137 7837 9171 7871
rect 9171 7837 9180 7871
rect 9128 7828 9180 7837
rect 10048 7760 10100 7812
rect 9036 7692 9088 7744
rect 11796 7828 11848 7880
rect 12164 7828 12216 7880
rect 12716 7828 12768 7880
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 14004 7871 14056 7880
rect 14004 7837 14013 7871
rect 14013 7837 14047 7871
rect 14047 7837 14056 7871
rect 14004 7828 14056 7837
rect 14096 7828 14148 7880
rect 15200 7896 15252 7948
rect 16304 7896 16356 7948
rect 19616 7896 19668 7948
rect 15292 7828 15344 7880
rect 15752 7871 15804 7880
rect 15752 7837 15761 7871
rect 15761 7837 15795 7871
rect 15795 7837 15804 7871
rect 15752 7828 15804 7837
rect 17592 7828 17644 7880
rect 19156 7828 19208 7880
rect 20720 7896 20772 7948
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 12808 7692 12860 7744
rect 15752 7692 15804 7744
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 17868 7692 17920 7744
rect 20444 7692 20496 7744
rect 4414 7590 4466 7642
rect 4478 7590 4530 7642
rect 4542 7590 4594 7642
rect 4606 7590 4658 7642
rect 11278 7590 11330 7642
rect 11342 7590 11394 7642
rect 11406 7590 11458 7642
rect 11470 7590 11522 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 18270 7590 18322 7642
rect 18334 7590 18386 7642
rect 2136 7531 2188 7540
rect 2136 7497 2145 7531
rect 2145 7497 2179 7531
rect 2179 7497 2188 7531
rect 2136 7488 2188 7497
rect 3056 7488 3108 7540
rect 4160 7488 4212 7540
rect 5724 7488 5776 7540
rect 6644 7488 6696 7540
rect 8852 7488 8904 7540
rect 9128 7488 9180 7540
rect 10140 7531 10192 7540
rect 3608 7420 3660 7472
rect 3792 7420 3844 7472
rect 2780 7395 2832 7404
rect 2780 7361 2789 7395
rect 2789 7361 2823 7395
rect 2823 7361 2832 7395
rect 2780 7352 2832 7361
rect 3056 7352 3108 7404
rect 3976 7352 4028 7404
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 5356 7352 5408 7404
rect 5632 7352 5684 7404
rect 7012 7352 7064 7404
rect 7104 7352 7156 7404
rect 8024 7352 8076 7404
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 14280 7488 14332 7540
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 19432 7488 19484 7540
rect 19800 7488 19852 7540
rect 20168 7488 20220 7540
rect 20352 7488 20404 7540
rect 14648 7420 14700 7472
rect 11152 7352 11204 7404
rect 12624 7352 12676 7404
rect 1952 7216 2004 7268
rect 3792 7216 3844 7268
rect 8208 7284 8260 7336
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 9036 7284 9088 7336
rect 9312 7284 9364 7336
rect 10232 7284 10284 7336
rect 12440 7284 12492 7336
rect 12808 7327 12860 7336
rect 12808 7293 12817 7327
rect 12817 7293 12851 7327
rect 12851 7293 12860 7327
rect 12808 7284 12860 7293
rect 12900 7284 12952 7336
rect 13176 7284 13228 7336
rect 19064 7352 19116 7404
rect 20536 7352 20588 7404
rect 4804 7148 4856 7200
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 6644 7148 6696 7200
rect 6920 7191 6972 7200
rect 6920 7157 6929 7191
rect 6929 7157 6963 7191
rect 6963 7157 6972 7191
rect 6920 7148 6972 7157
rect 7288 7191 7340 7200
rect 7288 7157 7297 7191
rect 7297 7157 7331 7191
rect 7331 7157 7340 7191
rect 7288 7148 7340 7157
rect 8300 7216 8352 7268
rect 11060 7216 11112 7268
rect 12716 7216 12768 7268
rect 13912 7259 13964 7268
rect 13912 7225 13946 7259
rect 13946 7225 13964 7259
rect 13912 7216 13964 7225
rect 14004 7216 14056 7268
rect 14832 7216 14884 7268
rect 15200 7216 15252 7268
rect 15844 7216 15896 7268
rect 9956 7148 10008 7200
rect 10508 7191 10560 7200
rect 10508 7157 10517 7191
rect 10517 7157 10551 7191
rect 10551 7157 10560 7191
rect 10508 7148 10560 7157
rect 11704 7148 11756 7200
rect 12532 7148 12584 7200
rect 12808 7148 12860 7200
rect 15108 7148 15160 7200
rect 15660 7191 15712 7200
rect 15660 7157 15669 7191
rect 15669 7157 15703 7191
rect 15703 7157 15712 7191
rect 15660 7148 15712 7157
rect 16672 7216 16724 7268
rect 19432 7284 19484 7336
rect 20720 7327 20772 7336
rect 20720 7293 20729 7327
rect 20729 7293 20763 7327
rect 20763 7293 20772 7327
rect 20720 7284 20772 7293
rect 18788 7216 18840 7268
rect 19524 7216 19576 7268
rect 17592 7148 17644 7200
rect 20076 7191 20128 7200
rect 20076 7157 20085 7191
rect 20085 7157 20119 7191
rect 20119 7157 20128 7191
rect 20076 7148 20128 7157
rect 20168 7191 20220 7200
rect 20168 7157 20177 7191
rect 20177 7157 20211 7191
rect 20211 7157 20220 7191
rect 20168 7148 20220 7157
rect 21088 7148 21140 7200
rect 7846 7046 7898 7098
rect 7910 7046 7962 7098
rect 7974 7046 8026 7098
rect 8038 7046 8090 7098
rect 14710 7046 14762 7098
rect 14774 7046 14826 7098
rect 14838 7046 14890 7098
rect 14902 7046 14954 7098
rect 3056 6987 3108 6996
rect 3056 6953 3065 6987
rect 3065 6953 3099 6987
rect 3099 6953 3108 6987
rect 3056 6944 3108 6953
rect 6920 6944 6972 6996
rect 10508 6944 10560 6996
rect 2412 6876 2464 6928
rect 5356 6876 5408 6928
rect 6368 6876 6420 6928
rect 9036 6876 9088 6928
rect 1676 6851 1728 6860
rect 1676 6817 1685 6851
rect 1685 6817 1719 6851
rect 1719 6817 1728 6851
rect 1676 6808 1728 6817
rect 2228 6808 2280 6860
rect 6000 6808 6052 6860
rect 6276 6808 6328 6860
rect 10232 6919 10284 6928
rect 10232 6885 10241 6919
rect 10241 6885 10275 6919
rect 10275 6885 10284 6919
rect 12256 6944 12308 6996
rect 17408 6944 17460 6996
rect 10232 6876 10284 6885
rect 13820 6876 13872 6928
rect 4160 6740 4212 6792
rect 6920 6740 6972 6792
rect 7196 6740 7248 6792
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 8300 6740 8352 6792
rect 11152 6808 11204 6860
rect 11796 6808 11848 6860
rect 7012 6672 7064 6724
rect 10140 6672 10192 6724
rect 5448 6604 5500 6656
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 9772 6604 9824 6656
rect 11060 6783 11112 6792
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 15476 6876 15528 6928
rect 19984 6876 20036 6928
rect 14648 6808 14700 6817
rect 15752 6808 15804 6860
rect 16396 6808 16448 6860
rect 18972 6851 19024 6860
rect 18972 6817 18981 6851
rect 18981 6817 19015 6851
rect 19015 6817 19024 6851
rect 18972 6808 19024 6817
rect 13636 6783 13688 6792
rect 10508 6672 10560 6724
rect 12624 6604 12676 6656
rect 12900 6604 12952 6656
rect 13636 6749 13645 6783
rect 13645 6749 13679 6783
rect 13679 6749 13688 6783
rect 13636 6740 13688 6749
rect 13912 6740 13964 6792
rect 14556 6740 14608 6792
rect 14740 6783 14792 6792
rect 14740 6749 14749 6783
rect 14749 6749 14783 6783
rect 14783 6749 14792 6783
rect 14740 6740 14792 6749
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 16948 6740 17000 6792
rect 14004 6672 14056 6724
rect 15660 6672 15712 6724
rect 15844 6715 15896 6724
rect 15844 6681 15853 6715
rect 15853 6681 15887 6715
rect 15887 6681 15896 6715
rect 15844 6672 15896 6681
rect 16120 6715 16172 6724
rect 16120 6681 16129 6715
rect 16129 6681 16163 6715
rect 16163 6681 16172 6715
rect 16120 6672 16172 6681
rect 15752 6604 15804 6656
rect 17224 6672 17276 6724
rect 17684 6604 17736 6656
rect 17868 6740 17920 6792
rect 19064 6783 19116 6792
rect 19064 6749 19073 6783
rect 19073 6749 19107 6783
rect 19107 6749 19116 6783
rect 19984 6783 20036 6792
rect 19064 6740 19116 6749
rect 19984 6749 19993 6783
rect 19993 6749 20027 6783
rect 20027 6749 20036 6783
rect 19984 6740 20036 6749
rect 20536 6740 20588 6792
rect 19340 6672 19392 6724
rect 19524 6715 19576 6724
rect 19524 6681 19533 6715
rect 19533 6681 19567 6715
rect 19567 6681 19576 6715
rect 19524 6672 19576 6681
rect 4414 6502 4466 6554
rect 4478 6502 4530 6554
rect 4542 6502 4594 6554
rect 4606 6502 4658 6554
rect 11278 6502 11330 6554
rect 11342 6502 11394 6554
rect 11406 6502 11458 6554
rect 11470 6502 11522 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 18270 6502 18322 6554
rect 18334 6502 18386 6554
rect 2780 6400 2832 6452
rect 4068 6400 4120 6452
rect 4804 6400 4856 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7196 6400 7248 6452
rect 8852 6400 8904 6452
rect 11888 6400 11940 6452
rect 12348 6400 12400 6452
rect 12624 6400 12676 6452
rect 16396 6400 16448 6452
rect 18696 6400 18748 6452
rect 20168 6400 20220 6452
rect 4160 6332 4212 6384
rect 6736 6332 6788 6384
rect 11152 6375 11204 6384
rect 1676 6264 1728 6316
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 2228 6196 2280 6248
rect 3608 6196 3660 6248
rect 5172 6264 5224 6316
rect 5448 6307 5500 6316
rect 5448 6273 5457 6307
rect 5457 6273 5491 6307
rect 5491 6273 5500 6307
rect 5448 6264 5500 6273
rect 7288 6264 7340 6316
rect 11152 6341 11161 6375
rect 11161 6341 11195 6375
rect 11195 6341 11204 6375
rect 11152 6332 11204 6341
rect 11336 6332 11388 6384
rect 11980 6332 12032 6384
rect 15660 6332 15712 6384
rect 19800 6332 19852 6384
rect 7564 6264 7616 6316
rect 9404 6264 9456 6316
rect 3056 6128 3108 6180
rect 5080 6128 5132 6180
rect 12072 6264 12124 6316
rect 16120 6264 16172 6316
rect 17132 6264 17184 6316
rect 17592 6264 17644 6316
rect 17868 6264 17920 6316
rect 20444 6264 20496 6316
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 3884 6060 3936 6112
rect 5264 6103 5316 6112
rect 5264 6069 5273 6103
rect 5273 6069 5307 6103
rect 5307 6069 5316 6103
rect 5264 6060 5316 6069
rect 8208 6128 8260 6180
rect 8300 6128 8352 6180
rect 8484 6128 8536 6180
rect 9404 6128 9456 6180
rect 9220 6060 9272 6112
rect 11060 6196 11112 6248
rect 12440 6239 12492 6248
rect 12440 6205 12449 6239
rect 12449 6205 12483 6239
rect 12483 6205 12492 6239
rect 12440 6196 12492 6205
rect 12716 6239 12768 6248
rect 12716 6205 12750 6239
rect 12750 6205 12768 6239
rect 12716 6196 12768 6205
rect 14280 6196 14332 6248
rect 12256 6128 12308 6180
rect 17224 6196 17276 6248
rect 19432 6239 19484 6248
rect 19432 6205 19441 6239
rect 19441 6205 19475 6239
rect 19475 6205 19484 6239
rect 19432 6196 19484 6205
rect 20628 6196 20680 6248
rect 10600 6060 10652 6112
rect 15108 6128 15160 6180
rect 12992 6060 13044 6112
rect 14556 6060 14608 6112
rect 18788 6128 18840 6180
rect 19248 6128 19300 6180
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 18328 6060 18380 6112
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 18696 6060 18748 6112
rect 19616 6060 19668 6112
rect 7846 5958 7898 6010
rect 7910 5958 7962 6010
rect 7974 5958 8026 6010
rect 8038 5958 8090 6010
rect 14710 5958 14762 6010
rect 14774 5958 14826 6010
rect 14838 5958 14890 6010
rect 14902 5958 14954 6010
rect 1952 5899 2004 5908
rect 1952 5865 1961 5899
rect 1961 5865 1995 5899
rect 1995 5865 2004 5899
rect 1952 5856 2004 5865
rect 3792 5856 3844 5908
rect 3976 5856 4028 5908
rect 4068 5788 4120 5840
rect 5264 5856 5316 5908
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 6460 5856 6512 5908
rect 6920 5788 6972 5840
rect 7104 5831 7156 5840
rect 7104 5797 7138 5831
rect 7138 5797 7156 5831
rect 7104 5788 7156 5797
rect 8852 5856 8904 5908
rect 10600 5856 10652 5908
rect 13084 5856 13136 5908
rect 3976 5720 4028 5772
rect 6736 5720 6788 5772
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 12164 5788 12216 5840
rect 12440 5788 12492 5840
rect 10048 5720 10100 5729
rect 12072 5720 12124 5772
rect 12900 5788 12952 5840
rect 13452 5788 13504 5840
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3056 5652 3108 5704
rect 4068 5695 4120 5704
rect 4068 5661 4084 5695
rect 4084 5661 4118 5695
rect 4118 5661 4120 5695
rect 4068 5652 4120 5661
rect 6000 5652 6052 5704
rect 6644 5652 6696 5704
rect 9036 5695 9088 5704
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 9956 5584 10008 5636
rect 10232 5695 10284 5704
rect 10232 5661 10241 5695
rect 10241 5661 10275 5695
rect 10275 5661 10284 5695
rect 10232 5652 10284 5661
rect 11244 5652 11296 5704
rect 11888 5652 11940 5704
rect 11980 5652 12032 5704
rect 12992 5763 13044 5772
rect 12992 5729 13026 5763
rect 13026 5729 13044 5763
rect 12992 5720 13044 5729
rect 14004 5720 14056 5772
rect 16120 5788 16172 5840
rect 17592 5856 17644 5908
rect 17868 5831 17920 5840
rect 17868 5797 17902 5831
rect 17902 5797 17920 5831
rect 17868 5788 17920 5797
rect 18512 5856 18564 5908
rect 18144 5720 18196 5772
rect 19156 5720 19208 5772
rect 13820 5652 13872 5704
rect 15660 5652 15712 5704
rect 15844 5652 15896 5704
rect 17592 5695 17644 5704
rect 10876 5584 10928 5636
rect 5540 5516 5592 5568
rect 8300 5516 8352 5568
rect 9404 5516 9456 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 11980 5516 12032 5568
rect 12440 5516 12492 5568
rect 12716 5584 12768 5636
rect 14280 5584 14332 5636
rect 13636 5516 13688 5568
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19708 5695 19760 5704
rect 19708 5661 19717 5695
rect 19717 5661 19751 5695
rect 19751 5661 19760 5695
rect 19708 5652 19760 5661
rect 19248 5584 19300 5636
rect 18972 5559 19024 5568
rect 18972 5525 18981 5559
rect 18981 5525 19015 5559
rect 19015 5525 19024 5559
rect 18972 5516 19024 5525
rect 20996 5516 21048 5568
rect 4414 5414 4466 5466
rect 4478 5414 4530 5466
rect 4542 5414 4594 5466
rect 4606 5414 4658 5466
rect 11278 5414 11330 5466
rect 11342 5414 11394 5466
rect 11406 5414 11458 5466
rect 11470 5414 11522 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 18270 5414 18322 5466
rect 18334 5414 18386 5466
rect 2412 5312 2464 5364
rect 4068 5312 4120 5364
rect 6092 5312 6144 5364
rect 7656 5312 7708 5364
rect 9036 5312 9088 5364
rect 12440 5312 12492 5364
rect 6736 5244 6788 5296
rect 7380 5244 7432 5296
rect 2228 5176 2280 5228
rect 4988 5176 5040 5228
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 6552 5176 6604 5228
rect 7104 5176 7156 5228
rect 7656 5176 7708 5228
rect 5448 5108 5500 5160
rect 5724 5108 5776 5160
rect 10600 5244 10652 5296
rect 8300 5176 8352 5228
rect 11796 5244 11848 5296
rect 12072 5244 12124 5296
rect 12716 5244 12768 5296
rect 17684 5312 17736 5364
rect 17868 5312 17920 5364
rect 17960 5312 18012 5364
rect 20536 5312 20588 5364
rect 13820 5244 13872 5296
rect 14464 5244 14516 5296
rect 19616 5244 19668 5296
rect 12992 5176 13044 5228
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 8208 5108 8260 5160
rect 9680 5108 9732 5160
rect 9956 5108 10008 5160
rect 13176 5108 13228 5160
rect 13544 5108 13596 5160
rect 2320 4972 2372 5024
rect 2964 5040 3016 5092
rect 3976 5040 4028 5092
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 4896 5015 4948 5024
rect 2504 4972 2556 4981
rect 4896 4981 4905 5015
rect 4905 4981 4939 5015
rect 4939 4981 4948 5015
rect 4896 4972 4948 4981
rect 6920 4972 6972 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 9680 4972 9732 5024
rect 10140 4972 10192 5024
rect 10692 4972 10744 5024
rect 10876 4972 10928 5024
rect 11888 5040 11940 5092
rect 13912 5040 13964 5092
rect 15844 5108 15896 5160
rect 18972 5176 19024 5228
rect 17960 5108 18012 5160
rect 18512 5151 18564 5160
rect 18512 5117 18521 5151
rect 18521 5117 18555 5151
rect 18555 5117 18564 5151
rect 18512 5108 18564 5117
rect 17592 5040 17644 5092
rect 18328 5040 18380 5092
rect 18696 5108 18748 5160
rect 19340 5108 19392 5160
rect 19524 5108 19576 5160
rect 21180 5108 21232 5160
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 12992 4972 13044 5024
rect 13360 4972 13412 5024
rect 14004 5015 14056 5024
rect 14004 4981 14013 5015
rect 14013 4981 14047 5015
rect 14047 4981 14056 5015
rect 14004 4972 14056 4981
rect 14280 4972 14332 5024
rect 19800 5040 19852 5092
rect 18788 4972 18840 5024
rect 7846 4870 7898 4922
rect 7910 4870 7962 4922
rect 7974 4870 8026 4922
rect 8038 4870 8090 4922
rect 14710 4870 14762 4922
rect 14774 4870 14826 4922
rect 14838 4870 14890 4922
rect 14902 4870 14954 4922
rect 3700 4811 3752 4820
rect 3700 4777 3709 4811
rect 3709 4777 3743 4811
rect 3743 4777 3752 4811
rect 3700 4768 3752 4777
rect 4068 4768 4120 4820
rect 2136 4632 2188 4684
rect 3240 4700 3292 4752
rect 4160 4700 4212 4752
rect 3148 4632 3200 4684
rect 5540 4700 5592 4752
rect 7472 4768 7524 4820
rect 8760 4768 8812 4820
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 10600 4768 10652 4820
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 11520 4700 11572 4752
rect 15200 4768 15252 4820
rect 19156 4768 19208 4820
rect 19800 4811 19852 4820
rect 19800 4777 19809 4811
rect 19809 4777 19843 4811
rect 19843 4777 19852 4811
rect 19800 4768 19852 4777
rect 13636 4743 13688 4752
rect 13636 4709 13670 4743
rect 13670 4709 13688 4743
rect 13636 4700 13688 4709
rect 17684 4700 17736 4752
rect 19340 4700 19392 4752
rect 5172 4632 5224 4684
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 9864 4632 9916 4684
rect 10048 4675 10100 4684
rect 10048 4641 10057 4675
rect 10057 4641 10091 4675
rect 10091 4641 10100 4675
rect 10048 4632 10100 4641
rect 11796 4632 11848 4684
rect 3424 4564 3476 4616
rect 4160 4564 4212 4616
rect 6276 4564 6328 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7472 4564 7524 4616
rect 8668 4607 8720 4616
rect 5356 4496 5408 4548
rect 6368 4496 6420 4548
rect 6828 4496 6880 4548
rect 7564 4496 7616 4548
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 10140 4607 10192 4616
rect 7932 4496 7984 4548
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 11060 4564 11112 4616
rect 12164 4564 12216 4616
rect 12716 4564 12768 4616
rect 9772 4496 9824 4548
rect 15292 4632 15344 4684
rect 17592 4632 17644 4684
rect 18512 4632 18564 4684
rect 18972 4632 19024 4684
rect 19432 4632 19484 4684
rect 19892 4632 19944 4684
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 16856 4607 16908 4616
rect 16856 4573 16865 4607
rect 16865 4573 16899 4607
rect 16899 4573 16908 4607
rect 16856 4564 16908 4573
rect 17868 4607 17920 4616
rect 17868 4573 17877 4607
rect 17877 4573 17911 4607
rect 17911 4573 17920 4607
rect 17868 4564 17920 4573
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 18328 4564 18380 4616
rect 5264 4428 5316 4480
rect 9680 4428 9732 4480
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 12900 4428 12952 4480
rect 13636 4428 13688 4480
rect 14556 4428 14608 4480
rect 16304 4428 16356 4480
rect 17408 4471 17460 4480
rect 17408 4437 17417 4471
rect 17417 4437 17451 4471
rect 17451 4437 17460 4471
rect 17408 4428 17460 4437
rect 17960 4428 18012 4480
rect 19524 4428 19576 4480
rect 4414 4326 4466 4378
rect 4478 4326 4530 4378
rect 4542 4326 4594 4378
rect 4606 4326 4658 4378
rect 11278 4326 11330 4378
rect 11342 4326 11394 4378
rect 11406 4326 11458 4378
rect 11470 4326 11522 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 18270 4326 18322 4378
rect 18334 4326 18386 4378
rect 2136 4224 2188 4276
rect 3148 4224 3200 4276
rect 3608 4224 3660 4276
rect 7656 4224 7708 4276
rect 10232 4224 10284 4276
rect 11612 4224 11664 4276
rect 12532 4224 12584 4276
rect 16856 4267 16908 4276
rect 3700 4156 3752 4208
rect 6276 4156 6328 4208
rect 4068 4131 4120 4140
rect 4068 4097 4077 4131
rect 4077 4097 4111 4131
rect 4111 4097 4120 4131
rect 4068 4088 4120 4097
rect 4896 4088 4948 4140
rect 5264 4088 5316 4140
rect 6644 4088 6696 4140
rect 6920 4088 6972 4140
rect 10048 4156 10100 4208
rect 3056 4020 3108 4072
rect 7932 4063 7984 4072
rect 1952 3952 2004 4004
rect 7932 4029 7966 4063
rect 7966 4029 7984 4063
rect 7932 4020 7984 4029
rect 8208 4020 8260 4072
rect 9772 4088 9824 4140
rect 11888 4131 11940 4140
rect 9404 4063 9456 4072
rect 9404 4029 9413 4063
rect 9413 4029 9447 4063
rect 9447 4029 9456 4063
rect 9404 4020 9456 4029
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 11060 4020 11112 4072
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 5356 3884 5408 3936
rect 8760 3952 8812 4004
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12440 4156 12492 4208
rect 12900 4131 12952 4140
rect 12900 4097 12909 4131
rect 12909 4097 12943 4131
rect 12943 4097 12952 4131
rect 12900 4088 12952 4097
rect 13360 4020 13412 4072
rect 16856 4233 16865 4267
rect 16865 4233 16899 4267
rect 16899 4233 16908 4267
rect 16856 4224 16908 4233
rect 17592 4224 17644 4276
rect 19524 4224 19576 4276
rect 20536 4156 20588 4208
rect 16672 4088 16724 4140
rect 19340 4088 19392 4140
rect 19800 4088 19852 4140
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 17316 4020 17368 4072
rect 17592 4020 17644 4072
rect 17960 4020 18012 4072
rect 20536 4020 20588 4072
rect 11520 3952 11572 4004
rect 5632 3884 5684 3936
rect 10048 3884 10100 3936
rect 11336 3884 11388 3936
rect 11612 3927 11664 3936
rect 11612 3893 11621 3927
rect 11621 3893 11655 3927
rect 11655 3893 11664 3927
rect 11612 3884 11664 3893
rect 12440 3927 12492 3936
rect 12440 3893 12449 3927
rect 12449 3893 12483 3927
rect 12483 3893 12492 3927
rect 14372 3952 14424 4004
rect 16948 3952 17000 4004
rect 18144 3952 18196 4004
rect 18604 3952 18656 4004
rect 12440 3884 12492 3893
rect 14556 3884 14608 3936
rect 15108 3927 15160 3936
rect 15108 3893 15117 3927
rect 15117 3893 15151 3927
rect 15151 3893 15160 3927
rect 15108 3884 15160 3893
rect 15660 3884 15712 3936
rect 17132 3884 17184 3936
rect 17316 3927 17368 3936
rect 17316 3893 17325 3927
rect 17325 3893 17359 3927
rect 17359 3893 17368 3927
rect 17316 3884 17368 3893
rect 17408 3884 17460 3936
rect 18512 3927 18564 3936
rect 18512 3893 18521 3927
rect 18521 3893 18555 3927
rect 18555 3893 18564 3927
rect 20260 3952 20312 4004
rect 18512 3884 18564 3893
rect 19340 3884 19392 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 20904 3884 20956 3936
rect 7846 3782 7898 3834
rect 7910 3782 7962 3834
rect 7974 3782 8026 3834
rect 8038 3782 8090 3834
rect 14710 3782 14762 3834
rect 14774 3782 14826 3834
rect 14838 3782 14890 3834
rect 14902 3782 14954 3834
rect 3516 3680 3568 3732
rect 204 3612 256 3664
rect 2872 3612 2924 3664
rect 10140 3680 10192 3732
rect 10692 3680 10744 3732
rect 11520 3723 11572 3732
rect 11520 3689 11529 3723
rect 11529 3689 11563 3723
rect 11563 3689 11572 3723
rect 11520 3680 11572 3689
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 12440 3680 12492 3732
rect 2412 3544 2464 3596
rect 1032 3476 1084 3528
rect 5540 3612 5592 3664
rect 7472 3612 7524 3664
rect 9956 3655 10008 3664
rect 5080 3544 5132 3596
rect 5172 3544 5224 3596
rect 6368 3544 6420 3596
rect 7012 3544 7064 3596
rect 8116 3544 8168 3596
rect 8576 3587 8628 3596
rect 8576 3553 8585 3587
rect 8585 3553 8619 3587
rect 8619 3553 8628 3587
rect 8576 3544 8628 3553
rect 8852 3544 8904 3596
rect 9680 3587 9732 3596
rect 9680 3553 9689 3587
rect 9689 3553 9723 3587
rect 9723 3553 9732 3587
rect 9680 3544 9732 3553
rect 3608 3476 3660 3528
rect 4252 3476 4304 3528
rect 4896 3476 4948 3528
rect 5264 3476 5316 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7564 3476 7616 3528
rect 8392 3476 8444 3528
rect 3332 3408 3384 3460
rect 7104 3408 7156 3460
rect 8944 3476 8996 3528
rect 9588 3476 9640 3528
rect 9956 3621 9965 3655
rect 9965 3621 9999 3655
rect 9999 3621 10008 3655
rect 9956 3612 10008 3621
rect 10876 3655 10928 3664
rect 10876 3621 10885 3655
rect 10885 3621 10919 3655
rect 10919 3621 10928 3655
rect 10876 3612 10928 3621
rect 14372 3680 14424 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15660 3680 15712 3689
rect 16488 3680 16540 3732
rect 14004 3612 14056 3664
rect 15844 3612 15896 3664
rect 16672 3655 16724 3664
rect 11612 3476 11664 3528
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 8852 3408 8904 3460
rect 2872 3340 2924 3392
rect 7012 3340 7064 3392
rect 9036 3340 9088 3392
rect 10232 3340 10284 3392
rect 13728 3544 13780 3596
rect 14556 3544 14608 3596
rect 16672 3621 16706 3655
rect 16706 3621 16724 3655
rect 16672 3612 16724 3621
rect 17684 3680 17736 3732
rect 18512 3723 18564 3732
rect 18512 3689 18521 3723
rect 18521 3689 18555 3723
rect 18555 3689 18564 3723
rect 18512 3680 18564 3689
rect 18972 3723 19024 3732
rect 18236 3612 18288 3664
rect 13084 3519 13136 3528
rect 13084 3485 13093 3519
rect 13093 3485 13127 3519
rect 13127 3485 13136 3519
rect 13084 3476 13136 3485
rect 15108 3476 15160 3528
rect 17868 3544 17920 3596
rect 18512 3544 18564 3596
rect 18972 3689 18981 3723
rect 18981 3689 19015 3723
rect 19015 3689 19024 3723
rect 18972 3680 19024 3689
rect 19064 3680 19116 3732
rect 19248 3680 19300 3732
rect 19984 3680 20036 3732
rect 19708 3612 19760 3664
rect 20536 3612 20588 3664
rect 19248 3544 19300 3596
rect 15016 3408 15068 3460
rect 19064 3519 19116 3528
rect 19064 3485 19073 3519
rect 19073 3485 19107 3519
rect 19107 3485 19116 3519
rect 19064 3476 19116 3485
rect 20444 3519 20496 3528
rect 19984 3408 20036 3460
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 20812 3408 20864 3460
rect 10600 3340 10652 3392
rect 12532 3383 12584 3392
rect 12532 3349 12541 3383
rect 12541 3349 12575 3383
rect 12575 3349 12584 3383
rect 12532 3340 12584 3349
rect 14096 3340 14148 3392
rect 17592 3340 17644 3392
rect 20904 3340 20956 3392
rect 4414 3238 4466 3290
rect 4478 3238 4530 3290
rect 4542 3238 4594 3290
rect 4606 3238 4658 3290
rect 11278 3238 11330 3290
rect 11342 3238 11394 3290
rect 11406 3238 11458 3290
rect 11470 3238 11522 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 18270 3238 18322 3290
rect 18334 3238 18386 3290
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 1492 3068 1544 3120
rect 572 3000 624 3052
rect 3148 3068 3200 3120
rect 2872 3000 2924 3052
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 4068 3136 4120 3188
rect 8208 3179 8260 3188
rect 6000 3068 6052 3120
rect 6736 3068 6788 3120
rect 5080 3043 5132 3052
rect 3056 3000 3108 3009
rect 5080 3009 5089 3043
rect 5089 3009 5123 3043
rect 5123 3009 5132 3043
rect 5080 3000 5132 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 8208 3145 8217 3179
rect 8217 3145 8251 3179
rect 8251 3145 8260 3179
rect 8208 3136 8260 3145
rect 12716 3136 12768 3188
rect 18972 3136 19024 3188
rect 8484 3068 8536 3120
rect 8944 3068 8996 3120
rect 11796 3068 11848 3120
rect 12256 3068 12308 3120
rect 17316 3068 17368 3120
rect 6368 3000 6420 3009
rect 3240 2932 3292 2984
rect 2412 2864 2464 2916
rect 6736 2932 6788 2984
rect 3608 2864 3660 2916
rect 3240 2796 3292 2848
rect 6644 2864 6696 2916
rect 7564 2932 7616 2984
rect 9036 2975 9088 2984
rect 6920 2864 6972 2916
rect 7012 2864 7064 2916
rect 5080 2796 5132 2848
rect 5816 2796 5868 2848
rect 6092 2839 6144 2848
rect 6092 2805 6101 2839
rect 6101 2805 6135 2839
rect 6135 2805 6144 2839
rect 6092 2796 6144 2805
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 9036 2941 9045 2975
rect 9045 2941 9079 2975
rect 9079 2941 9088 2975
rect 9036 2932 9088 2941
rect 15476 3000 15528 3052
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 17684 3000 17736 3052
rect 17868 3000 17920 3052
rect 10232 2932 10284 2984
rect 10324 2932 10376 2984
rect 12624 2975 12676 2984
rect 12624 2941 12633 2975
rect 12633 2941 12667 2975
rect 12667 2941 12676 2975
rect 12624 2932 12676 2941
rect 6184 2796 6236 2805
rect 10324 2796 10376 2848
rect 10600 2796 10652 2848
rect 11612 2864 11664 2916
rect 11980 2864 12032 2916
rect 14096 2975 14148 2984
rect 14096 2941 14105 2975
rect 14105 2941 14139 2975
rect 14139 2941 14148 2975
rect 14096 2932 14148 2941
rect 14924 2932 14976 2984
rect 15384 2932 15436 2984
rect 17040 2932 17092 2984
rect 17132 2932 17184 2984
rect 17500 2932 17552 2984
rect 18144 2932 18196 2984
rect 22100 3068 22152 3120
rect 20444 3043 20496 3052
rect 20444 3009 20453 3043
rect 20453 3009 20487 3043
rect 20487 3009 20496 3043
rect 20444 3000 20496 3009
rect 13544 2864 13596 2916
rect 13084 2796 13136 2848
rect 14464 2864 14516 2916
rect 15200 2864 15252 2916
rect 17868 2864 17920 2916
rect 22560 2932 22612 2984
rect 18788 2864 18840 2916
rect 18880 2864 18932 2916
rect 21640 2864 21692 2916
rect 15292 2796 15344 2848
rect 19340 2796 19392 2848
rect 19432 2839 19484 2848
rect 19432 2805 19441 2839
rect 19441 2805 19475 2839
rect 19475 2805 19484 2839
rect 19432 2796 19484 2805
rect 20168 2796 20220 2848
rect 7846 2694 7898 2746
rect 7910 2694 7962 2746
rect 7974 2694 8026 2746
rect 8038 2694 8090 2746
rect 14710 2694 14762 2746
rect 14774 2694 14826 2746
rect 14838 2694 14890 2746
rect 14902 2694 14954 2746
rect 3240 2592 3292 2644
rect 7104 2592 7156 2644
rect 7472 2592 7524 2644
rect 8576 2635 8628 2644
rect 3608 2524 3660 2576
rect 4896 2524 4948 2576
rect 8576 2601 8585 2635
rect 8585 2601 8619 2635
rect 8619 2601 8628 2635
rect 8576 2592 8628 2601
rect 9312 2592 9364 2644
rect 9864 2592 9916 2644
rect 10232 2635 10284 2644
rect 10232 2601 10241 2635
rect 10241 2601 10275 2635
rect 10275 2601 10284 2635
rect 10232 2592 10284 2601
rect 10324 2592 10376 2644
rect 3976 2456 4028 2508
rect 4804 2456 4856 2508
rect 2596 2388 2648 2440
rect 4068 2388 4120 2440
rect 7012 2456 7064 2508
rect 8484 2456 8536 2508
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 8852 2431 8904 2440
rect 7564 2388 7616 2397
rect 8852 2397 8861 2431
rect 8861 2397 8895 2431
rect 8895 2397 8904 2431
rect 8852 2388 8904 2397
rect 2872 2320 2924 2372
rect 5724 2320 5776 2372
rect 14004 2592 14056 2644
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 12532 2456 12584 2508
rect 16672 2524 16724 2576
rect 13268 2456 13320 2508
rect 13544 2456 13596 2508
rect 14464 2456 14516 2508
rect 15200 2456 15252 2508
rect 15476 2499 15528 2508
rect 15476 2465 15485 2499
rect 15485 2465 15519 2499
rect 15519 2465 15528 2499
rect 15476 2456 15528 2465
rect 16212 2456 16264 2508
rect 16580 2499 16632 2508
rect 16580 2465 16589 2499
rect 16589 2465 16623 2499
rect 16623 2465 16632 2499
rect 16580 2456 16632 2465
rect 17868 2635 17920 2644
rect 17868 2601 17877 2635
rect 17877 2601 17911 2635
rect 17911 2601 17920 2635
rect 17868 2592 17920 2601
rect 18604 2635 18656 2644
rect 18604 2601 18613 2635
rect 18613 2601 18647 2635
rect 18647 2601 18656 2635
rect 18604 2592 18656 2601
rect 19156 2592 19208 2644
rect 19524 2592 19576 2644
rect 19984 2635 20036 2644
rect 19984 2601 19993 2635
rect 19993 2601 20027 2635
rect 20027 2601 20036 2635
rect 19984 2592 20036 2601
rect 19432 2524 19484 2576
rect 17592 2456 17644 2508
rect 18880 2456 18932 2508
rect 19248 2456 19300 2508
rect 20076 2499 20128 2508
rect 20076 2465 20085 2499
rect 20085 2465 20119 2499
rect 20119 2465 20128 2499
rect 20076 2456 20128 2465
rect 17776 2388 17828 2440
rect 19156 2431 19208 2440
rect 19156 2397 19165 2431
rect 19165 2397 19199 2431
rect 19199 2397 19208 2431
rect 19156 2388 19208 2397
rect 20168 2431 20220 2440
rect 20168 2397 20177 2431
rect 20177 2397 20211 2431
rect 20211 2397 20220 2431
rect 20168 2388 20220 2397
rect 14372 2320 14424 2372
rect 17132 2320 17184 2372
rect 8668 2252 8720 2304
rect 15384 2252 15436 2304
rect 15844 2252 15896 2304
rect 17960 2320 18012 2372
rect 4414 2150 4466 2202
rect 4478 2150 4530 2202
rect 4542 2150 4594 2202
rect 4606 2150 4658 2202
rect 11278 2150 11330 2202
rect 11342 2150 11394 2202
rect 11406 2150 11458 2202
rect 11470 2150 11522 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 18270 2150 18322 2202
rect 18334 2150 18386 2202
rect 6644 2048 6696 2100
rect 8484 2048 8536 2100
rect 6736 1980 6788 2032
rect 8576 1980 8628 2032
rect 3976 1232 4028 1284
rect 4988 1232 5040 1284
rect 21088 620 21140 672
rect 20260 552 20312 604
rect 20720 552 20772 604
rect 20996 552 21048 604
<< metal2 >>
rect 2962 22536 3018 22545
rect 2962 22471 3018 22480
rect 2318 22128 2374 22137
rect 2318 22063 2374 22072
rect 1950 19816 2006 19825
rect 1950 19751 2006 19760
rect 1964 19514 1992 19751
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1950 19272 2006 19281
rect 1950 19207 2006 19216
rect 1964 18970 1992 19207
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 1950 18864 2006 18873
rect 1950 18799 2006 18808
rect 1964 18426 1992 18799
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1768 18216 1820 18222
rect 1768 18158 1820 18164
rect 1674 17912 1730 17921
rect 1674 17847 1730 17856
rect 1688 17338 1716 17847
rect 1780 17814 1808 18158
rect 1872 17882 1900 18255
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1768 17808 1820 17814
rect 1768 17750 1820 17756
rect 1950 17368 2006 17377
rect 1676 17332 1728 17338
rect 1950 17303 2006 17312
rect 1676 17274 1728 17280
rect 1964 16794 1992 17303
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1950 16552 2006 16561
rect 1950 16487 2006 16496
rect 1964 16250 1992 16487
rect 2332 16250 2360 22063
rect 2502 21176 2558 21185
rect 2502 21111 2558 21120
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 1950 16008 2006 16017
rect 1950 15943 2006 15952
rect 1964 15706 1992 15943
rect 2516 15706 2544 21111
rect 2778 20224 2834 20233
rect 2778 20159 2834 20168
rect 2792 19174 2820 20159
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2778 15600 2834 15609
rect 2778 15535 2834 15544
rect 2792 15162 2820 15535
rect 2780 15156 2832 15162
rect 2780 15098 2832 15104
rect 1952 15088 2004 15094
rect 1950 15056 1952 15065
rect 2004 15056 2006 15065
rect 1950 14991 2006 15000
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 2596 14952 2648 14958
rect 2596 14894 2648 14900
rect 2780 14952 2832 14958
rect 2780 14894 2832 14900
rect 1674 14648 1730 14657
rect 1674 14583 1676 14592
rect 1728 14583 1730 14592
rect 1676 14554 1728 14560
rect 1780 14550 1808 14894
rect 1768 14544 1820 14550
rect 1768 14486 1820 14492
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 9518 1440 12038
rect 1504 10713 1532 14418
rect 1582 14104 1638 14113
rect 1582 14039 1638 14048
rect 1596 13530 1624 14039
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1964 12850 1992 13330
rect 1952 12844 2004 12850
rect 1952 12786 2004 12792
rect 1768 12776 1820 12782
rect 1768 12718 1820 12724
rect 1780 10810 1808 12718
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 2056 11762 2084 12174
rect 2044 11756 2096 11762
rect 2044 11698 2096 11704
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 1490 10704 1546 10713
rect 1490 10639 1546 10648
rect 1872 9586 1900 11494
rect 2056 10130 2084 11698
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 2056 8634 2084 10066
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1688 6866 1716 8366
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1964 7993 1992 8026
rect 1950 7984 2006 7993
rect 1950 7919 2006 7928
rect 2148 7546 2176 13806
rect 2320 13388 2372 13394
rect 2320 13330 2372 13336
rect 2332 12442 2360 13330
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2424 12986 2452 13262
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2320 12436 2372 12442
rect 2320 12378 2372 12384
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2240 10606 2268 11494
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2332 9178 2360 11494
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 9722 2452 10406
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9178 2544 12582
rect 2608 10169 2636 14894
rect 2792 14074 2820 14894
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2884 13530 2912 14418
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 2976 12850 3004 22471
rect 5722 22320 5778 22800
rect 17130 22320 17186 22800
rect 19062 22536 19118 22545
rect 19062 22471 19118 22480
rect 3146 21584 3202 21593
rect 3146 21519 3202 21528
rect 3160 14618 3188 21519
rect 3698 20632 3754 20641
rect 3698 20567 3754 20576
rect 3712 19514 3740 20567
rect 4388 19612 4684 19632
rect 4444 19610 4468 19612
rect 4524 19610 4548 19612
rect 4604 19610 4628 19612
rect 4466 19558 4468 19610
rect 4530 19558 4542 19610
rect 4604 19558 4606 19610
rect 4444 19556 4468 19558
rect 4524 19556 4548 19558
rect 4604 19556 4628 19558
rect 4388 19536 4684 19556
rect 3700 19508 3752 19514
rect 3700 19450 3752 19456
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4388 18524 4684 18544
rect 4444 18522 4468 18524
rect 4524 18522 4548 18524
rect 4604 18522 4628 18524
rect 4466 18470 4468 18522
rect 4530 18470 4542 18522
rect 4604 18470 4606 18522
rect 4444 18468 4468 18470
rect 4524 18468 4548 18470
rect 4604 18468 4628 18470
rect 4388 18448 4684 18468
rect 4388 17436 4684 17456
rect 4444 17434 4468 17436
rect 4524 17434 4548 17436
rect 4604 17434 4628 17436
rect 4466 17382 4468 17434
rect 4530 17382 4542 17434
rect 4604 17382 4606 17434
rect 4444 17380 4468 17382
rect 4524 17380 4548 17382
rect 4604 17380 4628 17382
rect 4388 17360 4684 17380
rect 3422 16960 3478 16969
rect 3422 16895 3478 16904
rect 3436 16250 3464 16895
rect 4388 16348 4684 16368
rect 4444 16346 4468 16348
rect 4524 16346 4548 16348
rect 4604 16346 4628 16348
rect 4466 16294 4468 16346
rect 4530 16294 4542 16346
rect 4604 16294 4606 16346
rect 4444 16292 4468 16294
rect 4524 16292 4548 16294
rect 4604 16292 4628 16294
rect 4388 16272 4684 16292
rect 3424 16244 3476 16250
rect 3424 16186 3476 16192
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 15638 3280 15982
rect 3240 15632 3292 15638
rect 3240 15574 3292 15580
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4172 14906 4200 15370
rect 3792 14884 3844 14890
rect 3792 14826 3844 14832
rect 4080 14878 4200 14906
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3056 13796 3108 13802
rect 3056 13738 3108 13744
rect 3068 12850 3096 13738
rect 2964 12844 3016 12850
rect 2964 12786 3016 12792
rect 3056 12844 3108 12850
rect 3056 12786 3108 12792
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11354 2820 12242
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2594 10160 2650 10169
rect 2594 10095 2650 10104
rect 2700 9722 2728 11154
rect 2976 10810 3004 12310
rect 3068 12238 3096 12786
rect 3160 12306 3188 13806
rect 3252 13530 3280 14350
rect 3516 14068 3568 14074
rect 3516 14010 3568 14016
rect 3330 13696 3386 13705
rect 3330 13631 3386 13640
rect 3344 13530 3372 13631
rect 3240 13524 3292 13530
rect 3240 13466 3292 13472
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3436 12986 3464 13262
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3528 12918 3556 14010
rect 3804 13734 3832 14826
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 4080 13682 4108 14878
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14414 4200 14758
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 4172 13870 4200 14350
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 3804 13326 3832 13670
rect 4080 13654 4200 13682
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3792 13320 3844 13326
rect 3606 13288 3662 13297
rect 3792 13262 3844 13268
rect 3606 13223 3662 13232
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3528 12714 3556 12854
rect 3516 12708 3568 12714
rect 3516 12650 3568 12656
rect 3620 12442 3648 13223
rect 3896 12986 3924 13330
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3988 12850 4016 13194
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3974 12744 4030 12753
rect 3700 12708 3752 12714
rect 3700 12650 3752 12656
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 3148 12300 3200 12306
rect 3148 12242 3200 12248
rect 3516 12300 3568 12306
rect 3516 12242 3568 12248
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 10804 3016 10810
rect 2964 10746 3016 10752
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2884 9654 2912 10542
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1952 7268 2004 7274
rect 1952 7210 2004 7216
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6322 1716 6802
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1964 5914 1992 7210
rect 2424 6934 2452 7822
rect 2412 6928 2464 6934
rect 2412 6870 2464 6876
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2148 4690 2176 6258
rect 2240 6254 2268 6802
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 2240 5234 2268 6190
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2424 5370 2452 5646
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2516 5030 2544 9114
rect 2700 8974 2728 9454
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2148 4282 2176 4626
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 204 3664 256 3670
rect 204 3606 256 3612
rect 216 480 244 3606
rect 1032 3528 1084 3534
rect 1032 3470 1084 3476
rect 572 3052 624 3058
rect 572 2994 624 3000
rect 584 480 612 2994
rect 1044 480 1072 3470
rect 1492 3120 1544 3126
rect 1492 3062 1544 3068
rect 1504 480 1532 3062
rect 1964 480 1992 3946
rect 2332 2553 2360 4966
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2424 3194 2452 3538
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2412 2916 2464 2922
rect 2412 2858 2464 2864
rect 2318 2544 2374 2553
rect 2318 2479 2374 2488
rect 2424 480 2452 2858
rect 2516 1601 2544 4966
rect 2608 2446 2636 8910
rect 2700 8362 2728 8910
rect 2688 8356 2740 8362
rect 2688 8298 2740 8304
rect 2700 7886 2728 8298
rect 2688 7880 2740 7886
rect 2976 7857 3004 9318
rect 3068 9178 3096 12038
rect 3160 10606 3188 12106
rect 3332 11620 3384 11626
rect 3332 11562 3384 11568
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3252 10198 3280 11222
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9722 3188 9862
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3252 8294 3280 8570
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3056 8016 3108 8022
rect 3056 7958 3108 7964
rect 2688 7822 2740 7828
rect 2962 7848 3018 7857
rect 2962 7783 3018 7792
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2792 6458 2820 7346
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2870 5128 2926 5137
rect 2976 5098 3004 7783
rect 3068 7546 3096 7958
rect 3252 7818 3280 8230
rect 3240 7812 3292 7818
rect 3240 7754 3292 7760
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3068 7002 3096 7346
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 3068 6186 3096 6938
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3068 5710 3096 6122
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2870 5063 2926 5072
rect 2964 5092 3016 5098
rect 2884 3670 2912 5063
rect 2964 5034 3016 5040
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3160 4282 3188 4626
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2884 3058 2912 3334
rect 3068 3058 3096 4014
rect 3148 3120 3200 3126
rect 3146 3088 3148 3097
rect 3200 3088 3202 3097
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 3056 3052 3108 3058
rect 3146 3023 3202 3032
rect 3056 2994 3108 3000
rect 3252 2990 3280 4694
rect 3344 3466 3372 11562
rect 3528 11082 3556 12242
rect 3712 12238 3740 12650
rect 3896 12424 3924 12718
rect 3974 12679 3976 12688
rect 4028 12679 4030 12688
rect 3976 12650 4028 12656
rect 3804 12396 3924 12424
rect 3700 12232 3752 12238
rect 3700 12174 3752 12180
rect 3712 11218 3740 12174
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3528 10674 3556 11018
rect 3700 11008 3752 11014
rect 3700 10950 3752 10956
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3528 10130 3556 10406
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3620 9586 3648 10610
rect 3712 10033 3740 10950
rect 3698 10024 3754 10033
rect 3698 9959 3754 9968
rect 3804 9908 3832 12396
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 3896 12102 3924 12271
rect 3884 12096 3936 12102
rect 4080 12050 4108 13330
rect 4172 12374 4200 13654
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3884 12038 3936 12044
rect 3988 12022 4108 12050
rect 3988 11694 4016 12022
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4080 11801 4108 11834
rect 4066 11792 4122 11801
rect 4066 11727 4122 11736
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 3882 10840 3938 10849
rect 3882 10775 3938 10784
rect 3896 10674 3924 10775
rect 3884 10668 3936 10674
rect 3884 10610 3936 10616
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3712 9880 3832 9908
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3712 9518 3740 9880
rect 3700 9512 3752 9518
rect 3700 9454 3752 9460
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 3436 8022 3464 9046
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3424 8016 3476 8022
rect 3516 8016 3568 8022
rect 3424 7958 3476 7964
rect 3514 7984 3516 7993
rect 3568 7984 3570 7993
rect 3436 4622 3464 7958
rect 3514 7919 3570 7928
rect 3712 7886 3740 8434
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3792 7880 3844 7886
rect 3792 7822 3844 7828
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7342 3556 7686
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 3620 6254 3648 7414
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3712 4826 3740 7822
rect 3804 7478 3832 7822
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3792 7268 3844 7274
rect 3792 7210 3844 7216
rect 3804 7177 3832 7210
rect 3790 7168 3846 7177
rect 3790 7103 3846 7112
rect 3896 6118 3924 10474
rect 3988 8090 4016 11494
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4080 10606 4108 11154
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 9722 4108 10367
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4066 9480 4122 9489
rect 4066 9415 4122 9424
rect 4080 8838 4108 9415
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4172 8634 4200 11494
rect 4264 10266 4292 15506
rect 4388 15260 4684 15280
rect 4444 15258 4468 15260
rect 4524 15258 4548 15260
rect 4604 15258 4628 15260
rect 4466 15206 4468 15258
rect 4530 15206 4542 15258
rect 4604 15206 4606 15258
rect 4444 15204 4468 15206
rect 4524 15204 4548 15206
rect 4604 15204 4628 15206
rect 4388 15184 4684 15204
rect 4388 14172 4684 14192
rect 4444 14170 4468 14172
rect 4524 14170 4548 14172
rect 4604 14170 4628 14172
rect 4466 14118 4468 14170
rect 4530 14118 4542 14170
rect 4604 14118 4606 14170
rect 4444 14116 4468 14118
rect 4524 14116 4548 14118
rect 4604 14116 4628 14118
rect 4388 14096 4684 14116
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4388 13084 4684 13104
rect 4444 13082 4468 13084
rect 4524 13082 4548 13084
rect 4604 13082 4628 13084
rect 4466 13030 4468 13082
rect 4530 13030 4542 13082
rect 4604 13030 4606 13082
rect 4444 13028 4468 13030
rect 4524 13028 4548 13030
rect 4604 13028 4628 13030
rect 4388 13008 4684 13028
rect 4724 12782 4752 13126
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4388 11996 4684 12016
rect 4444 11994 4468 11996
rect 4524 11994 4548 11996
rect 4604 11994 4628 11996
rect 4466 11942 4468 11994
rect 4530 11942 4542 11994
rect 4604 11942 4606 11994
rect 4444 11940 4468 11942
rect 4524 11940 4548 11942
rect 4604 11940 4628 11942
rect 4388 11920 4684 11940
rect 4388 10908 4684 10928
rect 4444 10906 4468 10908
rect 4524 10906 4548 10908
rect 4604 10906 4628 10908
rect 4466 10854 4468 10906
rect 4530 10854 4542 10906
rect 4604 10854 4606 10906
rect 4444 10852 4468 10854
rect 4524 10852 4548 10854
rect 4604 10852 4628 10854
rect 4388 10832 4684 10852
rect 4618 10568 4674 10577
rect 4618 10503 4674 10512
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4264 9704 4292 10066
rect 4632 9994 4660 10503
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4388 9820 4684 9840
rect 4444 9818 4468 9820
rect 4524 9818 4548 9820
rect 4604 9818 4628 9820
rect 4466 9766 4468 9818
rect 4530 9766 4542 9818
rect 4604 9766 4606 9818
rect 4444 9764 4468 9766
rect 4524 9764 4548 9766
rect 4604 9764 4628 9766
rect 4388 9744 4684 9764
rect 4264 9676 4568 9704
rect 4448 9518 4476 9549
rect 4252 9512 4304 9518
rect 4436 9512 4488 9518
rect 4252 9454 4304 9460
rect 4356 9460 4436 9466
rect 4540 9466 4568 9676
rect 4488 9460 4568 9466
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4068 8560 4120 8566
rect 4066 8528 4068 8537
rect 4120 8528 4122 8537
rect 4066 8463 4122 8472
rect 4264 8090 4292 9454
rect 4356 9438 4568 9460
rect 4356 8888 4384 9438
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4448 8906 4476 9318
rect 4632 9042 4660 9318
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4325 8860 4384 8888
rect 4436 8900 4488 8906
rect 4325 8616 4353 8860
rect 4436 8842 4488 8848
rect 4388 8732 4684 8752
rect 4444 8730 4468 8732
rect 4524 8730 4548 8732
rect 4604 8730 4628 8732
rect 4466 8678 4468 8730
rect 4530 8678 4542 8730
rect 4604 8678 4606 8730
rect 4444 8676 4468 8678
rect 4524 8676 4548 8678
rect 4604 8676 4628 8678
rect 4388 8656 4684 8676
rect 4325 8588 4384 8616
rect 3976 8084 4028 8090
rect 3976 8026 4028 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 3974 7984 4030 7993
rect 4356 7970 4384 8588
rect 3974 7919 3976 7928
rect 4028 7919 4030 7928
rect 4160 7948 4212 7954
rect 3976 7890 4028 7896
rect 4160 7890 4212 7896
rect 4264 7942 4384 7970
rect 3974 7576 4030 7585
rect 4172 7546 4200 7890
rect 3974 7511 4030 7520
rect 4160 7540 4212 7546
rect 3988 7410 4016 7511
rect 4160 7482 4212 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3974 6216 4030 6225
rect 3974 6151 4030 6160
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3804 5914 3832 6054
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3608 4276 3660 4282
rect 3608 4218 3660 4224
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 3738 3556 3878
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 3620 3534 3648 4218
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3608 3528 3660 3534
rect 3608 3470 3660 3476
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 3330 2816 3386 2825
rect 3252 2650 3280 2790
rect 3330 2751 3386 2760
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2502 1592 2558 1601
rect 2502 1527 2558 1536
rect 2884 480 2912 2314
rect 3344 480 3372 2751
rect 3620 2582 3648 2858
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3712 480 3740 4150
rect 3896 3505 3924 6054
rect 3988 5914 4016 6151
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5846 4108 6394
rect 4172 6390 4200 6734
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4068 5840 4120 5846
rect 3974 5808 4030 5817
rect 4068 5782 4120 5788
rect 3974 5743 3976 5752
rect 4028 5743 4030 5752
rect 3976 5714 4028 5720
rect 4068 5704 4120 5710
rect 4172 5692 4200 6326
rect 4120 5664 4200 5692
rect 4068 5646 4120 5652
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4080 5273 4108 5306
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4865 4016 5034
rect 3974 4856 4030 4865
rect 3974 4791 4030 4800
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 4321 4108 4762
rect 4172 4758 4200 5664
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 4066 4312 4122 4321
rect 4066 4247 4122 4256
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3882 3496 3938 3505
rect 3882 3431 3938 3440
rect 4080 3194 4108 4082
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 3988 2009 4016 2450
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 3974 2000 4030 2009
rect 3974 1935 4030 1944
rect 3976 1284 4028 1290
rect 3976 1226 4028 1232
rect 3988 649 4016 1226
rect 4080 1057 4108 2382
rect 4066 1048 4122 1057
rect 4066 983 4122 992
rect 3974 640 4030 649
rect 3974 575 4030 584
rect 4172 480 4200 4558
rect 4264 3534 4292 7942
rect 4388 7644 4684 7664
rect 4444 7642 4468 7644
rect 4524 7642 4548 7644
rect 4604 7642 4628 7644
rect 4466 7590 4468 7642
rect 4530 7590 4542 7642
rect 4604 7590 4606 7642
rect 4444 7588 4468 7590
rect 4524 7588 4548 7590
rect 4604 7588 4628 7590
rect 4388 7568 4684 7588
rect 4388 6556 4684 6576
rect 4444 6554 4468 6556
rect 4524 6554 4548 6556
rect 4604 6554 4628 6556
rect 4466 6502 4468 6554
rect 4530 6502 4542 6554
rect 4604 6502 4606 6554
rect 4444 6500 4468 6502
rect 4524 6500 4548 6502
rect 4604 6500 4628 6502
rect 4388 6480 4684 6500
rect 4388 5468 4684 5488
rect 4444 5466 4468 5468
rect 4524 5466 4548 5468
rect 4604 5466 4628 5468
rect 4466 5414 4468 5466
rect 4530 5414 4542 5466
rect 4604 5414 4606 5466
rect 4444 5412 4468 5414
rect 4524 5412 4548 5414
rect 4604 5412 4628 5414
rect 4388 5392 4684 5412
rect 4388 4380 4684 4400
rect 4444 4378 4468 4380
rect 4524 4378 4548 4380
rect 4604 4378 4628 4380
rect 4466 4326 4468 4378
rect 4530 4326 4542 4378
rect 4604 4326 4606 4378
rect 4444 4324 4468 4326
rect 4524 4324 4548 4326
rect 4604 4324 4628 4326
rect 4388 4304 4684 4324
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 2961 4292 3470
rect 4388 3292 4684 3312
rect 4444 3290 4468 3292
rect 4524 3290 4548 3292
rect 4604 3290 4628 3292
rect 4466 3238 4468 3290
rect 4530 3238 4542 3290
rect 4604 3238 4606 3290
rect 4444 3236 4468 3238
rect 4524 3236 4548 3238
rect 4604 3236 4628 3238
rect 4388 3216 4684 3236
rect 4250 2952 4306 2961
rect 4250 2887 4306 2896
rect 4388 2204 4684 2224
rect 4444 2202 4468 2204
rect 4524 2202 4548 2204
rect 4604 2202 4628 2204
rect 4466 2150 4468 2202
rect 4530 2150 4542 2202
rect 4604 2150 4606 2202
rect 4444 2148 4468 2150
rect 4524 2148 4548 2150
rect 4604 2148 4628 2150
rect 4388 2128 4684 2148
rect 4724 1986 4752 12582
rect 4816 10282 4844 19246
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4908 10577 4936 19178
rect 5736 18222 5764 22320
rect 7820 20156 8116 20176
rect 7876 20154 7900 20156
rect 7956 20154 7980 20156
rect 8036 20154 8060 20156
rect 7898 20102 7900 20154
rect 7962 20102 7974 20154
rect 8036 20102 8038 20154
rect 7876 20100 7900 20102
rect 7956 20100 7980 20102
rect 8036 20100 8060 20102
rect 7820 20080 8116 20100
rect 14684 20156 14980 20176
rect 14740 20154 14764 20156
rect 14820 20154 14844 20156
rect 14900 20154 14924 20156
rect 14762 20102 14764 20154
rect 14826 20102 14838 20154
rect 14900 20102 14902 20154
rect 14740 20100 14764 20102
rect 14820 20100 14844 20102
rect 14900 20100 14924 20102
rect 14684 20080 14980 20100
rect 11252 19612 11548 19632
rect 11308 19610 11332 19612
rect 11388 19610 11412 19612
rect 11468 19610 11492 19612
rect 11330 19558 11332 19610
rect 11394 19558 11406 19610
rect 11468 19558 11470 19610
rect 11308 19556 11332 19558
rect 11388 19556 11412 19558
rect 11468 19556 11492 19558
rect 11252 19536 11548 19556
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5828 18902 5856 19246
rect 7820 19068 8116 19088
rect 7876 19066 7900 19068
rect 7956 19066 7980 19068
rect 8036 19066 8060 19068
rect 7898 19014 7900 19066
rect 7962 19014 7974 19066
rect 8036 19014 8038 19066
rect 7876 19012 7900 19014
rect 7956 19012 7980 19014
rect 8036 19012 8060 19014
rect 7820 18992 8116 19012
rect 14684 19068 14980 19088
rect 14740 19066 14764 19068
rect 14820 19066 14844 19068
rect 14900 19066 14924 19068
rect 14762 19014 14764 19066
rect 14826 19014 14838 19066
rect 14900 19014 14902 19066
rect 14740 19012 14764 19014
rect 14820 19012 14844 19014
rect 14900 19012 14924 19014
rect 14684 18992 14980 19012
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5080 15496 5132 15502
rect 5080 15438 5132 15444
rect 5092 14618 5120 15438
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5092 13530 5120 14554
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5080 13524 5132 13530
rect 5080 13466 5132 13472
rect 5080 12368 5132 12374
rect 5080 12310 5132 12316
rect 4894 10568 4950 10577
rect 4894 10503 4950 10512
rect 4816 10254 5028 10282
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9178 4844 10066
rect 5000 9654 5028 10254
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4908 8974 4936 9590
rect 4986 9480 5042 9489
rect 4986 9415 5042 9424
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 6458 4844 7142
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4908 6338 4936 8910
rect 4816 6310 4936 6338
rect 4816 2514 4844 6310
rect 5000 5273 5028 9415
rect 5092 8634 5120 12310
rect 5184 11762 5212 13942
rect 5276 12306 5304 14418
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5184 10538 5212 11698
rect 5276 11694 5304 12242
rect 5368 11778 5396 16594
rect 5448 15972 5500 15978
rect 5448 15914 5500 15920
rect 5460 13802 5488 15914
rect 5632 13864 5684 13870
rect 5632 13806 5684 13812
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5460 13530 5488 13738
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12714 5488 13262
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5460 12442 5488 12650
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5368 11750 5488 11778
rect 5460 11694 5488 11750
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5448 11688 5500 11694
rect 5448 11630 5500 11636
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5460 10810 5488 11154
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5356 10736 5408 10742
rect 5356 10678 5408 10684
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5184 8974 5212 10474
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5092 8362 5120 8570
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5080 7948 5132 7954
rect 5080 7890 5132 7896
rect 5092 6186 5120 7890
rect 5184 7818 5212 8910
rect 5276 8090 5304 10474
rect 5368 10266 5396 10678
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5354 10160 5410 10169
rect 5354 10095 5410 10104
rect 5368 9994 5396 10095
rect 5460 9994 5488 10746
rect 5552 10062 5580 11018
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5368 7886 5396 9930
rect 5460 9654 5488 9685
rect 5644 9654 5672 13806
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10198 5764 10406
rect 5724 10192 5776 10198
rect 5724 10134 5776 10140
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5448 9648 5500 9654
rect 5446 9616 5448 9625
rect 5632 9648 5684 9654
rect 5500 9616 5502 9625
rect 5632 9590 5684 9596
rect 5446 9551 5502 9560
rect 5460 8430 5488 9551
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5448 8288 5500 8294
rect 5540 8288 5592 8294
rect 5448 8230 5500 8236
rect 5538 8256 5540 8265
rect 5592 8256 5594 8265
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5184 7392 5212 7754
rect 5356 7404 5408 7410
rect 5184 7364 5356 7392
rect 5356 7346 5408 7352
rect 5460 7290 5488 8230
rect 5538 8191 5594 8200
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5184 7262 5488 7290
rect 5184 6322 5212 7262
rect 5264 7200 5316 7206
rect 5316 7160 5396 7188
rect 5264 7142 5316 7148
rect 5368 6934 5396 7160
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4986 5264 5042 5273
rect 4986 5199 4988 5208
rect 5040 5199 5042 5208
rect 4988 5170 5040 5176
rect 5000 5139 5028 5170
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4908 4146 4936 4966
rect 5092 4162 5120 6122
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5276 5914 5304 6054
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5012 5396 6870
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5460 6322 5488 6598
rect 5448 6316 5500 6322
rect 5448 6258 5500 6264
rect 5552 5658 5580 7822
rect 5644 7410 5672 8026
rect 5736 7546 5764 9998
rect 5828 8265 5856 18702
rect 6104 13530 6132 18770
rect 11252 18524 11548 18544
rect 11308 18522 11332 18524
rect 11388 18522 11412 18524
rect 11468 18522 11492 18524
rect 11330 18470 11332 18522
rect 11394 18470 11406 18522
rect 11468 18470 11470 18522
rect 11308 18468 11332 18470
rect 11388 18468 11412 18470
rect 11468 18468 11492 18470
rect 11252 18448 11548 18468
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7820 17980 8116 18000
rect 7876 17978 7900 17980
rect 7956 17978 7980 17980
rect 8036 17978 8060 17980
rect 7898 17926 7900 17978
rect 7962 17926 7974 17978
rect 8036 17926 8038 17978
rect 7876 17924 7900 17926
rect 7956 17924 7980 17926
rect 8036 17924 8060 17926
rect 7820 17904 8116 17924
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6184 13252 6236 13258
rect 6184 13194 6236 13200
rect 6196 12918 6224 13194
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5920 11558 5948 12174
rect 6184 11824 6236 11830
rect 6184 11766 6236 11772
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11286 5948 11494
rect 5998 11384 6054 11393
rect 5998 11319 6054 11328
rect 6012 11286 6040 11319
rect 5908 11280 5960 11286
rect 5908 11222 5960 11228
rect 6000 11280 6052 11286
rect 6000 11222 6052 11228
rect 5920 11150 5948 11222
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5920 10062 5948 11086
rect 6090 10704 6146 10713
rect 6196 10674 6224 11766
rect 6472 11558 6500 17070
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6090 10639 6146 10648
rect 6184 10668 6236 10674
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 6012 8498 6040 9454
rect 6000 8492 6052 8498
rect 6000 8434 6052 8440
rect 5814 8256 5870 8265
rect 5814 8191 5870 8200
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5460 5630 5580 5658
rect 5460 5166 5488 5630
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5552 5234 5580 5510
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5368 4984 5488 5012
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 4134 5120 4162
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4908 2582 4936 3470
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4632 1958 4752 1986
rect 4632 480 4660 1958
rect 5000 1290 5028 4134
rect 5184 3602 5212 4626
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 4146 5304 4422
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5092 3058 5120 3538
rect 5276 3534 5304 4082
rect 5368 3942 5396 4490
rect 5356 3936 5408 3942
rect 5460 3924 5488 4984
rect 5552 4758 5580 5170
rect 5724 5160 5776 5166
rect 5724 5102 5776 5108
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 5632 3936 5684 3942
rect 5460 3896 5632 3924
rect 5356 3878 5408 3884
rect 5632 3878 5684 3884
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 5080 2848 5132 2854
rect 5080 2790 5132 2796
rect 4988 1284 5040 1290
rect 4988 1226 5040 1232
rect 5092 480 5120 2790
rect 5552 480 5580 3606
rect 202 0 258 480
rect 570 0 626 480
rect 1030 0 1086 480
rect 1490 0 1546 480
rect 1950 0 2006 480
rect 2410 0 2466 480
rect 2870 0 2926 480
rect 3330 0 3386 480
rect 3698 0 3754 480
rect 4158 0 4214 480
rect 4618 0 4674 480
rect 5078 0 5134 480
rect 5538 0 5594 480
rect 5644 241 5672 3878
rect 5736 2378 5764 5102
rect 5828 2854 5856 7822
rect 6012 6866 6040 8434
rect 6104 8362 6132 10639
rect 6184 10610 6236 10616
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6196 9042 6224 9998
rect 6656 9654 6684 17682
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6840 13530 6868 13670
rect 6828 13524 6880 13530
rect 6828 13466 6880 13472
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6736 11348 6788 11354
rect 6736 11290 6788 11296
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6748 9042 6776 11290
rect 6840 10674 6868 13126
rect 7012 12368 7064 12374
rect 7012 12310 7064 12316
rect 7024 11801 7052 12310
rect 7010 11792 7066 11801
rect 7010 11727 7066 11736
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7116 11665 7144 11698
rect 7102 11656 7158 11665
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 7012 11620 7064 11626
rect 7102 11591 7158 11600
rect 7012 11562 7064 11568
rect 6932 11257 6960 11562
rect 6918 11248 6974 11257
rect 6918 11183 6974 11192
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 7024 10470 7052 11562
rect 7300 11218 7328 16050
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7392 12442 7420 13330
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7484 12374 7512 17614
rect 7820 16892 8116 16912
rect 7876 16890 7900 16892
rect 7956 16890 7980 16892
rect 8036 16890 8060 16892
rect 7898 16838 7900 16890
rect 7962 16838 7974 16890
rect 8036 16838 8038 16890
rect 7876 16836 7900 16838
rect 7956 16836 7980 16838
rect 8036 16836 8060 16838
rect 7820 16816 8116 16836
rect 7820 15804 8116 15824
rect 7876 15802 7900 15804
rect 7956 15802 7980 15804
rect 8036 15802 8060 15804
rect 7898 15750 7900 15802
rect 7962 15750 7974 15802
rect 8036 15750 8038 15802
rect 7876 15748 7900 15750
rect 7956 15748 7980 15750
rect 8036 15748 8060 15750
rect 7820 15728 8116 15748
rect 7820 14716 8116 14736
rect 7876 14714 7900 14716
rect 7956 14714 7980 14716
rect 8036 14714 8060 14716
rect 7898 14662 7900 14714
rect 7962 14662 7974 14714
rect 8036 14662 8038 14714
rect 7876 14660 7900 14662
rect 7956 14660 7980 14662
rect 8036 14660 8060 14662
rect 7820 14640 8116 14660
rect 8220 14550 8248 18158
rect 14684 17980 14980 18000
rect 14740 17978 14764 17980
rect 14820 17978 14844 17980
rect 14900 17978 14924 17980
rect 14762 17926 14764 17978
rect 14826 17926 14838 17978
rect 14900 17926 14902 17978
rect 14740 17924 14764 17926
rect 14820 17924 14844 17926
rect 14900 17924 14924 17926
rect 14684 17904 14980 17924
rect 11252 17436 11548 17456
rect 11308 17434 11332 17436
rect 11388 17434 11412 17436
rect 11468 17434 11492 17436
rect 11330 17382 11332 17434
rect 11394 17382 11406 17434
rect 11468 17382 11470 17434
rect 11308 17380 11332 17382
rect 11388 17380 11412 17382
rect 11468 17380 11492 17382
rect 11252 17360 11548 17380
rect 14684 16892 14980 16912
rect 14740 16890 14764 16892
rect 14820 16890 14844 16892
rect 14900 16890 14924 16892
rect 14762 16838 14764 16890
rect 14826 16838 14838 16890
rect 14900 16838 14902 16890
rect 14740 16836 14764 16838
rect 14820 16836 14844 16838
rect 14900 16836 14924 16838
rect 14684 16816 14980 16836
rect 11252 16348 11548 16368
rect 11308 16346 11332 16348
rect 11388 16346 11412 16348
rect 11468 16346 11492 16348
rect 11330 16294 11332 16346
rect 11394 16294 11406 16346
rect 11468 16294 11470 16346
rect 11308 16292 11332 16294
rect 11388 16292 11412 16294
rect 11468 16292 11492 16294
rect 11252 16272 11548 16292
rect 12808 16040 12860 16046
rect 12808 15982 12860 15988
rect 12820 15638 12848 15982
rect 14684 15804 14980 15824
rect 14740 15802 14764 15804
rect 14820 15802 14844 15804
rect 14900 15802 14924 15804
rect 14762 15750 14764 15802
rect 14826 15750 14838 15802
rect 14900 15750 14902 15802
rect 14740 15748 14764 15750
rect 14820 15748 14844 15750
rect 14900 15748 14924 15750
rect 14684 15728 14980 15748
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 11252 15260 11548 15280
rect 11308 15258 11332 15260
rect 11388 15258 11412 15260
rect 11468 15258 11492 15260
rect 11330 15206 11332 15258
rect 11394 15206 11406 15258
rect 11468 15206 11470 15258
rect 11308 15204 11332 15206
rect 11388 15204 11412 15206
rect 11468 15204 11492 15206
rect 11252 15184 11548 15204
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8404 13938 8432 14350
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 7576 13394 7604 13874
rect 7820 13628 8116 13648
rect 7876 13626 7900 13628
rect 7956 13626 7980 13628
rect 8036 13626 8060 13628
rect 7898 13574 7900 13626
rect 7962 13574 7974 13626
rect 8036 13574 8038 13626
rect 7876 13572 7900 13574
rect 7956 13572 7980 13574
rect 8036 13572 8060 13574
rect 7820 13552 8116 13572
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 12368 7524 12374
rect 7472 12310 7524 12316
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7484 11830 7512 12174
rect 7576 12170 7604 13330
rect 8404 13258 8432 13874
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8760 13796 8812 13802
rect 8760 13738 8812 13744
rect 8496 13258 8524 13738
rect 8772 13530 8800 13738
rect 9784 13734 9812 14418
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 10704 13938 10732 14350
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 9588 13728 9640 13734
rect 9586 13696 9588 13705
rect 9772 13728 9824 13734
rect 9640 13696 9642 13705
rect 9772 13670 9824 13676
rect 10416 13728 10468 13734
rect 10416 13670 10468 13676
rect 9586 13631 9642 13640
rect 8760 13524 8812 13530
rect 8760 13466 8812 13472
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8392 13252 8444 13258
rect 8392 13194 8444 13200
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 7656 12708 7708 12714
rect 7656 12650 7708 12656
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7562 11792 7618 11801
rect 7562 11727 7618 11736
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7576 10810 7604 11727
rect 7564 10804 7616 10810
rect 7300 10764 7564 10792
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 7012 10464 7064 10470
rect 7012 10406 7064 10412
rect 6932 9654 6960 10406
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6182 8936 6238 8945
rect 6182 8871 6184 8880
rect 6236 8871 6238 8880
rect 6184 8842 6236 8848
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6656 8537 6684 8570
rect 6642 8528 6698 8537
rect 6642 8463 6698 8472
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6550 8392 6606 8401
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6288 8090 6316 8230
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6380 7818 6408 8366
rect 6550 8327 6552 8336
rect 6604 8327 6606 8336
rect 6552 8298 6604 8304
rect 6644 8288 6696 8294
rect 6644 8230 6696 8236
rect 6656 7954 6684 8230
rect 6748 7954 6776 8978
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6736 7948 6788 7954
rect 6736 7890 6788 7896
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6368 7812 6420 7818
rect 6550 7783 6606 7792
rect 6368 7754 6420 7760
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6656 7206 6684 7482
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6012 5710 6040 6802
rect 6182 6216 6238 6225
rect 6182 6151 6238 6160
rect 6196 5914 6224 6151
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 6092 5364 6144 5370
rect 6092 5306 6144 5312
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 6012 480 6040 3062
rect 6104 2854 6132 5306
rect 6288 4622 6316 6802
rect 6380 4690 6408 6870
rect 6748 6390 6776 7890
rect 6840 6458 6868 8434
rect 7024 7834 7052 10406
rect 7300 9586 7328 10764
rect 7564 10746 7616 10752
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7116 7954 7144 9386
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8634 7236 9318
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7392 8090 7420 10134
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 7484 9722 7512 9862
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7576 9654 7604 10066
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7378 7984 7434 7993
rect 7104 7948 7156 7954
rect 7378 7919 7434 7928
rect 7104 7890 7156 7896
rect 7024 7806 7236 7834
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 7002 6960 7142
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6932 5930 6960 6734
rect 7024 6730 7052 7346
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6840 5902 6960 5930
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6288 4214 6316 4558
rect 6380 4554 6408 4626
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6182 4040 6238 4049
rect 6182 3975 6238 3984
rect 6196 2854 6224 3975
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6380 3058 6408 3538
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6092 2848 6144 2854
rect 6184 2848 6236 2854
rect 6092 2790 6144 2796
rect 6182 2816 6184 2825
rect 6236 2816 6238 2825
rect 6182 2751 6238 2760
rect 6472 480 6500 5850
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6564 4622 6592 5170
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6656 4146 6684 5646
rect 6748 5302 6776 5714
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6840 5114 6868 5902
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6748 5086 6868 5114
rect 6644 4140 6696 4146
rect 6644 4082 6696 4088
rect 6748 3126 6776 5086
rect 6932 5030 6960 5782
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6736 3120 6788 3126
rect 6736 3062 6788 3068
rect 6736 2984 6788 2990
rect 6736 2926 6788 2932
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6656 2106 6684 2858
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6748 2038 6776 2926
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6840 480 6868 4490
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6932 2961 6960 4082
rect 7024 3602 7052 6666
rect 7116 5846 7144 7346
rect 7208 6798 7236 7806
rect 7288 7200 7340 7206
rect 7288 7142 7340 7148
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6458 7236 6598
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 7300 6322 7328 7142
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7392 6066 7420 7919
rect 7300 6038 7420 6066
rect 7104 5840 7156 5846
rect 7104 5782 7156 5788
rect 7116 5234 7144 5782
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 7104 3460 7156 3466
rect 7104 3402 7156 3408
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6918 2952 6974 2961
rect 7024 2922 7052 3334
rect 6918 2887 6920 2896
rect 6972 2887 6974 2896
rect 7012 2916 7064 2922
rect 6920 2858 6972 2864
rect 7012 2858 7064 2864
rect 6932 2827 6960 2858
rect 7024 2514 7052 2858
rect 7116 2650 7144 3402
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7300 480 7328 6038
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7392 4185 7420 5238
rect 7484 4826 7512 9386
rect 7576 8906 7604 9590
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8498 7604 8842
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7576 8265 7604 8298
rect 7562 8256 7618 8265
rect 7562 8191 7618 8200
rect 7562 8120 7618 8129
rect 7562 8055 7564 8064
rect 7616 8055 7618 8064
rect 7564 8026 7616 8032
rect 7668 7562 7696 12650
rect 7820 12540 8116 12560
rect 7876 12538 7900 12540
rect 7956 12538 7980 12540
rect 8036 12538 8060 12540
rect 7898 12486 7900 12538
rect 7962 12486 7974 12538
rect 8036 12486 8038 12538
rect 7876 12484 7900 12486
rect 7956 12484 7980 12486
rect 8036 12484 8060 12486
rect 7820 12464 8116 12484
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 8208 12368 8260 12374
rect 8208 12310 8260 12316
rect 7748 11552 7800 11558
rect 7852 11540 7880 12310
rect 8022 11792 8078 11801
rect 8022 11727 8024 11736
rect 8076 11727 8078 11736
rect 8024 11698 8076 11704
rect 8220 11676 8248 12310
rect 8404 11830 8432 13194
rect 8496 12850 8524 13194
rect 9048 12986 9076 13330
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9036 12980 9088 12986
rect 9036 12922 9088 12928
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 9416 12714 9444 13126
rect 9784 12986 9812 13670
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12850 9812 12922
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9508 12628 9536 12786
rect 10324 12708 10376 12714
rect 10324 12650 10376 12656
rect 9588 12640 9640 12646
rect 9508 12600 9588 12628
rect 9588 12582 9640 12588
rect 8576 12300 8628 12306
rect 8576 12242 8628 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 8392 11824 8444 11830
rect 8392 11766 8444 11772
rect 8484 11688 8536 11694
rect 8220 11648 8340 11676
rect 8208 11552 8260 11558
rect 7852 11520 8208 11540
rect 8260 11520 8262 11529
rect 7852 11512 8206 11520
rect 7748 11494 7800 11500
rect 7760 11354 7788 11494
rect 7820 11452 8116 11472
rect 8206 11455 8262 11464
rect 7876 11450 7900 11452
rect 7956 11450 7980 11452
rect 8036 11450 8060 11452
rect 7898 11398 7900 11450
rect 7962 11398 7974 11450
rect 8036 11398 8038 11450
rect 7876 11396 7900 11398
rect 7956 11396 7980 11398
rect 8036 11396 8060 11398
rect 7820 11376 8116 11396
rect 8312 11354 8340 11648
rect 8484 11630 8536 11636
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8404 11286 8432 11494
rect 8392 11280 8444 11286
rect 8298 11248 8354 11257
rect 8392 11222 8444 11228
rect 8298 11183 8354 11192
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 7820 10364 8116 10384
rect 7876 10362 7900 10364
rect 7956 10362 7980 10364
rect 8036 10362 8060 10364
rect 7898 10310 7900 10362
rect 7962 10310 7974 10362
rect 8036 10310 8038 10362
rect 7876 10308 7900 10310
rect 7956 10308 7980 10310
rect 8036 10308 8060 10310
rect 7820 10288 8116 10308
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 7760 9586 7788 9930
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7852 9625 7880 9658
rect 7838 9616 7894 9625
rect 7748 9580 7800 9586
rect 7838 9551 7894 9560
rect 7748 9522 7800 9528
rect 7944 9364 7972 9930
rect 8220 9586 8248 11018
rect 8312 10266 8340 11183
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8404 9704 8432 10066
rect 8496 9994 8524 11630
rect 8588 11354 8616 12242
rect 10152 12209 10180 12242
rect 10232 12232 10284 12238
rect 10138 12200 10194 12209
rect 10232 12174 10284 12180
rect 10138 12135 10194 12144
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9496 11688 9548 11694
rect 8666 11656 8722 11665
rect 9496 11630 9548 11636
rect 8666 11591 8722 11600
rect 8680 11354 8708 11591
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 9036 11280 9088 11286
rect 9034 11248 9036 11257
rect 9088 11248 9090 11257
rect 8944 11212 8996 11218
rect 9034 11183 9090 11192
rect 8944 11154 8996 11160
rect 8956 11121 8984 11154
rect 8942 11112 8998 11121
rect 8942 11047 8998 11056
rect 8484 9988 8536 9994
rect 8484 9930 8536 9936
rect 8404 9676 8524 9704
rect 8496 9586 8524 9676
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 7760 9336 7972 9364
rect 8300 9376 8352 9382
rect 7760 8906 7788 9336
rect 8300 9318 8352 9324
rect 7820 9276 8116 9296
rect 7876 9274 7900 9276
rect 7956 9274 7980 9276
rect 8036 9274 8060 9276
rect 7898 9222 7900 9274
rect 7962 9222 7974 9274
rect 8036 9222 8038 9274
rect 7876 9220 7900 9222
rect 7956 9220 7980 9222
rect 8036 9220 8060 9222
rect 7820 9200 8116 9220
rect 8312 9110 8340 9318
rect 8300 9104 8352 9110
rect 8576 9104 8628 9110
rect 8300 9046 8352 9052
rect 8574 9072 8576 9081
rect 8628 9072 8630 9081
rect 9048 9058 9076 11183
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9324 10742 9352 11086
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9508 10130 9536 11630
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 10674 9628 11562
rect 10060 11558 10088 11698
rect 10244 11665 10272 12174
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10810 9720 11154
rect 10244 11150 10272 11494
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10152 10810 10180 11086
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9600 10266 9628 10610
rect 9864 10464 9916 10470
rect 9862 10432 9864 10441
rect 9956 10464 10008 10470
rect 9916 10432 9918 10441
rect 9956 10406 10008 10412
rect 9862 10367 9918 10376
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 8208 9036 8260 9042
rect 8574 9007 8630 9016
rect 8956 9030 9076 9058
rect 8208 8978 8260 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 8128 8498 8156 8910
rect 8220 8838 8248 8978
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7820 8188 8116 8208
rect 7876 8186 7900 8188
rect 7956 8186 7980 8188
rect 8036 8186 8060 8188
rect 7898 8134 7900 8186
rect 7962 8134 7974 8186
rect 8036 8134 8038 8186
rect 7876 8132 7900 8134
rect 7956 8132 7980 8134
rect 8036 8132 8060 8134
rect 7820 8112 8116 8132
rect 7668 7534 7788 7562
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 7378 4176 7434 4185
rect 7378 4111 7434 4120
rect 7392 2446 7420 4111
rect 7484 3670 7512 4558
rect 7576 4554 7604 6258
rect 7668 5370 7696 6734
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7668 4282 7696 5170
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 7562 3904 7618 3913
rect 7562 3839 7618 3848
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7576 3534 7604 3839
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7484 2650 7512 3470
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7576 2446 7604 2926
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7760 480 7788 7534
rect 8024 7404 8076 7410
rect 8076 7364 8156 7392
rect 8024 7346 8076 7352
rect 8128 7188 8156 7364
rect 8220 7342 8248 8774
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8312 7274 8340 8026
rect 8496 7342 8524 8366
rect 8588 8090 8616 8774
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8864 7546 8892 7958
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8128 7160 8248 7188
rect 7820 7100 8116 7120
rect 7876 7098 7900 7100
rect 7956 7098 7980 7100
rect 8036 7098 8060 7100
rect 7898 7046 7900 7098
rect 7962 7046 7974 7098
rect 8036 7046 8038 7098
rect 7876 7044 7900 7046
rect 7956 7044 7980 7046
rect 8036 7044 8060 7046
rect 7820 7024 8116 7044
rect 8220 6186 8248 7160
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8312 6186 8340 6734
rect 8496 6186 8524 7278
rect 8956 6746 8984 9030
rect 9036 8968 9088 8974
rect 9036 8910 9088 8916
rect 9048 7750 9076 8910
rect 9876 8906 9904 9386
rect 9864 8900 9916 8906
rect 9864 8842 9916 8848
rect 9876 8634 9904 8842
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 9312 8356 9364 8362
rect 9312 8298 9364 8304
rect 9140 7886 9168 8298
rect 9324 7993 9352 8298
rect 9692 8129 9720 8570
rect 9862 8528 9918 8537
rect 9862 8463 9918 8472
rect 9678 8120 9734 8129
rect 9678 8055 9734 8064
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9128 7880 9180 7886
rect 9128 7822 9180 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7342 9076 7686
rect 9140 7546 9168 7822
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9036 7336 9088 7342
rect 9036 7278 9088 7284
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9048 6934 9076 7278
rect 9036 6928 9088 6934
rect 9036 6870 9088 6876
rect 8956 6718 9168 6746
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8208 6180 8260 6186
rect 8208 6122 8260 6128
rect 8300 6180 8352 6186
rect 8484 6180 8536 6186
rect 8300 6122 8352 6128
rect 8404 6140 8484 6168
rect 7820 6012 8116 6032
rect 7876 6010 7900 6012
rect 7956 6010 7980 6012
rect 8036 6010 8060 6012
rect 7898 5958 7900 6010
rect 7962 5958 7974 6010
rect 8036 5958 8038 6010
rect 7876 5956 7900 5958
rect 7956 5956 7980 5958
rect 8036 5956 8060 5958
rect 7820 5936 8116 5956
rect 8220 5166 8248 6122
rect 8312 5574 8340 6122
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5234 8340 5510
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8300 5024 8352 5030
rect 8404 5012 8432 6140
rect 8484 6122 8536 6128
rect 8864 5914 8892 6394
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9048 5370 9076 5646
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 8850 5264 8906 5273
rect 8850 5199 8906 5208
rect 8352 4984 8432 5012
rect 8300 4966 8352 4972
rect 7820 4924 8116 4944
rect 7876 4922 7900 4924
rect 7956 4922 7980 4924
rect 8036 4922 8060 4924
rect 7898 4870 7900 4922
rect 7962 4870 7974 4922
rect 8036 4870 8038 4922
rect 7876 4868 7900 4870
rect 7956 4868 7980 4870
rect 8036 4868 8060 4870
rect 7820 4848 8116 4868
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 7944 4078 7972 4490
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 7820 3836 8116 3856
rect 7876 3834 7900 3836
rect 7956 3834 7980 3836
rect 8036 3834 8060 3836
rect 7898 3782 7900 3834
rect 7962 3782 7974 3834
rect 8036 3782 8038 3834
rect 7876 3780 7900 3782
rect 7956 3780 7980 3782
rect 8036 3780 8060 3782
rect 7820 3760 8116 3780
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3074 8156 3538
rect 8220 3194 8248 4014
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8128 3046 8248 3074
rect 7820 2748 8116 2768
rect 7876 2746 7900 2748
rect 7956 2746 7980 2748
rect 8036 2746 8060 2748
rect 7898 2694 7900 2746
rect 7962 2694 7974 2746
rect 8036 2694 8038 2746
rect 7876 2692 7900 2694
rect 7956 2692 7980 2694
rect 8036 2692 8060 2694
rect 7820 2672 8116 2692
rect 8220 480 8248 3046
rect 8312 2961 8340 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8390 3768 8446 3777
rect 8390 3703 8446 3712
rect 8404 3534 8432 3703
rect 8588 3602 8616 3839
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 8484 3120 8536 3126
rect 8588 3097 8616 3538
rect 8484 3062 8536 3068
rect 8574 3088 8630 3097
rect 8298 2952 8354 2961
rect 8298 2887 8354 2896
rect 8496 2514 8524 3062
rect 8574 3023 8630 3032
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8496 2106 8524 2450
rect 8484 2100 8536 2106
rect 8484 2042 8536 2048
rect 8588 2038 8616 2586
rect 8680 2310 8708 4558
rect 8772 4010 8800 4762
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8772 2122 8800 3946
rect 8864 3602 8892 5199
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8864 2446 8892 3402
rect 8956 3126 8984 3470
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9048 2990 9076 3334
rect 9036 2984 9088 2990
rect 9034 2952 9036 2961
rect 9088 2952 9090 2961
rect 9034 2887 9090 2896
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8680 2094 8800 2122
rect 8576 2032 8628 2038
rect 8576 1974 8628 1980
rect 8680 480 8708 2094
rect 9140 480 9168 6718
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9232 5710 9260 6054
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9324 2650 9352 7278
rect 9692 6769 9720 7890
rect 9770 7440 9826 7449
rect 9770 7375 9826 7384
rect 9678 6760 9734 6769
rect 9678 6695 9734 6704
rect 9784 6662 9812 7375
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9770 6352 9826 6361
rect 9404 6316 9456 6322
rect 9770 6287 9826 6296
rect 9404 6258 9456 6264
rect 9416 6186 9444 6258
rect 9494 6216 9550 6225
rect 9404 6180 9456 6186
rect 9494 6151 9550 6160
rect 9404 6122 9456 6128
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 4078 9444 5510
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9508 3380 9536 6151
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9586 5264 9642 5273
rect 9586 5199 9642 5208
rect 9600 5001 9628 5199
rect 9692 5166 9720 5510
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9680 5024 9732 5030
rect 9586 4992 9642 5001
rect 9680 4966 9732 4972
rect 9586 4927 9642 4936
rect 9692 4826 9720 4966
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4672 9812 6287
rect 9876 5930 9904 8463
rect 9968 7206 9996 10406
rect 10232 10124 10284 10130
rect 10232 10066 10284 10072
rect 10244 9722 10272 10066
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 7818 10088 8978
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10048 7812 10100 7818
rect 10048 7754 10100 7760
rect 10152 7546 10180 8910
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10244 7426 10272 9318
rect 10060 7398 10272 7426
rect 9956 7200 10008 7206
rect 9956 7142 10008 7148
rect 9876 5902 9996 5930
rect 9968 5642 9996 5902
rect 10060 5778 10088 7398
rect 10232 7336 10284 7342
rect 10232 7278 10284 7284
rect 10244 6934 10272 7278
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 10138 6760 10194 6769
rect 10138 6695 10140 6704
rect 10192 6695 10194 6704
rect 10140 6666 10192 6672
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9956 5160 10008 5166
rect 10060 5137 10088 5714
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 9956 5102 10008 5108
rect 10046 5128 10102 5137
rect 9692 4644 9812 4672
rect 9864 4684 9916 4690
rect 9692 4570 9720 4644
rect 9864 4626 9916 4632
rect 9600 4542 9720 4570
rect 9772 4548 9824 4554
rect 9600 3534 9628 4542
rect 9772 4490 9824 4496
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 3602 9720 4422
rect 9784 4146 9812 4490
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 3596 9732 3602
rect 9680 3538 9732 3544
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9508 3352 9628 3380
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9600 480 9628 3352
rect 9876 2650 9904 4626
rect 9968 3670 9996 5102
rect 10046 5063 10102 5072
rect 10140 5024 10192 5030
rect 10140 4966 10192 4972
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10060 4214 10088 4626
rect 10152 4622 10180 4966
rect 10244 4622 10272 5646
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 9956 3664 10008 3670
rect 9956 3606 10008 3612
rect 10060 3516 10088 3878
rect 10152 3738 10180 4558
rect 10244 4282 10272 4558
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 9968 3488 10088 3516
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9968 480 9996 3488
rect 10244 3398 10272 4014
rect 10336 3505 10364 12650
rect 10428 12646 10456 13670
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10520 12730 10548 12854
rect 10612 12850 10640 13194
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10520 12714 10640 12730
rect 10520 12708 10652 12714
rect 10520 12702 10600 12708
rect 10600 12650 10652 12656
rect 10416 12640 10468 12646
rect 10416 12582 10468 12588
rect 10428 7954 10456 12582
rect 10704 12306 10732 13874
rect 10980 13870 11008 14214
rect 11252 14172 11548 14192
rect 11308 14170 11332 14172
rect 11388 14170 11412 14172
rect 11468 14170 11492 14172
rect 11330 14118 11332 14170
rect 11394 14118 11406 14170
rect 11468 14118 11470 14170
rect 11308 14116 11332 14118
rect 11388 14116 11412 14118
rect 11468 14116 11492 14118
rect 11252 14096 11548 14116
rect 11808 13938 11836 14350
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10796 13326 10824 13806
rect 12070 13696 12126 13705
rect 12070 13631 12126 13640
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 10968 13388 11020 13394
rect 10968 13330 11020 13336
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10980 12986 11008 13330
rect 11252 13084 11548 13104
rect 11308 13082 11332 13084
rect 11388 13082 11412 13084
rect 11468 13082 11492 13084
rect 11330 13030 11332 13082
rect 11394 13030 11406 13082
rect 11468 13030 11470 13082
rect 11308 13028 11332 13030
rect 11388 13028 11412 13030
rect 11468 13028 11492 13030
rect 11252 13008 11548 13028
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10692 12300 10744 12306
rect 10612 12260 10692 12288
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11393 10548 12106
rect 10506 11384 10562 11393
rect 10506 11319 10562 11328
rect 10612 11150 10640 12260
rect 10692 12242 10744 12248
rect 11150 12200 11206 12209
rect 11150 12135 11206 12144
rect 10782 11792 10838 11801
rect 10782 11727 10838 11736
rect 10690 11520 10746 11529
rect 10690 11455 10746 11464
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10508 10464 10560 10470
rect 10508 10406 10560 10412
rect 10520 9722 10548 10406
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10520 8362 10548 8842
rect 10704 8537 10732 11455
rect 10796 11286 10824 11727
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10796 9586 10824 10134
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10888 9518 10916 11290
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10966 10024 11022 10033
rect 10966 9959 11022 9968
rect 10980 9926 11008 9959
rect 10968 9920 11020 9926
rect 10968 9862 11020 9868
rect 10966 9616 11022 9625
rect 10966 9551 11022 9560
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10888 8838 10916 9454
rect 10980 9382 11008 9551
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10690 8528 10746 8537
rect 10690 8463 10746 8472
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10508 8356 10560 8362
rect 10508 8298 10560 8304
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10416 7948 10468 7954
rect 10416 7890 10468 7896
rect 10520 7290 10548 8026
rect 10428 7262 10548 7290
rect 10428 4049 10456 7262
rect 10508 7200 10560 7206
rect 10612 7177 10640 8366
rect 10508 7142 10560 7148
rect 10598 7168 10654 7177
rect 10520 7002 10548 7142
rect 10598 7103 10654 7112
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10508 6724 10560 6730
rect 10508 6666 10560 6672
rect 10520 6361 10548 6666
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5914 10640 6054
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10612 4826 10640 5238
rect 10704 5030 10732 8463
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10414 4040 10470 4049
rect 10414 3975 10470 3984
rect 10414 3768 10470 3777
rect 10704 3738 10732 4422
rect 10414 3703 10470 3712
rect 10692 3732 10744 3738
rect 10322 3496 10378 3505
rect 10322 3431 10378 3440
rect 10232 3392 10284 3398
rect 10284 3352 10364 3380
rect 10232 3334 10284 3340
rect 10244 3269 10272 3334
rect 10336 2990 10364 3352
rect 10232 2984 10284 2990
rect 10232 2926 10284 2932
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 10244 2650 10272 2926
rect 10324 2848 10376 2854
rect 10324 2790 10376 2796
rect 10336 2650 10364 2790
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10428 480 10456 3703
rect 10692 3674 10744 3680
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 2854 10640 3334
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 10796 2514 10824 8774
rect 10876 8016 10928 8022
rect 10876 7958 10928 7964
rect 10888 6905 10916 7958
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10888 6089 10916 6831
rect 10874 6080 10930 6089
rect 10874 6015 10930 6024
rect 10874 5808 10930 5817
rect 10874 5743 10930 5752
rect 10888 5642 10916 5743
rect 10876 5636 10928 5642
rect 10876 5578 10928 5584
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10888 3670 10916 4966
rect 10876 3664 10928 3670
rect 10876 3606 10928 3612
rect 10874 3496 10930 3505
rect 10874 3431 10930 3440
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10888 480 10916 3431
rect 10980 2961 11008 8978
rect 11072 7274 11100 10066
rect 11164 8480 11192 12135
rect 11252 11996 11548 12016
rect 11308 11994 11332 11996
rect 11388 11994 11412 11996
rect 11468 11994 11492 11996
rect 11330 11942 11332 11994
rect 11394 11942 11406 11994
rect 11468 11942 11470 11994
rect 11308 11940 11332 11942
rect 11388 11940 11412 11942
rect 11468 11940 11492 11942
rect 11252 11920 11548 11940
rect 11624 11694 11652 13398
rect 11796 13320 11848 13326
rect 11794 13288 11796 13297
rect 11848 13288 11850 13297
rect 11794 13223 11850 13232
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11610 11112 11666 11121
rect 11610 11047 11666 11056
rect 11252 10908 11548 10928
rect 11308 10906 11332 10908
rect 11388 10906 11412 10908
rect 11468 10906 11492 10908
rect 11330 10854 11332 10906
rect 11394 10854 11406 10906
rect 11468 10854 11470 10906
rect 11308 10852 11332 10854
rect 11388 10852 11412 10854
rect 11468 10852 11492 10854
rect 11252 10832 11548 10852
rect 11624 10305 11652 11047
rect 11716 10606 11744 12038
rect 11808 11898 11836 12242
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11900 11286 11928 12106
rect 11888 11280 11940 11286
rect 11888 11222 11940 11228
rect 11900 10674 11928 11222
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11610 10296 11666 10305
rect 11610 10231 11666 10240
rect 11716 10130 11744 10406
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11252 9820 11548 9840
rect 11308 9818 11332 9820
rect 11388 9818 11412 9820
rect 11468 9818 11492 9820
rect 11330 9766 11332 9818
rect 11394 9766 11406 9818
rect 11468 9766 11470 9818
rect 11308 9764 11332 9766
rect 11388 9764 11412 9766
rect 11468 9764 11492 9766
rect 11252 9744 11548 9764
rect 11704 9376 11756 9382
rect 11704 9318 11756 9324
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11252 8732 11548 8752
rect 11308 8730 11332 8732
rect 11388 8730 11412 8732
rect 11468 8730 11492 8732
rect 11330 8678 11332 8730
rect 11394 8678 11406 8730
rect 11468 8678 11470 8730
rect 11308 8676 11332 8678
rect 11388 8676 11412 8678
rect 11468 8676 11492 8678
rect 11252 8656 11548 8676
rect 11164 8452 11284 8480
rect 11150 8392 11206 8401
rect 11150 8327 11206 8336
rect 11164 7954 11192 8327
rect 11256 8276 11284 8452
rect 11624 8401 11652 9046
rect 11716 8906 11744 9318
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11610 8392 11666 8401
rect 11610 8327 11666 8336
rect 11256 8248 11744 8276
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11252 7644 11548 7664
rect 11308 7642 11332 7644
rect 11388 7642 11412 7644
rect 11468 7642 11492 7644
rect 11330 7590 11332 7642
rect 11394 7590 11406 7642
rect 11468 7590 11470 7642
rect 11308 7588 11332 7590
rect 11388 7588 11412 7590
rect 11468 7588 11492 7590
rect 11252 7568 11548 7588
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11060 7268 11112 7274
rect 11060 7210 11112 7216
rect 11164 6866 11192 7346
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6254 11100 6734
rect 11164 6390 11192 6802
rect 11252 6556 11548 6576
rect 11308 6554 11332 6556
rect 11388 6554 11412 6556
rect 11468 6554 11492 6556
rect 11330 6502 11332 6554
rect 11394 6502 11406 6554
rect 11468 6502 11470 6554
rect 11308 6500 11332 6502
rect 11388 6500 11412 6502
rect 11468 6500 11492 6502
rect 11252 6480 11548 6500
rect 11152 6384 11204 6390
rect 11152 6326 11204 6332
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11058 6080 11114 6089
rect 11242 6080 11298 6089
rect 11058 6015 11114 6024
rect 11164 6038 11242 6066
rect 11072 4706 11100 6015
rect 11164 4826 11192 6038
rect 11242 6015 11298 6024
rect 11244 5704 11296 5710
rect 11348 5692 11376 6326
rect 11296 5664 11376 5692
rect 11244 5646 11296 5652
rect 11252 5468 11548 5488
rect 11308 5466 11332 5468
rect 11388 5466 11412 5468
rect 11468 5466 11492 5468
rect 11330 5414 11332 5466
rect 11394 5414 11406 5466
rect 11468 5414 11470 5466
rect 11308 5412 11332 5414
rect 11388 5412 11412 5414
rect 11468 5412 11492 5414
rect 11252 5392 11548 5412
rect 11624 5352 11652 7890
rect 11716 7206 11744 8248
rect 11808 7886 11836 10406
rect 11886 10296 11942 10305
rect 11992 10266 12020 12582
rect 11886 10231 11942 10240
rect 11980 10260 12032 10266
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11704 7200 11756 7206
rect 11704 7142 11756 7148
rect 11532 5324 11652 5352
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11532 4758 11560 5324
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11520 4752 11572 4758
rect 11072 4678 11192 4706
rect 11520 4694 11572 4700
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4078 11100 4558
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10966 2952 11022 2961
rect 10966 2887 11022 2896
rect 11164 2020 11192 4678
rect 11252 4380 11548 4400
rect 11308 4378 11332 4380
rect 11388 4378 11412 4380
rect 11468 4378 11492 4380
rect 11330 4326 11332 4378
rect 11394 4326 11406 4378
rect 11468 4326 11470 4378
rect 11308 4324 11332 4326
rect 11388 4324 11412 4326
rect 11468 4324 11492 4326
rect 11252 4304 11548 4324
rect 11624 4282 11652 4966
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11334 4040 11390 4049
rect 11334 3975 11390 3984
rect 11520 4004 11572 4010
rect 11348 3942 11376 3975
rect 11520 3946 11572 3952
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11532 3738 11560 3946
rect 11612 3936 11664 3942
rect 11716 3913 11744 7142
rect 11808 6866 11836 7822
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11808 5302 11836 6802
rect 11900 6458 11928 10231
rect 11980 10202 12032 10208
rect 12084 8906 12112 13631
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12442 12480 12718
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10577 12296 10950
rect 12360 10606 12388 11562
rect 12440 11280 12492 11286
rect 12438 11248 12440 11257
rect 12492 11248 12494 11257
rect 12438 11183 12494 11192
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12452 10674 12480 10950
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12348 10600 12400 10606
rect 12254 10568 12310 10577
rect 12348 10542 12400 10548
rect 12254 10503 12310 10512
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 12070 8664 12126 8673
rect 12176 8634 12204 9998
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 12348 9988 12400 9994
rect 12348 9930 12400 9936
rect 12070 8599 12126 8608
rect 12164 8628 12216 8634
rect 11980 8288 12032 8294
rect 11980 8230 12032 8236
rect 11992 7585 12020 8230
rect 12084 8090 12112 8599
rect 12164 8570 12216 8576
rect 12162 8392 12218 8401
rect 12162 8327 12218 8336
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12176 7970 12204 8327
rect 12268 8294 12296 9930
rect 12360 9722 12388 9930
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12348 9512 12400 9518
rect 12452 9466 12480 10610
rect 12544 10266 12572 15506
rect 15384 15088 15436 15094
rect 15384 15030 15436 15036
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14096 14884 14148 14890
rect 14096 14826 14148 14832
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 12716 14272 12768 14278
rect 12716 14214 12768 14220
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 12728 12646 12756 14214
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 12808 13320 12860 13326
rect 12808 13262 12860 13268
rect 12820 12782 12848 13262
rect 13004 12850 13032 13942
rect 13084 13932 13136 13938
rect 13084 13874 13136 13880
rect 13096 13394 13124 13874
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 13360 13388 13412 13394
rect 13412 13348 13492 13376
rect 13360 13330 13412 13336
rect 12992 12844 13044 12850
rect 12912 12804 12992 12832
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12728 11830 12756 12582
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12820 11694 12848 12038
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12820 11150 12848 11290
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10554 12848 10950
rect 12636 10538 12848 10554
rect 12624 10532 12848 10538
rect 12676 10526 12848 10532
rect 12624 10474 12676 10480
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12912 10146 12940 12804
rect 12992 12786 13044 12792
rect 13096 11898 13124 13330
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13004 11354 13032 11698
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 13004 10606 13032 11290
rect 13096 11218 13124 11834
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12992 10600 13044 10606
rect 12992 10542 13044 10548
rect 13188 10305 13216 12174
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13174 10296 13230 10305
rect 13084 10260 13136 10266
rect 13174 10231 13230 10240
rect 13084 10202 13136 10208
rect 12636 10118 12940 10146
rect 12636 9722 12664 10118
rect 12716 10056 12768 10062
rect 12716 9998 12768 10004
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12400 9460 12480 9466
rect 12348 9454 12480 9460
rect 12360 9438 12480 9454
rect 12728 9450 12756 9998
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12532 9444 12584 9450
rect 12532 9386 12584 9392
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8412 12388 8842
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12452 8537 12480 8570
rect 12438 8528 12494 8537
rect 12438 8463 12494 8472
rect 12360 8384 12480 8412
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12254 8120 12310 8129
rect 12310 8078 12388 8106
rect 12254 8055 12310 8064
rect 12360 8022 12388 8078
rect 12084 7942 12204 7970
rect 12348 8016 12400 8022
rect 12348 7958 12400 7964
rect 11978 7576 12034 7585
rect 11978 7511 12034 7520
rect 12084 7154 12112 7942
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 11992 7126 12112 7154
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 6390 12020 7126
rect 12176 6984 12204 7822
rect 12452 7342 12480 8384
rect 12544 8022 12572 9386
rect 12728 9178 12756 9386
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 8430 12664 8978
rect 12714 8936 12770 8945
rect 12714 8871 12770 8880
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12728 8362 12756 8871
rect 12820 8498 12848 9658
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12532 8016 12584 8022
rect 12532 7958 12584 7964
rect 12806 7984 12862 7993
rect 12806 7919 12808 7928
rect 12860 7919 12862 7928
rect 12808 7890 12860 7896
rect 12716 7880 12768 7886
rect 13004 7868 13032 8434
rect 13096 8090 13124 10202
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13188 8498 13216 8978
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13176 8356 13228 8362
rect 13176 8298 13228 8304
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13084 7880 13136 7886
rect 13004 7840 13084 7868
rect 12716 7822 12768 7828
rect 13084 7822 13136 7828
rect 12728 7721 12756 7822
rect 12808 7744 12860 7750
rect 12714 7712 12770 7721
rect 12808 7686 12860 7692
rect 12714 7647 12770 7656
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12084 6956 12204 6984
rect 12256 6996 12308 7002
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 12084 6322 12112 6956
rect 12256 6938 12308 6944
rect 12268 6769 12296 6938
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12070 5944 12126 5953
rect 12070 5879 12126 5888
rect 12084 5778 12112 5879
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11888 5704 11940 5710
rect 11886 5672 11888 5681
rect 11980 5704 12032 5710
rect 11940 5672 11942 5681
rect 12032 5652 12112 5658
rect 11980 5646 12112 5652
rect 11992 5630 12112 5646
rect 11886 5607 11942 5616
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11612 3878 11664 3884
rect 11702 3904 11758 3913
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11624 3534 11652 3878
rect 11702 3839 11758 3848
rect 11808 3754 11836 4626
rect 11900 4146 11928 5034
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 11886 3768 11942 3777
rect 11808 3726 11886 3754
rect 11886 3703 11888 3712
rect 11940 3703 11942 3712
rect 11888 3674 11940 3680
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11252 3292 11548 3312
rect 11308 3290 11332 3292
rect 11388 3290 11412 3292
rect 11468 3290 11492 3292
rect 11330 3238 11332 3290
rect 11394 3238 11406 3290
rect 11468 3238 11470 3290
rect 11308 3236 11332 3238
rect 11388 3236 11412 3238
rect 11468 3236 11492 3238
rect 11252 3216 11548 3236
rect 11624 2922 11652 3470
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11252 2204 11548 2224
rect 11308 2202 11332 2204
rect 11388 2202 11412 2204
rect 11468 2202 11492 2204
rect 11330 2150 11332 2202
rect 11394 2150 11406 2202
rect 11468 2150 11470 2202
rect 11308 2148 11332 2150
rect 11388 2148 11412 2150
rect 11468 2148 11492 2150
rect 11252 2128 11548 2148
rect 11164 1992 11376 2020
rect 11348 480 11376 1992
rect 11808 480 11836 3062
rect 11992 2922 12020 5510
rect 12084 5302 12112 5630
rect 12176 5545 12204 5782
rect 12162 5536 12218 5545
rect 12162 5471 12218 5480
rect 12072 5296 12124 5302
rect 12072 5238 12124 5244
rect 12070 5128 12126 5137
rect 12070 5063 12126 5072
rect 12084 4826 12112 5063
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 12176 3534 12204 4558
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12268 3126 12296 6122
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12360 2972 12388 6394
rect 12440 6248 12492 6254
rect 12440 6190 12492 6196
rect 12452 5846 12480 6190
rect 12440 5840 12492 5846
rect 12440 5782 12492 5788
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12452 5370 12480 5510
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12544 5080 12572 7142
rect 12636 6662 12664 7346
rect 12820 7342 12848 7686
rect 13188 7342 13216 8298
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 13176 7336 13228 7342
rect 13176 7278 13228 7284
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12728 6769 12756 7210
rect 12808 7200 12860 7206
rect 12808 7142 12860 7148
rect 12714 6760 12770 6769
rect 12714 6695 12770 6704
rect 12624 6656 12676 6662
rect 12676 6604 12756 6610
rect 12624 6598 12756 6604
rect 12636 6582 12756 6598
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12636 6225 12664 6394
rect 12728 6254 12756 6582
rect 12716 6248 12768 6254
rect 12622 6216 12678 6225
rect 12716 6190 12768 6196
rect 12622 6151 12678 6160
rect 12716 5636 12768 5642
rect 12820 5624 12848 7142
rect 12912 6662 12940 7278
rect 12900 6656 12952 6662
rect 12900 6598 12952 6604
rect 12912 5846 12940 6598
rect 13174 6352 13230 6361
rect 13174 6287 13230 6296
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12900 5840 12952 5846
rect 12900 5782 12952 5788
rect 13004 5778 13032 6054
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13096 5817 13124 5850
rect 13082 5808 13138 5817
rect 12992 5772 13044 5778
rect 13082 5743 13138 5752
rect 12992 5714 13044 5720
rect 13004 5681 13032 5714
rect 12768 5596 12848 5624
rect 12990 5672 13046 5681
rect 12990 5607 13046 5616
rect 12716 5578 12768 5584
rect 12716 5296 12768 5302
rect 12716 5238 12768 5244
rect 12544 5052 12664 5080
rect 12530 4312 12586 4321
rect 12530 4247 12532 4256
rect 12584 4247 12586 4256
rect 12532 4218 12584 4224
rect 12440 4208 12492 4214
rect 12438 4176 12440 4185
rect 12492 4176 12494 4185
rect 12438 4111 12494 4120
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12268 2944 12388 2972
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 12268 480 12296 2944
rect 12544 2514 12572 3334
rect 12636 2990 12664 5052
rect 12728 4622 12756 5238
rect 13004 5234 13032 5607
rect 12992 5228 13044 5234
rect 12992 5170 13044 5176
rect 13188 5166 13216 6287
rect 13176 5160 13228 5166
rect 13176 5102 13228 5108
rect 12992 5024 13044 5030
rect 12992 4966 13044 4972
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12900 4480 12952 4486
rect 12900 4422 12952 4428
rect 12912 4146 12940 4422
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12728 480 12756 3130
rect 13004 2122 13032 4966
rect 13084 3528 13136 3534
rect 13084 3470 13136 3476
rect 13096 2854 13124 3470
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13280 2514 13308 11086
rect 13372 10130 13400 11494
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13358 9480 13414 9489
rect 13464 9450 13492 13348
rect 13648 11218 13676 14214
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13820 11688 13872 11694
rect 13820 11630 13872 11636
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13544 11008 13596 11014
rect 13544 10950 13596 10956
rect 13358 9415 13414 9424
rect 13452 9444 13504 9450
rect 13372 7177 13400 9415
rect 13452 9386 13504 9392
rect 13556 8294 13584 10950
rect 13648 10674 13676 11154
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13832 10266 13860 11630
rect 13924 11218 13952 12135
rect 14016 11540 14044 14486
rect 14108 12986 14136 14826
rect 14188 14816 14240 14822
rect 14188 14758 14240 14764
rect 14200 14618 14228 14758
rect 14188 14612 14240 14618
rect 14188 14554 14240 14560
rect 14292 13462 14320 14826
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 13870 14504 14350
rect 14568 14074 14596 14962
rect 14684 14716 14980 14736
rect 14740 14714 14764 14716
rect 14820 14714 14844 14716
rect 14900 14714 14924 14716
rect 14762 14662 14764 14714
rect 14826 14662 14838 14714
rect 14900 14662 14902 14714
rect 14740 14660 14764 14662
rect 14820 14660 14844 14662
rect 14900 14660 14924 14662
rect 14684 14640 14980 14660
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12782 14228 13262
rect 14292 12850 14320 13398
rect 14476 13190 14504 13806
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 14568 13530 14596 13738
rect 14684 13628 14980 13648
rect 14740 13626 14764 13628
rect 14820 13626 14844 13628
rect 14900 13626 14924 13628
rect 14762 13574 14764 13626
rect 14826 13574 14838 13626
rect 14900 13574 14902 13626
rect 14740 13572 14764 13574
rect 14820 13572 14844 13574
rect 14900 13572 14924 13574
rect 14684 13552 14980 13572
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12850 14504 13126
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 15108 12708 15160 12714
rect 15108 12650 15160 12656
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 14684 12540 14980 12560
rect 14740 12538 14764 12540
rect 14820 12538 14844 12540
rect 14900 12538 14924 12540
rect 14762 12486 14764 12538
rect 14826 12486 14838 12538
rect 14900 12486 14902 12538
rect 14740 12484 14764 12486
rect 14820 12484 14844 12486
rect 14900 12484 14924 12486
rect 14684 12464 14980 12484
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14016 11512 14136 11540
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13912 10464 13964 10470
rect 13910 10432 13912 10441
rect 13964 10432 13966 10441
rect 13910 10367 13966 10376
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13358 7168 13414 7177
rect 13358 7103 13414 7112
rect 13372 5030 13400 7103
rect 13464 6089 13492 8026
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13556 6361 13584 7890
rect 13648 6798 13676 9862
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13542 6352 13598 6361
rect 13542 6287 13598 6296
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13360 4616 13412 4622
rect 13464 4604 13492 5782
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13412 4576 13492 4604
rect 13360 4558 13412 4564
rect 13372 4078 13400 4558
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13556 3777 13584 5102
rect 13648 4758 13676 5510
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13542 3768 13598 3777
rect 13542 3703 13598 3712
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 2514 13584 2858
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13648 2258 13676 4422
rect 13740 3602 13768 9998
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13832 9042 13860 9318
rect 14016 9110 14044 10066
rect 14004 9104 14056 9110
rect 14004 9046 14056 9052
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8362 13860 8978
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13832 7970 13860 8298
rect 13924 8090 13952 8910
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8084 13964 8090
rect 13912 8026 13964 8032
rect 13832 7954 13952 7970
rect 13832 7948 13964 7954
rect 13832 7942 13912 7948
rect 13832 6934 13860 7942
rect 13912 7890 13964 7896
rect 14016 7886 14044 8366
rect 14108 8022 14136 11512
rect 14476 11150 14504 12242
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11694 14780 12174
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14684 11452 14980 11472
rect 14740 11450 14764 11452
rect 14820 11450 14844 11452
rect 14900 11450 14924 11452
rect 14762 11398 14764 11450
rect 14826 11398 14838 11450
rect 14900 11398 14902 11450
rect 14740 11396 14764 11398
rect 14820 11396 14844 11398
rect 14900 11396 14924 11398
rect 14684 11376 14980 11396
rect 15028 11150 15056 11834
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14684 10364 14980 10384
rect 14740 10362 14764 10364
rect 14820 10362 14844 10364
rect 14900 10362 14924 10364
rect 14762 10310 14764 10362
rect 14826 10310 14838 10362
rect 14900 10310 14902 10362
rect 14740 10308 14764 10310
rect 14820 10308 14844 10310
rect 14900 10308 14924 10310
rect 14684 10288 14980 10308
rect 14464 10192 14516 10198
rect 14370 10160 14426 10169
rect 14464 10134 14516 10140
rect 14370 10095 14426 10104
rect 14278 10024 14334 10033
rect 14278 9959 14334 9968
rect 14188 9444 14240 9450
rect 14188 9386 14240 9392
rect 14096 8016 14148 8022
rect 14096 7958 14148 7964
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13820 6928 13872 6934
rect 13820 6870 13872 6876
rect 13924 6798 13952 7210
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 14016 6730 14044 7210
rect 14004 6724 14056 6730
rect 14004 6666 14056 6672
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13832 5710 13860 5879
rect 14004 5772 14056 5778
rect 14004 5714 14056 5720
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 14016 5545 14044 5714
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 13820 5296 13872 5302
rect 13820 5238 13872 5244
rect 13832 4321 13860 5238
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13818 4312 13874 4321
rect 13818 4247 13874 4256
rect 13924 3641 13952 5034
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 14016 3670 14044 4966
rect 14108 4049 14136 7822
rect 14200 7528 14228 9386
rect 14292 7857 14320 9959
rect 14278 7848 14334 7857
rect 14278 7783 14334 7792
rect 14280 7540 14332 7546
rect 14200 7500 14280 7528
rect 14280 7482 14332 7488
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14186 5808 14242 5817
rect 14186 5743 14242 5752
rect 14200 5001 14228 5743
rect 14292 5642 14320 6190
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14384 5114 14412 10095
rect 14476 8378 14504 10134
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 9178 14596 9318
rect 14684 9276 14980 9296
rect 14740 9274 14764 9276
rect 14820 9274 14844 9276
rect 14900 9274 14924 9276
rect 14762 9222 14764 9274
rect 14826 9222 14838 9274
rect 14900 9222 14902 9274
rect 14740 9220 14764 9222
rect 14820 9220 14844 9222
rect 14900 9220 14924 9222
rect 14684 9200 14980 9220
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8566 14872 8910
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 14554 8392 14610 8401
rect 14476 8350 14554 8378
rect 14554 8327 14610 8336
rect 14568 8090 14596 8327
rect 14684 8188 14980 8208
rect 14740 8186 14764 8188
rect 14820 8186 14844 8188
rect 14900 8186 14924 8188
rect 14762 8134 14764 8186
rect 14826 8134 14838 8186
rect 14900 8134 14902 8186
rect 14740 8132 14764 8134
rect 14820 8132 14844 8134
rect 14900 8132 14924 8134
rect 14684 8112 14980 8132
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 15028 7970 15056 11086
rect 15120 10742 15148 12650
rect 15212 12442 15240 12650
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 10266 15148 10542
rect 15304 10266 15332 11290
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15108 9444 15160 9450
rect 15108 9386 15160 9392
rect 15120 8566 15148 9386
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 14476 7942 15056 7970
rect 15212 7954 15240 10066
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9178 15332 9318
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15200 7948 15252 7954
rect 14476 5302 14504 7942
rect 15200 7890 15252 7896
rect 15304 7886 15332 8910
rect 15292 7880 15344 7886
rect 14554 7848 14610 7857
rect 15292 7822 15344 7828
rect 14554 7783 14610 7792
rect 14568 6882 14596 7783
rect 14646 7712 14702 7721
rect 14646 7647 14702 7656
rect 14660 7478 14688 7647
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14844 7274 15240 7290
rect 14832 7268 15252 7274
rect 14884 7262 15200 7268
rect 14832 7210 14884 7216
rect 15200 7210 15252 7216
rect 15108 7200 15160 7206
rect 15028 7160 15108 7188
rect 14684 7100 14980 7120
rect 14740 7098 14764 7100
rect 14820 7098 14844 7100
rect 14900 7098 14924 7100
rect 14762 7046 14764 7098
rect 14826 7046 14838 7098
rect 14900 7046 14902 7098
rect 14740 7044 14764 7046
rect 14820 7044 14844 7046
rect 14900 7044 14924 7046
rect 14684 7024 14980 7044
rect 14568 6866 14688 6882
rect 14568 6860 14700 6866
rect 14568 6854 14648 6860
rect 14648 6802 14700 6808
rect 14556 6792 14608 6798
rect 14740 6792 14792 6798
rect 14608 6740 14740 6746
rect 14556 6734 14792 6740
rect 14568 6718 14780 6734
rect 14556 6112 14608 6118
rect 14752 6100 14780 6718
rect 14608 6072 14780 6100
rect 14556 6054 14608 6060
rect 14684 6012 14980 6032
rect 14740 6010 14764 6012
rect 14820 6010 14844 6012
rect 14900 6010 14924 6012
rect 14762 5958 14764 6010
rect 14826 5958 14838 6010
rect 14900 5958 14902 6010
rect 14740 5956 14764 5958
rect 14820 5956 14844 5958
rect 14900 5956 14924 5958
rect 14684 5936 14980 5956
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14292 5086 14412 5114
rect 14292 5030 14320 5086
rect 14280 5024 14332 5030
rect 14186 4992 14242 5001
rect 14280 4966 14332 4972
rect 14186 4927 14242 4936
rect 14568 4486 14596 5170
rect 14684 4924 14980 4944
rect 14740 4922 14764 4924
rect 14820 4922 14844 4924
rect 14900 4922 14924 4924
rect 14762 4870 14764 4922
rect 14826 4870 14838 4922
rect 14900 4870 14902 4922
rect 14740 4868 14764 4870
rect 14820 4868 14844 4870
rect 14900 4868 14924 4870
rect 14684 4848 14980 4868
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14384 3738 14412 3946
rect 14568 3942 14596 4422
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14004 3664 14056 3670
rect 13910 3632 13966 3641
rect 13728 3596 13780 3602
rect 14004 3606 14056 3612
rect 14568 3602 14596 3878
rect 14684 3836 14980 3856
rect 14740 3834 14764 3836
rect 14820 3834 14844 3836
rect 14900 3834 14924 3836
rect 14762 3782 14764 3834
rect 14826 3782 14838 3834
rect 14900 3782 14902 3834
rect 14740 3780 14764 3782
rect 14820 3780 14844 3782
rect 14900 3780 14924 3782
rect 14684 3760 14980 3780
rect 15028 3618 15056 7160
rect 15108 7142 15160 7148
rect 15108 6180 15160 6186
rect 15108 6122 15160 6128
rect 15120 3942 15148 6122
rect 15198 4856 15254 4865
rect 15198 4791 15200 4800
rect 15252 4791 15254 4800
rect 15200 4762 15252 4768
rect 15292 4684 15344 4690
rect 15292 4626 15344 4632
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 13910 3567 13966 3576
rect 14556 3596 14608 3602
rect 13728 3538 13780 3544
rect 14556 3538 14608 3544
rect 14936 3590 15056 3618
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 2990 14136 3334
rect 14936 2990 14964 3590
rect 15120 3534 15148 3878
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15016 3460 15068 3466
rect 15016 3402 15068 3408
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14464 2916 14516 2922
rect 14464 2858 14516 2864
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13556 2230 13676 2258
rect 13004 2094 13216 2122
rect 13188 480 13216 2094
rect 13556 480 13584 2230
rect 14016 480 14044 2586
rect 14476 2514 14504 2858
rect 14684 2748 14980 2768
rect 14740 2746 14764 2748
rect 14820 2746 14844 2748
rect 14900 2746 14924 2748
rect 14762 2694 14764 2746
rect 14826 2694 14838 2746
rect 14900 2694 14902 2746
rect 14740 2692 14764 2694
rect 14820 2692 14844 2694
rect 14900 2692 14924 2694
rect 14684 2672 14980 2692
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 1170 14412 2314
rect 15028 1714 15056 3402
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 15212 2514 15240 2858
rect 15304 2854 15332 4626
rect 15396 2990 15424 15030
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14550 16252 14758
rect 16212 14544 16264 14550
rect 16212 14486 16264 14492
rect 16948 14544 17000 14550
rect 16948 14486 17000 14492
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 13802 15608 14282
rect 16316 13818 16344 14350
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 16224 13790 16344 13818
rect 16776 13802 16804 14214
rect 16960 13938 16988 14486
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16764 13796 16816 13802
rect 15580 13394 15608 13738
rect 16224 13734 16252 13790
rect 16764 13738 16816 13744
rect 15936 13728 15988 13734
rect 15936 13670 15988 13676
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 11762 15608 13330
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15856 11626 15884 12786
rect 15948 12782 15976 13670
rect 16224 13462 16252 13670
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 16224 12850 16252 13398
rect 16592 12986 16620 13670
rect 16960 13530 16988 13874
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17144 13462 17172 22320
rect 18116 19612 18412 19632
rect 18172 19610 18196 19612
rect 18252 19610 18276 19612
rect 18332 19610 18356 19612
rect 18194 19558 18196 19610
rect 18258 19558 18270 19610
rect 18332 19558 18334 19610
rect 18172 19556 18196 19558
rect 18252 19556 18276 19558
rect 18332 19556 18356 19558
rect 18116 19536 18412 19556
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18432 18902 18460 19246
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17866 16960 17922 16969
rect 17866 16895 17922 16904
rect 17880 16250 17908 16895
rect 17868 16244 17920 16250
rect 17868 16186 17920 16192
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17512 13802 17540 14418
rect 17500 13796 17552 13802
rect 17500 13738 17552 13744
rect 17592 13796 17644 13802
rect 17592 13738 17644 13744
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17130 13288 17186 13297
rect 17130 13223 17186 13232
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 15936 12776 15988 12782
rect 15936 12718 15988 12724
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 15948 12442 15976 12582
rect 15936 12436 15988 12442
rect 15936 12378 15988 12384
rect 16028 12436 16080 12442
rect 16028 12378 16080 12384
rect 16040 12322 16068 12378
rect 15948 12294 16068 12322
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16120 12300 16172 12306
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15566 11248 15622 11257
rect 15566 11183 15622 11192
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 10198 15516 10406
rect 15476 10192 15528 10198
rect 15476 10134 15528 10140
rect 15580 9602 15608 11183
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15764 10810 15792 11086
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15672 10130 15700 10610
rect 15750 10568 15806 10577
rect 15750 10503 15752 10512
rect 15804 10503 15806 10512
rect 15752 10474 15804 10480
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15856 10062 15884 11562
rect 15948 11286 15976 12294
rect 16120 12242 16172 12248
rect 16132 11354 16160 12242
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15844 10056 15896 10062
rect 15844 9998 15896 10004
rect 15488 9574 15608 9602
rect 15660 9580 15712 9586
rect 15488 9382 15516 9574
rect 15660 9522 15712 9528
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15672 9178 15700 9522
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15764 9110 15792 9522
rect 15752 9104 15804 9110
rect 15752 9046 15804 9052
rect 15948 8537 15976 11222
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 16040 10674 16068 11086
rect 16028 10668 16080 10674
rect 16028 10610 16080 10616
rect 16028 9172 16080 9178
rect 16028 9114 16080 9120
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15568 8356 15620 8362
rect 15568 8298 15620 8304
rect 15474 7576 15530 7585
rect 15474 7511 15530 7520
rect 15488 6934 15516 7511
rect 15580 7449 15608 8298
rect 16040 8022 16068 9114
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16028 8016 16080 8022
rect 16028 7958 16080 7964
rect 15752 7880 15804 7886
rect 15804 7840 15884 7868
rect 15752 7822 15804 7828
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15566 7440 15622 7449
rect 15566 7375 15622 7384
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15672 6730 15700 7142
rect 15764 6866 15792 7686
rect 15856 7274 15884 7840
rect 15844 7268 15896 7274
rect 15844 7210 15896 7216
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15764 6662 15792 6802
rect 15856 6730 15884 7210
rect 16132 6730 16160 8366
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15660 6384 15712 6390
rect 15660 6326 15712 6332
rect 15672 5710 15700 6326
rect 15856 5710 15884 6666
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 16132 5846 16160 6258
rect 16120 5840 16172 5846
rect 16120 5782 16172 5788
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15856 5166 15884 5646
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3738 15700 3878
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15856 3670 15884 5102
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15488 2514 15516 2994
rect 16224 2514 16252 11494
rect 16500 11150 16528 12174
rect 16592 11801 16620 12310
rect 16578 11792 16634 11801
rect 16578 11727 16634 11736
rect 16580 11620 16632 11626
rect 16580 11562 16632 11568
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16486 10704 16542 10713
rect 16486 10639 16542 10648
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10266 16436 10406
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16302 7984 16358 7993
rect 16302 7919 16304 7928
rect 16356 7919 16358 7928
rect 16304 7890 16356 7896
rect 16394 6896 16450 6905
rect 16394 6831 16396 6840
rect 16448 6831 16450 6840
rect 16396 6802 16448 6808
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16408 6118 16436 6394
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 4480 16356 4486
rect 16304 4422 16356 4428
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 14936 1686 15056 1714
rect 14384 1142 14504 1170
rect 14476 480 14504 1142
rect 14936 480 14964 1686
rect 15396 480 15424 2246
rect 15856 480 15884 2246
rect 16316 480 16344 4422
rect 16500 3738 16528 10639
rect 16488 3732 16540 3738
rect 16488 3674 16540 3680
rect 16592 2514 16620 11562
rect 16684 8673 16712 12582
rect 17052 12442 17080 12582
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16854 12200 16910 12209
rect 16854 12135 16910 12144
rect 16868 11898 16896 12135
rect 16856 11892 16908 11898
rect 16856 11834 16908 11840
rect 17052 11801 17080 12378
rect 17038 11792 17094 11801
rect 17038 11727 17094 11736
rect 16856 11688 16908 11694
rect 16856 11630 16908 11636
rect 16868 11150 16896 11630
rect 16856 11144 16908 11150
rect 16908 11104 17080 11132
rect 16856 11086 16908 11092
rect 17052 10690 17080 11104
rect 17144 10810 17172 13223
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17328 12442 17356 12854
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11694 17264 12038
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17224 10736 17276 10742
rect 17052 10684 17224 10690
rect 17052 10678 17276 10684
rect 17052 10662 17264 10678
rect 16854 10568 16910 10577
rect 16764 10532 16816 10538
rect 16854 10503 16910 10512
rect 16764 10474 16816 10480
rect 16776 9654 16804 10474
rect 16868 10470 16896 10503
rect 16856 10464 16908 10470
rect 16856 10406 16908 10412
rect 16764 9648 16816 9654
rect 16764 9590 16816 9596
rect 16670 8664 16726 8673
rect 16670 8599 16726 8608
rect 16868 7800 16896 10406
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 17052 9586 17080 9998
rect 17132 9716 17184 9722
rect 17132 9658 17184 9664
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8566 16988 8774
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 16868 7772 16988 7800
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16684 6798 16712 7210
rect 16960 6798 16988 7772
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16856 4616 16908 4622
rect 16856 4558 16908 4564
rect 16868 4282 16896 4558
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16684 3670 16712 4082
rect 16960 4010 16988 6734
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16672 3664 16724 3670
rect 16672 3606 16724 3612
rect 17052 2990 17080 8502
rect 17144 8401 17172 9658
rect 17236 8956 17264 10202
rect 17420 9994 17448 12174
rect 17512 11898 17540 12174
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17512 11286 17540 11834
rect 17604 11558 17632 13738
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17788 12850 17816 13330
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17972 12322 18000 18770
rect 18116 18524 18412 18544
rect 18172 18522 18196 18524
rect 18252 18522 18276 18524
rect 18332 18522 18356 18524
rect 18194 18470 18196 18522
rect 18258 18470 18270 18522
rect 18332 18470 18334 18522
rect 18172 18468 18196 18470
rect 18252 18468 18276 18470
rect 18332 18468 18356 18470
rect 18116 18448 18412 18468
rect 18116 17436 18412 17456
rect 18172 17434 18196 17436
rect 18252 17434 18276 17436
rect 18332 17434 18356 17436
rect 18194 17382 18196 17434
rect 18258 17382 18270 17434
rect 18332 17382 18334 17434
rect 18172 17380 18196 17382
rect 18252 17380 18276 17382
rect 18332 17380 18356 17382
rect 18116 17360 18412 17380
rect 18116 16348 18412 16368
rect 18172 16346 18196 16348
rect 18252 16346 18276 16348
rect 18332 16346 18356 16348
rect 18194 16294 18196 16346
rect 18258 16294 18270 16346
rect 18332 16294 18334 16346
rect 18172 16292 18196 16294
rect 18252 16292 18276 16294
rect 18332 16292 18356 16294
rect 18116 16272 18412 16292
rect 18694 15600 18750 15609
rect 18694 15535 18750 15544
rect 18116 15260 18412 15280
rect 18172 15258 18196 15260
rect 18252 15258 18276 15260
rect 18332 15258 18356 15260
rect 18194 15206 18196 15258
rect 18258 15206 18270 15258
rect 18332 15206 18334 15258
rect 18172 15204 18196 15206
rect 18252 15204 18276 15206
rect 18332 15204 18356 15206
rect 18116 15184 18412 15204
rect 18512 14272 18564 14278
rect 18512 14214 18564 14220
rect 18116 14172 18412 14192
rect 18172 14170 18196 14172
rect 18252 14170 18276 14172
rect 18332 14170 18356 14172
rect 18194 14118 18196 14170
rect 18258 14118 18270 14170
rect 18332 14118 18334 14170
rect 18172 14116 18196 14118
rect 18252 14116 18276 14118
rect 18332 14116 18356 14118
rect 18116 14096 18412 14116
rect 18524 13394 18552 14214
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18116 13084 18412 13104
rect 18172 13082 18196 13084
rect 18252 13082 18276 13084
rect 18332 13082 18356 13084
rect 18194 13030 18196 13082
rect 18258 13030 18270 13082
rect 18332 13030 18334 13082
rect 18172 13028 18196 13030
rect 18252 13028 18276 13030
rect 18332 13028 18356 13030
rect 18116 13008 18412 13028
rect 18524 12782 18552 13126
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17880 12294 18000 12322
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17500 11280 17552 11286
rect 17788 11257 17816 12242
rect 17880 11778 17908 12294
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 17972 11898 18000 12174
rect 18524 12102 18552 12718
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18116 11996 18412 12016
rect 18172 11994 18196 11996
rect 18252 11994 18276 11996
rect 18332 11994 18356 11996
rect 18194 11942 18196 11994
rect 18258 11942 18270 11994
rect 18332 11942 18334 11994
rect 18172 11940 18196 11942
rect 18252 11940 18276 11942
rect 18332 11940 18356 11942
rect 18116 11920 18412 11940
rect 17960 11892 18012 11898
rect 17960 11834 18012 11840
rect 17880 11750 18000 11778
rect 17500 11222 17552 11228
rect 17774 11248 17830 11257
rect 17774 11183 17830 11192
rect 17500 10464 17552 10470
rect 17500 10406 17552 10412
rect 17512 10266 17540 10406
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17512 9382 17540 10066
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17328 9110 17356 9318
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 17316 8968 17368 8974
rect 17236 8928 17316 8956
rect 17316 8910 17368 8916
rect 17130 8392 17186 8401
rect 17130 8327 17186 8336
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 6322 17172 7686
rect 17236 6730 17264 8298
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17236 4078 17264 6190
rect 17328 4078 17356 8910
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17420 4486 17448 6938
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17144 2990 17172 3878
rect 17328 3126 17356 3878
rect 17316 3120 17368 3126
rect 17316 3062 17368 3068
rect 17420 3058 17448 3878
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17512 2990 17540 9318
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17604 7886 17632 8910
rect 17972 8786 18000 11750
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 18116 10908 18412 10928
rect 18172 10906 18196 10908
rect 18252 10906 18276 10908
rect 18332 10906 18356 10908
rect 18194 10854 18196 10906
rect 18258 10854 18270 10906
rect 18332 10854 18334 10906
rect 18172 10852 18196 10854
rect 18252 10852 18276 10854
rect 18332 10852 18356 10854
rect 18116 10832 18412 10852
rect 18328 10532 18380 10538
rect 18328 10474 18380 10480
rect 18050 10432 18106 10441
rect 18050 10367 18106 10376
rect 18064 9994 18092 10367
rect 18340 10062 18368 10474
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 18116 9820 18412 9840
rect 18172 9818 18196 9820
rect 18252 9818 18276 9820
rect 18332 9818 18356 9820
rect 18194 9766 18196 9818
rect 18258 9766 18270 9818
rect 18332 9766 18334 9818
rect 18172 9764 18196 9766
rect 18252 9764 18276 9766
rect 18332 9764 18356 9766
rect 18116 9744 18412 9764
rect 18524 9625 18552 11494
rect 18604 10600 18656 10606
rect 18604 10542 18656 10548
rect 18616 10130 18644 10542
rect 18604 10124 18656 10130
rect 18604 10066 18656 10072
rect 18510 9616 18566 9625
rect 18510 9551 18566 9560
rect 18604 9104 18656 9110
rect 18510 9072 18566 9081
rect 18604 9046 18656 9052
rect 18510 9007 18566 9016
rect 17880 8758 18000 8786
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17696 8022 17724 8434
rect 17880 8378 17908 8758
rect 18116 8732 18412 8752
rect 18172 8730 18196 8732
rect 18252 8730 18276 8732
rect 18332 8730 18356 8732
rect 18194 8678 18196 8730
rect 18258 8678 18270 8730
rect 18332 8678 18334 8730
rect 18172 8676 18196 8678
rect 18252 8676 18276 8678
rect 18332 8676 18356 8678
rect 18116 8656 18412 8676
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17972 8537 18000 8570
rect 18524 8566 18552 9007
rect 18512 8560 18564 8566
rect 17958 8528 18014 8537
rect 18512 8502 18564 8508
rect 17958 8463 18014 8472
rect 17880 8350 18000 8378
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7206 17632 7822
rect 17696 7546 17724 7958
rect 17868 7744 17920 7750
rect 17868 7686 17920 7692
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17774 7168 17830 7177
rect 17774 7103 17830 7112
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17604 5914 17632 6258
rect 17592 5908 17644 5914
rect 17592 5850 17644 5856
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 17604 5098 17632 5646
rect 17696 5370 17724 6598
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17684 4752 17736 4758
rect 17684 4694 17736 4700
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17604 4282 17632 4626
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17592 4072 17644 4078
rect 17592 4014 17644 4020
rect 17604 3398 17632 4014
rect 17696 3738 17724 4694
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17696 3058 17724 3674
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 17040 2984 17092 2990
rect 17040 2926 17092 2932
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17590 2816 17646 2825
rect 17590 2751 17646 2760
rect 17604 2689 17632 2751
rect 17590 2680 17646 2689
rect 17590 2615 17646 2624
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 16684 480 16712 2518
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 17144 480 17172 2314
rect 17604 480 17632 2450
rect 17788 2446 17816 7103
rect 17880 6798 17908 7686
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5846 17908 6258
rect 17868 5840 17920 5846
rect 17868 5782 17920 5788
rect 17972 5370 18000 8350
rect 18116 7644 18412 7664
rect 18172 7642 18196 7644
rect 18252 7642 18276 7644
rect 18332 7642 18356 7644
rect 18194 7590 18196 7642
rect 18258 7590 18270 7642
rect 18332 7590 18334 7642
rect 18172 7588 18196 7590
rect 18252 7588 18276 7590
rect 18332 7588 18356 7590
rect 18116 7568 18412 7588
rect 18116 6556 18412 6576
rect 18172 6554 18196 6556
rect 18252 6554 18276 6556
rect 18332 6554 18356 6556
rect 18194 6502 18196 6554
rect 18258 6502 18270 6554
rect 18332 6502 18334 6554
rect 18172 6500 18196 6502
rect 18252 6500 18276 6502
rect 18332 6500 18356 6502
rect 18116 6480 18412 6500
rect 18142 6216 18198 6225
rect 18142 6151 18198 6160
rect 18156 5778 18184 6151
rect 18328 6112 18380 6118
rect 18512 6112 18564 6118
rect 18380 6072 18460 6100
rect 18328 6054 18380 6060
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18432 5658 18460 6072
rect 18512 6054 18564 6060
rect 18524 5914 18552 6054
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18432 5630 18552 5658
rect 18116 5468 18412 5488
rect 18172 5466 18196 5468
rect 18252 5466 18276 5468
rect 18332 5466 18356 5468
rect 18194 5414 18196 5466
rect 18258 5414 18270 5466
rect 18332 5414 18334 5466
rect 18172 5412 18196 5414
rect 18252 5412 18276 5414
rect 18332 5412 18356 5414
rect 18116 5392 18412 5412
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17880 5012 17908 5306
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 17972 5166 18000 5199
rect 18524 5166 18552 5630
rect 17960 5160 18012 5166
rect 17960 5102 18012 5108
rect 18512 5160 18564 5166
rect 18512 5102 18564 5108
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 17880 4984 18000 5012
rect 17972 4622 18000 4984
rect 18340 4622 18368 5034
rect 18616 4978 18644 9046
rect 18708 6458 18736 15535
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18800 12170 18828 12718
rect 18892 12322 18920 14554
rect 18970 14104 19026 14113
rect 18970 14039 18972 14048
rect 19024 14039 19026 14048
rect 18972 14010 19024 14016
rect 18892 12294 19012 12322
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18880 12164 18932 12170
rect 18880 12106 18932 12112
rect 18892 11762 18920 12106
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 18984 11393 19012 12294
rect 18970 11384 19026 11393
rect 18970 11319 19026 11328
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 7585 18828 8774
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18788 7268 18840 7274
rect 18788 7210 18840 7216
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18800 6186 18828 7210
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5166 18736 6054
rect 18696 5160 18748 5166
rect 18696 5102 18748 5108
rect 18524 4950 18644 4978
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18524 4690 18552 4950
rect 18512 4684 18564 4690
rect 18512 4626 18564 4632
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 17880 3890 17908 4558
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17972 4078 18000 4422
rect 18116 4380 18412 4400
rect 18172 4378 18196 4380
rect 18252 4378 18276 4380
rect 18332 4378 18356 4380
rect 18194 4326 18196 4378
rect 18258 4326 18270 4378
rect 18332 4326 18334 4378
rect 18172 4324 18196 4326
rect 18252 4324 18276 4326
rect 18332 4324 18356 4326
rect 18116 4304 18412 4324
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 18144 4004 18196 4010
rect 18144 3946 18196 3952
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 17880 3862 18000 3890
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17880 3058 17908 3538
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17868 2916 17920 2922
rect 17868 2858 17920 2864
rect 17880 2650 17908 2858
rect 17972 2825 18000 3862
rect 18156 3505 18184 3946
rect 18512 3936 18564 3942
rect 18512 3878 18564 3884
rect 18524 3738 18552 3878
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18236 3664 18288 3670
rect 18234 3632 18236 3641
rect 18288 3632 18290 3641
rect 18234 3567 18290 3576
rect 18512 3596 18564 3602
rect 18512 3538 18564 3544
rect 18142 3496 18198 3505
rect 18142 3431 18198 3440
rect 18116 3292 18412 3312
rect 18172 3290 18196 3292
rect 18252 3290 18276 3292
rect 18332 3290 18356 3292
rect 18194 3238 18196 3290
rect 18258 3238 18270 3290
rect 18332 3238 18334 3290
rect 18172 3236 18196 3238
rect 18252 3236 18276 3238
rect 18332 3236 18356 3238
rect 18116 3216 18412 3236
rect 18144 2984 18196 2990
rect 18144 2926 18196 2932
rect 17958 2816 18014 2825
rect 17958 2751 18014 2760
rect 18156 2666 18184 2926
rect 18524 2825 18552 3538
rect 18510 2816 18566 2825
rect 18510 2751 18566 2760
rect 18234 2680 18290 2689
rect 17868 2644 17920 2650
rect 18156 2638 18234 2666
rect 18616 2650 18644 3946
rect 18800 3890 18828 4966
rect 18708 3862 18828 3890
rect 18234 2615 18290 2624
rect 18604 2644 18656 2650
rect 17868 2586 17920 2592
rect 18604 2586 18656 2592
rect 18708 2530 18736 3862
rect 18892 3516 18920 11018
rect 19076 10198 19104 22471
rect 20902 22128 20958 22137
rect 20902 22063 20958 22072
rect 20626 21584 20682 21593
rect 20626 21519 20682 21528
rect 20258 21176 20314 21185
rect 20258 21111 20314 21120
rect 19154 20632 19210 20641
rect 19154 20567 19210 20576
rect 19168 19514 19196 20567
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19616 15088 19668 15094
rect 19614 15056 19616 15065
rect 19668 15056 19670 15065
rect 19614 14991 19670 15000
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19246 14648 19302 14657
rect 19246 14583 19302 14592
rect 19260 14074 19288 14583
rect 19444 14550 19472 14894
rect 19432 14544 19484 14550
rect 19432 14486 19484 14492
rect 19616 14476 19668 14482
rect 19616 14418 19668 14424
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19248 14068 19300 14074
rect 19248 14010 19300 14016
rect 19156 14000 19208 14006
rect 19156 13942 19208 13948
rect 19064 10192 19116 10198
rect 19064 10134 19116 10140
rect 19064 9036 19116 9042
rect 19064 8978 19116 8984
rect 18972 8356 19024 8362
rect 18972 8298 19024 8304
rect 18984 6866 19012 8298
rect 19076 8090 19104 8978
rect 19168 8634 19196 13942
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 12753 19288 13330
rect 19352 13297 19380 14214
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19338 13288 19394 13297
rect 19338 13223 19394 13232
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19246 12744 19302 12753
rect 19246 12679 19302 12688
rect 19352 11898 19380 13126
rect 19444 12209 19472 13806
rect 19536 13462 19564 14350
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19628 12850 19656 14418
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19524 12232 19576 12238
rect 19430 12200 19486 12209
rect 19628 12186 19656 12582
rect 19576 12180 19656 12186
rect 19524 12174 19656 12180
rect 19536 12158 19656 12174
rect 19430 12135 19486 12144
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19628 11694 19656 12158
rect 19616 11688 19668 11694
rect 19246 11656 19302 11665
rect 19616 11630 19668 11636
rect 19246 11591 19302 11600
rect 19260 11234 19288 11591
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 19260 11206 19380 11234
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10849 19288 11086
rect 19246 10840 19302 10849
rect 19246 10775 19302 10784
rect 19352 10690 19380 11206
rect 19444 11150 19472 11494
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19260 10662 19380 10690
rect 19444 10674 19472 11086
rect 19720 10690 19748 17682
rect 19984 17128 20036 17134
rect 19984 17070 20036 17076
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19812 11218 19840 15914
rect 19904 12714 19932 15982
rect 19892 12708 19944 12714
rect 19892 12650 19944 12656
rect 19890 12608 19946 12617
rect 19890 12543 19946 12552
rect 19904 11234 19932 12543
rect 19996 11370 20024 17070
rect 20166 16552 20222 16561
rect 20166 16487 20222 16496
rect 20180 16250 20208 16487
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 20088 11694 20116 15506
rect 20272 15162 20300 21111
rect 20536 19304 20588 19310
rect 20442 19272 20498 19281
rect 20536 19246 20588 19252
rect 20442 19207 20498 19216
rect 20350 18184 20406 18193
rect 20350 18119 20406 18128
rect 20260 15156 20312 15162
rect 20260 15098 20312 15104
rect 20364 15026 20392 18119
rect 20456 16794 20484 19207
rect 20548 18329 20576 19246
rect 20534 18320 20590 18329
rect 20534 18255 20590 18264
rect 20536 18216 20588 18222
rect 20536 18158 20588 18164
rect 20548 17814 20576 18158
rect 20536 17808 20588 17814
rect 20536 17750 20588 17756
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20442 16008 20498 16017
rect 20442 15943 20498 15952
rect 20456 15706 20484 15943
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20168 13864 20220 13870
rect 20168 13806 20220 13812
rect 20180 12306 20208 13806
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 20076 11688 20128 11694
rect 20076 11630 20128 11636
rect 19996 11342 20116 11370
rect 19800 11212 19852 11218
rect 19904 11206 20024 11234
rect 19800 11154 19852 11160
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19432 10668 19484 10674
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19260 8129 19288 10662
rect 19432 10610 19484 10616
rect 19628 10662 19748 10690
rect 19628 9654 19656 10662
rect 19708 10600 19760 10606
rect 19708 10542 19760 10548
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19720 9586 19748 10542
rect 19800 10124 19852 10130
rect 19800 10066 19852 10072
rect 19708 9580 19760 9586
rect 19708 9522 19760 9528
rect 19812 9178 19840 10066
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19340 8356 19392 8362
rect 19340 8298 19392 8304
rect 19246 8120 19302 8129
rect 19064 8084 19116 8090
rect 19246 8055 19302 8064
rect 19064 8026 19116 8032
rect 19076 7410 19104 8026
rect 19156 7880 19208 7886
rect 19154 7848 19156 7857
rect 19208 7848 19210 7857
rect 19154 7783 19210 7792
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 19076 6798 19104 7346
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 19352 6730 19380 8298
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19444 7546 19472 8230
rect 19628 7954 19656 8978
rect 19812 8498 19840 9114
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19432 7540 19484 7546
rect 19432 7482 19484 7488
rect 19432 7336 19484 7342
rect 19432 7278 19484 7284
rect 19340 6724 19392 6730
rect 19340 6666 19392 6672
rect 19062 6352 19118 6361
rect 19062 6287 19118 6296
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 5234 19012 5510
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18984 3738 19012 4626
rect 19076 3738 19104 6287
rect 19444 6254 19472 7278
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19536 6730 19564 7210
rect 19524 6724 19576 6730
rect 19524 6666 19576 6672
rect 19432 6248 19484 6254
rect 19432 6190 19484 6196
rect 19248 6180 19300 6186
rect 19248 6122 19300 6128
rect 19156 5772 19208 5778
rect 19260 5760 19288 6122
rect 19628 6118 19656 7890
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19812 6390 19840 7482
rect 19800 6384 19852 6390
rect 19800 6326 19852 6332
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19260 5732 19472 5760
rect 19156 5714 19208 5720
rect 19168 4826 19196 5714
rect 19248 5636 19300 5642
rect 19248 5578 19300 5584
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19064 3528 19116 3534
rect 18800 3488 19064 3516
rect 18800 2922 18828 3488
rect 19064 3470 19116 3476
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18880 2916 18932 2922
rect 18880 2858 18932 2864
rect 18786 2816 18842 2825
rect 18786 2751 18842 2760
rect 18524 2502 18736 2530
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17960 2372 18012 2378
rect 17960 2314 18012 2320
rect 17972 1170 18000 2314
rect 18116 2204 18412 2224
rect 18172 2202 18196 2204
rect 18252 2202 18276 2204
rect 18332 2202 18356 2204
rect 18194 2150 18196 2202
rect 18258 2150 18270 2202
rect 18332 2150 18334 2202
rect 18172 2148 18196 2150
rect 18252 2148 18276 2150
rect 18332 2148 18356 2150
rect 18116 2128 18412 2148
rect 17972 1142 18092 1170
rect 18064 480 18092 1142
rect 18524 480 18552 2502
rect 5630 232 5686 241
rect 5630 167 5686 176
rect 5998 0 6054 480
rect 6458 0 6514 480
rect 6826 0 6882 480
rect 7286 0 7342 480
rect 7746 0 7802 480
rect 8206 0 8262 480
rect 8666 0 8722 480
rect 9126 0 9182 480
rect 9586 0 9642 480
rect 9954 0 10010 480
rect 10414 0 10470 480
rect 10874 0 10930 480
rect 11334 0 11390 480
rect 11794 0 11850 480
rect 12254 0 12310 480
rect 12714 0 12770 480
rect 13174 0 13230 480
rect 13542 0 13598 480
rect 14002 0 14058 480
rect 14462 0 14518 480
rect 14922 0 14978 480
rect 15382 0 15438 480
rect 15842 0 15898 480
rect 16302 0 16358 480
rect 16670 0 16726 480
rect 17130 0 17186 480
rect 17590 0 17646 480
rect 18050 0 18106 480
rect 18510 0 18566 480
rect 18800 241 18828 2751
rect 18892 2514 18920 2858
rect 18880 2508 18932 2514
rect 18880 2450 18932 2456
rect 18984 480 19012 3130
rect 19076 2530 19104 3470
rect 19168 2825 19196 4762
rect 19260 3913 19288 5578
rect 19340 5160 19392 5166
rect 19340 5102 19392 5108
rect 19352 4758 19380 5102
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19444 4690 19472 5732
rect 19708 5704 19760 5710
rect 19708 5646 19760 5652
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19432 4684 19484 4690
rect 19432 4626 19484 4632
rect 19536 4486 19564 5102
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19340 4140 19392 4146
rect 19340 4082 19392 4088
rect 19352 4026 19380 4082
rect 19352 3998 19472 4026
rect 19340 3936 19392 3942
rect 19246 3904 19302 3913
rect 19340 3878 19392 3884
rect 19246 3839 19302 3848
rect 19248 3732 19300 3738
rect 19248 3674 19300 3680
rect 19260 3602 19288 3674
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19154 2816 19210 2825
rect 19154 2751 19210 2760
rect 19168 2650 19196 2751
rect 19156 2644 19208 2650
rect 19156 2586 19208 2592
rect 19076 2502 19196 2530
rect 19260 2514 19288 3538
rect 19352 2854 19380 3878
rect 19444 2854 19472 3998
rect 19340 2848 19392 2854
rect 19340 2790 19392 2796
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19536 2650 19564 4218
rect 19524 2644 19576 2650
rect 19524 2586 19576 2592
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19628 2530 19656 5238
rect 19720 3670 19748 5646
rect 19800 5092 19852 5098
rect 19800 5034 19852 5040
rect 19812 4826 19840 5034
rect 19800 4820 19852 4826
rect 19800 4762 19852 4768
rect 19812 4146 19840 4762
rect 19904 4690 19932 11018
rect 19996 9178 20024 11206
rect 20088 9722 20116 11342
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20180 10266 20208 11154
rect 20168 10260 20220 10266
rect 20168 10202 20220 10208
rect 20076 9716 20128 9722
rect 20076 9658 20128 9664
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 19996 6934 20024 8230
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20180 7546 20208 7822
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20168 7200 20220 7206
rect 20168 7142 20220 7148
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19800 4140 19852 4146
rect 19800 4082 19852 4088
rect 19996 3738 20024 6734
rect 20088 3942 20116 7142
rect 20180 6458 20208 7142
rect 20168 6452 20220 6458
rect 20168 6394 20220 6400
rect 20272 4010 20300 13738
rect 20442 13696 20498 13705
rect 20442 13631 20498 13640
rect 20352 13388 20404 13394
rect 20352 13330 20404 13336
rect 20364 12442 20392 13330
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20364 12345 20392 12378
rect 20350 12336 20406 12345
rect 20350 12271 20406 12280
rect 20456 12170 20484 13631
rect 20444 12164 20496 12170
rect 20444 12106 20496 12112
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20352 11144 20404 11150
rect 20352 11086 20404 11092
rect 20364 10470 20392 11086
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 9518 20392 10406
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20456 9330 20484 11630
rect 20548 11286 20576 16594
rect 20640 15162 20668 21519
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19514 20760 19751
rect 20720 19508 20772 19514
rect 20720 19450 20772 19456
rect 20718 18864 20774 18873
rect 20718 18799 20774 18808
rect 20732 18426 20760 18799
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20718 17912 20774 17921
rect 20718 17847 20774 17856
rect 20732 17338 20760 17847
rect 20810 17368 20866 17377
rect 20720 17332 20772 17338
rect 20810 17303 20866 17312
rect 20720 17274 20772 17280
rect 20824 16250 20852 17303
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20640 12866 20668 14962
rect 20916 12986 20944 22063
rect 20994 20224 21050 20233
rect 20994 20159 21050 20168
rect 20904 12980 20956 12986
rect 20904 12922 20956 12928
rect 20640 12838 20760 12866
rect 20628 12776 20680 12782
rect 20628 12718 20680 12724
rect 20640 12238 20668 12718
rect 20732 12617 20760 12838
rect 20718 12608 20774 12617
rect 20718 12543 20774 12552
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 21008 11898 21036 20159
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20536 11280 20588 11286
rect 20536 11222 20588 11228
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20364 9302 20484 9330
rect 20364 7546 20392 9302
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20456 8090 20484 8230
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20548 8022 20576 8434
rect 20536 8016 20588 8022
rect 20536 7958 20588 7964
rect 20444 7744 20496 7750
rect 20444 7686 20496 7692
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20456 6322 20484 7686
rect 20548 7410 20576 7958
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 6798 20576 7346
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 20456 5386 20484 6258
rect 20640 6254 20668 10134
rect 20732 7954 20760 11630
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20916 8090 20944 8298
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20720 7948 20772 7954
rect 20720 7890 20772 7896
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20456 5370 20576 5386
rect 20456 5364 20588 5370
rect 20456 5358 20536 5364
rect 20536 5306 20588 5312
rect 20548 4214 20576 5306
rect 20732 4321 20760 7278
rect 21088 7200 21140 7206
rect 21088 7142 21140 7148
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 20718 4312 20774 4321
rect 20718 4247 20774 4256
rect 20536 4208 20588 4214
rect 20456 4156 20536 4162
rect 20456 4150 20588 4156
rect 20456 4134 20576 4150
rect 20260 4004 20312 4010
rect 20260 3946 20312 3952
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 20074 3632 20130 3641
rect 20074 3567 20130 3576
rect 19984 3460 20036 3466
rect 19984 3402 20036 3408
rect 19996 2650 20024 3402
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 19168 2446 19196 2502
rect 19248 2508 19300 2514
rect 19248 2450 19300 2456
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 19260 2009 19288 2450
rect 19246 2000 19302 2009
rect 19246 1935 19302 1944
rect 19444 480 19472 2518
rect 19628 2502 19840 2530
rect 20088 2514 20116 3567
rect 20456 3534 20484 4134
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3670 20576 4014
rect 20904 3936 20956 3942
rect 20904 3878 20956 3884
rect 20536 3664 20588 3670
rect 20536 3606 20588 3612
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20456 2961 20484 2994
rect 20442 2952 20498 2961
rect 20442 2887 20498 2896
rect 20168 2848 20220 2854
rect 20168 2790 20220 2796
rect 19812 480 19840 2502
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20180 2446 20208 2790
rect 20168 2440 20220 2446
rect 20168 2382 20220 2388
rect 20548 1057 20576 3606
rect 20812 3460 20864 3466
rect 20812 3402 20864 3408
rect 20824 2689 20852 3402
rect 20916 3398 20944 3878
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20810 2680 20866 2689
rect 20810 2615 20866 2624
rect 20824 1601 20852 2615
rect 20810 1592 20866 1601
rect 20810 1527 20866 1536
rect 20534 1048 20590 1057
rect 20534 983 20590 992
rect 20916 649 20944 3334
rect 20902 640 20958 649
rect 20260 604 20312 610
rect 20260 546 20312 552
rect 20720 604 20772 610
rect 21008 610 21036 5510
rect 21100 678 21128 7142
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21088 672 21140 678
rect 21088 614 21140 620
rect 20902 575 20958 584
rect 20996 604 21048 610
rect 20720 546 20772 552
rect 20996 546 21048 552
rect 20272 480 20300 546
rect 20732 480 20760 546
rect 21192 480 21220 5102
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21640 2916 21692 2922
rect 21640 2858 21692 2864
rect 21652 480 21680 2858
rect 22112 480 22140 3062
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22572 480 22600 2926
rect 18786 232 18842 241
rect 18786 167 18842 176
rect 18970 0 19026 480
rect 19430 0 19486 480
rect 19798 0 19854 480
rect 20258 0 20314 480
rect 20718 0 20774 480
rect 21178 0 21234 480
rect 21638 0 21694 480
rect 22098 0 22154 480
rect 22558 0 22614 480
<< via2 >>
rect 2962 22480 3018 22536
rect 2318 22072 2374 22128
rect 1950 19760 2006 19816
rect 1950 19216 2006 19272
rect 1950 18808 2006 18864
rect 1858 18264 1914 18320
rect 1674 17856 1730 17912
rect 1950 17312 2006 17368
rect 1950 16496 2006 16552
rect 2502 21120 2558 21176
rect 1950 15952 2006 16008
rect 2778 20168 2834 20224
rect 2778 15544 2834 15600
rect 1950 15036 1952 15056
rect 1952 15036 2004 15056
rect 2004 15036 2006 15056
rect 1950 15000 2006 15036
rect 1674 14612 1730 14648
rect 1674 14592 1676 14612
rect 1676 14592 1728 14612
rect 1728 14592 1730 14612
rect 1582 14048 1638 14104
rect 1490 10648 1546 10704
rect 1950 7928 2006 7984
rect 19062 22480 19118 22536
rect 3146 21528 3202 21584
rect 3698 20576 3754 20632
rect 4388 19610 4444 19612
rect 4468 19610 4524 19612
rect 4548 19610 4604 19612
rect 4628 19610 4684 19612
rect 4388 19558 4414 19610
rect 4414 19558 4444 19610
rect 4468 19558 4478 19610
rect 4478 19558 4524 19610
rect 4548 19558 4594 19610
rect 4594 19558 4604 19610
rect 4628 19558 4658 19610
rect 4658 19558 4684 19610
rect 4388 19556 4444 19558
rect 4468 19556 4524 19558
rect 4548 19556 4604 19558
rect 4628 19556 4684 19558
rect 4388 18522 4444 18524
rect 4468 18522 4524 18524
rect 4548 18522 4604 18524
rect 4628 18522 4684 18524
rect 4388 18470 4414 18522
rect 4414 18470 4444 18522
rect 4468 18470 4478 18522
rect 4478 18470 4524 18522
rect 4548 18470 4594 18522
rect 4594 18470 4604 18522
rect 4628 18470 4658 18522
rect 4658 18470 4684 18522
rect 4388 18468 4444 18470
rect 4468 18468 4524 18470
rect 4548 18468 4604 18470
rect 4628 18468 4684 18470
rect 4388 17434 4444 17436
rect 4468 17434 4524 17436
rect 4548 17434 4604 17436
rect 4628 17434 4684 17436
rect 4388 17382 4414 17434
rect 4414 17382 4444 17434
rect 4468 17382 4478 17434
rect 4478 17382 4524 17434
rect 4548 17382 4594 17434
rect 4594 17382 4604 17434
rect 4628 17382 4658 17434
rect 4658 17382 4684 17434
rect 4388 17380 4444 17382
rect 4468 17380 4524 17382
rect 4548 17380 4604 17382
rect 4628 17380 4684 17382
rect 3422 16904 3478 16960
rect 4388 16346 4444 16348
rect 4468 16346 4524 16348
rect 4548 16346 4604 16348
rect 4628 16346 4684 16348
rect 4388 16294 4414 16346
rect 4414 16294 4444 16346
rect 4468 16294 4478 16346
rect 4478 16294 4524 16346
rect 4548 16294 4594 16346
rect 4594 16294 4604 16346
rect 4628 16294 4658 16346
rect 4658 16294 4684 16346
rect 4388 16292 4444 16294
rect 4468 16292 4524 16294
rect 4548 16292 4604 16294
rect 4628 16292 4684 16294
rect 2594 10104 2650 10160
rect 3330 13640 3386 13696
rect 3606 13232 3662 13288
rect 2318 2488 2374 2544
rect 2962 7792 3018 7848
rect 2870 5072 2926 5128
rect 3146 3068 3148 3088
rect 3148 3068 3200 3088
rect 3200 3068 3202 3088
rect 3146 3032 3202 3068
rect 3974 12708 4030 12744
rect 3974 12688 3976 12708
rect 3976 12688 4028 12708
rect 4028 12688 4030 12708
rect 3698 9968 3754 10024
rect 3882 12280 3938 12336
rect 4066 11736 4122 11792
rect 3882 10784 3938 10840
rect 3514 7964 3516 7984
rect 3516 7964 3568 7984
rect 3568 7964 3570 7984
rect 3514 7928 3570 7964
rect 3790 7112 3846 7168
rect 4066 10376 4122 10432
rect 4066 9424 4122 9480
rect 4388 15258 4444 15260
rect 4468 15258 4524 15260
rect 4548 15258 4604 15260
rect 4628 15258 4684 15260
rect 4388 15206 4414 15258
rect 4414 15206 4444 15258
rect 4468 15206 4478 15258
rect 4478 15206 4524 15258
rect 4548 15206 4594 15258
rect 4594 15206 4604 15258
rect 4628 15206 4658 15258
rect 4658 15206 4684 15258
rect 4388 15204 4444 15206
rect 4468 15204 4524 15206
rect 4548 15204 4604 15206
rect 4628 15204 4684 15206
rect 4388 14170 4444 14172
rect 4468 14170 4524 14172
rect 4548 14170 4604 14172
rect 4628 14170 4684 14172
rect 4388 14118 4414 14170
rect 4414 14118 4444 14170
rect 4468 14118 4478 14170
rect 4478 14118 4524 14170
rect 4548 14118 4594 14170
rect 4594 14118 4604 14170
rect 4628 14118 4658 14170
rect 4658 14118 4684 14170
rect 4388 14116 4444 14118
rect 4468 14116 4524 14118
rect 4548 14116 4604 14118
rect 4628 14116 4684 14118
rect 4388 13082 4444 13084
rect 4468 13082 4524 13084
rect 4548 13082 4604 13084
rect 4628 13082 4684 13084
rect 4388 13030 4414 13082
rect 4414 13030 4444 13082
rect 4468 13030 4478 13082
rect 4478 13030 4524 13082
rect 4548 13030 4594 13082
rect 4594 13030 4604 13082
rect 4628 13030 4658 13082
rect 4658 13030 4684 13082
rect 4388 13028 4444 13030
rect 4468 13028 4524 13030
rect 4548 13028 4604 13030
rect 4628 13028 4684 13030
rect 4388 11994 4444 11996
rect 4468 11994 4524 11996
rect 4548 11994 4604 11996
rect 4628 11994 4684 11996
rect 4388 11942 4414 11994
rect 4414 11942 4444 11994
rect 4468 11942 4478 11994
rect 4478 11942 4524 11994
rect 4548 11942 4594 11994
rect 4594 11942 4604 11994
rect 4628 11942 4658 11994
rect 4658 11942 4684 11994
rect 4388 11940 4444 11942
rect 4468 11940 4524 11942
rect 4548 11940 4604 11942
rect 4628 11940 4684 11942
rect 4388 10906 4444 10908
rect 4468 10906 4524 10908
rect 4548 10906 4604 10908
rect 4628 10906 4684 10908
rect 4388 10854 4414 10906
rect 4414 10854 4444 10906
rect 4468 10854 4478 10906
rect 4478 10854 4524 10906
rect 4548 10854 4594 10906
rect 4594 10854 4604 10906
rect 4628 10854 4658 10906
rect 4658 10854 4684 10906
rect 4388 10852 4444 10854
rect 4468 10852 4524 10854
rect 4548 10852 4604 10854
rect 4628 10852 4684 10854
rect 4618 10512 4674 10568
rect 4388 9818 4444 9820
rect 4468 9818 4524 9820
rect 4548 9818 4604 9820
rect 4628 9818 4684 9820
rect 4388 9766 4414 9818
rect 4414 9766 4444 9818
rect 4468 9766 4478 9818
rect 4478 9766 4524 9818
rect 4548 9766 4594 9818
rect 4594 9766 4604 9818
rect 4628 9766 4658 9818
rect 4658 9766 4684 9818
rect 4388 9764 4444 9766
rect 4468 9764 4524 9766
rect 4548 9764 4604 9766
rect 4628 9764 4684 9766
rect 4066 8508 4068 8528
rect 4068 8508 4120 8528
rect 4120 8508 4122 8528
rect 4066 8472 4122 8508
rect 4388 8730 4444 8732
rect 4468 8730 4524 8732
rect 4548 8730 4604 8732
rect 4628 8730 4684 8732
rect 4388 8678 4414 8730
rect 4414 8678 4444 8730
rect 4468 8678 4478 8730
rect 4478 8678 4524 8730
rect 4548 8678 4594 8730
rect 4594 8678 4604 8730
rect 4628 8678 4658 8730
rect 4658 8678 4684 8730
rect 4388 8676 4444 8678
rect 4468 8676 4524 8678
rect 4548 8676 4604 8678
rect 4628 8676 4684 8678
rect 3974 7948 4030 7984
rect 3974 7928 3976 7948
rect 3976 7928 4028 7948
rect 4028 7928 4030 7948
rect 3974 7520 4030 7576
rect 3974 6160 4030 6216
rect 3330 2760 3386 2816
rect 2502 1536 2558 1592
rect 3974 5772 4030 5808
rect 3974 5752 3976 5772
rect 3976 5752 4028 5772
rect 4028 5752 4030 5772
rect 4066 5208 4122 5264
rect 3974 4800 4030 4856
rect 4066 4256 4122 4312
rect 3882 3440 3938 3496
rect 3974 1944 4030 2000
rect 4066 992 4122 1048
rect 3974 584 4030 640
rect 4388 7642 4444 7644
rect 4468 7642 4524 7644
rect 4548 7642 4604 7644
rect 4628 7642 4684 7644
rect 4388 7590 4414 7642
rect 4414 7590 4444 7642
rect 4468 7590 4478 7642
rect 4478 7590 4524 7642
rect 4548 7590 4594 7642
rect 4594 7590 4604 7642
rect 4628 7590 4658 7642
rect 4658 7590 4684 7642
rect 4388 7588 4444 7590
rect 4468 7588 4524 7590
rect 4548 7588 4604 7590
rect 4628 7588 4684 7590
rect 4388 6554 4444 6556
rect 4468 6554 4524 6556
rect 4548 6554 4604 6556
rect 4628 6554 4684 6556
rect 4388 6502 4414 6554
rect 4414 6502 4444 6554
rect 4468 6502 4478 6554
rect 4478 6502 4524 6554
rect 4548 6502 4594 6554
rect 4594 6502 4604 6554
rect 4628 6502 4658 6554
rect 4658 6502 4684 6554
rect 4388 6500 4444 6502
rect 4468 6500 4524 6502
rect 4548 6500 4604 6502
rect 4628 6500 4684 6502
rect 4388 5466 4444 5468
rect 4468 5466 4524 5468
rect 4548 5466 4604 5468
rect 4628 5466 4684 5468
rect 4388 5414 4414 5466
rect 4414 5414 4444 5466
rect 4468 5414 4478 5466
rect 4478 5414 4524 5466
rect 4548 5414 4594 5466
rect 4594 5414 4604 5466
rect 4628 5414 4658 5466
rect 4658 5414 4684 5466
rect 4388 5412 4444 5414
rect 4468 5412 4524 5414
rect 4548 5412 4604 5414
rect 4628 5412 4684 5414
rect 4388 4378 4444 4380
rect 4468 4378 4524 4380
rect 4548 4378 4604 4380
rect 4628 4378 4684 4380
rect 4388 4326 4414 4378
rect 4414 4326 4444 4378
rect 4468 4326 4478 4378
rect 4478 4326 4524 4378
rect 4548 4326 4594 4378
rect 4594 4326 4604 4378
rect 4628 4326 4658 4378
rect 4658 4326 4684 4378
rect 4388 4324 4444 4326
rect 4468 4324 4524 4326
rect 4548 4324 4604 4326
rect 4628 4324 4684 4326
rect 4388 3290 4444 3292
rect 4468 3290 4524 3292
rect 4548 3290 4604 3292
rect 4628 3290 4684 3292
rect 4388 3238 4414 3290
rect 4414 3238 4444 3290
rect 4468 3238 4478 3290
rect 4478 3238 4524 3290
rect 4548 3238 4594 3290
rect 4594 3238 4604 3290
rect 4628 3238 4658 3290
rect 4658 3238 4684 3290
rect 4388 3236 4444 3238
rect 4468 3236 4524 3238
rect 4548 3236 4604 3238
rect 4628 3236 4684 3238
rect 4250 2896 4306 2952
rect 4388 2202 4444 2204
rect 4468 2202 4524 2204
rect 4548 2202 4604 2204
rect 4628 2202 4684 2204
rect 4388 2150 4414 2202
rect 4414 2150 4444 2202
rect 4468 2150 4478 2202
rect 4478 2150 4524 2202
rect 4548 2150 4594 2202
rect 4594 2150 4604 2202
rect 4628 2150 4658 2202
rect 4658 2150 4684 2202
rect 4388 2148 4444 2150
rect 4468 2148 4524 2150
rect 4548 2148 4604 2150
rect 4628 2148 4684 2150
rect 7820 20154 7876 20156
rect 7900 20154 7956 20156
rect 7980 20154 8036 20156
rect 8060 20154 8116 20156
rect 7820 20102 7846 20154
rect 7846 20102 7876 20154
rect 7900 20102 7910 20154
rect 7910 20102 7956 20154
rect 7980 20102 8026 20154
rect 8026 20102 8036 20154
rect 8060 20102 8090 20154
rect 8090 20102 8116 20154
rect 7820 20100 7876 20102
rect 7900 20100 7956 20102
rect 7980 20100 8036 20102
rect 8060 20100 8116 20102
rect 14684 20154 14740 20156
rect 14764 20154 14820 20156
rect 14844 20154 14900 20156
rect 14924 20154 14980 20156
rect 14684 20102 14710 20154
rect 14710 20102 14740 20154
rect 14764 20102 14774 20154
rect 14774 20102 14820 20154
rect 14844 20102 14890 20154
rect 14890 20102 14900 20154
rect 14924 20102 14954 20154
rect 14954 20102 14980 20154
rect 14684 20100 14740 20102
rect 14764 20100 14820 20102
rect 14844 20100 14900 20102
rect 14924 20100 14980 20102
rect 11252 19610 11308 19612
rect 11332 19610 11388 19612
rect 11412 19610 11468 19612
rect 11492 19610 11548 19612
rect 11252 19558 11278 19610
rect 11278 19558 11308 19610
rect 11332 19558 11342 19610
rect 11342 19558 11388 19610
rect 11412 19558 11458 19610
rect 11458 19558 11468 19610
rect 11492 19558 11522 19610
rect 11522 19558 11548 19610
rect 11252 19556 11308 19558
rect 11332 19556 11388 19558
rect 11412 19556 11468 19558
rect 11492 19556 11548 19558
rect 7820 19066 7876 19068
rect 7900 19066 7956 19068
rect 7980 19066 8036 19068
rect 8060 19066 8116 19068
rect 7820 19014 7846 19066
rect 7846 19014 7876 19066
rect 7900 19014 7910 19066
rect 7910 19014 7956 19066
rect 7980 19014 8026 19066
rect 8026 19014 8036 19066
rect 8060 19014 8090 19066
rect 8090 19014 8116 19066
rect 7820 19012 7876 19014
rect 7900 19012 7956 19014
rect 7980 19012 8036 19014
rect 8060 19012 8116 19014
rect 14684 19066 14740 19068
rect 14764 19066 14820 19068
rect 14844 19066 14900 19068
rect 14924 19066 14980 19068
rect 14684 19014 14710 19066
rect 14710 19014 14740 19066
rect 14764 19014 14774 19066
rect 14774 19014 14820 19066
rect 14844 19014 14890 19066
rect 14890 19014 14900 19066
rect 14924 19014 14954 19066
rect 14954 19014 14980 19066
rect 14684 19012 14740 19014
rect 14764 19012 14820 19014
rect 14844 19012 14900 19014
rect 14924 19012 14980 19014
rect 4894 10512 4950 10568
rect 4986 9424 5042 9480
rect 5354 10104 5410 10160
rect 5446 9596 5448 9616
rect 5448 9596 5500 9616
rect 5500 9596 5502 9616
rect 5446 9560 5502 9596
rect 5538 8236 5540 8256
rect 5540 8236 5592 8256
rect 5592 8236 5594 8256
rect 5538 8200 5594 8236
rect 4986 5228 5042 5264
rect 4986 5208 4988 5228
rect 4988 5208 5040 5228
rect 5040 5208 5042 5228
rect 11252 18522 11308 18524
rect 11332 18522 11388 18524
rect 11412 18522 11468 18524
rect 11492 18522 11548 18524
rect 11252 18470 11278 18522
rect 11278 18470 11308 18522
rect 11332 18470 11342 18522
rect 11342 18470 11388 18522
rect 11412 18470 11458 18522
rect 11458 18470 11468 18522
rect 11492 18470 11522 18522
rect 11522 18470 11548 18522
rect 11252 18468 11308 18470
rect 11332 18468 11388 18470
rect 11412 18468 11468 18470
rect 11492 18468 11548 18470
rect 7820 17978 7876 17980
rect 7900 17978 7956 17980
rect 7980 17978 8036 17980
rect 8060 17978 8116 17980
rect 7820 17926 7846 17978
rect 7846 17926 7876 17978
rect 7900 17926 7910 17978
rect 7910 17926 7956 17978
rect 7980 17926 8026 17978
rect 8026 17926 8036 17978
rect 8060 17926 8090 17978
rect 8090 17926 8116 17978
rect 7820 17924 7876 17926
rect 7900 17924 7956 17926
rect 7980 17924 8036 17926
rect 8060 17924 8116 17926
rect 5998 11328 6054 11384
rect 6090 10648 6146 10704
rect 5814 8200 5870 8256
rect 7010 11736 7066 11792
rect 7102 11600 7158 11656
rect 6918 11192 6974 11248
rect 7820 16890 7876 16892
rect 7900 16890 7956 16892
rect 7980 16890 8036 16892
rect 8060 16890 8116 16892
rect 7820 16838 7846 16890
rect 7846 16838 7876 16890
rect 7900 16838 7910 16890
rect 7910 16838 7956 16890
rect 7980 16838 8026 16890
rect 8026 16838 8036 16890
rect 8060 16838 8090 16890
rect 8090 16838 8116 16890
rect 7820 16836 7876 16838
rect 7900 16836 7956 16838
rect 7980 16836 8036 16838
rect 8060 16836 8116 16838
rect 7820 15802 7876 15804
rect 7900 15802 7956 15804
rect 7980 15802 8036 15804
rect 8060 15802 8116 15804
rect 7820 15750 7846 15802
rect 7846 15750 7876 15802
rect 7900 15750 7910 15802
rect 7910 15750 7956 15802
rect 7980 15750 8026 15802
rect 8026 15750 8036 15802
rect 8060 15750 8090 15802
rect 8090 15750 8116 15802
rect 7820 15748 7876 15750
rect 7900 15748 7956 15750
rect 7980 15748 8036 15750
rect 8060 15748 8116 15750
rect 7820 14714 7876 14716
rect 7900 14714 7956 14716
rect 7980 14714 8036 14716
rect 8060 14714 8116 14716
rect 7820 14662 7846 14714
rect 7846 14662 7876 14714
rect 7900 14662 7910 14714
rect 7910 14662 7956 14714
rect 7980 14662 8026 14714
rect 8026 14662 8036 14714
rect 8060 14662 8090 14714
rect 8090 14662 8116 14714
rect 7820 14660 7876 14662
rect 7900 14660 7956 14662
rect 7980 14660 8036 14662
rect 8060 14660 8116 14662
rect 14684 17978 14740 17980
rect 14764 17978 14820 17980
rect 14844 17978 14900 17980
rect 14924 17978 14980 17980
rect 14684 17926 14710 17978
rect 14710 17926 14740 17978
rect 14764 17926 14774 17978
rect 14774 17926 14820 17978
rect 14844 17926 14890 17978
rect 14890 17926 14900 17978
rect 14924 17926 14954 17978
rect 14954 17926 14980 17978
rect 14684 17924 14740 17926
rect 14764 17924 14820 17926
rect 14844 17924 14900 17926
rect 14924 17924 14980 17926
rect 11252 17434 11308 17436
rect 11332 17434 11388 17436
rect 11412 17434 11468 17436
rect 11492 17434 11548 17436
rect 11252 17382 11278 17434
rect 11278 17382 11308 17434
rect 11332 17382 11342 17434
rect 11342 17382 11388 17434
rect 11412 17382 11458 17434
rect 11458 17382 11468 17434
rect 11492 17382 11522 17434
rect 11522 17382 11548 17434
rect 11252 17380 11308 17382
rect 11332 17380 11388 17382
rect 11412 17380 11468 17382
rect 11492 17380 11548 17382
rect 14684 16890 14740 16892
rect 14764 16890 14820 16892
rect 14844 16890 14900 16892
rect 14924 16890 14980 16892
rect 14684 16838 14710 16890
rect 14710 16838 14740 16890
rect 14764 16838 14774 16890
rect 14774 16838 14820 16890
rect 14844 16838 14890 16890
rect 14890 16838 14900 16890
rect 14924 16838 14954 16890
rect 14954 16838 14980 16890
rect 14684 16836 14740 16838
rect 14764 16836 14820 16838
rect 14844 16836 14900 16838
rect 14924 16836 14980 16838
rect 11252 16346 11308 16348
rect 11332 16346 11388 16348
rect 11412 16346 11468 16348
rect 11492 16346 11548 16348
rect 11252 16294 11278 16346
rect 11278 16294 11308 16346
rect 11332 16294 11342 16346
rect 11342 16294 11388 16346
rect 11412 16294 11458 16346
rect 11458 16294 11468 16346
rect 11492 16294 11522 16346
rect 11522 16294 11548 16346
rect 11252 16292 11308 16294
rect 11332 16292 11388 16294
rect 11412 16292 11468 16294
rect 11492 16292 11548 16294
rect 14684 15802 14740 15804
rect 14764 15802 14820 15804
rect 14844 15802 14900 15804
rect 14924 15802 14980 15804
rect 14684 15750 14710 15802
rect 14710 15750 14740 15802
rect 14764 15750 14774 15802
rect 14774 15750 14820 15802
rect 14844 15750 14890 15802
rect 14890 15750 14900 15802
rect 14924 15750 14954 15802
rect 14954 15750 14980 15802
rect 14684 15748 14740 15750
rect 14764 15748 14820 15750
rect 14844 15748 14900 15750
rect 14924 15748 14980 15750
rect 11252 15258 11308 15260
rect 11332 15258 11388 15260
rect 11412 15258 11468 15260
rect 11492 15258 11548 15260
rect 11252 15206 11278 15258
rect 11278 15206 11308 15258
rect 11332 15206 11342 15258
rect 11342 15206 11388 15258
rect 11412 15206 11458 15258
rect 11458 15206 11468 15258
rect 11492 15206 11522 15258
rect 11522 15206 11548 15258
rect 11252 15204 11308 15206
rect 11332 15204 11388 15206
rect 11412 15204 11468 15206
rect 11492 15204 11548 15206
rect 7820 13626 7876 13628
rect 7900 13626 7956 13628
rect 7980 13626 8036 13628
rect 8060 13626 8116 13628
rect 7820 13574 7846 13626
rect 7846 13574 7876 13626
rect 7900 13574 7910 13626
rect 7910 13574 7956 13626
rect 7980 13574 8026 13626
rect 8026 13574 8036 13626
rect 8060 13574 8090 13626
rect 8090 13574 8116 13626
rect 7820 13572 7876 13574
rect 7900 13572 7956 13574
rect 7980 13572 8036 13574
rect 8060 13572 8116 13574
rect 9586 13676 9588 13696
rect 9588 13676 9640 13696
rect 9640 13676 9642 13696
rect 9586 13640 9642 13676
rect 7562 11736 7618 11792
rect 6182 8900 6238 8936
rect 6182 8880 6184 8900
rect 6184 8880 6236 8900
rect 6236 8880 6238 8900
rect 6642 8472 6698 8528
rect 6550 8356 6606 8392
rect 6550 8336 6552 8356
rect 6552 8336 6604 8356
rect 6604 8336 6606 8356
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 6182 6160 6238 6216
rect 7378 7928 7434 7984
rect 6182 3984 6238 4040
rect 6182 2796 6184 2816
rect 6184 2796 6236 2816
rect 6236 2796 6238 2816
rect 6182 2760 6238 2796
rect 6918 2916 6974 2952
rect 6918 2896 6920 2916
rect 6920 2896 6972 2916
rect 6972 2896 6974 2916
rect 7562 8200 7618 8256
rect 7562 8084 7618 8120
rect 7562 8064 7564 8084
rect 7564 8064 7616 8084
rect 7616 8064 7618 8084
rect 7820 12538 7876 12540
rect 7900 12538 7956 12540
rect 7980 12538 8036 12540
rect 8060 12538 8116 12540
rect 7820 12486 7846 12538
rect 7846 12486 7876 12538
rect 7900 12486 7910 12538
rect 7910 12486 7956 12538
rect 7980 12486 8026 12538
rect 8026 12486 8036 12538
rect 8060 12486 8090 12538
rect 8090 12486 8116 12538
rect 7820 12484 7876 12486
rect 7900 12484 7956 12486
rect 7980 12484 8036 12486
rect 8060 12484 8116 12486
rect 8022 11756 8078 11792
rect 8022 11736 8024 11756
rect 8024 11736 8076 11756
rect 8076 11736 8078 11756
rect 8206 11500 8208 11520
rect 8208 11500 8260 11520
rect 8260 11500 8262 11520
rect 8206 11464 8262 11500
rect 7820 11450 7876 11452
rect 7900 11450 7956 11452
rect 7980 11450 8036 11452
rect 8060 11450 8116 11452
rect 7820 11398 7846 11450
rect 7846 11398 7876 11450
rect 7900 11398 7910 11450
rect 7910 11398 7956 11450
rect 7980 11398 8026 11450
rect 8026 11398 8036 11450
rect 8060 11398 8090 11450
rect 8090 11398 8116 11450
rect 7820 11396 7876 11398
rect 7900 11396 7956 11398
rect 7980 11396 8036 11398
rect 8060 11396 8116 11398
rect 8298 11192 8354 11248
rect 7820 10362 7876 10364
rect 7900 10362 7956 10364
rect 7980 10362 8036 10364
rect 8060 10362 8116 10364
rect 7820 10310 7846 10362
rect 7846 10310 7876 10362
rect 7900 10310 7910 10362
rect 7910 10310 7956 10362
rect 7980 10310 8026 10362
rect 8026 10310 8036 10362
rect 8060 10310 8090 10362
rect 8090 10310 8116 10362
rect 7820 10308 7876 10310
rect 7900 10308 7956 10310
rect 7980 10308 8036 10310
rect 8060 10308 8116 10310
rect 7838 9560 7894 9616
rect 10138 12144 10194 12200
rect 8666 11600 8722 11656
rect 9034 11228 9036 11248
rect 9036 11228 9088 11248
rect 9088 11228 9090 11248
rect 9034 11192 9090 11228
rect 8942 11056 8998 11112
rect 7820 9274 7876 9276
rect 7900 9274 7956 9276
rect 7980 9274 8036 9276
rect 8060 9274 8116 9276
rect 7820 9222 7846 9274
rect 7846 9222 7876 9274
rect 7900 9222 7910 9274
rect 7910 9222 7956 9274
rect 7980 9222 8026 9274
rect 8026 9222 8036 9274
rect 8060 9222 8090 9274
rect 8090 9222 8116 9274
rect 7820 9220 7876 9222
rect 7900 9220 7956 9222
rect 7980 9220 8036 9222
rect 8060 9220 8116 9222
rect 8574 9052 8576 9072
rect 8576 9052 8628 9072
rect 8628 9052 8630 9072
rect 10230 11600 10286 11656
rect 9862 10412 9864 10432
rect 9864 10412 9916 10432
rect 9916 10412 9918 10432
rect 9862 10376 9918 10412
rect 8574 9016 8630 9052
rect 7820 8186 7876 8188
rect 7900 8186 7956 8188
rect 7980 8186 8036 8188
rect 8060 8186 8116 8188
rect 7820 8134 7846 8186
rect 7846 8134 7876 8186
rect 7900 8134 7910 8186
rect 7910 8134 7956 8186
rect 7980 8134 8026 8186
rect 8026 8134 8036 8186
rect 8060 8134 8090 8186
rect 8090 8134 8116 8186
rect 7820 8132 7876 8134
rect 7900 8132 7956 8134
rect 7980 8132 8036 8134
rect 8060 8132 8116 8134
rect 7378 4120 7434 4176
rect 7562 3848 7618 3904
rect 7820 7098 7876 7100
rect 7900 7098 7956 7100
rect 7980 7098 8036 7100
rect 8060 7098 8116 7100
rect 7820 7046 7846 7098
rect 7846 7046 7876 7098
rect 7900 7046 7910 7098
rect 7910 7046 7956 7098
rect 7980 7046 8026 7098
rect 8026 7046 8036 7098
rect 8060 7046 8090 7098
rect 8090 7046 8116 7098
rect 7820 7044 7876 7046
rect 7900 7044 7956 7046
rect 7980 7044 8036 7046
rect 8060 7044 8116 7046
rect 9862 8472 9918 8528
rect 9678 8064 9734 8120
rect 9310 7928 9366 7984
rect 7820 6010 7876 6012
rect 7900 6010 7956 6012
rect 7980 6010 8036 6012
rect 8060 6010 8116 6012
rect 7820 5958 7846 6010
rect 7846 5958 7876 6010
rect 7900 5958 7910 6010
rect 7910 5958 7956 6010
rect 7980 5958 8026 6010
rect 8026 5958 8036 6010
rect 8060 5958 8090 6010
rect 8090 5958 8116 6010
rect 7820 5956 7876 5958
rect 7900 5956 7956 5958
rect 7980 5956 8036 5958
rect 8060 5956 8116 5958
rect 8850 5208 8906 5264
rect 7820 4922 7876 4924
rect 7900 4922 7956 4924
rect 7980 4922 8036 4924
rect 8060 4922 8116 4924
rect 7820 4870 7846 4922
rect 7846 4870 7876 4922
rect 7900 4870 7910 4922
rect 7910 4870 7956 4922
rect 7980 4870 8026 4922
rect 8026 4870 8036 4922
rect 8060 4870 8090 4922
rect 8090 4870 8116 4922
rect 7820 4868 7876 4870
rect 7900 4868 7956 4870
rect 7980 4868 8036 4870
rect 8060 4868 8116 4870
rect 7820 3834 7876 3836
rect 7900 3834 7956 3836
rect 7980 3834 8036 3836
rect 8060 3834 8116 3836
rect 7820 3782 7846 3834
rect 7846 3782 7876 3834
rect 7900 3782 7910 3834
rect 7910 3782 7956 3834
rect 7980 3782 8026 3834
rect 8026 3782 8036 3834
rect 8060 3782 8090 3834
rect 8090 3782 8116 3834
rect 7820 3780 7876 3782
rect 7900 3780 7956 3782
rect 7980 3780 8036 3782
rect 8060 3780 8116 3782
rect 7820 2746 7876 2748
rect 7900 2746 7956 2748
rect 7980 2746 8036 2748
rect 8060 2746 8116 2748
rect 7820 2694 7846 2746
rect 7846 2694 7876 2746
rect 7900 2694 7910 2746
rect 7910 2694 7956 2746
rect 7980 2694 8026 2746
rect 8026 2694 8036 2746
rect 8060 2694 8090 2746
rect 8090 2694 8116 2746
rect 7820 2692 7876 2694
rect 7900 2692 7956 2694
rect 7980 2692 8036 2694
rect 8060 2692 8116 2694
rect 8574 3848 8630 3904
rect 8390 3712 8446 3768
rect 8298 2896 8354 2952
rect 8574 3032 8630 3088
rect 9034 2932 9036 2952
rect 9036 2932 9088 2952
rect 9088 2932 9090 2952
rect 9034 2896 9090 2932
rect 9770 7384 9826 7440
rect 9678 6704 9734 6760
rect 9770 6296 9826 6352
rect 9494 6160 9550 6216
rect 9586 5208 9642 5264
rect 9586 4936 9642 4992
rect 10138 6724 10194 6760
rect 10138 6704 10140 6724
rect 10140 6704 10192 6724
rect 10192 6704 10194 6724
rect 10046 5072 10102 5128
rect 11252 14170 11308 14172
rect 11332 14170 11388 14172
rect 11412 14170 11468 14172
rect 11492 14170 11548 14172
rect 11252 14118 11278 14170
rect 11278 14118 11308 14170
rect 11332 14118 11342 14170
rect 11342 14118 11388 14170
rect 11412 14118 11458 14170
rect 11458 14118 11468 14170
rect 11492 14118 11522 14170
rect 11522 14118 11548 14170
rect 11252 14116 11308 14118
rect 11332 14116 11388 14118
rect 11412 14116 11468 14118
rect 11492 14116 11548 14118
rect 12070 13640 12126 13696
rect 11252 13082 11308 13084
rect 11332 13082 11388 13084
rect 11412 13082 11468 13084
rect 11492 13082 11548 13084
rect 11252 13030 11278 13082
rect 11278 13030 11308 13082
rect 11332 13030 11342 13082
rect 11342 13030 11388 13082
rect 11412 13030 11458 13082
rect 11458 13030 11468 13082
rect 11492 13030 11522 13082
rect 11522 13030 11548 13082
rect 11252 13028 11308 13030
rect 11332 13028 11388 13030
rect 11412 13028 11468 13030
rect 11492 13028 11548 13030
rect 10506 11328 10562 11384
rect 11150 12144 11206 12200
rect 10782 11736 10838 11792
rect 10690 11464 10746 11520
rect 10966 9968 11022 10024
rect 10966 9560 11022 9616
rect 10690 8472 10746 8528
rect 10598 7112 10654 7168
rect 10506 6296 10562 6352
rect 10414 3984 10470 4040
rect 10414 3712 10470 3768
rect 10322 3440 10378 3496
rect 10874 6840 10930 6896
rect 10874 6024 10930 6080
rect 10874 5752 10930 5808
rect 10874 3440 10930 3496
rect 11252 11994 11308 11996
rect 11332 11994 11388 11996
rect 11412 11994 11468 11996
rect 11492 11994 11548 11996
rect 11252 11942 11278 11994
rect 11278 11942 11308 11994
rect 11332 11942 11342 11994
rect 11342 11942 11388 11994
rect 11412 11942 11458 11994
rect 11458 11942 11468 11994
rect 11492 11942 11522 11994
rect 11522 11942 11548 11994
rect 11252 11940 11308 11942
rect 11332 11940 11388 11942
rect 11412 11940 11468 11942
rect 11492 11940 11548 11942
rect 11794 13268 11796 13288
rect 11796 13268 11848 13288
rect 11848 13268 11850 13288
rect 11794 13232 11850 13268
rect 11610 11056 11666 11112
rect 11252 10906 11308 10908
rect 11332 10906 11388 10908
rect 11412 10906 11468 10908
rect 11492 10906 11548 10908
rect 11252 10854 11278 10906
rect 11278 10854 11308 10906
rect 11332 10854 11342 10906
rect 11342 10854 11388 10906
rect 11412 10854 11458 10906
rect 11458 10854 11468 10906
rect 11492 10854 11522 10906
rect 11522 10854 11548 10906
rect 11252 10852 11308 10854
rect 11332 10852 11388 10854
rect 11412 10852 11468 10854
rect 11492 10852 11548 10854
rect 11610 10240 11666 10296
rect 11252 9818 11308 9820
rect 11332 9818 11388 9820
rect 11412 9818 11468 9820
rect 11492 9818 11548 9820
rect 11252 9766 11278 9818
rect 11278 9766 11308 9818
rect 11332 9766 11342 9818
rect 11342 9766 11388 9818
rect 11412 9766 11458 9818
rect 11458 9766 11468 9818
rect 11492 9766 11522 9818
rect 11522 9766 11548 9818
rect 11252 9764 11308 9766
rect 11332 9764 11388 9766
rect 11412 9764 11468 9766
rect 11492 9764 11548 9766
rect 11252 8730 11308 8732
rect 11332 8730 11388 8732
rect 11412 8730 11468 8732
rect 11492 8730 11548 8732
rect 11252 8678 11278 8730
rect 11278 8678 11308 8730
rect 11332 8678 11342 8730
rect 11342 8678 11388 8730
rect 11412 8678 11458 8730
rect 11458 8678 11468 8730
rect 11492 8678 11522 8730
rect 11522 8678 11548 8730
rect 11252 8676 11308 8678
rect 11332 8676 11388 8678
rect 11412 8676 11468 8678
rect 11492 8676 11548 8678
rect 11150 8336 11206 8392
rect 11610 8336 11666 8392
rect 11252 7642 11308 7644
rect 11332 7642 11388 7644
rect 11412 7642 11468 7644
rect 11492 7642 11548 7644
rect 11252 7590 11278 7642
rect 11278 7590 11308 7642
rect 11332 7590 11342 7642
rect 11342 7590 11388 7642
rect 11412 7590 11458 7642
rect 11458 7590 11468 7642
rect 11492 7590 11522 7642
rect 11522 7590 11548 7642
rect 11252 7588 11308 7590
rect 11332 7588 11388 7590
rect 11412 7588 11468 7590
rect 11492 7588 11548 7590
rect 11252 6554 11308 6556
rect 11332 6554 11388 6556
rect 11412 6554 11468 6556
rect 11492 6554 11548 6556
rect 11252 6502 11278 6554
rect 11278 6502 11308 6554
rect 11332 6502 11342 6554
rect 11342 6502 11388 6554
rect 11412 6502 11458 6554
rect 11458 6502 11468 6554
rect 11492 6502 11522 6554
rect 11522 6502 11548 6554
rect 11252 6500 11308 6502
rect 11332 6500 11388 6502
rect 11412 6500 11468 6502
rect 11492 6500 11548 6502
rect 11058 6024 11114 6080
rect 11242 6024 11298 6080
rect 11252 5466 11308 5468
rect 11332 5466 11388 5468
rect 11412 5466 11468 5468
rect 11492 5466 11548 5468
rect 11252 5414 11278 5466
rect 11278 5414 11308 5466
rect 11332 5414 11342 5466
rect 11342 5414 11388 5466
rect 11412 5414 11458 5466
rect 11458 5414 11468 5466
rect 11492 5414 11522 5466
rect 11522 5414 11548 5466
rect 11252 5412 11308 5414
rect 11332 5412 11388 5414
rect 11412 5412 11468 5414
rect 11492 5412 11548 5414
rect 11886 10240 11942 10296
rect 10966 2896 11022 2952
rect 11252 4378 11308 4380
rect 11332 4378 11388 4380
rect 11412 4378 11468 4380
rect 11492 4378 11548 4380
rect 11252 4326 11278 4378
rect 11278 4326 11308 4378
rect 11332 4326 11342 4378
rect 11342 4326 11388 4378
rect 11412 4326 11458 4378
rect 11458 4326 11468 4378
rect 11492 4326 11522 4378
rect 11522 4326 11548 4378
rect 11252 4324 11308 4326
rect 11332 4324 11388 4326
rect 11412 4324 11468 4326
rect 11492 4324 11548 4326
rect 11334 3984 11390 4040
rect 12438 11228 12440 11248
rect 12440 11228 12492 11248
rect 12492 11228 12494 11248
rect 12438 11192 12494 11228
rect 12254 10512 12310 10568
rect 12070 8608 12126 8664
rect 12162 8336 12218 8392
rect 13174 10240 13230 10296
rect 12438 8472 12494 8528
rect 12254 8064 12310 8120
rect 11978 7520 12034 7576
rect 12714 8880 12770 8936
rect 12806 7948 12862 7984
rect 12806 7928 12808 7948
rect 12808 7928 12860 7948
rect 12860 7928 12862 7948
rect 12714 7656 12770 7712
rect 12254 6704 12310 6760
rect 12070 5888 12126 5944
rect 11886 5652 11888 5672
rect 11888 5652 11940 5672
rect 11940 5652 11942 5672
rect 11886 5616 11942 5652
rect 11702 3848 11758 3904
rect 11886 3732 11942 3768
rect 11886 3712 11888 3732
rect 11888 3712 11940 3732
rect 11940 3712 11942 3732
rect 11252 3290 11308 3292
rect 11332 3290 11388 3292
rect 11412 3290 11468 3292
rect 11492 3290 11548 3292
rect 11252 3238 11278 3290
rect 11278 3238 11308 3290
rect 11332 3238 11342 3290
rect 11342 3238 11388 3290
rect 11412 3238 11458 3290
rect 11458 3238 11468 3290
rect 11492 3238 11522 3290
rect 11522 3238 11548 3290
rect 11252 3236 11308 3238
rect 11332 3236 11388 3238
rect 11412 3236 11468 3238
rect 11492 3236 11548 3238
rect 11252 2202 11308 2204
rect 11332 2202 11388 2204
rect 11412 2202 11468 2204
rect 11492 2202 11548 2204
rect 11252 2150 11278 2202
rect 11278 2150 11308 2202
rect 11332 2150 11342 2202
rect 11342 2150 11388 2202
rect 11412 2150 11458 2202
rect 11458 2150 11468 2202
rect 11492 2150 11522 2202
rect 11522 2150 11548 2202
rect 11252 2148 11308 2150
rect 11332 2148 11388 2150
rect 11412 2148 11468 2150
rect 11492 2148 11548 2150
rect 12162 5480 12218 5536
rect 12070 5072 12126 5128
rect 12714 6704 12770 6760
rect 12622 6160 12678 6216
rect 13174 6296 13230 6352
rect 13082 5752 13138 5808
rect 12990 5616 13046 5672
rect 12530 4276 12586 4312
rect 12530 4256 12532 4276
rect 12532 4256 12584 4276
rect 12584 4256 12586 4276
rect 12438 4156 12440 4176
rect 12440 4156 12492 4176
rect 12492 4156 12494 4176
rect 12438 4120 12494 4156
rect 13358 9424 13414 9480
rect 13910 12144 13966 12200
rect 14684 14714 14740 14716
rect 14764 14714 14820 14716
rect 14844 14714 14900 14716
rect 14924 14714 14980 14716
rect 14684 14662 14710 14714
rect 14710 14662 14740 14714
rect 14764 14662 14774 14714
rect 14774 14662 14820 14714
rect 14844 14662 14890 14714
rect 14890 14662 14900 14714
rect 14924 14662 14954 14714
rect 14954 14662 14980 14714
rect 14684 14660 14740 14662
rect 14764 14660 14820 14662
rect 14844 14660 14900 14662
rect 14924 14660 14980 14662
rect 14684 13626 14740 13628
rect 14764 13626 14820 13628
rect 14844 13626 14900 13628
rect 14924 13626 14980 13628
rect 14684 13574 14710 13626
rect 14710 13574 14740 13626
rect 14764 13574 14774 13626
rect 14774 13574 14820 13626
rect 14844 13574 14890 13626
rect 14890 13574 14900 13626
rect 14924 13574 14954 13626
rect 14954 13574 14980 13626
rect 14684 13572 14740 13574
rect 14764 13572 14820 13574
rect 14844 13572 14900 13574
rect 14924 13572 14980 13574
rect 14684 12538 14740 12540
rect 14764 12538 14820 12540
rect 14844 12538 14900 12540
rect 14924 12538 14980 12540
rect 14684 12486 14710 12538
rect 14710 12486 14740 12538
rect 14764 12486 14774 12538
rect 14774 12486 14820 12538
rect 14844 12486 14890 12538
rect 14890 12486 14900 12538
rect 14924 12486 14954 12538
rect 14954 12486 14980 12538
rect 14684 12484 14740 12486
rect 14764 12484 14820 12486
rect 14844 12484 14900 12486
rect 14924 12484 14980 12486
rect 13910 10412 13912 10432
rect 13912 10412 13964 10432
rect 13964 10412 13966 10432
rect 13910 10376 13966 10412
rect 13358 7112 13414 7168
rect 13542 6296 13598 6352
rect 13450 6024 13506 6080
rect 13542 3712 13598 3768
rect 14684 11450 14740 11452
rect 14764 11450 14820 11452
rect 14844 11450 14900 11452
rect 14924 11450 14980 11452
rect 14684 11398 14710 11450
rect 14710 11398 14740 11450
rect 14764 11398 14774 11450
rect 14774 11398 14820 11450
rect 14844 11398 14890 11450
rect 14890 11398 14900 11450
rect 14924 11398 14954 11450
rect 14954 11398 14980 11450
rect 14684 11396 14740 11398
rect 14764 11396 14820 11398
rect 14844 11396 14900 11398
rect 14924 11396 14980 11398
rect 14684 10362 14740 10364
rect 14764 10362 14820 10364
rect 14844 10362 14900 10364
rect 14924 10362 14980 10364
rect 14684 10310 14710 10362
rect 14710 10310 14740 10362
rect 14764 10310 14774 10362
rect 14774 10310 14820 10362
rect 14844 10310 14890 10362
rect 14890 10310 14900 10362
rect 14924 10310 14954 10362
rect 14954 10310 14980 10362
rect 14684 10308 14740 10310
rect 14764 10308 14820 10310
rect 14844 10308 14900 10310
rect 14924 10308 14980 10310
rect 14370 10104 14426 10160
rect 14278 9968 14334 10024
rect 13818 5888 13874 5944
rect 14002 5480 14058 5536
rect 13818 4256 13874 4312
rect 14278 7792 14334 7848
rect 14186 5752 14242 5808
rect 14684 9274 14740 9276
rect 14764 9274 14820 9276
rect 14844 9274 14900 9276
rect 14924 9274 14980 9276
rect 14684 9222 14710 9274
rect 14710 9222 14740 9274
rect 14764 9222 14774 9274
rect 14774 9222 14820 9274
rect 14844 9222 14890 9274
rect 14890 9222 14900 9274
rect 14924 9222 14954 9274
rect 14954 9222 14980 9274
rect 14684 9220 14740 9222
rect 14764 9220 14820 9222
rect 14844 9220 14900 9222
rect 14924 9220 14980 9222
rect 14554 8336 14610 8392
rect 14684 8186 14740 8188
rect 14764 8186 14820 8188
rect 14844 8186 14900 8188
rect 14924 8186 14980 8188
rect 14684 8134 14710 8186
rect 14710 8134 14740 8186
rect 14764 8134 14774 8186
rect 14774 8134 14820 8186
rect 14844 8134 14890 8186
rect 14890 8134 14900 8186
rect 14924 8134 14954 8186
rect 14954 8134 14980 8186
rect 14684 8132 14740 8134
rect 14764 8132 14820 8134
rect 14844 8132 14900 8134
rect 14924 8132 14980 8134
rect 14554 7792 14610 7848
rect 14646 7656 14702 7712
rect 14684 7098 14740 7100
rect 14764 7098 14820 7100
rect 14844 7098 14900 7100
rect 14924 7098 14980 7100
rect 14684 7046 14710 7098
rect 14710 7046 14740 7098
rect 14764 7046 14774 7098
rect 14774 7046 14820 7098
rect 14844 7046 14890 7098
rect 14890 7046 14900 7098
rect 14924 7046 14954 7098
rect 14954 7046 14980 7098
rect 14684 7044 14740 7046
rect 14764 7044 14820 7046
rect 14844 7044 14900 7046
rect 14924 7044 14980 7046
rect 14684 6010 14740 6012
rect 14764 6010 14820 6012
rect 14844 6010 14900 6012
rect 14924 6010 14980 6012
rect 14684 5958 14710 6010
rect 14710 5958 14740 6010
rect 14764 5958 14774 6010
rect 14774 5958 14820 6010
rect 14844 5958 14890 6010
rect 14890 5958 14900 6010
rect 14924 5958 14954 6010
rect 14954 5958 14980 6010
rect 14684 5956 14740 5958
rect 14764 5956 14820 5958
rect 14844 5956 14900 5958
rect 14924 5956 14980 5958
rect 14186 4936 14242 4992
rect 14684 4922 14740 4924
rect 14764 4922 14820 4924
rect 14844 4922 14900 4924
rect 14924 4922 14980 4924
rect 14684 4870 14710 4922
rect 14710 4870 14740 4922
rect 14764 4870 14774 4922
rect 14774 4870 14820 4922
rect 14844 4870 14890 4922
rect 14890 4870 14900 4922
rect 14924 4870 14954 4922
rect 14954 4870 14980 4922
rect 14684 4868 14740 4870
rect 14764 4868 14820 4870
rect 14844 4868 14900 4870
rect 14924 4868 14980 4870
rect 14094 3984 14150 4040
rect 13910 3576 13966 3632
rect 14684 3834 14740 3836
rect 14764 3834 14820 3836
rect 14844 3834 14900 3836
rect 14924 3834 14980 3836
rect 14684 3782 14710 3834
rect 14710 3782 14740 3834
rect 14764 3782 14774 3834
rect 14774 3782 14820 3834
rect 14844 3782 14890 3834
rect 14890 3782 14900 3834
rect 14924 3782 14954 3834
rect 14954 3782 14980 3834
rect 14684 3780 14740 3782
rect 14764 3780 14820 3782
rect 14844 3780 14900 3782
rect 14924 3780 14980 3782
rect 15198 4820 15254 4856
rect 15198 4800 15200 4820
rect 15200 4800 15252 4820
rect 15252 4800 15254 4820
rect 14684 2746 14740 2748
rect 14764 2746 14820 2748
rect 14844 2746 14900 2748
rect 14924 2746 14980 2748
rect 14684 2694 14710 2746
rect 14710 2694 14740 2746
rect 14764 2694 14774 2746
rect 14774 2694 14820 2746
rect 14844 2694 14890 2746
rect 14890 2694 14900 2746
rect 14924 2694 14954 2746
rect 14954 2694 14980 2746
rect 14684 2692 14740 2694
rect 14764 2692 14820 2694
rect 14844 2692 14900 2694
rect 14924 2692 14980 2694
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 18276 19610 18332 19612
rect 18356 19610 18412 19612
rect 18116 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 18276 19558 18322 19610
rect 18322 19558 18332 19610
rect 18356 19558 18386 19610
rect 18386 19558 18412 19610
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 18276 19556 18332 19558
rect 18356 19556 18412 19558
rect 17866 16904 17922 16960
rect 17130 13232 17186 13288
rect 15566 11192 15622 11248
rect 15750 10532 15806 10568
rect 15750 10512 15752 10532
rect 15752 10512 15804 10532
rect 15804 10512 15806 10532
rect 15934 8472 15990 8528
rect 15474 7520 15530 7576
rect 15566 7384 15622 7440
rect 16578 11736 16634 11792
rect 16486 10648 16542 10704
rect 16302 7948 16358 7984
rect 16302 7928 16304 7948
rect 16304 7928 16356 7948
rect 16356 7928 16358 7948
rect 16394 6860 16450 6896
rect 16394 6840 16396 6860
rect 16396 6840 16448 6860
rect 16448 6840 16450 6860
rect 16854 12144 16910 12200
rect 17038 11736 17094 11792
rect 16854 10512 16910 10568
rect 16670 8608 16726 8664
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 18276 18522 18332 18524
rect 18356 18522 18412 18524
rect 18116 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 18276 18470 18322 18522
rect 18322 18470 18332 18522
rect 18356 18470 18386 18522
rect 18386 18470 18412 18522
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 18276 18468 18332 18470
rect 18356 18468 18412 18470
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 18276 17434 18332 17436
rect 18356 17434 18412 17436
rect 18116 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 18276 17382 18322 17434
rect 18322 17382 18332 17434
rect 18356 17382 18386 17434
rect 18386 17382 18412 17434
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18276 17380 18332 17382
rect 18356 17380 18412 17382
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 18276 16346 18332 16348
rect 18356 16346 18412 16348
rect 18116 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 18276 16294 18322 16346
rect 18322 16294 18332 16346
rect 18356 16294 18386 16346
rect 18386 16294 18412 16346
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 18276 16292 18332 16294
rect 18356 16292 18412 16294
rect 18694 15544 18750 15600
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 18276 15258 18332 15260
rect 18356 15258 18412 15260
rect 18116 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 18276 15206 18322 15258
rect 18322 15206 18332 15258
rect 18356 15206 18386 15258
rect 18386 15206 18412 15258
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18276 15204 18332 15206
rect 18356 15204 18412 15206
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 18276 14170 18332 14172
rect 18356 14170 18412 14172
rect 18116 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 18276 14118 18322 14170
rect 18322 14118 18332 14170
rect 18356 14118 18386 14170
rect 18386 14118 18412 14170
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18276 14116 18332 14118
rect 18356 14116 18412 14118
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 18276 13082 18332 13084
rect 18356 13082 18412 13084
rect 18116 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 18276 13030 18322 13082
rect 18322 13030 18332 13082
rect 18356 13030 18386 13082
rect 18386 13030 18412 13082
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18276 13028 18332 13030
rect 18356 13028 18412 13030
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 18276 11994 18332 11996
rect 18356 11994 18412 11996
rect 18116 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 18276 11942 18322 11994
rect 18322 11942 18332 11994
rect 18356 11942 18386 11994
rect 18386 11942 18412 11994
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 18276 11940 18332 11942
rect 18356 11940 18412 11942
rect 17774 11192 17830 11248
rect 17130 8336 17186 8392
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 18276 10906 18332 10908
rect 18356 10906 18412 10908
rect 18116 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 18276 10854 18322 10906
rect 18322 10854 18332 10906
rect 18356 10854 18386 10906
rect 18386 10854 18412 10906
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18276 10852 18332 10854
rect 18356 10852 18412 10854
rect 18050 10376 18106 10432
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 18276 9818 18332 9820
rect 18356 9818 18412 9820
rect 18116 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 18276 9766 18322 9818
rect 18322 9766 18332 9818
rect 18356 9766 18386 9818
rect 18386 9766 18412 9818
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 18276 9764 18332 9766
rect 18356 9764 18412 9766
rect 18510 9560 18566 9616
rect 18510 9016 18566 9072
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 18276 8730 18332 8732
rect 18356 8730 18412 8732
rect 18116 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 18276 8678 18322 8730
rect 18322 8678 18332 8730
rect 18356 8678 18386 8730
rect 18386 8678 18412 8730
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18276 8676 18332 8678
rect 18356 8676 18412 8678
rect 17958 8472 18014 8528
rect 17774 7112 17830 7168
rect 17590 2760 17646 2816
rect 17590 2624 17646 2680
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 18276 7642 18332 7644
rect 18356 7642 18412 7644
rect 18116 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 18276 7590 18322 7642
rect 18322 7590 18332 7642
rect 18356 7590 18386 7642
rect 18386 7590 18412 7642
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18276 7588 18332 7590
rect 18356 7588 18412 7590
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 18276 6554 18332 6556
rect 18356 6554 18412 6556
rect 18116 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 18276 6502 18322 6554
rect 18322 6502 18332 6554
rect 18356 6502 18386 6554
rect 18386 6502 18412 6554
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18276 6500 18332 6502
rect 18356 6500 18412 6502
rect 18142 6160 18198 6216
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 18276 5466 18332 5468
rect 18356 5466 18412 5468
rect 18116 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 18276 5414 18322 5466
rect 18322 5414 18332 5466
rect 18356 5414 18386 5466
rect 18386 5414 18412 5466
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18276 5412 18332 5414
rect 18356 5412 18412 5414
rect 17958 5208 18014 5264
rect 18970 14068 19026 14104
rect 18970 14048 18972 14068
rect 18972 14048 19024 14068
rect 19024 14048 19026 14068
rect 18970 11328 19026 11384
rect 18786 7520 18842 7576
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 18276 4378 18332 4380
rect 18356 4378 18412 4380
rect 18116 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 18276 4326 18322 4378
rect 18322 4326 18332 4378
rect 18356 4326 18386 4378
rect 18386 4326 18412 4378
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18276 4324 18332 4326
rect 18356 4324 18412 4326
rect 18234 3612 18236 3632
rect 18236 3612 18288 3632
rect 18288 3612 18290 3632
rect 18234 3576 18290 3612
rect 18142 3440 18198 3496
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 18276 3290 18332 3292
rect 18356 3290 18412 3292
rect 18116 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 18276 3238 18322 3290
rect 18322 3238 18332 3290
rect 18356 3238 18386 3290
rect 18386 3238 18412 3290
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 18276 3236 18332 3238
rect 18356 3236 18412 3238
rect 17958 2760 18014 2816
rect 18510 2760 18566 2816
rect 18234 2624 18290 2680
rect 20902 22072 20958 22128
rect 20626 21528 20682 21584
rect 20258 21120 20314 21176
rect 19154 20576 19210 20632
rect 19614 15036 19616 15056
rect 19616 15036 19668 15056
rect 19668 15036 19670 15056
rect 19614 15000 19670 15036
rect 19246 14592 19302 14648
rect 19338 13232 19394 13288
rect 19246 12688 19302 12744
rect 19430 12144 19486 12200
rect 19246 11600 19302 11656
rect 19246 10784 19302 10840
rect 19890 12552 19946 12608
rect 20166 16496 20222 16552
rect 20442 19216 20498 19272
rect 20350 18128 20406 18184
rect 20534 18264 20590 18320
rect 20442 15952 20498 16008
rect 19246 8064 19302 8120
rect 19154 7828 19156 7848
rect 19156 7828 19208 7848
rect 19208 7828 19210 7848
rect 19154 7792 19210 7828
rect 19062 6296 19118 6352
rect 18786 2760 18842 2816
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 18276 2202 18332 2204
rect 18356 2202 18412 2204
rect 18116 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 18276 2150 18322 2202
rect 18322 2150 18332 2202
rect 18356 2150 18386 2202
rect 18386 2150 18412 2202
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 18276 2148 18332 2150
rect 18356 2148 18412 2150
rect 5630 176 5686 232
rect 19246 3848 19302 3904
rect 19154 2760 19210 2816
rect 20442 13640 20498 13696
rect 20350 12280 20406 12336
rect 20718 19760 20774 19816
rect 20718 18808 20774 18864
rect 20718 17856 20774 17912
rect 20810 17312 20866 17368
rect 20994 20168 21050 20224
rect 20718 12552 20774 12608
rect 20718 4256 20774 4312
rect 20074 3576 20130 3632
rect 19246 1944 19302 2000
rect 20442 2896 20498 2952
rect 20810 2624 20866 2680
rect 20810 1536 20866 1592
rect 20534 992 20590 1048
rect 20902 584 20958 640
rect 18786 176 18842 232
<< metal3 >>
rect 0 22538 480 22568
rect 2957 22538 3023 22541
rect 0 22536 3023 22538
rect 0 22480 2962 22536
rect 3018 22480 3023 22536
rect 0 22478 3023 22480
rect 0 22448 480 22478
rect 2957 22475 3023 22478
rect 19057 22538 19123 22541
rect 22320 22538 22800 22568
rect 19057 22536 22800 22538
rect 19057 22480 19062 22536
rect 19118 22480 22800 22536
rect 19057 22478 22800 22480
rect 19057 22475 19123 22478
rect 22320 22448 22800 22478
rect 0 22130 480 22160
rect 2313 22130 2379 22133
rect 0 22128 2379 22130
rect 0 22072 2318 22128
rect 2374 22072 2379 22128
rect 0 22070 2379 22072
rect 0 22040 480 22070
rect 2313 22067 2379 22070
rect 20897 22130 20963 22133
rect 22320 22130 22800 22160
rect 20897 22128 22800 22130
rect 20897 22072 20902 22128
rect 20958 22072 22800 22128
rect 20897 22070 22800 22072
rect 20897 22067 20963 22070
rect 22320 22040 22800 22070
rect 0 21586 480 21616
rect 3141 21586 3207 21589
rect 0 21584 3207 21586
rect 0 21528 3146 21584
rect 3202 21528 3207 21584
rect 0 21526 3207 21528
rect 0 21496 480 21526
rect 3141 21523 3207 21526
rect 20621 21586 20687 21589
rect 22320 21586 22800 21616
rect 20621 21584 22800 21586
rect 20621 21528 20626 21584
rect 20682 21528 22800 21584
rect 20621 21526 22800 21528
rect 20621 21523 20687 21526
rect 22320 21496 22800 21526
rect 0 21178 480 21208
rect 2497 21178 2563 21181
rect 0 21176 2563 21178
rect 0 21120 2502 21176
rect 2558 21120 2563 21176
rect 0 21118 2563 21120
rect 0 21088 480 21118
rect 2497 21115 2563 21118
rect 20253 21178 20319 21181
rect 22320 21178 22800 21208
rect 20253 21176 22800 21178
rect 20253 21120 20258 21176
rect 20314 21120 22800 21176
rect 20253 21118 22800 21120
rect 20253 21115 20319 21118
rect 22320 21088 22800 21118
rect 0 20634 480 20664
rect 3693 20634 3759 20637
rect 0 20632 3759 20634
rect 0 20576 3698 20632
rect 3754 20576 3759 20632
rect 0 20574 3759 20576
rect 0 20544 480 20574
rect 3693 20571 3759 20574
rect 19149 20634 19215 20637
rect 22320 20634 22800 20664
rect 19149 20632 22800 20634
rect 19149 20576 19154 20632
rect 19210 20576 22800 20632
rect 19149 20574 22800 20576
rect 19149 20571 19215 20574
rect 22320 20544 22800 20574
rect 0 20226 480 20256
rect 2773 20226 2839 20229
rect 0 20224 2839 20226
rect 0 20168 2778 20224
rect 2834 20168 2839 20224
rect 0 20166 2839 20168
rect 0 20136 480 20166
rect 2773 20163 2839 20166
rect 20989 20226 21055 20229
rect 22320 20226 22800 20256
rect 20989 20224 22800 20226
rect 20989 20168 20994 20224
rect 21050 20168 22800 20224
rect 20989 20166 22800 20168
rect 20989 20163 21055 20166
rect 7808 20160 8128 20161
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 20095 8128 20096
rect 14672 20160 14992 20161
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 22320 20136 22800 20166
rect 14672 20095 14992 20096
rect 0 19818 480 19848
rect 1945 19818 2011 19821
rect 0 19816 2011 19818
rect 0 19760 1950 19816
rect 2006 19760 2011 19816
rect 0 19758 2011 19760
rect 0 19728 480 19758
rect 1945 19755 2011 19758
rect 20713 19818 20779 19821
rect 22320 19818 22800 19848
rect 20713 19816 22800 19818
rect 20713 19760 20718 19816
rect 20774 19760 22800 19816
rect 20713 19758 22800 19760
rect 20713 19755 20779 19758
rect 22320 19728 22800 19758
rect 4376 19616 4696 19617
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 19551 4696 19552
rect 11240 19616 11560 19617
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 19551 11560 19552
rect 18104 19616 18424 19617
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 19551 18424 19552
rect 0 19274 480 19304
rect 1945 19274 2011 19277
rect 0 19272 2011 19274
rect 0 19216 1950 19272
rect 2006 19216 2011 19272
rect 0 19214 2011 19216
rect 0 19184 480 19214
rect 1945 19211 2011 19214
rect 20437 19274 20503 19277
rect 22320 19274 22800 19304
rect 20437 19272 22800 19274
rect 20437 19216 20442 19272
rect 20498 19216 22800 19272
rect 20437 19214 22800 19216
rect 20437 19211 20503 19214
rect 22320 19184 22800 19214
rect 7808 19072 8128 19073
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 19007 8128 19008
rect 14672 19072 14992 19073
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 19007 14992 19008
rect 0 18866 480 18896
rect 1945 18866 2011 18869
rect 0 18864 2011 18866
rect 0 18808 1950 18864
rect 2006 18808 2011 18864
rect 0 18806 2011 18808
rect 0 18776 480 18806
rect 1945 18803 2011 18806
rect 20713 18866 20779 18869
rect 22320 18866 22800 18896
rect 20713 18864 22800 18866
rect 20713 18808 20718 18864
rect 20774 18808 22800 18864
rect 20713 18806 22800 18808
rect 20713 18803 20779 18806
rect 22320 18776 22800 18806
rect 4376 18528 4696 18529
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 18463 4696 18464
rect 11240 18528 11560 18529
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 18463 11560 18464
rect 18104 18528 18424 18529
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 18463 18424 18464
rect 0 18322 480 18352
rect 1853 18322 1919 18325
rect 0 18320 1919 18322
rect 0 18264 1858 18320
rect 1914 18264 1919 18320
rect 0 18262 1919 18264
rect 0 18232 480 18262
rect 1853 18259 1919 18262
rect 19926 18260 19932 18324
rect 19996 18322 20002 18324
rect 20529 18322 20595 18325
rect 22320 18322 22800 18352
rect 19996 18320 20595 18322
rect 19996 18264 20534 18320
rect 20590 18264 20595 18320
rect 19996 18262 20595 18264
rect 19996 18260 20002 18262
rect 20529 18259 20595 18262
rect 20854 18262 22800 18322
rect 20345 18186 20411 18189
rect 20854 18186 20914 18262
rect 22320 18232 22800 18262
rect 20345 18184 20914 18186
rect 20345 18128 20350 18184
rect 20406 18128 20914 18184
rect 20345 18126 20914 18128
rect 20345 18123 20411 18126
rect 7808 17984 8128 17985
rect 0 17914 480 17944
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 17919 8128 17920
rect 14672 17984 14992 17985
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 17919 14992 17920
rect 1669 17914 1735 17917
rect 0 17912 1735 17914
rect 0 17856 1674 17912
rect 1730 17856 1735 17912
rect 0 17854 1735 17856
rect 0 17824 480 17854
rect 1669 17851 1735 17854
rect 20713 17914 20779 17917
rect 22320 17914 22800 17944
rect 20713 17912 22800 17914
rect 20713 17856 20718 17912
rect 20774 17856 22800 17912
rect 20713 17854 22800 17856
rect 20713 17851 20779 17854
rect 22320 17824 22800 17854
rect 4376 17440 4696 17441
rect 0 17370 480 17400
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 17375 4696 17376
rect 11240 17440 11560 17441
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 17375 11560 17376
rect 18104 17440 18424 17441
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 17375 18424 17376
rect 1945 17370 2011 17373
rect 0 17368 2011 17370
rect 0 17312 1950 17368
rect 2006 17312 2011 17368
rect 0 17310 2011 17312
rect 0 17280 480 17310
rect 1945 17307 2011 17310
rect 20805 17370 20871 17373
rect 22320 17370 22800 17400
rect 20805 17368 22800 17370
rect 20805 17312 20810 17368
rect 20866 17312 22800 17368
rect 20805 17310 22800 17312
rect 20805 17307 20871 17310
rect 22320 17280 22800 17310
rect 0 16962 480 16992
rect 3417 16962 3483 16965
rect 0 16960 3483 16962
rect 0 16904 3422 16960
rect 3478 16904 3483 16960
rect 0 16902 3483 16904
rect 0 16872 480 16902
rect 3417 16899 3483 16902
rect 17861 16962 17927 16965
rect 22320 16962 22800 16992
rect 17861 16960 22800 16962
rect 17861 16904 17866 16960
rect 17922 16904 22800 16960
rect 17861 16902 22800 16904
rect 17861 16899 17927 16902
rect 7808 16896 8128 16897
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 16831 8128 16832
rect 14672 16896 14992 16897
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 22320 16872 22800 16902
rect 14672 16831 14992 16832
rect 0 16554 480 16584
rect 1945 16554 2011 16557
rect 0 16552 2011 16554
rect 0 16496 1950 16552
rect 2006 16496 2011 16552
rect 0 16494 2011 16496
rect 0 16464 480 16494
rect 1945 16491 2011 16494
rect 20161 16554 20227 16557
rect 22320 16554 22800 16584
rect 20161 16552 22800 16554
rect 20161 16496 20166 16552
rect 20222 16496 22800 16552
rect 20161 16494 22800 16496
rect 20161 16491 20227 16494
rect 22320 16464 22800 16494
rect 4376 16352 4696 16353
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 16287 4696 16288
rect 11240 16352 11560 16353
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 16287 11560 16288
rect 18104 16352 18424 16353
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 16287 18424 16288
rect 0 16010 480 16040
rect 1945 16010 2011 16013
rect 0 16008 2011 16010
rect 0 15952 1950 16008
rect 2006 15952 2011 16008
rect 0 15950 2011 15952
rect 0 15920 480 15950
rect 1945 15947 2011 15950
rect 20437 16010 20503 16013
rect 22320 16010 22800 16040
rect 20437 16008 22800 16010
rect 20437 15952 20442 16008
rect 20498 15952 22800 16008
rect 20437 15950 22800 15952
rect 20437 15947 20503 15950
rect 22320 15920 22800 15950
rect 7808 15808 8128 15809
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 15743 8128 15744
rect 14672 15808 14992 15809
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 15743 14992 15744
rect 0 15602 480 15632
rect 2773 15602 2839 15605
rect 0 15600 2839 15602
rect 0 15544 2778 15600
rect 2834 15544 2839 15600
rect 0 15542 2839 15544
rect 0 15512 480 15542
rect 2773 15539 2839 15542
rect 18689 15602 18755 15605
rect 22320 15602 22800 15632
rect 18689 15600 22800 15602
rect 18689 15544 18694 15600
rect 18750 15544 22800 15600
rect 18689 15542 22800 15544
rect 18689 15539 18755 15542
rect 22320 15512 22800 15542
rect 4376 15264 4696 15265
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 15199 4696 15200
rect 11240 15264 11560 15265
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 15199 11560 15200
rect 18104 15264 18424 15265
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 15199 18424 15200
rect 0 15058 480 15088
rect 1945 15058 2011 15061
rect 0 15056 2011 15058
rect 0 15000 1950 15056
rect 2006 15000 2011 15056
rect 0 14998 2011 15000
rect 0 14968 480 14998
rect 1945 14995 2011 14998
rect 19609 15058 19675 15061
rect 22320 15058 22800 15088
rect 19609 15056 22800 15058
rect 19609 15000 19614 15056
rect 19670 15000 22800 15056
rect 19609 14998 22800 15000
rect 19609 14995 19675 14998
rect 22320 14968 22800 14998
rect 7808 14720 8128 14721
rect 0 14650 480 14680
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 14655 8128 14656
rect 14672 14720 14992 14721
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 14655 14992 14656
rect 1669 14650 1735 14653
rect 0 14648 1735 14650
rect 0 14592 1674 14648
rect 1730 14592 1735 14648
rect 0 14590 1735 14592
rect 0 14560 480 14590
rect 1669 14587 1735 14590
rect 19241 14650 19307 14653
rect 22320 14650 22800 14680
rect 19241 14648 22800 14650
rect 19241 14592 19246 14648
rect 19302 14592 22800 14648
rect 19241 14590 22800 14592
rect 19241 14587 19307 14590
rect 22320 14560 22800 14590
rect 4376 14176 4696 14177
rect 0 14106 480 14136
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 14111 4696 14112
rect 11240 14176 11560 14177
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 14111 11560 14112
rect 18104 14176 18424 14177
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 14111 18424 14112
rect 1577 14106 1643 14109
rect 0 14104 1643 14106
rect 0 14048 1582 14104
rect 1638 14048 1643 14104
rect 0 14046 1643 14048
rect 0 14016 480 14046
rect 1577 14043 1643 14046
rect 18965 14106 19031 14109
rect 22320 14106 22800 14136
rect 18965 14104 22800 14106
rect 18965 14048 18970 14104
rect 19026 14048 22800 14104
rect 18965 14046 22800 14048
rect 18965 14043 19031 14046
rect 22320 14016 22800 14046
rect 0 13698 480 13728
rect 3325 13698 3391 13701
rect 0 13696 3391 13698
rect 0 13640 3330 13696
rect 3386 13640 3391 13696
rect 0 13638 3391 13640
rect 0 13608 480 13638
rect 3325 13635 3391 13638
rect 9581 13698 9647 13701
rect 12065 13698 12131 13701
rect 9581 13696 12131 13698
rect 9581 13640 9586 13696
rect 9642 13640 12070 13696
rect 12126 13640 12131 13696
rect 9581 13638 12131 13640
rect 9581 13635 9647 13638
rect 12065 13635 12131 13638
rect 20437 13698 20503 13701
rect 22320 13698 22800 13728
rect 20437 13696 22800 13698
rect 20437 13640 20442 13696
rect 20498 13640 22800 13696
rect 20437 13638 22800 13640
rect 20437 13635 20503 13638
rect 7808 13632 8128 13633
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 13567 8128 13568
rect 14672 13632 14992 13633
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 22320 13608 22800 13638
rect 14672 13567 14992 13568
rect 0 13290 480 13320
rect 3601 13290 3667 13293
rect 0 13288 3667 13290
rect 0 13232 3606 13288
rect 3662 13232 3667 13288
rect 0 13230 3667 13232
rect 0 13200 480 13230
rect 3601 13227 3667 13230
rect 11789 13290 11855 13293
rect 17125 13290 17191 13293
rect 11789 13288 17191 13290
rect 11789 13232 11794 13288
rect 11850 13232 17130 13288
rect 17186 13232 17191 13288
rect 11789 13230 17191 13232
rect 11789 13227 11855 13230
rect 17125 13227 17191 13230
rect 19333 13290 19399 13293
rect 22320 13290 22800 13320
rect 19333 13288 22800 13290
rect 19333 13232 19338 13288
rect 19394 13232 22800 13288
rect 19333 13230 22800 13232
rect 19333 13227 19399 13230
rect 22320 13200 22800 13230
rect 4376 13088 4696 13089
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 13023 4696 13024
rect 11240 13088 11560 13089
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 13023 11560 13024
rect 18104 13088 18424 13089
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 13023 18424 13024
rect 0 12746 480 12776
rect 3969 12746 4035 12749
rect 0 12744 4035 12746
rect 0 12688 3974 12744
rect 4030 12688 4035 12744
rect 0 12686 4035 12688
rect 0 12656 480 12686
rect 3969 12683 4035 12686
rect 19241 12746 19307 12749
rect 22320 12746 22800 12776
rect 19241 12744 22800 12746
rect 19241 12688 19246 12744
rect 19302 12688 22800 12744
rect 19241 12686 22800 12688
rect 19241 12683 19307 12686
rect 22320 12656 22800 12686
rect 19885 12610 19951 12613
rect 20713 12610 20779 12613
rect 19885 12608 20779 12610
rect 19885 12552 19890 12608
rect 19946 12552 20718 12608
rect 20774 12552 20779 12608
rect 19885 12550 20779 12552
rect 19885 12547 19951 12550
rect 20713 12547 20779 12550
rect 7808 12544 8128 12545
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 12479 8128 12480
rect 14672 12544 14992 12545
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 12479 14992 12480
rect 0 12338 480 12368
rect 3877 12338 3943 12341
rect 0 12336 3943 12338
rect 0 12280 3882 12336
rect 3938 12280 3943 12336
rect 0 12278 3943 12280
rect 0 12248 480 12278
rect 3877 12275 3943 12278
rect 20345 12338 20411 12341
rect 22320 12338 22800 12368
rect 20345 12336 22800 12338
rect 20345 12280 20350 12336
rect 20406 12280 22800 12336
rect 20345 12278 22800 12280
rect 20345 12275 20411 12278
rect 22320 12248 22800 12278
rect 10133 12202 10199 12205
rect 11145 12202 11211 12205
rect 13905 12202 13971 12205
rect 10133 12200 13971 12202
rect 10133 12144 10138 12200
rect 10194 12144 11150 12200
rect 11206 12144 13910 12200
rect 13966 12144 13971 12200
rect 10133 12142 13971 12144
rect 10133 12139 10199 12142
rect 11145 12139 11211 12142
rect 13905 12139 13971 12142
rect 16849 12202 16915 12205
rect 19425 12202 19491 12205
rect 16849 12200 19491 12202
rect 16849 12144 16854 12200
rect 16910 12144 19430 12200
rect 19486 12144 19491 12200
rect 16849 12142 19491 12144
rect 16849 12139 16915 12142
rect 19425 12139 19491 12142
rect 4376 12000 4696 12001
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 11935 4696 11936
rect 11240 12000 11560 12001
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 11935 11560 11936
rect 18104 12000 18424 12001
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 11935 18424 11936
rect 0 11794 480 11824
rect 4061 11794 4127 11797
rect 0 11792 4127 11794
rect 0 11736 4066 11792
rect 4122 11736 4127 11792
rect 0 11734 4127 11736
rect 0 11704 480 11734
rect 4061 11731 4127 11734
rect 7005 11794 7071 11797
rect 7557 11794 7623 11797
rect 8017 11794 8083 11797
rect 7005 11792 8083 11794
rect 7005 11736 7010 11792
rect 7066 11736 7562 11792
rect 7618 11736 8022 11792
rect 8078 11736 8083 11792
rect 7005 11734 8083 11736
rect 7005 11731 7071 11734
rect 7557 11731 7623 11734
rect 8017 11731 8083 11734
rect 10777 11794 10843 11797
rect 16573 11794 16639 11797
rect 10777 11792 16639 11794
rect 10777 11736 10782 11792
rect 10838 11736 16578 11792
rect 16634 11736 16639 11792
rect 10777 11734 16639 11736
rect 10777 11731 10843 11734
rect 16573 11731 16639 11734
rect 17033 11794 17099 11797
rect 22320 11794 22800 11824
rect 17033 11792 22800 11794
rect 17033 11736 17038 11792
rect 17094 11736 22800 11792
rect 17033 11734 22800 11736
rect 17033 11731 17099 11734
rect 22320 11704 22800 11734
rect 7097 11658 7163 11661
rect 8661 11658 8727 11661
rect 7097 11656 8727 11658
rect 7097 11600 7102 11656
rect 7158 11600 8666 11656
rect 8722 11600 8727 11656
rect 7097 11598 8727 11600
rect 7097 11595 7163 11598
rect 8661 11595 8727 11598
rect 10225 11658 10291 11661
rect 19241 11658 19307 11661
rect 10225 11656 19307 11658
rect 10225 11600 10230 11656
rect 10286 11600 19246 11656
rect 19302 11600 19307 11656
rect 10225 11598 19307 11600
rect 10225 11595 10291 11598
rect 19241 11595 19307 11598
rect 8201 11522 8267 11525
rect 10685 11522 10751 11525
rect 8201 11520 10751 11522
rect 8201 11464 8206 11520
rect 8262 11464 10690 11520
rect 10746 11464 10751 11520
rect 8201 11462 10751 11464
rect 8201 11459 8267 11462
rect 10685 11459 10751 11462
rect 7808 11456 8128 11457
rect 0 11386 480 11416
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 11391 8128 11392
rect 14672 11456 14992 11457
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 11391 14992 11392
rect 5993 11386 6059 11389
rect 0 11384 6059 11386
rect 0 11328 5998 11384
rect 6054 11328 6059 11384
rect 0 11326 6059 11328
rect 0 11296 480 11326
rect 5993 11323 6059 11326
rect 10501 11386 10567 11389
rect 18965 11386 19031 11389
rect 22320 11386 22800 11416
rect 10501 11384 14474 11386
rect 10501 11328 10506 11384
rect 10562 11328 14474 11384
rect 10501 11326 14474 11328
rect 10501 11323 10567 11326
rect 6913 11250 6979 11253
rect 8293 11250 8359 11253
rect 6913 11248 8359 11250
rect 6913 11192 6918 11248
rect 6974 11192 8298 11248
rect 8354 11192 8359 11248
rect 6913 11190 8359 11192
rect 6913 11187 6979 11190
rect 8293 11187 8359 11190
rect 9029 11250 9095 11253
rect 12433 11250 12499 11253
rect 9029 11248 12499 11250
rect 9029 11192 9034 11248
rect 9090 11192 12438 11248
rect 12494 11192 12499 11248
rect 9029 11190 12499 11192
rect 14414 11250 14474 11326
rect 18965 11384 22800 11386
rect 18965 11328 18970 11384
rect 19026 11328 22800 11384
rect 18965 11326 22800 11328
rect 18965 11323 19031 11326
rect 22320 11296 22800 11326
rect 15561 11250 15627 11253
rect 17769 11250 17835 11253
rect 14414 11248 17835 11250
rect 14414 11192 15566 11248
rect 15622 11192 17774 11248
rect 17830 11192 17835 11248
rect 14414 11190 17835 11192
rect 9029 11187 9095 11190
rect 12433 11187 12499 11190
rect 15561 11187 15627 11190
rect 17769 11187 17835 11190
rect 8937 11114 9003 11117
rect 11605 11114 11671 11117
rect 8937 11112 11671 11114
rect 8937 11056 8942 11112
rect 8998 11056 11610 11112
rect 11666 11056 11671 11112
rect 8937 11054 11671 11056
rect 8937 11051 9003 11054
rect 11605 11051 11671 11054
rect 4376 10912 4696 10913
rect 0 10842 480 10872
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 10847 4696 10848
rect 11240 10912 11560 10913
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 10847 11560 10848
rect 18104 10912 18424 10913
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 10847 18424 10848
rect 3877 10842 3943 10845
rect 0 10840 3943 10842
rect 0 10784 3882 10840
rect 3938 10784 3943 10840
rect 0 10782 3943 10784
rect 0 10752 480 10782
rect 3877 10779 3943 10782
rect 19241 10842 19307 10845
rect 22320 10842 22800 10872
rect 19241 10840 22800 10842
rect 19241 10784 19246 10840
rect 19302 10784 22800 10840
rect 19241 10782 22800 10784
rect 19241 10779 19307 10782
rect 22320 10752 22800 10782
rect 1485 10706 1551 10709
rect 6085 10706 6151 10709
rect 16481 10706 16547 10709
rect 19926 10706 19932 10708
rect 1485 10704 6151 10706
rect 1485 10648 1490 10704
rect 1546 10648 6090 10704
rect 6146 10648 6151 10704
rect 1485 10646 6151 10648
rect 1485 10643 1551 10646
rect 6085 10643 6151 10646
rect 15518 10704 19932 10706
rect 15518 10648 16486 10704
rect 16542 10648 19932 10704
rect 15518 10646 19932 10648
rect 4613 10570 4679 10573
rect 4889 10570 4955 10573
rect 4613 10568 4955 10570
rect 4613 10512 4618 10568
rect 4674 10512 4894 10568
rect 4950 10512 4955 10568
rect 4613 10510 4955 10512
rect 4613 10507 4679 10510
rect 4889 10507 4955 10510
rect 12249 10570 12315 10573
rect 15518 10570 15578 10646
rect 16481 10643 16547 10646
rect 19926 10644 19932 10646
rect 19996 10644 20002 10708
rect 12249 10568 15578 10570
rect 12249 10512 12254 10568
rect 12310 10512 15578 10568
rect 12249 10510 15578 10512
rect 15745 10570 15811 10573
rect 16849 10570 16915 10573
rect 15745 10568 16915 10570
rect 15745 10512 15750 10568
rect 15806 10512 16854 10568
rect 16910 10512 16915 10568
rect 15745 10510 16915 10512
rect 12249 10507 12315 10510
rect 15745 10507 15811 10510
rect 16849 10507 16915 10510
rect 0 10434 480 10464
rect 4061 10434 4127 10437
rect 0 10432 4127 10434
rect 0 10376 4066 10432
rect 4122 10376 4127 10432
rect 0 10374 4127 10376
rect 0 10344 480 10374
rect 4061 10371 4127 10374
rect 9857 10434 9923 10437
rect 13905 10434 13971 10437
rect 9857 10432 13971 10434
rect 9857 10376 9862 10432
rect 9918 10376 13910 10432
rect 13966 10376 13971 10432
rect 9857 10374 13971 10376
rect 9857 10371 9923 10374
rect 13905 10371 13971 10374
rect 18045 10434 18111 10437
rect 22320 10434 22800 10464
rect 18045 10432 22800 10434
rect 18045 10376 18050 10432
rect 18106 10376 22800 10432
rect 18045 10374 22800 10376
rect 18045 10371 18111 10374
rect 7808 10368 8128 10369
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 10303 8128 10304
rect 14672 10368 14992 10369
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 22320 10344 22800 10374
rect 14672 10303 14992 10304
rect 11605 10298 11671 10301
rect 11881 10298 11947 10301
rect 13169 10298 13235 10301
rect 11605 10296 13235 10298
rect 11605 10240 11610 10296
rect 11666 10240 11886 10296
rect 11942 10240 13174 10296
rect 13230 10240 13235 10296
rect 11605 10238 13235 10240
rect 11605 10235 11671 10238
rect 11881 10235 11947 10238
rect 13169 10235 13235 10238
rect 2589 10162 2655 10165
rect 5349 10162 5415 10165
rect 14365 10162 14431 10165
rect 2589 10160 4906 10162
rect 2589 10104 2594 10160
rect 2650 10104 4906 10160
rect 2589 10102 4906 10104
rect 2589 10099 2655 10102
rect 0 10026 480 10056
rect 3693 10026 3759 10029
rect 0 10024 3759 10026
rect 0 9968 3698 10024
rect 3754 9968 3759 10024
rect 0 9966 3759 9968
rect 0 9936 480 9966
rect 3693 9963 3759 9966
rect 4376 9824 4696 9825
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 9759 4696 9760
rect 0 9482 480 9512
rect 4061 9482 4127 9485
rect 0 9480 4127 9482
rect 0 9424 4066 9480
rect 4122 9424 4127 9480
rect 0 9422 4127 9424
rect 4846 9482 4906 10102
rect 5349 10160 18154 10162
rect 5349 10104 5354 10160
rect 5410 10104 14370 10160
rect 14426 10104 18154 10160
rect 5349 10102 18154 10104
rect 5349 10099 5415 10102
rect 14365 10099 14431 10102
rect 10961 10026 11027 10029
rect 14273 10026 14339 10029
rect 10961 10024 14339 10026
rect 10961 9968 10966 10024
rect 11022 9968 14278 10024
rect 14334 9968 14339 10024
rect 10961 9966 14339 9968
rect 18094 10026 18154 10102
rect 22320 10026 22800 10056
rect 18094 9966 22800 10026
rect 10961 9963 11027 9966
rect 14273 9963 14339 9966
rect 22320 9936 22800 9966
rect 11240 9824 11560 9825
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 11240 9759 11560 9760
rect 18104 9824 18424 9825
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 9759 18424 9760
rect 5441 9618 5507 9621
rect 7833 9618 7899 9621
rect 5441 9616 7899 9618
rect 5441 9560 5446 9616
rect 5502 9560 7838 9616
rect 7894 9560 7899 9616
rect 5441 9558 7899 9560
rect 5441 9555 5507 9558
rect 7833 9555 7899 9558
rect 10961 9618 11027 9621
rect 18505 9618 18571 9621
rect 10961 9616 18571 9618
rect 10961 9560 10966 9616
rect 11022 9560 18510 9616
rect 18566 9560 18571 9616
rect 10961 9558 18571 9560
rect 10961 9555 11027 9558
rect 18505 9555 18571 9558
rect 4981 9482 5047 9485
rect 4846 9480 5047 9482
rect 4846 9424 4986 9480
rect 5042 9424 5047 9480
rect 4846 9422 5047 9424
rect 0 9392 480 9422
rect 4061 9419 4127 9422
rect 4981 9419 5047 9422
rect 13353 9482 13419 9485
rect 22320 9482 22800 9512
rect 13353 9480 22800 9482
rect 13353 9424 13358 9480
rect 13414 9424 22800 9480
rect 13353 9422 22800 9424
rect 13353 9419 13419 9422
rect 22320 9392 22800 9422
rect 7808 9280 8128 9281
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 9215 8128 9216
rect 14672 9280 14992 9281
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 9215 14992 9216
rect 0 9074 480 9104
rect 8569 9074 8635 9077
rect 0 9014 4538 9074
rect 0 8984 480 9014
rect 4478 8938 4538 9014
rect 5030 9072 8635 9074
rect 5030 9016 8574 9072
rect 8630 9016 8635 9072
rect 5030 9014 8635 9016
rect 5030 8938 5090 9014
rect 8569 9011 8635 9014
rect 18505 9074 18571 9077
rect 22320 9074 22800 9104
rect 18505 9072 22800 9074
rect 18505 9016 18510 9072
rect 18566 9016 22800 9072
rect 18505 9014 22800 9016
rect 18505 9011 18571 9014
rect 22320 8984 22800 9014
rect 4478 8878 5090 8938
rect 6177 8938 6243 8941
rect 10358 8938 10364 8940
rect 6177 8936 10364 8938
rect 6177 8880 6182 8936
rect 6238 8880 10364 8936
rect 6177 8878 10364 8880
rect 6177 8875 6243 8878
rect 10358 8876 10364 8878
rect 10428 8938 10434 8940
rect 12709 8938 12775 8941
rect 10428 8936 12775 8938
rect 10428 8880 12714 8936
rect 12770 8880 12775 8936
rect 10428 8878 12775 8880
rect 10428 8876 10434 8878
rect 12709 8875 12775 8878
rect 4376 8736 4696 8737
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 8671 4696 8672
rect 11240 8736 11560 8737
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 8671 11560 8672
rect 18104 8736 18424 8737
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 8671 18424 8672
rect 12065 8666 12131 8669
rect 16665 8666 16731 8669
rect 12065 8664 16731 8666
rect 12065 8608 12070 8664
rect 12126 8608 16670 8664
rect 16726 8608 16731 8664
rect 12065 8606 16731 8608
rect 12065 8603 12131 8606
rect 16665 8603 16731 8606
rect 0 8530 480 8560
rect 4061 8530 4127 8533
rect 0 8528 4127 8530
rect 0 8472 4066 8528
rect 4122 8472 4127 8528
rect 0 8470 4127 8472
rect 0 8440 480 8470
rect 4061 8467 4127 8470
rect 6637 8530 6703 8533
rect 9857 8530 9923 8533
rect 6637 8528 9923 8530
rect 6637 8472 6642 8528
rect 6698 8472 9862 8528
rect 9918 8472 9923 8528
rect 6637 8470 9923 8472
rect 6637 8467 6703 8470
rect 9857 8467 9923 8470
rect 10685 8530 10751 8533
rect 12433 8530 12499 8533
rect 15929 8530 15995 8533
rect 10685 8528 12499 8530
rect 10685 8472 10690 8528
rect 10746 8472 12438 8528
rect 12494 8472 12499 8528
rect 10685 8470 12499 8472
rect 10685 8467 10751 8470
rect 12433 8467 12499 8470
rect 14230 8528 15995 8530
rect 14230 8472 15934 8528
rect 15990 8472 15995 8528
rect 14230 8470 15995 8472
rect 6545 8394 6611 8397
rect 11145 8394 11211 8397
rect 6545 8392 11211 8394
rect 6545 8336 6550 8392
rect 6606 8336 11150 8392
rect 11206 8336 11211 8392
rect 6545 8334 11211 8336
rect 6545 8331 6611 8334
rect 11145 8331 11211 8334
rect 11605 8394 11671 8397
rect 12157 8394 12223 8397
rect 14230 8394 14290 8470
rect 15929 8467 15995 8470
rect 17953 8530 18019 8533
rect 22320 8530 22800 8560
rect 17953 8528 22800 8530
rect 17953 8472 17958 8528
rect 18014 8472 22800 8528
rect 17953 8470 22800 8472
rect 17953 8467 18019 8470
rect 22320 8440 22800 8470
rect 11605 8392 14290 8394
rect 11605 8336 11610 8392
rect 11666 8336 12162 8392
rect 12218 8336 14290 8392
rect 11605 8334 14290 8336
rect 14549 8394 14615 8397
rect 17125 8394 17191 8397
rect 14549 8392 17191 8394
rect 14549 8336 14554 8392
rect 14610 8336 17130 8392
rect 17186 8336 17191 8392
rect 14549 8334 17191 8336
rect 11605 8331 11671 8334
rect 12157 8331 12223 8334
rect 14549 8331 14615 8334
rect 17125 8331 17191 8334
rect 5533 8258 5599 8261
rect 5809 8258 5875 8261
rect 7557 8258 7623 8261
rect 5533 8256 7623 8258
rect 5533 8200 5538 8256
rect 5594 8200 5814 8256
rect 5870 8200 7562 8256
rect 7618 8200 7623 8256
rect 5533 8198 7623 8200
rect 5533 8195 5599 8198
rect 5809 8195 5875 8198
rect 7557 8195 7623 8198
rect 7808 8192 8128 8193
rect 0 8122 480 8152
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 8127 8128 8128
rect 14672 8192 14992 8193
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 8127 14992 8128
rect 7557 8122 7623 8125
rect 0 8120 7623 8122
rect 0 8064 7562 8120
rect 7618 8064 7623 8120
rect 0 8062 7623 8064
rect 0 8032 480 8062
rect 7557 8059 7623 8062
rect 9673 8122 9739 8125
rect 12249 8122 12315 8125
rect 9673 8120 12315 8122
rect 9673 8064 9678 8120
rect 9734 8064 12254 8120
rect 12310 8064 12315 8120
rect 9673 8062 12315 8064
rect 9673 8059 9739 8062
rect 12249 8059 12315 8062
rect 19241 8122 19307 8125
rect 22320 8122 22800 8152
rect 19241 8120 22800 8122
rect 19241 8064 19246 8120
rect 19302 8064 22800 8120
rect 19241 8062 22800 8064
rect 19241 8059 19307 8062
rect 22320 8032 22800 8062
rect 1945 7986 2011 7989
rect 3509 7986 3575 7989
rect 1945 7984 3575 7986
rect 1945 7928 1950 7984
rect 2006 7928 3514 7984
rect 3570 7928 3575 7984
rect 1945 7926 3575 7928
rect 1945 7923 2011 7926
rect 3509 7923 3575 7926
rect 3969 7986 4035 7989
rect 7373 7986 7439 7989
rect 9305 7986 9371 7989
rect 3969 7984 9371 7986
rect 3969 7928 3974 7984
rect 4030 7928 7378 7984
rect 7434 7928 9310 7984
rect 9366 7928 9371 7984
rect 3969 7926 9371 7928
rect 3969 7923 4035 7926
rect 7373 7923 7439 7926
rect 9305 7923 9371 7926
rect 12801 7986 12867 7989
rect 16297 7986 16363 7989
rect 12801 7984 16363 7986
rect 12801 7928 12806 7984
rect 12862 7928 16302 7984
rect 16358 7928 16363 7984
rect 12801 7926 16363 7928
rect 12801 7923 12867 7926
rect 16297 7923 16363 7926
rect 2957 7850 3023 7853
rect 6545 7850 6611 7853
rect 2957 7848 6611 7850
rect 2957 7792 2962 7848
rect 3018 7792 6550 7848
rect 6606 7792 6611 7848
rect 2957 7790 6611 7792
rect 2957 7787 3023 7790
rect 6545 7787 6611 7790
rect 14273 7850 14339 7853
rect 14549 7850 14615 7853
rect 19149 7850 19215 7853
rect 14273 7848 19215 7850
rect 14273 7792 14278 7848
rect 14334 7792 14554 7848
rect 14610 7792 19154 7848
rect 19210 7792 19215 7848
rect 14273 7790 19215 7792
rect 14273 7787 14339 7790
rect 14549 7787 14615 7790
rect 19149 7787 19215 7790
rect 12709 7714 12775 7717
rect 14641 7714 14707 7717
rect 12709 7712 14707 7714
rect 12709 7656 12714 7712
rect 12770 7656 14646 7712
rect 14702 7656 14707 7712
rect 12709 7654 14707 7656
rect 12709 7651 12775 7654
rect 14641 7651 14707 7654
rect 4376 7648 4696 7649
rect 0 7578 480 7608
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 7583 4696 7584
rect 11240 7648 11560 7649
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 7583 11560 7584
rect 18104 7648 18424 7649
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 7583 18424 7584
rect 3969 7578 4035 7581
rect 0 7576 4035 7578
rect 0 7520 3974 7576
rect 4030 7520 4035 7576
rect 0 7518 4035 7520
rect 0 7488 480 7518
rect 3969 7515 4035 7518
rect 11973 7578 12039 7581
rect 15469 7578 15535 7581
rect 11973 7576 15535 7578
rect 11973 7520 11978 7576
rect 12034 7520 15474 7576
rect 15530 7520 15535 7576
rect 11973 7518 15535 7520
rect 11973 7515 12039 7518
rect 15469 7515 15535 7518
rect 18781 7578 18847 7581
rect 22320 7578 22800 7608
rect 18781 7576 22800 7578
rect 18781 7520 18786 7576
rect 18842 7520 22800 7576
rect 18781 7518 22800 7520
rect 18781 7515 18847 7518
rect 22320 7488 22800 7518
rect 9765 7442 9831 7445
rect 15561 7442 15627 7445
rect 9765 7440 15627 7442
rect 9765 7384 9770 7440
rect 9826 7384 15566 7440
rect 15622 7384 15627 7440
rect 9765 7382 15627 7384
rect 9765 7379 9831 7382
rect 15561 7379 15627 7382
rect 0 7170 480 7200
rect 3785 7170 3851 7173
rect 0 7168 3851 7170
rect 0 7112 3790 7168
rect 3846 7112 3851 7168
rect 0 7110 3851 7112
rect 0 7080 480 7110
rect 3785 7107 3851 7110
rect 10593 7170 10659 7173
rect 13353 7170 13419 7173
rect 10593 7168 13419 7170
rect 10593 7112 10598 7168
rect 10654 7112 13358 7168
rect 13414 7112 13419 7168
rect 10593 7110 13419 7112
rect 10593 7107 10659 7110
rect 13353 7107 13419 7110
rect 17769 7170 17835 7173
rect 22320 7170 22800 7200
rect 17769 7168 22800 7170
rect 17769 7112 17774 7168
rect 17830 7112 22800 7168
rect 17769 7110 22800 7112
rect 17769 7107 17835 7110
rect 7808 7104 8128 7105
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 7039 8128 7040
rect 14672 7104 14992 7105
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 22320 7080 22800 7110
rect 14672 7039 14992 7040
rect 10869 6898 10935 6901
rect 16389 6898 16455 6901
rect 10869 6896 16455 6898
rect 10869 6840 10874 6896
rect 10930 6840 16394 6896
rect 16450 6840 16455 6896
rect 10869 6838 16455 6840
rect 10869 6835 10935 6838
rect 16389 6835 16455 6838
rect 0 6762 480 6792
rect 9673 6762 9739 6765
rect 0 6760 9739 6762
rect 0 6704 9678 6760
rect 9734 6704 9739 6760
rect 0 6702 9739 6704
rect 0 6672 480 6702
rect 9673 6699 9739 6702
rect 10133 6762 10199 6765
rect 12249 6762 12315 6765
rect 10133 6760 12315 6762
rect 10133 6704 10138 6760
rect 10194 6704 12254 6760
rect 12310 6704 12315 6760
rect 10133 6702 12315 6704
rect 10133 6699 10199 6702
rect 12249 6699 12315 6702
rect 12709 6762 12775 6765
rect 22320 6762 22800 6792
rect 12709 6760 22800 6762
rect 12709 6704 12714 6760
rect 12770 6704 22800 6760
rect 12709 6702 22800 6704
rect 12709 6699 12775 6702
rect 22320 6672 22800 6702
rect 4376 6560 4696 6561
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 6495 4696 6496
rect 11240 6560 11560 6561
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 6495 11560 6496
rect 18104 6560 18424 6561
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 6495 18424 6496
rect 9765 6354 9831 6357
rect 10501 6354 10567 6357
rect 13169 6354 13235 6357
rect 9765 6352 13235 6354
rect 9765 6296 9770 6352
rect 9826 6296 10506 6352
rect 10562 6296 13174 6352
rect 13230 6296 13235 6352
rect 9765 6294 13235 6296
rect 9765 6291 9831 6294
rect 10501 6291 10567 6294
rect 13169 6291 13235 6294
rect 13537 6354 13603 6357
rect 19057 6354 19123 6357
rect 13537 6352 19123 6354
rect 13537 6296 13542 6352
rect 13598 6296 19062 6352
rect 19118 6296 19123 6352
rect 13537 6294 19123 6296
rect 13537 6291 13603 6294
rect 19057 6291 19123 6294
rect 0 6218 480 6248
rect 3969 6218 4035 6221
rect 0 6216 4035 6218
rect 0 6160 3974 6216
rect 4030 6160 4035 6216
rect 0 6158 4035 6160
rect 0 6128 480 6158
rect 3969 6155 4035 6158
rect 6177 6218 6243 6221
rect 9489 6218 9555 6221
rect 12617 6218 12683 6221
rect 6177 6216 12683 6218
rect 6177 6160 6182 6216
rect 6238 6160 9494 6216
rect 9550 6160 12622 6216
rect 12678 6160 12683 6216
rect 6177 6158 12683 6160
rect 6177 6155 6243 6158
rect 9489 6155 9555 6158
rect 12617 6155 12683 6158
rect 18137 6218 18203 6221
rect 22320 6218 22800 6248
rect 18137 6216 22800 6218
rect 18137 6160 18142 6216
rect 18198 6160 22800 6216
rect 18137 6158 22800 6160
rect 18137 6155 18203 6158
rect 22320 6128 22800 6158
rect 10869 6082 10935 6085
rect 11053 6082 11119 6085
rect 10869 6080 11119 6082
rect 10869 6024 10874 6080
rect 10930 6024 11058 6080
rect 11114 6024 11119 6080
rect 10869 6022 11119 6024
rect 10869 6019 10935 6022
rect 11053 6019 11119 6022
rect 11237 6082 11303 6085
rect 13445 6082 13511 6085
rect 11237 6080 13511 6082
rect 11237 6024 11242 6080
rect 11298 6024 13450 6080
rect 13506 6024 13511 6080
rect 11237 6022 13511 6024
rect 11237 6019 11303 6022
rect 13445 6019 13511 6022
rect 7808 6016 8128 6017
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 5951 8128 5952
rect 14672 6016 14992 6017
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 5951 14992 5952
rect 12065 5946 12131 5949
rect 13813 5946 13879 5949
rect 12065 5944 13879 5946
rect 12065 5888 12070 5944
rect 12126 5888 13818 5944
rect 13874 5888 13879 5944
rect 12065 5886 13879 5888
rect 12065 5883 12131 5886
rect 13813 5883 13879 5886
rect 0 5810 480 5840
rect 3969 5810 4035 5813
rect 0 5808 4035 5810
rect 0 5752 3974 5808
rect 4030 5752 4035 5808
rect 0 5750 4035 5752
rect 0 5720 480 5750
rect 3969 5747 4035 5750
rect 10869 5810 10935 5813
rect 13077 5810 13143 5813
rect 10869 5808 13143 5810
rect 10869 5752 10874 5808
rect 10930 5752 13082 5808
rect 13138 5752 13143 5808
rect 10869 5750 13143 5752
rect 10869 5747 10935 5750
rect 13077 5747 13143 5750
rect 14181 5810 14247 5813
rect 22320 5810 22800 5840
rect 14181 5808 22800 5810
rect 14181 5752 14186 5808
rect 14242 5752 22800 5808
rect 14181 5750 22800 5752
rect 14181 5747 14247 5750
rect 22320 5720 22800 5750
rect 11881 5674 11947 5677
rect 12985 5674 13051 5677
rect 11881 5672 13051 5674
rect 11881 5616 11886 5672
rect 11942 5616 12990 5672
rect 13046 5616 13051 5672
rect 11881 5614 13051 5616
rect 11881 5611 11947 5614
rect 12985 5611 13051 5614
rect 12157 5538 12223 5541
rect 13997 5538 14063 5541
rect 12157 5536 14063 5538
rect 12157 5480 12162 5536
rect 12218 5480 14002 5536
rect 14058 5480 14063 5536
rect 12157 5478 14063 5480
rect 12157 5475 12223 5478
rect 13997 5475 14063 5478
rect 4376 5472 4696 5473
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 5407 4696 5408
rect 11240 5472 11560 5473
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 5407 11560 5408
rect 18104 5472 18424 5473
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 5407 18424 5408
rect 0 5266 480 5296
rect 4061 5266 4127 5269
rect 0 5264 4127 5266
rect 0 5208 4066 5264
rect 4122 5208 4127 5264
rect 0 5206 4127 5208
rect 0 5176 480 5206
rect 4061 5203 4127 5206
rect 4981 5266 5047 5269
rect 8845 5266 8911 5269
rect 9581 5266 9647 5269
rect 4981 5264 9647 5266
rect 4981 5208 4986 5264
rect 5042 5208 8850 5264
rect 8906 5208 9586 5264
rect 9642 5208 9647 5264
rect 4981 5206 9647 5208
rect 4981 5203 5047 5206
rect 8845 5203 8911 5206
rect 9581 5203 9647 5206
rect 17953 5266 18019 5269
rect 22320 5266 22800 5296
rect 17953 5264 22800 5266
rect 17953 5208 17958 5264
rect 18014 5208 22800 5264
rect 17953 5206 22800 5208
rect 17953 5203 18019 5206
rect 22320 5176 22800 5206
rect 2865 5130 2931 5133
rect 10041 5130 10107 5133
rect 12065 5130 12131 5133
rect 2865 5128 12131 5130
rect 2865 5072 2870 5128
rect 2926 5072 10046 5128
rect 10102 5072 12070 5128
rect 12126 5072 12131 5128
rect 2865 5070 12131 5072
rect 2865 5067 2931 5070
rect 10041 5067 10107 5070
rect 12065 5067 12131 5070
rect 9581 4994 9647 4997
rect 14181 4994 14247 4997
rect 9581 4992 14247 4994
rect 9581 4936 9586 4992
rect 9642 4936 14186 4992
rect 14242 4936 14247 4992
rect 9581 4934 14247 4936
rect 9581 4931 9647 4934
rect 14181 4931 14247 4934
rect 7808 4928 8128 4929
rect 0 4858 480 4888
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 4863 8128 4864
rect 14672 4928 14992 4929
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 4863 14992 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4768 480 4798
rect 3969 4795 4035 4798
rect 15193 4858 15259 4861
rect 22320 4858 22800 4888
rect 15193 4856 22800 4858
rect 15193 4800 15198 4856
rect 15254 4800 22800 4856
rect 15193 4798 22800 4800
rect 15193 4795 15259 4798
rect 22320 4768 22800 4798
rect 4376 4384 4696 4385
rect 0 4314 480 4344
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 4319 4696 4320
rect 11240 4384 11560 4385
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 11240 4319 11560 4320
rect 18104 4384 18424 4385
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 4319 18424 4320
rect 4061 4314 4127 4317
rect 0 4312 4127 4314
rect 0 4256 4066 4312
rect 4122 4256 4127 4312
rect 0 4254 4127 4256
rect 0 4224 480 4254
rect 4061 4251 4127 4254
rect 12525 4314 12591 4317
rect 13813 4314 13879 4317
rect 12525 4312 13879 4314
rect 12525 4256 12530 4312
rect 12586 4256 13818 4312
rect 13874 4256 13879 4312
rect 12525 4254 13879 4256
rect 12525 4251 12591 4254
rect 13813 4251 13879 4254
rect 20713 4314 20779 4317
rect 22320 4314 22800 4344
rect 20713 4312 22800 4314
rect 20713 4256 20718 4312
rect 20774 4256 22800 4312
rect 20713 4254 22800 4256
rect 20713 4251 20779 4254
rect 22320 4224 22800 4254
rect 7373 4178 7439 4181
rect 12433 4178 12499 4181
rect 7373 4176 12499 4178
rect 7373 4120 7378 4176
rect 7434 4120 12438 4176
rect 12494 4120 12499 4176
rect 7373 4118 12499 4120
rect 7373 4115 7439 4118
rect 12433 4115 12499 4118
rect 6177 4042 6243 4045
rect 10409 4042 10475 4045
rect 6177 4040 10475 4042
rect 6177 3984 6182 4040
rect 6238 3984 10414 4040
rect 10470 3984 10475 4040
rect 6177 3982 10475 3984
rect 6177 3979 6243 3982
rect 10409 3979 10475 3982
rect 11329 4042 11395 4045
rect 14089 4042 14155 4045
rect 11329 4040 14155 4042
rect 11329 3984 11334 4040
rect 11390 3984 14094 4040
rect 14150 3984 14155 4040
rect 11329 3982 14155 3984
rect 11329 3979 11395 3982
rect 14089 3979 14155 3982
rect 0 3906 480 3936
rect 7557 3906 7623 3909
rect 0 3904 7623 3906
rect 0 3848 7562 3904
rect 7618 3848 7623 3904
rect 0 3846 7623 3848
rect 0 3816 480 3846
rect 7557 3843 7623 3846
rect 8569 3906 8635 3909
rect 11697 3906 11763 3909
rect 8569 3904 11763 3906
rect 8569 3848 8574 3904
rect 8630 3848 11702 3904
rect 11758 3848 11763 3904
rect 8569 3846 11763 3848
rect 8569 3843 8635 3846
rect 11697 3843 11763 3846
rect 19241 3906 19307 3909
rect 22320 3906 22800 3936
rect 19241 3904 22800 3906
rect 19241 3848 19246 3904
rect 19302 3848 22800 3904
rect 19241 3846 22800 3848
rect 19241 3843 19307 3846
rect 7808 3840 8128 3841
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 3775 8128 3776
rect 14672 3840 14992 3841
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 22320 3816 22800 3846
rect 14672 3775 14992 3776
rect 8385 3770 8451 3773
rect 10409 3772 10475 3773
rect 10358 3770 10364 3772
rect 8385 3768 9552 3770
rect 8385 3712 8390 3768
rect 8446 3736 9552 3768
rect 8446 3712 9690 3736
rect 8385 3710 9690 3712
rect 10318 3710 10364 3770
rect 10428 3768 10475 3772
rect 10470 3712 10475 3768
rect 8385 3707 8451 3710
rect 9492 3676 9690 3710
rect 10358 3708 10364 3710
rect 10428 3708 10475 3712
rect 10409 3707 10475 3708
rect 11881 3770 11947 3773
rect 13537 3770 13603 3773
rect 11881 3768 13603 3770
rect 11881 3712 11886 3768
rect 11942 3712 13542 3768
rect 13598 3712 13603 3768
rect 11881 3710 13603 3712
rect 11881 3707 11947 3710
rect 13537 3707 13603 3710
rect 9630 3634 9690 3676
rect 13905 3634 13971 3637
rect 9630 3632 13971 3634
rect 9630 3576 13910 3632
rect 13966 3576 13971 3632
rect 9630 3574 13971 3576
rect 13905 3571 13971 3574
rect 18229 3634 18295 3637
rect 20069 3634 20135 3637
rect 18229 3632 20135 3634
rect 18229 3576 18234 3632
rect 18290 3576 20074 3632
rect 20130 3576 20135 3632
rect 18229 3574 20135 3576
rect 18229 3571 18295 3574
rect 20069 3571 20135 3574
rect 0 3498 480 3528
rect 3877 3498 3943 3501
rect 0 3496 3943 3498
rect 0 3440 3882 3496
rect 3938 3440 3943 3496
rect 0 3438 3943 3440
rect 0 3408 480 3438
rect 3877 3435 3943 3438
rect 10317 3498 10383 3501
rect 10869 3498 10935 3501
rect 10317 3496 10935 3498
rect 10317 3440 10322 3496
rect 10378 3440 10874 3496
rect 10930 3440 10935 3496
rect 10317 3438 10935 3440
rect 10317 3435 10383 3438
rect 10869 3435 10935 3438
rect 18137 3498 18203 3501
rect 22320 3498 22800 3528
rect 18137 3496 22800 3498
rect 18137 3440 18142 3496
rect 18198 3440 22800 3496
rect 18137 3438 22800 3440
rect 18137 3435 18203 3438
rect 22320 3408 22800 3438
rect 4376 3296 4696 3297
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 3231 4696 3232
rect 11240 3296 11560 3297
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 3231 11560 3232
rect 18104 3296 18424 3297
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 3231 18424 3232
rect 3141 3090 3207 3093
rect 8569 3090 8635 3093
rect 3141 3088 8635 3090
rect 3141 3032 3146 3088
rect 3202 3032 8574 3088
rect 8630 3032 8635 3088
rect 3141 3030 8635 3032
rect 3141 3027 3207 3030
rect 8569 3027 8635 3030
rect 0 2954 480 2984
rect 4245 2954 4311 2957
rect 0 2952 4311 2954
rect 0 2896 4250 2952
rect 4306 2896 4311 2952
rect 0 2894 4311 2896
rect 0 2864 480 2894
rect 4245 2891 4311 2894
rect 6913 2954 6979 2957
rect 8293 2954 8359 2957
rect 9029 2954 9095 2957
rect 6913 2952 9095 2954
rect 6913 2896 6918 2952
rect 6974 2896 8298 2952
rect 8354 2896 9034 2952
rect 9090 2896 9095 2952
rect 6913 2894 9095 2896
rect 6913 2891 6979 2894
rect 8293 2891 8359 2894
rect 9029 2891 9095 2894
rect 10961 2954 11027 2957
rect 20437 2954 20503 2957
rect 22320 2954 22800 2984
rect 10961 2952 20503 2954
rect 10961 2896 10966 2952
rect 11022 2896 20442 2952
rect 20498 2896 20503 2952
rect 10961 2894 20503 2896
rect 10961 2891 11027 2894
rect 20437 2891 20503 2894
rect 20670 2894 22800 2954
rect 3325 2818 3391 2821
rect 6177 2818 6243 2821
rect 3325 2816 6243 2818
rect 3325 2760 3330 2816
rect 3386 2760 6182 2816
rect 6238 2760 6243 2816
rect 3325 2758 6243 2760
rect 3325 2755 3391 2758
rect 6177 2755 6243 2758
rect 17585 2818 17651 2821
rect 17953 2818 18019 2821
rect 17585 2816 18019 2818
rect 17585 2760 17590 2816
rect 17646 2760 17958 2816
rect 18014 2760 18019 2816
rect 17585 2758 18019 2760
rect 17585 2755 17651 2758
rect 17953 2755 18019 2758
rect 18505 2818 18571 2821
rect 18781 2818 18847 2821
rect 18505 2816 18847 2818
rect 18505 2760 18510 2816
rect 18566 2760 18786 2816
rect 18842 2760 18847 2816
rect 18505 2758 18847 2760
rect 18505 2755 18571 2758
rect 18781 2755 18847 2758
rect 19149 2818 19215 2821
rect 20670 2818 20730 2894
rect 22320 2864 22800 2894
rect 19149 2816 20730 2818
rect 19149 2760 19154 2816
rect 19210 2760 20730 2816
rect 19149 2758 20730 2760
rect 19149 2755 19215 2758
rect 7808 2752 8128 2753
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2687 8128 2688
rect 14672 2752 14992 2753
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2687 14992 2688
rect 17585 2682 17651 2685
rect 18229 2682 18295 2685
rect 20805 2682 20871 2685
rect 17585 2680 18154 2682
rect 17585 2624 17590 2680
rect 17646 2624 18154 2680
rect 17585 2622 18154 2624
rect 17585 2619 17651 2622
rect 0 2546 480 2576
rect 2313 2546 2379 2549
rect 0 2544 2379 2546
rect 0 2488 2318 2544
rect 2374 2488 2379 2544
rect 0 2486 2379 2488
rect 18094 2546 18154 2622
rect 18229 2680 20871 2682
rect 18229 2624 18234 2680
rect 18290 2624 20810 2680
rect 20866 2624 20871 2680
rect 18229 2622 20871 2624
rect 18229 2619 18295 2622
rect 20805 2619 20871 2622
rect 22320 2546 22800 2576
rect 18094 2486 22800 2546
rect 0 2456 480 2486
rect 2313 2483 2379 2486
rect 22320 2456 22800 2486
rect 4376 2208 4696 2209
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2143 4696 2144
rect 11240 2208 11560 2209
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2143 11560 2144
rect 18104 2208 18424 2209
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2143 18424 2144
rect 0 2002 480 2032
rect 3969 2002 4035 2005
rect 0 2000 4035 2002
rect 0 1944 3974 2000
rect 4030 1944 4035 2000
rect 0 1942 4035 1944
rect 0 1912 480 1942
rect 3969 1939 4035 1942
rect 19241 2002 19307 2005
rect 22320 2002 22800 2032
rect 19241 2000 22800 2002
rect 19241 1944 19246 2000
rect 19302 1944 22800 2000
rect 19241 1942 22800 1944
rect 19241 1939 19307 1942
rect 22320 1912 22800 1942
rect 0 1594 480 1624
rect 2497 1594 2563 1597
rect 0 1592 2563 1594
rect 0 1536 2502 1592
rect 2558 1536 2563 1592
rect 0 1534 2563 1536
rect 0 1504 480 1534
rect 2497 1531 2563 1534
rect 20805 1594 20871 1597
rect 22320 1594 22800 1624
rect 20805 1592 22800 1594
rect 20805 1536 20810 1592
rect 20866 1536 22800 1592
rect 20805 1534 22800 1536
rect 20805 1531 20871 1534
rect 22320 1504 22800 1534
rect 0 1050 480 1080
rect 4061 1050 4127 1053
rect 0 1048 4127 1050
rect 0 992 4066 1048
rect 4122 992 4127 1048
rect 0 990 4127 992
rect 0 960 480 990
rect 4061 987 4127 990
rect 20529 1050 20595 1053
rect 22320 1050 22800 1080
rect 20529 1048 22800 1050
rect 20529 992 20534 1048
rect 20590 992 22800 1048
rect 20529 990 22800 992
rect 20529 987 20595 990
rect 22320 960 22800 990
rect 0 642 480 672
rect 3969 642 4035 645
rect 0 640 4035 642
rect 0 584 3974 640
rect 4030 584 4035 640
rect 0 582 4035 584
rect 0 552 480 582
rect 3969 579 4035 582
rect 20897 642 20963 645
rect 22320 642 22800 672
rect 20897 640 22800 642
rect 20897 584 20902 640
rect 20958 584 22800 640
rect 20897 582 22800 584
rect 20897 579 20963 582
rect 22320 552 22800 582
rect 0 234 480 264
rect 5625 234 5691 237
rect 0 232 5691 234
rect 0 176 5630 232
rect 5686 176 5691 232
rect 0 174 5691 176
rect 0 144 480 174
rect 5625 171 5691 174
rect 18781 234 18847 237
rect 22320 234 22800 264
rect 18781 232 22800 234
rect 18781 176 18786 232
rect 18842 176 22800 232
rect 18781 174 22800 176
rect 18781 171 18847 174
rect 22320 144 22800 174
<< via3 >>
rect 7816 20156 7880 20160
rect 7816 20100 7820 20156
rect 7820 20100 7876 20156
rect 7876 20100 7880 20156
rect 7816 20096 7880 20100
rect 7896 20156 7960 20160
rect 7896 20100 7900 20156
rect 7900 20100 7956 20156
rect 7956 20100 7960 20156
rect 7896 20096 7960 20100
rect 7976 20156 8040 20160
rect 7976 20100 7980 20156
rect 7980 20100 8036 20156
rect 8036 20100 8040 20156
rect 7976 20096 8040 20100
rect 8056 20156 8120 20160
rect 8056 20100 8060 20156
rect 8060 20100 8116 20156
rect 8116 20100 8120 20156
rect 8056 20096 8120 20100
rect 14680 20156 14744 20160
rect 14680 20100 14684 20156
rect 14684 20100 14740 20156
rect 14740 20100 14744 20156
rect 14680 20096 14744 20100
rect 14760 20156 14824 20160
rect 14760 20100 14764 20156
rect 14764 20100 14820 20156
rect 14820 20100 14824 20156
rect 14760 20096 14824 20100
rect 14840 20156 14904 20160
rect 14840 20100 14844 20156
rect 14844 20100 14900 20156
rect 14900 20100 14904 20156
rect 14840 20096 14904 20100
rect 14920 20156 14984 20160
rect 14920 20100 14924 20156
rect 14924 20100 14980 20156
rect 14980 20100 14984 20156
rect 14920 20096 14984 20100
rect 4384 19612 4448 19616
rect 4384 19556 4388 19612
rect 4388 19556 4444 19612
rect 4444 19556 4448 19612
rect 4384 19552 4448 19556
rect 4464 19612 4528 19616
rect 4464 19556 4468 19612
rect 4468 19556 4524 19612
rect 4524 19556 4528 19612
rect 4464 19552 4528 19556
rect 4544 19612 4608 19616
rect 4544 19556 4548 19612
rect 4548 19556 4604 19612
rect 4604 19556 4608 19612
rect 4544 19552 4608 19556
rect 4624 19612 4688 19616
rect 4624 19556 4628 19612
rect 4628 19556 4684 19612
rect 4684 19556 4688 19612
rect 4624 19552 4688 19556
rect 11248 19612 11312 19616
rect 11248 19556 11252 19612
rect 11252 19556 11308 19612
rect 11308 19556 11312 19612
rect 11248 19552 11312 19556
rect 11328 19612 11392 19616
rect 11328 19556 11332 19612
rect 11332 19556 11388 19612
rect 11388 19556 11392 19612
rect 11328 19552 11392 19556
rect 11408 19612 11472 19616
rect 11408 19556 11412 19612
rect 11412 19556 11468 19612
rect 11468 19556 11472 19612
rect 11408 19552 11472 19556
rect 11488 19612 11552 19616
rect 11488 19556 11492 19612
rect 11492 19556 11548 19612
rect 11548 19556 11552 19612
rect 11488 19552 11552 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 18272 19612 18336 19616
rect 18272 19556 18276 19612
rect 18276 19556 18332 19612
rect 18332 19556 18336 19612
rect 18272 19552 18336 19556
rect 18352 19612 18416 19616
rect 18352 19556 18356 19612
rect 18356 19556 18412 19612
rect 18412 19556 18416 19612
rect 18352 19552 18416 19556
rect 7816 19068 7880 19072
rect 7816 19012 7820 19068
rect 7820 19012 7876 19068
rect 7876 19012 7880 19068
rect 7816 19008 7880 19012
rect 7896 19068 7960 19072
rect 7896 19012 7900 19068
rect 7900 19012 7956 19068
rect 7956 19012 7960 19068
rect 7896 19008 7960 19012
rect 7976 19068 8040 19072
rect 7976 19012 7980 19068
rect 7980 19012 8036 19068
rect 8036 19012 8040 19068
rect 7976 19008 8040 19012
rect 8056 19068 8120 19072
rect 8056 19012 8060 19068
rect 8060 19012 8116 19068
rect 8116 19012 8120 19068
rect 8056 19008 8120 19012
rect 14680 19068 14744 19072
rect 14680 19012 14684 19068
rect 14684 19012 14740 19068
rect 14740 19012 14744 19068
rect 14680 19008 14744 19012
rect 14760 19068 14824 19072
rect 14760 19012 14764 19068
rect 14764 19012 14820 19068
rect 14820 19012 14824 19068
rect 14760 19008 14824 19012
rect 14840 19068 14904 19072
rect 14840 19012 14844 19068
rect 14844 19012 14900 19068
rect 14900 19012 14904 19068
rect 14840 19008 14904 19012
rect 14920 19068 14984 19072
rect 14920 19012 14924 19068
rect 14924 19012 14980 19068
rect 14980 19012 14984 19068
rect 14920 19008 14984 19012
rect 4384 18524 4448 18528
rect 4384 18468 4388 18524
rect 4388 18468 4444 18524
rect 4444 18468 4448 18524
rect 4384 18464 4448 18468
rect 4464 18524 4528 18528
rect 4464 18468 4468 18524
rect 4468 18468 4524 18524
rect 4524 18468 4528 18524
rect 4464 18464 4528 18468
rect 4544 18524 4608 18528
rect 4544 18468 4548 18524
rect 4548 18468 4604 18524
rect 4604 18468 4608 18524
rect 4544 18464 4608 18468
rect 4624 18524 4688 18528
rect 4624 18468 4628 18524
rect 4628 18468 4684 18524
rect 4684 18468 4688 18524
rect 4624 18464 4688 18468
rect 11248 18524 11312 18528
rect 11248 18468 11252 18524
rect 11252 18468 11308 18524
rect 11308 18468 11312 18524
rect 11248 18464 11312 18468
rect 11328 18524 11392 18528
rect 11328 18468 11332 18524
rect 11332 18468 11388 18524
rect 11388 18468 11392 18524
rect 11328 18464 11392 18468
rect 11408 18524 11472 18528
rect 11408 18468 11412 18524
rect 11412 18468 11468 18524
rect 11468 18468 11472 18524
rect 11408 18464 11472 18468
rect 11488 18524 11552 18528
rect 11488 18468 11492 18524
rect 11492 18468 11548 18524
rect 11548 18468 11552 18524
rect 11488 18464 11552 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 18272 18524 18336 18528
rect 18272 18468 18276 18524
rect 18276 18468 18332 18524
rect 18332 18468 18336 18524
rect 18272 18464 18336 18468
rect 18352 18524 18416 18528
rect 18352 18468 18356 18524
rect 18356 18468 18412 18524
rect 18412 18468 18416 18524
rect 18352 18464 18416 18468
rect 19932 18260 19996 18324
rect 7816 17980 7880 17984
rect 7816 17924 7820 17980
rect 7820 17924 7876 17980
rect 7876 17924 7880 17980
rect 7816 17920 7880 17924
rect 7896 17980 7960 17984
rect 7896 17924 7900 17980
rect 7900 17924 7956 17980
rect 7956 17924 7960 17980
rect 7896 17920 7960 17924
rect 7976 17980 8040 17984
rect 7976 17924 7980 17980
rect 7980 17924 8036 17980
rect 8036 17924 8040 17980
rect 7976 17920 8040 17924
rect 8056 17980 8120 17984
rect 8056 17924 8060 17980
rect 8060 17924 8116 17980
rect 8116 17924 8120 17980
rect 8056 17920 8120 17924
rect 14680 17980 14744 17984
rect 14680 17924 14684 17980
rect 14684 17924 14740 17980
rect 14740 17924 14744 17980
rect 14680 17920 14744 17924
rect 14760 17980 14824 17984
rect 14760 17924 14764 17980
rect 14764 17924 14820 17980
rect 14820 17924 14824 17980
rect 14760 17920 14824 17924
rect 14840 17980 14904 17984
rect 14840 17924 14844 17980
rect 14844 17924 14900 17980
rect 14900 17924 14904 17980
rect 14840 17920 14904 17924
rect 14920 17980 14984 17984
rect 14920 17924 14924 17980
rect 14924 17924 14980 17980
rect 14980 17924 14984 17980
rect 14920 17920 14984 17924
rect 4384 17436 4448 17440
rect 4384 17380 4388 17436
rect 4388 17380 4444 17436
rect 4444 17380 4448 17436
rect 4384 17376 4448 17380
rect 4464 17436 4528 17440
rect 4464 17380 4468 17436
rect 4468 17380 4524 17436
rect 4524 17380 4528 17436
rect 4464 17376 4528 17380
rect 4544 17436 4608 17440
rect 4544 17380 4548 17436
rect 4548 17380 4604 17436
rect 4604 17380 4608 17436
rect 4544 17376 4608 17380
rect 4624 17436 4688 17440
rect 4624 17380 4628 17436
rect 4628 17380 4684 17436
rect 4684 17380 4688 17436
rect 4624 17376 4688 17380
rect 11248 17436 11312 17440
rect 11248 17380 11252 17436
rect 11252 17380 11308 17436
rect 11308 17380 11312 17436
rect 11248 17376 11312 17380
rect 11328 17436 11392 17440
rect 11328 17380 11332 17436
rect 11332 17380 11388 17436
rect 11388 17380 11392 17436
rect 11328 17376 11392 17380
rect 11408 17436 11472 17440
rect 11408 17380 11412 17436
rect 11412 17380 11468 17436
rect 11468 17380 11472 17436
rect 11408 17376 11472 17380
rect 11488 17436 11552 17440
rect 11488 17380 11492 17436
rect 11492 17380 11548 17436
rect 11548 17380 11552 17436
rect 11488 17376 11552 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 18272 17436 18336 17440
rect 18272 17380 18276 17436
rect 18276 17380 18332 17436
rect 18332 17380 18336 17436
rect 18272 17376 18336 17380
rect 18352 17436 18416 17440
rect 18352 17380 18356 17436
rect 18356 17380 18412 17436
rect 18412 17380 18416 17436
rect 18352 17376 18416 17380
rect 7816 16892 7880 16896
rect 7816 16836 7820 16892
rect 7820 16836 7876 16892
rect 7876 16836 7880 16892
rect 7816 16832 7880 16836
rect 7896 16892 7960 16896
rect 7896 16836 7900 16892
rect 7900 16836 7956 16892
rect 7956 16836 7960 16892
rect 7896 16832 7960 16836
rect 7976 16892 8040 16896
rect 7976 16836 7980 16892
rect 7980 16836 8036 16892
rect 8036 16836 8040 16892
rect 7976 16832 8040 16836
rect 8056 16892 8120 16896
rect 8056 16836 8060 16892
rect 8060 16836 8116 16892
rect 8116 16836 8120 16892
rect 8056 16832 8120 16836
rect 14680 16892 14744 16896
rect 14680 16836 14684 16892
rect 14684 16836 14740 16892
rect 14740 16836 14744 16892
rect 14680 16832 14744 16836
rect 14760 16892 14824 16896
rect 14760 16836 14764 16892
rect 14764 16836 14820 16892
rect 14820 16836 14824 16892
rect 14760 16832 14824 16836
rect 14840 16892 14904 16896
rect 14840 16836 14844 16892
rect 14844 16836 14900 16892
rect 14900 16836 14904 16892
rect 14840 16832 14904 16836
rect 14920 16892 14984 16896
rect 14920 16836 14924 16892
rect 14924 16836 14980 16892
rect 14980 16836 14984 16892
rect 14920 16832 14984 16836
rect 4384 16348 4448 16352
rect 4384 16292 4388 16348
rect 4388 16292 4444 16348
rect 4444 16292 4448 16348
rect 4384 16288 4448 16292
rect 4464 16348 4528 16352
rect 4464 16292 4468 16348
rect 4468 16292 4524 16348
rect 4524 16292 4528 16348
rect 4464 16288 4528 16292
rect 4544 16348 4608 16352
rect 4544 16292 4548 16348
rect 4548 16292 4604 16348
rect 4604 16292 4608 16348
rect 4544 16288 4608 16292
rect 4624 16348 4688 16352
rect 4624 16292 4628 16348
rect 4628 16292 4684 16348
rect 4684 16292 4688 16348
rect 4624 16288 4688 16292
rect 11248 16348 11312 16352
rect 11248 16292 11252 16348
rect 11252 16292 11308 16348
rect 11308 16292 11312 16348
rect 11248 16288 11312 16292
rect 11328 16348 11392 16352
rect 11328 16292 11332 16348
rect 11332 16292 11388 16348
rect 11388 16292 11392 16348
rect 11328 16288 11392 16292
rect 11408 16348 11472 16352
rect 11408 16292 11412 16348
rect 11412 16292 11468 16348
rect 11468 16292 11472 16348
rect 11408 16288 11472 16292
rect 11488 16348 11552 16352
rect 11488 16292 11492 16348
rect 11492 16292 11548 16348
rect 11548 16292 11552 16348
rect 11488 16288 11552 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 18272 16348 18336 16352
rect 18272 16292 18276 16348
rect 18276 16292 18332 16348
rect 18332 16292 18336 16348
rect 18272 16288 18336 16292
rect 18352 16348 18416 16352
rect 18352 16292 18356 16348
rect 18356 16292 18412 16348
rect 18412 16292 18416 16348
rect 18352 16288 18416 16292
rect 7816 15804 7880 15808
rect 7816 15748 7820 15804
rect 7820 15748 7876 15804
rect 7876 15748 7880 15804
rect 7816 15744 7880 15748
rect 7896 15804 7960 15808
rect 7896 15748 7900 15804
rect 7900 15748 7956 15804
rect 7956 15748 7960 15804
rect 7896 15744 7960 15748
rect 7976 15804 8040 15808
rect 7976 15748 7980 15804
rect 7980 15748 8036 15804
rect 8036 15748 8040 15804
rect 7976 15744 8040 15748
rect 8056 15804 8120 15808
rect 8056 15748 8060 15804
rect 8060 15748 8116 15804
rect 8116 15748 8120 15804
rect 8056 15744 8120 15748
rect 14680 15804 14744 15808
rect 14680 15748 14684 15804
rect 14684 15748 14740 15804
rect 14740 15748 14744 15804
rect 14680 15744 14744 15748
rect 14760 15804 14824 15808
rect 14760 15748 14764 15804
rect 14764 15748 14820 15804
rect 14820 15748 14824 15804
rect 14760 15744 14824 15748
rect 14840 15804 14904 15808
rect 14840 15748 14844 15804
rect 14844 15748 14900 15804
rect 14900 15748 14904 15804
rect 14840 15744 14904 15748
rect 14920 15804 14984 15808
rect 14920 15748 14924 15804
rect 14924 15748 14980 15804
rect 14980 15748 14984 15804
rect 14920 15744 14984 15748
rect 4384 15260 4448 15264
rect 4384 15204 4388 15260
rect 4388 15204 4444 15260
rect 4444 15204 4448 15260
rect 4384 15200 4448 15204
rect 4464 15260 4528 15264
rect 4464 15204 4468 15260
rect 4468 15204 4524 15260
rect 4524 15204 4528 15260
rect 4464 15200 4528 15204
rect 4544 15260 4608 15264
rect 4544 15204 4548 15260
rect 4548 15204 4604 15260
rect 4604 15204 4608 15260
rect 4544 15200 4608 15204
rect 4624 15260 4688 15264
rect 4624 15204 4628 15260
rect 4628 15204 4684 15260
rect 4684 15204 4688 15260
rect 4624 15200 4688 15204
rect 11248 15260 11312 15264
rect 11248 15204 11252 15260
rect 11252 15204 11308 15260
rect 11308 15204 11312 15260
rect 11248 15200 11312 15204
rect 11328 15260 11392 15264
rect 11328 15204 11332 15260
rect 11332 15204 11388 15260
rect 11388 15204 11392 15260
rect 11328 15200 11392 15204
rect 11408 15260 11472 15264
rect 11408 15204 11412 15260
rect 11412 15204 11468 15260
rect 11468 15204 11472 15260
rect 11408 15200 11472 15204
rect 11488 15260 11552 15264
rect 11488 15204 11492 15260
rect 11492 15204 11548 15260
rect 11548 15204 11552 15260
rect 11488 15200 11552 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 18272 15260 18336 15264
rect 18272 15204 18276 15260
rect 18276 15204 18332 15260
rect 18332 15204 18336 15260
rect 18272 15200 18336 15204
rect 18352 15260 18416 15264
rect 18352 15204 18356 15260
rect 18356 15204 18412 15260
rect 18412 15204 18416 15260
rect 18352 15200 18416 15204
rect 7816 14716 7880 14720
rect 7816 14660 7820 14716
rect 7820 14660 7876 14716
rect 7876 14660 7880 14716
rect 7816 14656 7880 14660
rect 7896 14716 7960 14720
rect 7896 14660 7900 14716
rect 7900 14660 7956 14716
rect 7956 14660 7960 14716
rect 7896 14656 7960 14660
rect 7976 14716 8040 14720
rect 7976 14660 7980 14716
rect 7980 14660 8036 14716
rect 8036 14660 8040 14716
rect 7976 14656 8040 14660
rect 8056 14716 8120 14720
rect 8056 14660 8060 14716
rect 8060 14660 8116 14716
rect 8116 14660 8120 14716
rect 8056 14656 8120 14660
rect 14680 14716 14744 14720
rect 14680 14660 14684 14716
rect 14684 14660 14740 14716
rect 14740 14660 14744 14716
rect 14680 14656 14744 14660
rect 14760 14716 14824 14720
rect 14760 14660 14764 14716
rect 14764 14660 14820 14716
rect 14820 14660 14824 14716
rect 14760 14656 14824 14660
rect 14840 14716 14904 14720
rect 14840 14660 14844 14716
rect 14844 14660 14900 14716
rect 14900 14660 14904 14716
rect 14840 14656 14904 14660
rect 14920 14716 14984 14720
rect 14920 14660 14924 14716
rect 14924 14660 14980 14716
rect 14980 14660 14984 14716
rect 14920 14656 14984 14660
rect 4384 14172 4448 14176
rect 4384 14116 4388 14172
rect 4388 14116 4444 14172
rect 4444 14116 4448 14172
rect 4384 14112 4448 14116
rect 4464 14172 4528 14176
rect 4464 14116 4468 14172
rect 4468 14116 4524 14172
rect 4524 14116 4528 14172
rect 4464 14112 4528 14116
rect 4544 14172 4608 14176
rect 4544 14116 4548 14172
rect 4548 14116 4604 14172
rect 4604 14116 4608 14172
rect 4544 14112 4608 14116
rect 4624 14172 4688 14176
rect 4624 14116 4628 14172
rect 4628 14116 4684 14172
rect 4684 14116 4688 14172
rect 4624 14112 4688 14116
rect 11248 14172 11312 14176
rect 11248 14116 11252 14172
rect 11252 14116 11308 14172
rect 11308 14116 11312 14172
rect 11248 14112 11312 14116
rect 11328 14172 11392 14176
rect 11328 14116 11332 14172
rect 11332 14116 11388 14172
rect 11388 14116 11392 14172
rect 11328 14112 11392 14116
rect 11408 14172 11472 14176
rect 11408 14116 11412 14172
rect 11412 14116 11468 14172
rect 11468 14116 11472 14172
rect 11408 14112 11472 14116
rect 11488 14172 11552 14176
rect 11488 14116 11492 14172
rect 11492 14116 11548 14172
rect 11548 14116 11552 14172
rect 11488 14112 11552 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 18272 14172 18336 14176
rect 18272 14116 18276 14172
rect 18276 14116 18332 14172
rect 18332 14116 18336 14172
rect 18272 14112 18336 14116
rect 18352 14172 18416 14176
rect 18352 14116 18356 14172
rect 18356 14116 18412 14172
rect 18412 14116 18416 14172
rect 18352 14112 18416 14116
rect 7816 13628 7880 13632
rect 7816 13572 7820 13628
rect 7820 13572 7876 13628
rect 7876 13572 7880 13628
rect 7816 13568 7880 13572
rect 7896 13628 7960 13632
rect 7896 13572 7900 13628
rect 7900 13572 7956 13628
rect 7956 13572 7960 13628
rect 7896 13568 7960 13572
rect 7976 13628 8040 13632
rect 7976 13572 7980 13628
rect 7980 13572 8036 13628
rect 8036 13572 8040 13628
rect 7976 13568 8040 13572
rect 8056 13628 8120 13632
rect 8056 13572 8060 13628
rect 8060 13572 8116 13628
rect 8116 13572 8120 13628
rect 8056 13568 8120 13572
rect 14680 13628 14744 13632
rect 14680 13572 14684 13628
rect 14684 13572 14740 13628
rect 14740 13572 14744 13628
rect 14680 13568 14744 13572
rect 14760 13628 14824 13632
rect 14760 13572 14764 13628
rect 14764 13572 14820 13628
rect 14820 13572 14824 13628
rect 14760 13568 14824 13572
rect 14840 13628 14904 13632
rect 14840 13572 14844 13628
rect 14844 13572 14900 13628
rect 14900 13572 14904 13628
rect 14840 13568 14904 13572
rect 14920 13628 14984 13632
rect 14920 13572 14924 13628
rect 14924 13572 14980 13628
rect 14980 13572 14984 13628
rect 14920 13568 14984 13572
rect 4384 13084 4448 13088
rect 4384 13028 4388 13084
rect 4388 13028 4444 13084
rect 4444 13028 4448 13084
rect 4384 13024 4448 13028
rect 4464 13084 4528 13088
rect 4464 13028 4468 13084
rect 4468 13028 4524 13084
rect 4524 13028 4528 13084
rect 4464 13024 4528 13028
rect 4544 13084 4608 13088
rect 4544 13028 4548 13084
rect 4548 13028 4604 13084
rect 4604 13028 4608 13084
rect 4544 13024 4608 13028
rect 4624 13084 4688 13088
rect 4624 13028 4628 13084
rect 4628 13028 4684 13084
rect 4684 13028 4688 13084
rect 4624 13024 4688 13028
rect 11248 13084 11312 13088
rect 11248 13028 11252 13084
rect 11252 13028 11308 13084
rect 11308 13028 11312 13084
rect 11248 13024 11312 13028
rect 11328 13084 11392 13088
rect 11328 13028 11332 13084
rect 11332 13028 11388 13084
rect 11388 13028 11392 13084
rect 11328 13024 11392 13028
rect 11408 13084 11472 13088
rect 11408 13028 11412 13084
rect 11412 13028 11468 13084
rect 11468 13028 11472 13084
rect 11408 13024 11472 13028
rect 11488 13084 11552 13088
rect 11488 13028 11492 13084
rect 11492 13028 11548 13084
rect 11548 13028 11552 13084
rect 11488 13024 11552 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 18272 13084 18336 13088
rect 18272 13028 18276 13084
rect 18276 13028 18332 13084
rect 18332 13028 18336 13084
rect 18272 13024 18336 13028
rect 18352 13084 18416 13088
rect 18352 13028 18356 13084
rect 18356 13028 18412 13084
rect 18412 13028 18416 13084
rect 18352 13024 18416 13028
rect 7816 12540 7880 12544
rect 7816 12484 7820 12540
rect 7820 12484 7876 12540
rect 7876 12484 7880 12540
rect 7816 12480 7880 12484
rect 7896 12540 7960 12544
rect 7896 12484 7900 12540
rect 7900 12484 7956 12540
rect 7956 12484 7960 12540
rect 7896 12480 7960 12484
rect 7976 12540 8040 12544
rect 7976 12484 7980 12540
rect 7980 12484 8036 12540
rect 8036 12484 8040 12540
rect 7976 12480 8040 12484
rect 8056 12540 8120 12544
rect 8056 12484 8060 12540
rect 8060 12484 8116 12540
rect 8116 12484 8120 12540
rect 8056 12480 8120 12484
rect 14680 12540 14744 12544
rect 14680 12484 14684 12540
rect 14684 12484 14740 12540
rect 14740 12484 14744 12540
rect 14680 12480 14744 12484
rect 14760 12540 14824 12544
rect 14760 12484 14764 12540
rect 14764 12484 14820 12540
rect 14820 12484 14824 12540
rect 14760 12480 14824 12484
rect 14840 12540 14904 12544
rect 14840 12484 14844 12540
rect 14844 12484 14900 12540
rect 14900 12484 14904 12540
rect 14840 12480 14904 12484
rect 14920 12540 14984 12544
rect 14920 12484 14924 12540
rect 14924 12484 14980 12540
rect 14980 12484 14984 12540
rect 14920 12480 14984 12484
rect 4384 11996 4448 12000
rect 4384 11940 4388 11996
rect 4388 11940 4444 11996
rect 4444 11940 4448 11996
rect 4384 11936 4448 11940
rect 4464 11996 4528 12000
rect 4464 11940 4468 11996
rect 4468 11940 4524 11996
rect 4524 11940 4528 11996
rect 4464 11936 4528 11940
rect 4544 11996 4608 12000
rect 4544 11940 4548 11996
rect 4548 11940 4604 11996
rect 4604 11940 4608 11996
rect 4544 11936 4608 11940
rect 4624 11996 4688 12000
rect 4624 11940 4628 11996
rect 4628 11940 4684 11996
rect 4684 11940 4688 11996
rect 4624 11936 4688 11940
rect 11248 11996 11312 12000
rect 11248 11940 11252 11996
rect 11252 11940 11308 11996
rect 11308 11940 11312 11996
rect 11248 11936 11312 11940
rect 11328 11996 11392 12000
rect 11328 11940 11332 11996
rect 11332 11940 11388 11996
rect 11388 11940 11392 11996
rect 11328 11936 11392 11940
rect 11408 11996 11472 12000
rect 11408 11940 11412 11996
rect 11412 11940 11468 11996
rect 11468 11940 11472 11996
rect 11408 11936 11472 11940
rect 11488 11996 11552 12000
rect 11488 11940 11492 11996
rect 11492 11940 11548 11996
rect 11548 11940 11552 11996
rect 11488 11936 11552 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 18272 11996 18336 12000
rect 18272 11940 18276 11996
rect 18276 11940 18332 11996
rect 18332 11940 18336 11996
rect 18272 11936 18336 11940
rect 18352 11996 18416 12000
rect 18352 11940 18356 11996
rect 18356 11940 18412 11996
rect 18412 11940 18416 11996
rect 18352 11936 18416 11940
rect 7816 11452 7880 11456
rect 7816 11396 7820 11452
rect 7820 11396 7876 11452
rect 7876 11396 7880 11452
rect 7816 11392 7880 11396
rect 7896 11452 7960 11456
rect 7896 11396 7900 11452
rect 7900 11396 7956 11452
rect 7956 11396 7960 11452
rect 7896 11392 7960 11396
rect 7976 11452 8040 11456
rect 7976 11396 7980 11452
rect 7980 11396 8036 11452
rect 8036 11396 8040 11452
rect 7976 11392 8040 11396
rect 8056 11452 8120 11456
rect 8056 11396 8060 11452
rect 8060 11396 8116 11452
rect 8116 11396 8120 11452
rect 8056 11392 8120 11396
rect 14680 11452 14744 11456
rect 14680 11396 14684 11452
rect 14684 11396 14740 11452
rect 14740 11396 14744 11452
rect 14680 11392 14744 11396
rect 14760 11452 14824 11456
rect 14760 11396 14764 11452
rect 14764 11396 14820 11452
rect 14820 11396 14824 11452
rect 14760 11392 14824 11396
rect 14840 11452 14904 11456
rect 14840 11396 14844 11452
rect 14844 11396 14900 11452
rect 14900 11396 14904 11452
rect 14840 11392 14904 11396
rect 14920 11452 14984 11456
rect 14920 11396 14924 11452
rect 14924 11396 14980 11452
rect 14980 11396 14984 11452
rect 14920 11392 14984 11396
rect 4384 10908 4448 10912
rect 4384 10852 4388 10908
rect 4388 10852 4444 10908
rect 4444 10852 4448 10908
rect 4384 10848 4448 10852
rect 4464 10908 4528 10912
rect 4464 10852 4468 10908
rect 4468 10852 4524 10908
rect 4524 10852 4528 10908
rect 4464 10848 4528 10852
rect 4544 10908 4608 10912
rect 4544 10852 4548 10908
rect 4548 10852 4604 10908
rect 4604 10852 4608 10908
rect 4544 10848 4608 10852
rect 4624 10908 4688 10912
rect 4624 10852 4628 10908
rect 4628 10852 4684 10908
rect 4684 10852 4688 10908
rect 4624 10848 4688 10852
rect 11248 10908 11312 10912
rect 11248 10852 11252 10908
rect 11252 10852 11308 10908
rect 11308 10852 11312 10908
rect 11248 10848 11312 10852
rect 11328 10908 11392 10912
rect 11328 10852 11332 10908
rect 11332 10852 11388 10908
rect 11388 10852 11392 10908
rect 11328 10848 11392 10852
rect 11408 10908 11472 10912
rect 11408 10852 11412 10908
rect 11412 10852 11468 10908
rect 11468 10852 11472 10908
rect 11408 10848 11472 10852
rect 11488 10908 11552 10912
rect 11488 10852 11492 10908
rect 11492 10852 11548 10908
rect 11548 10852 11552 10908
rect 11488 10848 11552 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 18272 10908 18336 10912
rect 18272 10852 18276 10908
rect 18276 10852 18332 10908
rect 18332 10852 18336 10908
rect 18272 10848 18336 10852
rect 18352 10908 18416 10912
rect 18352 10852 18356 10908
rect 18356 10852 18412 10908
rect 18412 10852 18416 10908
rect 18352 10848 18416 10852
rect 19932 10644 19996 10708
rect 7816 10364 7880 10368
rect 7816 10308 7820 10364
rect 7820 10308 7876 10364
rect 7876 10308 7880 10364
rect 7816 10304 7880 10308
rect 7896 10364 7960 10368
rect 7896 10308 7900 10364
rect 7900 10308 7956 10364
rect 7956 10308 7960 10364
rect 7896 10304 7960 10308
rect 7976 10364 8040 10368
rect 7976 10308 7980 10364
rect 7980 10308 8036 10364
rect 8036 10308 8040 10364
rect 7976 10304 8040 10308
rect 8056 10364 8120 10368
rect 8056 10308 8060 10364
rect 8060 10308 8116 10364
rect 8116 10308 8120 10364
rect 8056 10304 8120 10308
rect 14680 10364 14744 10368
rect 14680 10308 14684 10364
rect 14684 10308 14740 10364
rect 14740 10308 14744 10364
rect 14680 10304 14744 10308
rect 14760 10364 14824 10368
rect 14760 10308 14764 10364
rect 14764 10308 14820 10364
rect 14820 10308 14824 10364
rect 14760 10304 14824 10308
rect 14840 10364 14904 10368
rect 14840 10308 14844 10364
rect 14844 10308 14900 10364
rect 14900 10308 14904 10364
rect 14840 10304 14904 10308
rect 14920 10364 14984 10368
rect 14920 10308 14924 10364
rect 14924 10308 14980 10364
rect 14980 10308 14984 10364
rect 14920 10304 14984 10308
rect 4384 9820 4448 9824
rect 4384 9764 4388 9820
rect 4388 9764 4444 9820
rect 4444 9764 4448 9820
rect 4384 9760 4448 9764
rect 4464 9820 4528 9824
rect 4464 9764 4468 9820
rect 4468 9764 4524 9820
rect 4524 9764 4528 9820
rect 4464 9760 4528 9764
rect 4544 9820 4608 9824
rect 4544 9764 4548 9820
rect 4548 9764 4604 9820
rect 4604 9764 4608 9820
rect 4544 9760 4608 9764
rect 4624 9820 4688 9824
rect 4624 9764 4628 9820
rect 4628 9764 4684 9820
rect 4684 9764 4688 9820
rect 4624 9760 4688 9764
rect 11248 9820 11312 9824
rect 11248 9764 11252 9820
rect 11252 9764 11308 9820
rect 11308 9764 11312 9820
rect 11248 9760 11312 9764
rect 11328 9820 11392 9824
rect 11328 9764 11332 9820
rect 11332 9764 11388 9820
rect 11388 9764 11392 9820
rect 11328 9760 11392 9764
rect 11408 9820 11472 9824
rect 11408 9764 11412 9820
rect 11412 9764 11468 9820
rect 11468 9764 11472 9820
rect 11408 9760 11472 9764
rect 11488 9820 11552 9824
rect 11488 9764 11492 9820
rect 11492 9764 11548 9820
rect 11548 9764 11552 9820
rect 11488 9760 11552 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 18272 9820 18336 9824
rect 18272 9764 18276 9820
rect 18276 9764 18332 9820
rect 18332 9764 18336 9820
rect 18272 9760 18336 9764
rect 18352 9820 18416 9824
rect 18352 9764 18356 9820
rect 18356 9764 18412 9820
rect 18412 9764 18416 9820
rect 18352 9760 18416 9764
rect 7816 9276 7880 9280
rect 7816 9220 7820 9276
rect 7820 9220 7876 9276
rect 7876 9220 7880 9276
rect 7816 9216 7880 9220
rect 7896 9276 7960 9280
rect 7896 9220 7900 9276
rect 7900 9220 7956 9276
rect 7956 9220 7960 9276
rect 7896 9216 7960 9220
rect 7976 9276 8040 9280
rect 7976 9220 7980 9276
rect 7980 9220 8036 9276
rect 8036 9220 8040 9276
rect 7976 9216 8040 9220
rect 8056 9276 8120 9280
rect 8056 9220 8060 9276
rect 8060 9220 8116 9276
rect 8116 9220 8120 9276
rect 8056 9216 8120 9220
rect 14680 9276 14744 9280
rect 14680 9220 14684 9276
rect 14684 9220 14740 9276
rect 14740 9220 14744 9276
rect 14680 9216 14744 9220
rect 14760 9276 14824 9280
rect 14760 9220 14764 9276
rect 14764 9220 14820 9276
rect 14820 9220 14824 9276
rect 14760 9216 14824 9220
rect 14840 9276 14904 9280
rect 14840 9220 14844 9276
rect 14844 9220 14900 9276
rect 14900 9220 14904 9276
rect 14840 9216 14904 9220
rect 14920 9276 14984 9280
rect 14920 9220 14924 9276
rect 14924 9220 14980 9276
rect 14980 9220 14984 9276
rect 14920 9216 14984 9220
rect 10364 8876 10428 8940
rect 4384 8732 4448 8736
rect 4384 8676 4388 8732
rect 4388 8676 4444 8732
rect 4444 8676 4448 8732
rect 4384 8672 4448 8676
rect 4464 8732 4528 8736
rect 4464 8676 4468 8732
rect 4468 8676 4524 8732
rect 4524 8676 4528 8732
rect 4464 8672 4528 8676
rect 4544 8732 4608 8736
rect 4544 8676 4548 8732
rect 4548 8676 4604 8732
rect 4604 8676 4608 8732
rect 4544 8672 4608 8676
rect 4624 8732 4688 8736
rect 4624 8676 4628 8732
rect 4628 8676 4684 8732
rect 4684 8676 4688 8732
rect 4624 8672 4688 8676
rect 11248 8732 11312 8736
rect 11248 8676 11252 8732
rect 11252 8676 11308 8732
rect 11308 8676 11312 8732
rect 11248 8672 11312 8676
rect 11328 8732 11392 8736
rect 11328 8676 11332 8732
rect 11332 8676 11388 8732
rect 11388 8676 11392 8732
rect 11328 8672 11392 8676
rect 11408 8732 11472 8736
rect 11408 8676 11412 8732
rect 11412 8676 11468 8732
rect 11468 8676 11472 8732
rect 11408 8672 11472 8676
rect 11488 8732 11552 8736
rect 11488 8676 11492 8732
rect 11492 8676 11548 8732
rect 11548 8676 11552 8732
rect 11488 8672 11552 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 18272 8732 18336 8736
rect 18272 8676 18276 8732
rect 18276 8676 18332 8732
rect 18332 8676 18336 8732
rect 18272 8672 18336 8676
rect 18352 8732 18416 8736
rect 18352 8676 18356 8732
rect 18356 8676 18412 8732
rect 18412 8676 18416 8732
rect 18352 8672 18416 8676
rect 7816 8188 7880 8192
rect 7816 8132 7820 8188
rect 7820 8132 7876 8188
rect 7876 8132 7880 8188
rect 7816 8128 7880 8132
rect 7896 8188 7960 8192
rect 7896 8132 7900 8188
rect 7900 8132 7956 8188
rect 7956 8132 7960 8188
rect 7896 8128 7960 8132
rect 7976 8188 8040 8192
rect 7976 8132 7980 8188
rect 7980 8132 8036 8188
rect 8036 8132 8040 8188
rect 7976 8128 8040 8132
rect 8056 8188 8120 8192
rect 8056 8132 8060 8188
rect 8060 8132 8116 8188
rect 8116 8132 8120 8188
rect 8056 8128 8120 8132
rect 14680 8188 14744 8192
rect 14680 8132 14684 8188
rect 14684 8132 14740 8188
rect 14740 8132 14744 8188
rect 14680 8128 14744 8132
rect 14760 8188 14824 8192
rect 14760 8132 14764 8188
rect 14764 8132 14820 8188
rect 14820 8132 14824 8188
rect 14760 8128 14824 8132
rect 14840 8188 14904 8192
rect 14840 8132 14844 8188
rect 14844 8132 14900 8188
rect 14900 8132 14904 8188
rect 14840 8128 14904 8132
rect 14920 8188 14984 8192
rect 14920 8132 14924 8188
rect 14924 8132 14980 8188
rect 14980 8132 14984 8188
rect 14920 8128 14984 8132
rect 4384 7644 4448 7648
rect 4384 7588 4388 7644
rect 4388 7588 4444 7644
rect 4444 7588 4448 7644
rect 4384 7584 4448 7588
rect 4464 7644 4528 7648
rect 4464 7588 4468 7644
rect 4468 7588 4524 7644
rect 4524 7588 4528 7644
rect 4464 7584 4528 7588
rect 4544 7644 4608 7648
rect 4544 7588 4548 7644
rect 4548 7588 4604 7644
rect 4604 7588 4608 7644
rect 4544 7584 4608 7588
rect 4624 7644 4688 7648
rect 4624 7588 4628 7644
rect 4628 7588 4684 7644
rect 4684 7588 4688 7644
rect 4624 7584 4688 7588
rect 11248 7644 11312 7648
rect 11248 7588 11252 7644
rect 11252 7588 11308 7644
rect 11308 7588 11312 7644
rect 11248 7584 11312 7588
rect 11328 7644 11392 7648
rect 11328 7588 11332 7644
rect 11332 7588 11388 7644
rect 11388 7588 11392 7644
rect 11328 7584 11392 7588
rect 11408 7644 11472 7648
rect 11408 7588 11412 7644
rect 11412 7588 11468 7644
rect 11468 7588 11472 7644
rect 11408 7584 11472 7588
rect 11488 7644 11552 7648
rect 11488 7588 11492 7644
rect 11492 7588 11548 7644
rect 11548 7588 11552 7644
rect 11488 7584 11552 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 18272 7644 18336 7648
rect 18272 7588 18276 7644
rect 18276 7588 18332 7644
rect 18332 7588 18336 7644
rect 18272 7584 18336 7588
rect 18352 7644 18416 7648
rect 18352 7588 18356 7644
rect 18356 7588 18412 7644
rect 18412 7588 18416 7644
rect 18352 7584 18416 7588
rect 7816 7100 7880 7104
rect 7816 7044 7820 7100
rect 7820 7044 7876 7100
rect 7876 7044 7880 7100
rect 7816 7040 7880 7044
rect 7896 7100 7960 7104
rect 7896 7044 7900 7100
rect 7900 7044 7956 7100
rect 7956 7044 7960 7100
rect 7896 7040 7960 7044
rect 7976 7100 8040 7104
rect 7976 7044 7980 7100
rect 7980 7044 8036 7100
rect 8036 7044 8040 7100
rect 7976 7040 8040 7044
rect 8056 7100 8120 7104
rect 8056 7044 8060 7100
rect 8060 7044 8116 7100
rect 8116 7044 8120 7100
rect 8056 7040 8120 7044
rect 14680 7100 14744 7104
rect 14680 7044 14684 7100
rect 14684 7044 14740 7100
rect 14740 7044 14744 7100
rect 14680 7040 14744 7044
rect 14760 7100 14824 7104
rect 14760 7044 14764 7100
rect 14764 7044 14820 7100
rect 14820 7044 14824 7100
rect 14760 7040 14824 7044
rect 14840 7100 14904 7104
rect 14840 7044 14844 7100
rect 14844 7044 14900 7100
rect 14900 7044 14904 7100
rect 14840 7040 14904 7044
rect 14920 7100 14984 7104
rect 14920 7044 14924 7100
rect 14924 7044 14980 7100
rect 14980 7044 14984 7100
rect 14920 7040 14984 7044
rect 4384 6556 4448 6560
rect 4384 6500 4388 6556
rect 4388 6500 4444 6556
rect 4444 6500 4448 6556
rect 4384 6496 4448 6500
rect 4464 6556 4528 6560
rect 4464 6500 4468 6556
rect 4468 6500 4524 6556
rect 4524 6500 4528 6556
rect 4464 6496 4528 6500
rect 4544 6556 4608 6560
rect 4544 6500 4548 6556
rect 4548 6500 4604 6556
rect 4604 6500 4608 6556
rect 4544 6496 4608 6500
rect 4624 6556 4688 6560
rect 4624 6500 4628 6556
rect 4628 6500 4684 6556
rect 4684 6500 4688 6556
rect 4624 6496 4688 6500
rect 11248 6556 11312 6560
rect 11248 6500 11252 6556
rect 11252 6500 11308 6556
rect 11308 6500 11312 6556
rect 11248 6496 11312 6500
rect 11328 6556 11392 6560
rect 11328 6500 11332 6556
rect 11332 6500 11388 6556
rect 11388 6500 11392 6556
rect 11328 6496 11392 6500
rect 11408 6556 11472 6560
rect 11408 6500 11412 6556
rect 11412 6500 11468 6556
rect 11468 6500 11472 6556
rect 11408 6496 11472 6500
rect 11488 6556 11552 6560
rect 11488 6500 11492 6556
rect 11492 6500 11548 6556
rect 11548 6500 11552 6556
rect 11488 6496 11552 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 18272 6556 18336 6560
rect 18272 6500 18276 6556
rect 18276 6500 18332 6556
rect 18332 6500 18336 6556
rect 18272 6496 18336 6500
rect 18352 6556 18416 6560
rect 18352 6500 18356 6556
rect 18356 6500 18412 6556
rect 18412 6500 18416 6556
rect 18352 6496 18416 6500
rect 7816 6012 7880 6016
rect 7816 5956 7820 6012
rect 7820 5956 7876 6012
rect 7876 5956 7880 6012
rect 7816 5952 7880 5956
rect 7896 6012 7960 6016
rect 7896 5956 7900 6012
rect 7900 5956 7956 6012
rect 7956 5956 7960 6012
rect 7896 5952 7960 5956
rect 7976 6012 8040 6016
rect 7976 5956 7980 6012
rect 7980 5956 8036 6012
rect 8036 5956 8040 6012
rect 7976 5952 8040 5956
rect 8056 6012 8120 6016
rect 8056 5956 8060 6012
rect 8060 5956 8116 6012
rect 8116 5956 8120 6012
rect 8056 5952 8120 5956
rect 14680 6012 14744 6016
rect 14680 5956 14684 6012
rect 14684 5956 14740 6012
rect 14740 5956 14744 6012
rect 14680 5952 14744 5956
rect 14760 6012 14824 6016
rect 14760 5956 14764 6012
rect 14764 5956 14820 6012
rect 14820 5956 14824 6012
rect 14760 5952 14824 5956
rect 14840 6012 14904 6016
rect 14840 5956 14844 6012
rect 14844 5956 14900 6012
rect 14900 5956 14904 6012
rect 14840 5952 14904 5956
rect 14920 6012 14984 6016
rect 14920 5956 14924 6012
rect 14924 5956 14980 6012
rect 14980 5956 14984 6012
rect 14920 5952 14984 5956
rect 4384 5468 4448 5472
rect 4384 5412 4388 5468
rect 4388 5412 4444 5468
rect 4444 5412 4448 5468
rect 4384 5408 4448 5412
rect 4464 5468 4528 5472
rect 4464 5412 4468 5468
rect 4468 5412 4524 5468
rect 4524 5412 4528 5468
rect 4464 5408 4528 5412
rect 4544 5468 4608 5472
rect 4544 5412 4548 5468
rect 4548 5412 4604 5468
rect 4604 5412 4608 5468
rect 4544 5408 4608 5412
rect 4624 5468 4688 5472
rect 4624 5412 4628 5468
rect 4628 5412 4684 5468
rect 4684 5412 4688 5468
rect 4624 5408 4688 5412
rect 11248 5468 11312 5472
rect 11248 5412 11252 5468
rect 11252 5412 11308 5468
rect 11308 5412 11312 5468
rect 11248 5408 11312 5412
rect 11328 5468 11392 5472
rect 11328 5412 11332 5468
rect 11332 5412 11388 5468
rect 11388 5412 11392 5468
rect 11328 5408 11392 5412
rect 11408 5468 11472 5472
rect 11408 5412 11412 5468
rect 11412 5412 11468 5468
rect 11468 5412 11472 5468
rect 11408 5408 11472 5412
rect 11488 5468 11552 5472
rect 11488 5412 11492 5468
rect 11492 5412 11548 5468
rect 11548 5412 11552 5468
rect 11488 5408 11552 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 18272 5468 18336 5472
rect 18272 5412 18276 5468
rect 18276 5412 18332 5468
rect 18332 5412 18336 5468
rect 18272 5408 18336 5412
rect 18352 5468 18416 5472
rect 18352 5412 18356 5468
rect 18356 5412 18412 5468
rect 18412 5412 18416 5468
rect 18352 5408 18416 5412
rect 7816 4924 7880 4928
rect 7816 4868 7820 4924
rect 7820 4868 7876 4924
rect 7876 4868 7880 4924
rect 7816 4864 7880 4868
rect 7896 4924 7960 4928
rect 7896 4868 7900 4924
rect 7900 4868 7956 4924
rect 7956 4868 7960 4924
rect 7896 4864 7960 4868
rect 7976 4924 8040 4928
rect 7976 4868 7980 4924
rect 7980 4868 8036 4924
rect 8036 4868 8040 4924
rect 7976 4864 8040 4868
rect 8056 4924 8120 4928
rect 8056 4868 8060 4924
rect 8060 4868 8116 4924
rect 8116 4868 8120 4924
rect 8056 4864 8120 4868
rect 14680 4924 14744 4928
rect 14680 4868 14684 4924
rect 14684 4868 14740 4924
rect 14740 4868 14744 4924
rect 14680 4864 14744 4868
rect 14760 4924 14824 4928
rect 14760 4868 14764 4924
rect 14764 4868 14820 4924
rect 14820 4868 14824 4924
rect 14760 4864 14824 4868
rect 14840 4924 14904 4928
rect 14840 4868 14844 4924
rect 14844 4868 14900 4924
rect 14900 4868 14904 4924
rect 14840 4864 14904 4868
rect 14920 4924 14984 4928
rect 14920 4868 14924 4924
rect 14924 4868 14980 4924
rect 14980 4868 14984 4924
rect 14920 4864 14984 4868
rect 4384 4380 4448 4384
rect 4384 4324 4388 4380
rect 4388 4324 4444 4380
rect 4444 4324 4448 4380
rect 4384 4320 4448 4324
rect 4464 4380 4528 4384
rect 4464 4324 4468 4380
rect 4468 4324 4524 4380
rect 4524 4324 4528 4380
rect 4464 4320 4528 4324
rect 4544 4380 4608 4384
rect 4544 4324 4548 4380
rect 4548 4324 4604 4380
rect 4604 4324 4608 4380
rect 4544 4320 4608 4324
rect 4624 4380 4688 4384
rect 4624 4324 4628 4380
rect 4628 4324 4684 4380
rect 4684 4324 4688 4380
rect 4624 4320 4688 4324
rect 11248 4380 11312 4384
rect 11248 4324 11252 4380
rect 11252 4324 11308 4380
rect 11308 4324 11312 4380
rect 11248 4320 11312 4324
rect 11328 4380 11392 4384
rect 11328 4324 11332 4380
rect 11332 4324 11388 4380
rect 11388 4324 11392 4380
rect 11328 4320 11392 4324
rect 11408 4380 11472 4384
rect 11408 4324 11412 4380
rect 11412 4324 11468 4380
rect 11468 4324 11472 4380
rect 11408 4320 11472 4324
rect 11488 4380 11552 4384
rect 11488 4324 11492 4380
rect 11492 4324 11548 4380
rect 11548 4324 11552 4380
rect 11488 4320 11552 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 18272 4380 18336 4384
rect 18272 4324 18276 4380
rect 18276 4324 18332 4380
rect 18332 4324 18336 4380
rect 18272 4320 18336 4324
rect 18352 4380 18416 4384
rect 18352 4324 18356 4380
rect 18356 4324 18412 4380
rect 18412 4324 18416 4380
rect 18352 4320 18416 4324
rect 7816 3836 7880 3840
rect 7816 3780 7820 3836
rect 7820 3780 7876 3836
rect 7876 3780 7880 3836
rect 7816 3776 7880 3780
rect 7896 3836 7960 3840
rect 7896 3780 7900 3836
rect 7900 3780 7956 3836
rect 7956 3780 7960 3836
rect 7896 3776 7960 3780
rect 7976 3836 8040 3840
rect 7976 3780 7980 3836
rect 7980 3780 8036 3836
rect 8036 3780 8040 3836
rect 7976 3776 8040 3780
rect 8056 3836 8120 3840
rect 8056 3780 8060 3836
rect 8060 3780 8116 3836
rect 8116 3780 8120 3836
rect 8056 3776 8120 3780
rect 14680 3836 14744 3840
rect 14680 3780 14684 3836
rect 14684 3780 14740 3836
rect 14740 3780 14744 3836
rect 14680 3776 14744 3780
rect 14760 3836 14824 3840
rect 14760 3780 14764 3836
rect 14764 3780 14820 3836
rect 14820 3780 14824 3836
rect 14760 3776 14824 3780
rect 14840 3836 14904 3840
rect 14840 3780 14844 3836
rect 14844 3780 14900 3836
rect 14900 3780 14904 3836
rect 14840 3776 14904 3780
rect 14920 3836 14984 3840
rect 14920 3780 14924 3836
rect 14924 3780 14980 3836
rect 14980 3780 14984 3836
rect 14920 3776 14984 3780
rect 10364 3768 10428 3772
rect 10364 3712 10414 3768
rect 10414 3712 10428 3768
rect 10364 3708 10428 3712
rect 4384 3292 4448 3296
rect 4384 3236 4388 3292
rect 4388 3236 4444 3292
rect 4444 3236 4448 3292
rect 4384 3232 4448 3236
rect 4464 3292 4528 3296
rect 4464 3236 4468 3292
rect 4468 3236 4524 3292
rect 4524 3236 4528 3292
rect 4464 3232 4528 3236
rect 4544 3292 4608 3296
rect 4544 3236 4548 3292
rect 4548 3236 4604 3292
rect 4604 3236 4608 3292
rect 4544 3232 4608 3236
rect 4624 3292 4688 3296
rect 4624 3236 4628 3292
rect 4628 3236 4684 3292
rect 4684 3236 4688 3292
rect 4624 3232 4688 3236
rect 11248 3292 11312 3296
rect 11248 3236 11252 3292
rect 11252 3236 11308 3292
rect 11308 3236 11312 3292
rect 11248 3232 11312 3236
rect 11328 3292 11392 3296
rect 11328 3236 11332 3292
rect 11332 3236 11388 3292
rect 11388 3236 11392 3292
rect 11328 3232 11392 3236
rect 11408 3292 11472 3296
rect 11408 3236 11412 3292
rect 11412 3236 11468 3292
rect 11468 3236 11472 3292
rect 11408 3232 11472 3236
rect 11488 3292 11552 3296
rect 11488 3236 11492 3292
rect 11492 3236 11548 3292
rect 11548 3236 11552 3292
rect 11488 3232 11552 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 18272 3292 18336 3296
rect 18272 3236 18276 3292
rect 18276 3236 18332 3292
rect 18332 3236 18336 3292
rect 18272 3232 18336 3236
rect 18352 3292 18416 3296
rect 18352 3236 18356 3292
rect 18356 3236 18412 3292
rect 18412 3236 18416 3292
rect 18352 3232 18416 3236
rect 7816 2748 7880 2752
rect 7816 2692 7820 2748
rect 7820 2692 7876 2748
rect 7876 2692 7880 2748
rect 7816 2688 7880 2692
rect 7896 2748 7960 2752
rect 7896 2692 7900 2748
rect 7900 2692 7956 2748
rect 7956 2692 7960 2748
rect 7896 2688 7960 2692
rect 7976 2748 8040 2752
rect 7976 2692 7980 2748
rect 7980 2692 8036 2748
rect 8036 2692 8040 2748
rect 7976 2688 8040 2692
rect 8056 2748 8120 2752
rect 8056 2692 8060 2748
rect 8060 2692 8116 2748
rect 8116 2692 8120 2748
rect 8056 2688 8120 2692
rect 14680 2748 14744 2752
rect 14680 2692 14684 2748
rect 14684 2692 14740 2748
rect 14740 2692 14744 2748
rect 14680 2688 14744 2692
rect 14760 2748 14824 2752
rect 14760 2692 14764 2748
rect 14764 2692 14820 2748
rect 14820 2692 14824 2748
rect 14760 2688 14824 2692
rect 14840 2748 14904 2752
rect 14840 2692 14844 2748
rect 14844 2692 14900 2748
rect 14900 2692 14904 2748
rect 14840 2688 14904 2692
rect 14920 2748 14984 2752
rect 14920 2692 14924 2748
rect 14924 2692 14980 2748
rect 14980 2692 14984 2748
rect 14920 2688 14984 2692
rect 4384 2204 4448 2208
rect 4384 2148 4388 2204
rect 4388 2148 4444 2204
rect 4444 2148 4448 2204
rect 4384 2144 4448 2148
rect 4464 2204 4528 2208
rect 4464 2148 4468 2204
rect 4468 2148 4524 2204
rect 4524 2148 4528 2204
rect 4464 2144 4528 2148
rect 4544 2204 4608 2208
rect 4544 2148 4548 2204
rect 4548 2148 4604 2204
rect 4604 2148 4608 2204
rect 4544 2144 4608 2148
rect 4624 2204 4688 2208
rect 4624 2148 4628 2204
rect 4628 2148 4684 2204
rect 4684 2148 4688 2204
rect 4624 2144 4688 2148
rect 11248 2204 11312 2208
rect 11248 2148 11252 2204
rect 11252 2148 11308 2204
rect 11308 2148 11312 2204
rect 11248 2144 11312 2148
rect 11328 2204 11392 2208
rect 11328 2148 11332 2204
rect 11332 2148 11388 2204
rect 11388 2148 11392 2204
rect 11328 2144 11392 2148
rect 11408 2204 11472 2208
rect 11408 2148 11412 2204
rect 11412 2148 11468 2204
rect 11468 2148 11472 2204
rect 11408 2144 11472 2148
rect 11488 2204 11552 2208
rect 11488 2148 11492 2204
rect 11492 2148 11548 2204
rect 11548 2148 11552 2204
rect 11488 2144 11552 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 18272 2204 18336 2208
rect 18272 2148 18276 2204
rect 18276 2148 18332 2204
rect 18332 2148 18336 2204
rect 18272 2144 18336 2148
rect 18352 2204 18416 2208
rect 18352 2148 18356 2204
rect 18356 2148 18412 2204
rect 18412 2148 18416 2204
rect 18352 2144 18416 2148
<< metal4 >>
rect 4376 19616 4696 20176
rect 4376 19552 4384 19616
rect 4448 19552 4464 19616
rect 4528 19552 4544 19616
rect 4608 19552 4624 19616
rect 4688 19552 4696 19616
rect 4376 18528 4696 19552
rect 4376 18464 4384 18528
rect 4448 18464 4464 18528
rect 4528 18464 4544 18528
rect 4608 18464 4624 18528
rect 4688 18464 4696 18528
rect 4376 17440 4696 18464
rect 4376 17376 4384 17440
rect 4448 17376 4464 17440
rect 4528 17376 4544 17440
rect 4608 17376 4624 17440
rect 4688 17376 4696 17440
rect 4376 16352 4696 17376
rect 4376 16288 4384 16352
rect 4448 16288 4464 16352
rect 4528 16288 4544 16352
rect 4608 16288 4624 16352
rect 4688 16288 4696 16352
rect 4376 15264 4696 16288
rect 4376 15200 4384 15264
rect 4448 15200 4464 15264
rect 4528 15200 4544 15264
rect 4608 15200 4624 15264
rect 4688 15200 4696 15264
rect 4376 14176 4696 15200
rect 4376 14112 4384 14176
rect 4448 14112 4464 14176
rect 4528 14112 4544 14176
rect 4608 14112 4624 14176
rect 4688 14112 4696 14176
rect 4376 13088 4696 14112
rect 4376 13024 4384 13088
rect 4448 13024 4464 13088
rect 4528 13024 4544 13088
rect 4608 13024 4624 13088
rect 4688 13024 4696 13088
rect 4376 12000 4696 13024
rect 4376 11936 4384 12000
rect 4448 11936 4464 12000
rect 4528 11936 4544 12000
rect 4608 11936 4624 12000
rect 4688 11936 4696 12000
rect 4376 10912 4696 11936
rect 4376 10848 4384 10912
rect 4448 10848 4464 10912
rect 4528 10848 4544 10912
rect 4608 10848 4624 10912
rect 4688 10848 4696 10912
rect 4376 9824 4696 10848
rect 4376 9760 4384 9824
rect 4448 9760 4464 9824
rect 4528 9760 4544 9824
rect 4608 9760 4624 9824
rect 4688 9760 4696 9824
rect 4376 8736 4696 9760
rect 4376 8672 4384 8736
rect 4448 8672 4464 8736
rect 4528 8672 4544 8736
rect 4608 8672 4624 8736
rect 4688 8672 4696 8736
rect 4376 7648 4696 8672
rect 4376 7584 4384 7648
rect 4448 7584 4464 7648
rect 4528 7584 4544 7648
rect 4608 7584 4624 7648
rect 4688 7584 4696 7648
rect 4376 6560 4696 7584
rect 4376 6496 4384 6560
rect 4448 6496 4464 6560
rect 4528 6496 4544 6560
rect 4608 6496 4624 6560
rect 4688 6496 4696 6560
rect 4376 5472 4696 6496
rect 4376 5408 4384 5472
rect 4448 5408 4464 5472
rect 4528 5408 4544 5472
rect 4608 5408 4624 5472
rect 4688 5408 4696 5472
rect 4376 4384 4696 5408
rect 4376 4320 4384 4384
rect 4448 4320 4464 4384
rect 4528 4320 4544 4384
rect 4608 4320 4624 4384
rect 4688 4320 4696 4384
rect 4376 3296 4696 4320
rect 4376 3232 4384 3296
rect 4448 3232 4464 3296
rect 4528 3232 4544 3296
rect 4608 3232 4624 3296
rect 4688 3232 4696 3296
rect 4376 2208 4696 3232
rect 4376 2144 4384 2208
rect 4448 2144 4464 2208
rect 4528 2144 4544 2208
rect 4608 2144 4624 2208
rect 4688 2144 4696 2208
rect 4376 2128 4696 2144
rect 7808 20160 8128 20176
rect 7808 20096 7816 20160
rect 7880 20096 7896 20160
rect 7960 20096 7976 20160
rect 8040 20096 8056 20160
rect 8120 20096 8128 20160
rect 7808 19072 8128 20096
rect 7808 19008 7816 19072
rect 7880 19008 7896 19072
rect 7960 19008 7976 19072
rect 8040 19008 8056 19072
rect 8120 19008 8128 19072
rect 7808 17984 8128 19008
rect 7808 17920 7816 17984
rect 7880 17920 7896 17984
rect 7960 17920 7976 17984
rect 8040 17920 8056 17984
rect 8120 17920 8128 17984
rect 7808 16896 8128 17920
rect 7808 16832 7816 16896
rect 7880 16832 7896 16896
rect 7960 16832 7976 16896
rect 8040 16832 8056 16896
rect 8120 16832 8128 16896
rect 7808 15808 8128 16832
rect 7808 15744 7816 15808
rect 7880 15744 7896 15808
rect 7960 15744 7976 15808
rect 8040 15744 8056 15808
rect 8120 15744 8128 15808
rect 7808 14720 8128 15744
rect 7808 14656 7816 14720
rect 7880 14656 7896 14720
rect 7960 14656 7976 14720
rect 8040 14656 8056 14720
rect 8120 14656 8128 14720
rect 7808 13632 8128 14656
rect 7808 13568 7816 13632
rect 7880 13568 7896 13632
rect 7960 13568 7976 13632
rect 8040 13568 8056 13632
rect 8120 13568 8128 13632
rect 7808 12544 8128 13568
rect 7808 12480 7816 12544
rect 7880 12480 7896 12544
rect 7960 12480 7976 12544
rect 8040 12480 8056 12544
rect 8120 12480 8128 12544
rect 7808 11456 8128 12480
rect 7808 11392 7816 11456
rect 7880 11392 7896 11456
rect 7960 11392 7976 11456
rect 8040 11392 8056 11456
rect 8120 11392 8128 11456
rect 7808 10368 8128 11392
rect 7808 10304 7816 10368
rect 7880 10304 7896 10368
rect 7960 10304 7976 10368
rect 8040 10304 8056 10368
rect 8120 10304 8128 10368
rect 7808 9280 8128 10304
rect 7808 9216 7816 9280
rect 7880 9216 7896 9280
rect 7960 9216 7976 9280
rect 8040 9216 8056 9280
rect 8120 9216 8128 9280
rect 7808 8192 8128 9216
rect 11240 19616 11560 20176
rect 11240 19552 11248 19616
rect 11312 19552 11328 19616
rect 11392 19552 11408 19616
rect 11472 19552 11488 19616
rect 11552 19552 11560 19616
rect 11240 18528 11560 19552
rect 11240 18464 11248 18528
rect 11312 18464 11328 18528
rect 11392 18464 11408 18528
rect 11472 18464 11488 18528
rect 11552 18464 11560 18528
rect 11240 17440 11560 18464
rect 11240 17376 11248 17440
rect 11312 17376 11328 17440
rect 11392 17376 11408 17440
rect 11472 17376 11488 17440
rect 11552 17376 11560 17440
rect 11240 16352 11560 17376
rect 11240 16288 11248 16352
rect 11312 16288 11328 16352
rect 11392 16288 11408 16352
rect 11472 16288 11488 16352
rect 11552 16288 11560 16352
rect 11240 15264 11560 16288
rect 11240 15200 11248 15264
rect 11312 15200 11328 15264
rect 11392 15200 11408 15264
rect 11472 15200 11488 15264
rect 11552 15200 11560 15264
rect 11240 14176 11560 15200
rect 11240 14112 11248 14176
rect 11312 14112 11328 14176
rect 11392 14112 11408 14176
rect 11472 14112 11488 14176
rect 11552 14112 11560 14176
rect 11240 13088 11560 14112
rect 11240 13024 11248 13088
rect 11312 13024 11328 13088
rect 11392 13024 11408 13088
rect 11472 13024 11488 13088
rect 11552 13024 11560 13088
rect 11240 12000 11560 13024
rect 11240 11936 11248 12000
rect 11312 11936 11328 12000
rect 11392 11936 11408 12000
rect 11472 11936 11488 12000
rect 11552 11936 11560 12000
rect 11240 10912 11560 11936
rect 11240 10848 11248 10912
rect 11312 10848 11328 10912
rect 11392 10848 11408 10912
rect 11472 10848 11488 10912
rect 11552 10848 11560 10912
rect 11240 9824 11560 10848
rect 11240 9760 11248 9824
rect 11312 9760 11328 9824
rect 11392 9760 11408 9824
rect 11472 9760 11488 9824
rect 11552 9760 11560 9824
rect 10363 8940 10429 8941
rect 10363 8876 10364 8940
rect 10428 8876 10429 8940
rect 10363 8875 10429 8876
rect 7808 8128 7816 8192
rect 7880 8128 7896 8192
rect 7960 8128 7976 8192
rect 8040 8128 8056 8192
rect 8120 8128 8128 8192
rect 7808 7104 8128 8128
rect 7808 7040 7816 7104
rect 7880 7040 7896 7104
rect 7960 7040 7976 7104
rect 8040 7040 8056 7104
rect 8120 7040 8128 7104
rect 7808 6016 8128 7040
rect 7808 5952 7816 6016
rect 7880 5952 7896 6016
rect 7960 5952 7976 6016
rect 8040 5952 8056 6016
rect 8120 5952 8128 6016
rect 7808 4928 8128 5952
rect 7808 4864 7816 4928
rect 7880 4864 7896 4928
rect 7960 4864 7976 4928
rect 8040 4864 8056 4928
rect 8120 4864 8128 4928
rect 7808 3840 8128 4864
rect 7808 3776 7816 3840
rect 7880 3776 7896 3840
rect 7960 3776 7976 3840
rect 8040 3776 8056 3840
rect 8120 3776 8128 3840
rect 7808 2752 8128 3776
rect 10366 3773 10426 8875
rect 11240 8736 11560 9760
rect 11240 8672 11248 8736
rect 11312 8672 11328 8736
rect 11392 8672 11408 8736
rect 11472 8672 11488 8736
rect 11552 8672 11560 8736
rect 11240 7648 11560 8672
rect 11240 7584 11248 7648
rect 11312 7584 11328 7648
rect 11392 7584 11408 7648
rect 11472 7584 11488 7648
rect 11552 7584 11560 7648
rect 11240 6560 11560 7584
rect 11240 6496 11248 6560
rect 11312 6496 11328 6560
rect 11392 6496 11408 6560
rect 11472 6496 11488 6560
rect 11552 6496 11560 6560
rect 11240 5472 11560 6496
rect 11240 5408 11248 5472
rect 11312 5408 11328 5472
rect 11392 5408 11408 5472
rect 11472 5408 11488 5472
rect 11552 5408 11560 5472
rect 11240 4384 11560 5408
rect 11240 4320 11248 4384
rect 11312 4320 11328 4384
rect 11392 4320 11408 4384
rect 11472 4320 11488 4384
rect 11552 4320 11560 4384
rect 10363 3772 10429 3773
rect 10363 3708 10364 3772
rect 10428 3708 10429 3772
rect 10363 3707 10429 3708
rect 7808 2688 7816 2752
rect 7880 2688 7896 2752
rect 7960 2688 7976 2752
rect 8040 2688 8056 2752
rect 8120 2688 8128 2752
rect 7808 2128 8128 2688
rect 11240 3296 11560 4320
rect 11240 3232 11248 3296
rect 11312 3232 11328 3296
rect 11392 3232 11408 3296
rect 11472 3232 11488 3296
rect 11552 3232 11560 3296
rect 11240 2208 11560 3232
rect 11240 2144 11248 2208
rect 11312 2144 11328 2208
rect 11392 2144 11408 2208
rect 11472 2144 11488 2208
rect 11552 2144 11560 2208
rect 11240 2128 11560 2144
rect 14672 20160 14992 20176
rect 14672 20096 14680 20160
rect 14744 20096 14760 20160
rect 14824 20096 14840 20160
rect 14904 20096 14920 20160
rect 14984 20096 14992 20160
rect 14672 19072 14992 20096
rect 14672 19008 14680 19072
rect 14744 19008 14760 19072
rect 14824 19008 14840 19072
rect 14904 19008 14920 19072
rect 14984 19008 14992 19072
rect 14672 17984 14992 19008
rect 14672 17920 14680 17984
rect 14744 17920 14760 17984
rect 14824 17920 14840 17984
rect 14904 17920 14920 17984
rect 14984 17920 14992 17984
rect 14672 16896 14992 17920
rect 14672 16832 14680 16896
rect 14744 16832 14760 16896
rect 14824 16832 14840 16896
rect 14904 16832 14920 16896
rect 14984 16832 14992 16896
rect 14672 15808 14992 16832
rect 14672 15744 14680 15808
rect 14744 15744 14760 15808
rect 14824 15744 14840 15808
rect 14904 15744 14920 15808
rect 14984 15744 14992 15808
rect 14672 14720 14992 15744
rect 14672 14656 14680 14720
rect 14744 14656 14760 14720
rect 14824 14656 14840 14720
rect 14904 14656 14920 14720
rect 14984 14656 14992 14720
rect 14672 13632 14992 14656
rect 14672 13568 14680 13632
rect 14744 13568 14760 13632
rect 14824 13568 14840 13632
rect 14904 13568 14920 13632
rect 14984 13568 14992 13632
rect 14672 12544 14992 13568
rect 14672 12480 14680 12544
rect 14744 12480 14760 12544
rect 14824 12480 14840 12544
rect 14904 12480 14920 12544
rect 14984 12480 14992 12544
rect 14672 11456 14992 12480
rect 14672 11392 14680 11456
rect 14744 11392 14760 11456
rect 14824 11392 14840 11456
rect 14904 11392 14920 11456
rect 14984 11392 14992 11456
rect 14672 10368 14992 11392
rect 14672 10304 14680 10368
rect 14744 10304 14760 10368
rect 14824 10304 14840 10368
rect 14904 10304 14920 10368
rect 14984 10304 14992 10368
rect 14672 9280 14992 10304
rect 14672 9216 14680 9280
rect 14744 9216 14760 9280
rect 14824 9216 14840 9280
rect 14904 9216 14920 9280
rect 14984 9216 14992 9280
rect 14672 8192 14992 9216
rect 14672 8128 14680 8192
rect 14744 8128 14760 8192
rect 14824 8128 14840 8192
rect 14904 8128 14920 8192
rect 14984 8128 14992 8192
rect 14672 7104 14992 8128
rect 14672 7040 14680 7104
rect 14744 7040 14760 7104
rect 14824 7040 14840 7104
rect 14904 7040 14920 7104
rect 14984 7040 14992 7104
rect 14672 6016 14992 7040
rect 14672 5952 14680 6016
rect 14744 5952 14760 6016
rect 14824 5952 14840 6016
rect 14904 5952 14920 6016
rect 14984 5952 14992 6016
rect 14672 4928 14992 5952
rect 14672 4864 14680 4928
rect 14744 4864 14760 4928
rect 14824 4864 14840 4928
rect 14904 4864 14920 4928
rect 14984 4864 14992 4928
rect 14672 3840 14992 4864
rect 14672 3776 14680 3840
rect 14744 3776 14760 3840
rect 14824 3776 14840 3840
rect 14904 3776 14920 3840
rect 14984 3776 14992 3840
rect 14672 2752 14992 3776
rect 14672 2688 14680 2752
rect 14744 2688 14760 2752
rect 14824 2688 14840 2752
rect 14904 2688 14920 2752
rect 14984 2688 14992 2752
rect 14672 2128 14992 2688
rect 18104 19616 18424 20176
rect 18104 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18272 19616
rect 18336 19552 18352 19616
rect 18416 19552 18424 19616
rect 18104 18528 18424 19552
rect 18104 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18272 18528
rect 18336 18464 18352 18528
rect 18416 18464 18424 18528
rect 18104 17440 18424 18464
rect 19931 18324 19997 18325
rect 19931 18260 19932 18324
rect 19996 18260 19997 18324
rect 19931 18259 19997 18260
rect 18104 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18272 17440
rect 18336 17376 18352 17440
rect 18416 17376 18424 17440
rect 18104 16352 18424 17376
rect 18104 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18272 16352
rect 18336 16288 18352 16352
rect 18416 16288 18424 16352
rect 18104 15264 18424 16288
rect 18104 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18272 15264
rect 18336 15200 18352 15264
rect 18416 15200 18424 15264
rect 18104 14176 18424 15200
rect 18104 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18272 14176
rect 18336 14112 18352 14176
rect 18416 14112 18424 14176
rect 18104 13088 18424 14112
rect 18104 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18272 13088
rect 18336 13024 18352 13088
rect 18416 13024 18424 13088
rect 18104 12000 18424 13024
rect 18104 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18272 12000
rect 18336 11936 18352 12000
rect 18416 11936 18424 12000
rect 18104 10912 18424 11936
rect 18104 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18272 10912
rect 18336 10848 18352 10912
rect 18416 10848 18424 10912
rect 18104 9824 18424 10848
rect 19934 10709 19994 18259
rect 19931 10708 19997 10709
rect 19931 10644 19932 10708
rect 19996 10644 19997 10708
rect 19931 10643 19997 10644
rect 18104 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18272 9824
rect 18336 9760 18352 9824
rect 18416 9760 18424 9824
rect 18104 8736 18424 9760
rect 18104 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18272 8736
rect 18336 8672 18352 8736
rect 18416 8672 18424 8736
rect 18104 7648 18424 8672
rect 18104 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18272 7648
rect 18336 7584 18352 7648
rect 18416 7584 18424 7648
rect 18104 6560 18424 7584
rect 18104 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18272 6560
rect 18336 6496 18352 6560
rect 18416 6496 18424 6560
rect 18104 5472 18424 6496
rect 18104 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18272 5472
rect 18336 5408 18352 5472
rect 18416 5408 18424 5472
rect 18104 4384 18424 5408
rect 18104 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18272 4384
rect 18336 4320 18352 4384
rect 18416 4320 18424 4384
rect 18104 3296 18424 4320
rect 18104 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18272 3296
rect 18336 3232 18352 3296
rect 18416 3232 18424 3296
rect 18104 2208 18424 3232
rect 18104 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18272 2208
rect 18336 2144 18352 2208
rect 18416 2144 18424 2208
rect 18104 2128 18424 2144
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 2392 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606821651
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606821651
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 1380 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_11
timestamp 1606821651
transform 1 0 2116 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3404 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1606821651
transform 1 0 4048 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_66 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp 1606821651
transform 1 0 4876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_41
timestamp 1606821651
transform 1 0 4876 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1606821651
transform 1 0 5336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1606821651
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5796 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5704 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _033_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 5060 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1606821651
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60
timestamp 1606821651
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606821651
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_67
timestamp 1606821651
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6808 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _116_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8464 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6900 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1606821651
transform 1 0 7728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8096 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78
timestamp 1606821651
transform 1 0 8280 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 10672 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9016 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9752 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68
timestamp 1606821651
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 9016 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1606821651
transform 1 0 9568 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606821651
transform 1 0 10580 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_84
timestamp 1606821651
transform 1 0 8832 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1606821651
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_111
timestamp 1606821651
transform 1 0 11316 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10764 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 11500 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_123
timestamp 1606821651
transform 1 0 12420 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1606821651
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_123
timestamp 1606821651
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1606821651
transform 1 0 12052 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606821651
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1606821651
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12604 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _113_
timestamp 1606821651
transform 1 0 12604 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1606821651
transform 1 0 13156 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 1606821651
transform 1 0 12972 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _112_
timestamp 1606821651
transform 1 0 13156 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 1606821651
transform 1 0 13524 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13340 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _110_
timestamp 1606821651
transform 1 0 13708 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_139
timestamp 1606821651
transform 1 0 13892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_141
timestamp 1606821651
transform 1 0 14076 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14076 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _107_
timestamp 1606821651
transform 1 0 14260 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1606821651
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_147
timestamp 1606821651
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 14812 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _106_
timestamp 1606821651
transform 1 0 14812 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_155
timestamp 1606821651
transform 1 0 15364 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1606821651
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606821651
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 15548 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _109_
timestamp 1606821651
transform 1 0 15456 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_163
timestamp 1606821651
transform 1 0 16100 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1606821651
transform 1 0 16376 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_160
timestamp 1606821651
transform 1 0 15824 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _105_
timestamp 1606821651
transform 1 0 16008 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _102_
timestamp 1606821651
transform 1 0 16376 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_170
timestamp 1606821651
transform 1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1606821651
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1606821651
transform 1 0 16928 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _104_
timestamp 1606821651
transform 1 0 16560 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _101_
timestamp 1606821651
transform 1 0 17112 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1606821651
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606821651
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606821651
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1606821651
transform 1 0 17480 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606821651
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606821651
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _056_
timestamp 1606821651
transform 1 0 17664 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1606821651
transform 1 0 18584 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19596 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 20056 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_199
timestamp 1606821651
transform 1 0 19412 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_200
timestamp 1606821651
transform 1 0 19504 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606821651
transform -1 0 21620 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606821651
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606821651
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_210
timestamp 1606821651
transform 1 0 20424 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_216
timestamp 1606821651
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_218
timestamp 1606821651
transform 1 0 21160 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_218
timestamp 1606821651
transform 1 0 21160 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2576 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606821651
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606821651
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_15
timestamp 1606821651
transform 1 0 2484 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1606821651
transform 1 0 4048 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606821651
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_25
timestamp 1606821651
transform 1 0 3404 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_41
timestamp 1606821651
transform 1 0 4876 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 5796 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1606821651
transform 1 0 5612 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1606821651
transform 1 0 7452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1606821651
transform 1 0 7268 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72
timestamp 1606821651
transform 1 0 7728 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_76
timestamp 1606821651
transform 1 0 8096 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 10488 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9660 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606821651
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_86
timestamp 1606821651
transform 1 0 9016 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_2_99
timestamp 1606821651
transform 1 0 10212 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_111
timestamp 1606821651
transform 1 0 11316 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_122
timestamp 1606821651
transform 1 0 12328 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _111_
timestamp 1606821651
transform 1 0 13616 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_133
timestamp 1606821651
transform 1 0 13340 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1606821651
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 16376 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606821651
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1606821651
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_163
timestamp 1606821651
transform 1 0 16100 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1606821651
transform 1 0 18032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1606821651
transform 1 0 17848 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 1606821651
transform 1 0 18308 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18492 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1606821651
transform 1 0 19780 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_2_198
timestamp 1606821651
transform 1 0 19320 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_202
timestamp 1606821651
transform 1 0 19688 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606821651
transform -1 0 21620 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606821651
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1606821651
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_215
timestamp 1606821651
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_219
timestamp 1606821651
transform 1 0 21252 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1840 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606821651
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 1606821651
transform 1 0 1380 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 1606821651
transform 1 0 1748 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4508 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3496 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1606821651
transform 1 0 3312 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1606821651
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5520 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606821651
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_46
timestamp 1606821651
transform 1 0 5336 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1606821651
transform 1 0 6348 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_62
timestamp 1606821651
transform 1 0 6808 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 7636 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_3_70
timestamp 1606821651
transform 1 0 7544 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10212 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 9384 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_87
timestamp 1606821651
transform 1 0 9108 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp 1606821651
transform 1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1606821651
transform 1 0 11868 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606821651
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1606821651
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1606821651
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13708 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_132
timestamp 1606821651
transform 1 0 13248 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_136
timestamp 1606821651
transform 1 0 13616 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1606821651
transform 1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15824 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_153
timestamp 1606821651
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1606821651
transform 1 0 15640 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16836 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606821651
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1606821651
transform 1 0 16652 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_180
timestamp 1606821651
transform 1 0 17664 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1606821651
transform 1 0 19044 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1606821651
transform 1 0 20056 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1606821651
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1606821651
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606821651
transform -1 0 21620 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_215
timestamp 1606821651
transform 1 0 20884 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_219
timestamp 1606821651
transform 1 0 21252 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 2300 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606821651
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1606821651
transform 1 0 1380 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1606821651
transform 1 0 2116 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4324 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606821651
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1606821651
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 1606821651
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5980 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_51
timestamp 1606821651
transform 1 0 5796 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1606821651
transform 1 0 6808 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8188 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1606821651
transform 1 0 7176 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_75
timestamp 1606821651
transform 1 0 8004 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10672 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9660 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606821651
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_86
timestamp 1606821651
transform 1 0 9016 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_102
timestamp 1606821651
transform 1 0 10488 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11684 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_113
timestamp 1606821651
transform 1 0 11500 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_124
timestamp 1606821651
transform 1 0 12512 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _114_
timestamp 1606821651
transform 1 0 12788 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13340 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1606821651
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _108_
timestamp 1606821651
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1606821651
transform 1 0 16376 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606821651
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606821651
transform 1 0 14812 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1606821651
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1606821651
transform 1 0 16008 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1606821651
transform 1 0 17388 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_175
timestamp 1606821651
transform 1 0 17204 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_186
timestamp 1606821651
transform 1 0 18216 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18400 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20056 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_204
timestamp 1606821651
transform 1 0 19872 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606821651
transform -1 0 21620 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606821651
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_212
timestamp 1606821651
transform 1 0 20608 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_215
timestamp 1606821651
transform 1 0 20884 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_219
timestamp 1606821651
transform 1 0 21252 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2024 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606821651
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_3
timestamp 1606821651
transform 1 0 1380 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_9
timestamp 1606821651
transform 1 0 1932 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1606821651
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4876 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_31
timestamp 1606821651
transform 1 0 3956 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_39
timestamp 1606821651
transform 1 0 4692 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606821651
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_50
timestamp 1606821651
transform 1 0 5704 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_58
timestamp 1606821651
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1606821651
transform 1 0 6808 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 7268 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 8556 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 8280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1606821651
transform 1 0 7176 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_76
timestamp 1606821651
transform 1 0 8096 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10120 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_5_90
timestamp 1606821651
transform 1 0 9384 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _115_
timestamp 1606821651
transform 1 0 12420 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1606821651
transform 1 0 11132 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606821651
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_107
timestamp 1606821651
transform 1 0 10948 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_118
timestamp 1606821651
transform 1 0 11960 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13064 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13984 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_5_127
timestamp 1606821651
transform 1 0 12788 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_139
timestamp 1606821651
transform 1 0 13892 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _097_
timestamp 1606821651
transform 1 0 15180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15732 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 14996 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1606821651
transform 1 0 14812 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1606821651
transform 1 0 15548 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _100_
timestamp 1606821651
transform 1 0 17388 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606821651
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_175
timestamp 1606821651
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1606821651
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _103_
timestamp 1606821651
transform 1 0 19044 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19596 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1606821651
transform 1 0 18860 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1606821651
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606821651
transform -1 0 21620 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 1606821651
transform 1 0 21068 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1606821651
transform 1 0 1656 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2116 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606821651
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606821651
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_3
timestamp 1606821651
transform 1 0 1380 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_18
timestamp 1606821651
transform 1 0 2760 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 1606821651
transform 1 0 1380 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_9
timestamp 1606821651
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1606821651
transform 1 0 4876 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1606821651
transform 1 0 3772 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606821651
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1606821651
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1606821651
transform 1 0 3588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_38
timestamp 1606821651
transform 1 0 4600 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_50
timestamp 1606821651
transform 1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_48
timestamp 1606821651
transform 1 0 5520 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 5888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5796 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606821651
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1606821651
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1606821651
transform 1 0 6624 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606821651
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1606821651
transform 1 0 6808 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1606821651
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6808 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8096 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8556 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_6_78
timestamp 1606821651
transform 1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_71
timestamp 1606821651
transform 1 0 7636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_75
timestamp 1606821651
transform 1 0 8004 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 9752 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1606821651
transform 1 0 10672 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606821651
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1606821651
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_102
timestamp 1606821651
transform 1 0 10488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_92
timestamp 1606821651
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1606821651
transform 1 0 11868 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11684 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606821651
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_113
timestamp 1606821651
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1606821651
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_110
timestamp 1606821651
transform 1 0 11224 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_116
timestamp 1606821651
transform 1 0 11776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 1606821651
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1606821651
transform 1 0 14352 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 12696 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14352 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_142
timestamp 1606821651
transform 1 0 14168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1606821651
transform 1 0 13892 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_143
timestamp 1606821651
transform 1 0 14260 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15916 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606821651
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_147
timestamp 1606821651
transform 1 0 14628 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_6_154
timestamp 1606821651
transform 1 0 15272 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_160
timestamp 1606821651
transform 1 0 15824 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_160
timestamp 1606821651
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _091_
timestamp 1606821651
transform 1 0 17388 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 17572 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606821651
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_177
timestamp 1606821651
transform 1 0 17388 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_171
timestamp 1606821651
transform 1 0 16836 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1606821651
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _098_
timestamp 1606821651
transform 1 0 20240 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19228 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19044 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1606821651
transform 1 0 20240 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_6_195
timestamp 1606821651
transform 1 0 19044 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1606821651
transform 1 0 20056 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1606821651
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_204
timestamp 1606821651
transform 1 0 19872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606821651
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606821651
transform -1 0 21620 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606821651
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606821651
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_215
timestamp 1606821651
transform 1 0 20884 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_219
timestamp 1606821651
transform 1 0 21252 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 1606821651
transform 1 0 21068 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1656 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606821651
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1606821651
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4692 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606821651
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_22
timestamp 1606821651
transform 1 0 3128 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_30
timestamp 1606821651
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1606821651
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1606821651
transform 1 0 4600 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_55
timestamp 1606821651
transform 1 0 6164 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7176 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8188 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_8_63
timestamp 1606821651
transform 1 0 6900 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 1606821651
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1606821651
transform 1 0 9844 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606821651
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_86
timestamp 1606821651
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_8_93
timestamp 1606821651
transform 1 0 9660 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_104
timestamp 1606821651
transform 1 0 10672 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 11040 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1606821651
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13156 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1606821651
transform 1 0 14168 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 12696 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 1606821651
transform 1 0 12972 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_140
timestamp 1606821651
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1606821651
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1606821651
transform 1 0 16100 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606821651
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1606821651
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_157
timestamp 1606821651
transform 1 0 15548 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1606821651
transform 1 0 17112 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_172
timestamp 1606821651
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_183
timestamp 1606821651
transform 1 0 17940 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19504 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1606821651
transform 1 0 18492 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1606821651
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606821651
transform -1 0 21620 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606821651
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_209
timestamp 1606821651
transform 1 0 20332 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1606821651
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_215
timestamp 1606821651
transform 1 0 20884 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_219
timestamp 1606821651
transform 1 0 21252 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2116 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606821651
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp 1606821651
transform 1 0 1380 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_20
timestamp 1606821651
transform 1 0 2944 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1606821651
transform 1 0 3128 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1606821651
transform 1 0 4876 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_31
timestamp 1606821651
transform 1 0 3956 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_39
timestamp 1606821651
transform 1 0 4692 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606821651
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_50
timestamp 1606821651
transform 1 0 5704 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_58
timestamp 1606821651
transform 1 0 6440 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1606821651
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 8464 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6900 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7912 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_72
timestamp 1606821651
transform 1 0 7728 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_77
timestamp 1606821651
transform 1 0 8188 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10120 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1606821651
transform 1 0 9936 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1606821651
transform 1 0 11132 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606821651
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_107
timestamp 1606821651
transform 1 0 10948 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_118
timestamp 1606821651
transform 1 0 11960 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13616 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_9_132
timestamp 1606821651
transform 1 0 13248 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 16284 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15272 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1606821651
transform 1 0 15088 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_163
timestamp 1606821651
transform 1 0 16100 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1606821651
transform 1 0 18124 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606821651
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1606821651
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1606821651
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19688 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1606821651
transform 1 0 18676 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_9_188
timestamp 1606821651
transform 1 0 18400 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1606821651
transform 1 0 19504 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _099_
timestamp 1606821651
transform 1 0 20700 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606821651
transform -1 0 21620 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_211
timestamp 1606821651
transform 1 0 20516 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp 1606821651
transform 1 0 21068 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1606821651
transform 1 0 2944 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1606821651
transform 1 0 1932 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606821651
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_3
timestamp 1606821651
transform 1 0 1380 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_18
timestamp 1606821651
transform 1 0 2760 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1606821651
transform 1 0 4048 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606821651
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1606821651
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1606821651
transform 1 0 4876 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1606821651
transform 1 0 5244 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1606821651
transform 1 0 6348 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_10_54
timestamp 1606821651
transform 1 0 6072 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1606821651
transform 1 0 8556 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7360 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1606821651
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_77
timestamp 1606821651
transform 1 0 8188 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1606821651
transform 1 0 10120 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606821651
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1606821651
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_93
timestamp 1606821651
transform 1 0 9660 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_97
timestamp 1606821651
transform 1 0 10028 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11500 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1606821651
transform 1 0 12512 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_107
timestamp 1606821651
transform 1 0 10948 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1606821651
transform 1 0 12328 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13340 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14168 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 15732 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606821651
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 15456 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606821651
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_154
timestamp 1606821651
transform 1 0 15272 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 17664 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_175
timestamp 1606821651
transform 1 0 17204 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_179
timestamp 1606821651
transform 1 0 17572 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1606821651
transform 1 0 19688 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_10_196
timestamp 1606821651
transform 1 0 19136 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1606821651
transform 1 0 20884 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606821651
transform -1 0 21620 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606821651
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1606821651
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_218
timestamp 1606821651
transform 1 0 21160 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 1840 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606821651
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1606821651
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp 1606821651
transform 1 0 1748 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4140 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_11_24
timestamp 1606821651
transform 1 0 3312 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_32
timestamp 1606821651
transform 1 0 4048 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1606821651
transform 1 0 6256 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1606821651
transform 1 0 5152 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606821651
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 1606821651
transform 1 0 4968 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_53
timestamp 1606821651
transform 1 0 5980 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606821651
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1606821651
transform 1 0 8004 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8464 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1606821651
transform 1 0 7636 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_78
timestamp 1606821651
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10672 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_11_96
timestamp 1606821651
transform 1 0 9936 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1606821651
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606821651
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1606821651
transform 1 0 12144 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13432 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1606821651
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15180 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_11_150
timestamp 1606821651
transform 1 0 14904 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_162
timestamp 1606821651
transform 1 0 16008 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1606821651
transform 1 0 16744 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606821651
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1606821651
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_184
timestamp 1606821651
transform 1 0 18032 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1606821651
transform 1 0 19964 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1606821651
transform 1 0 18952 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_192
timestamp 1606821651
transform 1 0 18768 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_203
timestamp 1606821651
transform 1 0 19780 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606821651
transform -1 0 21620 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_214
timestamp 1606821651
transform 1 0 20792 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1606821651
transform 1 0 2024 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606821651
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1606821651
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1606821651
transform 1 0 1932 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1606821651
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1606821651
transform 1 0 3036 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1606821651
transform 1 0 4416 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606821651
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_24
timestamp 1606821651
transform 1 0 3312 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1606821651
transform 1 0 3864 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_32
timestamp 1606821651
transform 1 0 4048 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1606821651
transform 1 0 5428 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6164 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_45
timestamp 1606821651
transform 1 0 5244 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_50
timestamp 1606821651
transform 1 0 5704 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_54
timestamp 1606821651
transform 1 0 6072 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1606821651
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 7820 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_71
timestamp 1606821651
transform 1 0 7636 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1606821651
transform 1 0 8096 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606821651
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606821651
transform 1 0 10672 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1606821651
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1606821651
transform 1 0 10488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 12512 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1606821651
transform 1 0 14168 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_140
timestamp 1606821651
transform 1 0 13984 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 15272 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606821651
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1606821651
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_170
timestamp 1606821651
transform 1 0 16744 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_181
timestamp 1606821651
transform 1 0 17756 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_187
timestamp 1606821651
transform 1 0 18308 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _085_
timestamp 1606821651
transform 1 0 20240 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 18400 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_12_204
timestamp 1606821651
transform 1 0 19872 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606821651
transform -1 0 21620 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606821651
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1606821651
transform 1 0 20608 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1606821651
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1606821651
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 1748 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1606821651
transform 1 0 2852 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1840 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606821651
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606821651
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1606821651
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1606821651
transform 1 0 1748 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_17
timestamp 1606821651
transform 1 0 2668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1606821651
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1606821651
transform 1 0 4232 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1606821651
transform 1 0 3956 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606821651
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_28
timestamp 1606821651
transform 1 0 3680 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_40
timestamp 1606821651
transform 1 0 4784 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1606821651
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1606821651
transform 1 0 4048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 6440 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1606821651
transform 1 0 5244 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1606821651
transform 1 0 5520 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606821651
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1606821651
transform 1 0 6348 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1606821651
transform 1 0 5060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1606821651
transform 1 0 6072 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7820 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1606821651
transform 1 0 8096 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_71
timestamp 1606821651
transform 1 0 7636 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_82
timestamp 1606821651
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_74
timestamp 1606821651
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 8832 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 9660 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 10488 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606821651
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp 1606821651
transform 1 0 10304 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1606821651
transform 1 0 8924 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1606821651
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1606821651
transform 1 0 11316 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1606821651
transform 1 0 11592 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12604 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606821651
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1606821651
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_109
timestamp 1606821651
transform 1 0 11132 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_113
timestamp 1606821651
transform 1 0 11500 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1606821651
transform 1 0 12420 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 13616 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1606821651
transform 1 0 14168 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14352 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1606821651
transform 1 0 13892 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1606821651
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_142
timestamp 1606821651
transform 1 0 14168 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_154
timestamp 1606821651
transform 1 0 15272 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606821651
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_147
timestamp 1606821651
transform 1 0 14628 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1606821651
transform 1 0 14996 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 14812 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606821651
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1606821651
transform 1 0 15180 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1606821651
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1606821651
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1606821651
transform 1 0 15456 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1606821651
transform 1 0 16192 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_176
timestamp 1606821651
transform 1 0 17296 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_171
timestamp 1606821651
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_167
timestamp 1606821651
transform 1 0 16468 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1606821651
transform 1 0 16928 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16468 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_187
timestamp 1606821651
transform 1 0 18308 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_181
timestamp 1606821651
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606821651
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1606821651
transform 1 0 17480 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606821651
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19688 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 18676 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_13_196
timestamp 1606821651
transform 1 0 19136 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1606821651
transform 1 0 20148 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1606821651
transform 1 0 20332 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606821651
transform -1 0 21620 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606821651
transform -1 0 21620 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606821651
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1606821651
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1606821651
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_215
timestamp 1606821651
transform 1 0 20884 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 1606821651
transform 1 0 21252 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606821651
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_3
timestamp 1606821651
transform 1 0 1380 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_9
timestamp 1606821651
transform 1 0 1932 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1606821651
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4048 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1606821651
transform 1 0 3036 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_30
timestamp 1606821651
transform 1 0 3864 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1606821651
transform 1 0 5704 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606821651
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1606821651
transform 1 0 5520 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606821651
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1606821651
transform 1 0 8556 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_78
timestamp 1606821651
transform 1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 10028 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 9016 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1606821651
transform 1 0 8832 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_95
timestamp 1606821651
transform 1 0 9844 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 12420 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1606821651
transform 1 0 11316 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606821651
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_106
timestamp 1606821651
transform 1 0 10856 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_110
timestamp 1606821651
transform 1 0 11224 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606821651
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1606821651
transform 1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_139
timestamp 1606821651
transform 1 0 13892 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1606821651
transform 1 0 15456 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1606821651
transform 1 0 15088 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_165
timestamp 1606821651
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 18032 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606821651
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 17480 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1606821651
transform 1 0 17296 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606821651
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 19688 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 1606821651
transform 1 0 19504 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606821651
transform -1 0 21620 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1606821651
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 1840 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606821651
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1606821651
transform 1 0 1380 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1606821651
transform 1 0 1748 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1606821651
transform 1 0 3496 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 4232 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606821651
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_24
timestamp 1606821651
transform 1 0 3312 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1606821651
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1606821651
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 5888 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_50
timestamp 1606821651
transform 1 0 5704 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7544 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1606821651
transform 1 0 8556 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_68
timestamp 1606821651
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1606821651
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 9660 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 10672 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606821651
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 1606821651
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_102
timestamp 1606821651
transform 1 0 10488 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 11500 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_110
timestamp 1606821651
transform 1 0 11224 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13340 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_129
timestamp 1606821651
transform 1 0 12972 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1606821651
transform 1 0 16284 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1606821651
transform 1 0 15272 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606821651
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606821651
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 1606821651
transform 1 0 16100 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16836 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 1606821651
transform 1 0 16560 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_187
timestamp 1606821651
transform 1 0 18308 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1606821651
transform 1 0 18768 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1606821651
transform 1 0 19780 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_16_191
timestamp 1606821651
transform 1 0 18676 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1606821651
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606821651
transform -1 0 21620 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606821651
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1606821651
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_215
timestamp 1606821651
transform 1 0 20884 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_219
timestamp 1606821651
transform 1 0 21252 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2852 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1606821651
transform 1 0 1840 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606821651
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606821651
transform 1 0 1380 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_7
timestamp 1606821651
transform 1 0 1748 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_17
timestamp 1606821651
transform 1 0 2668 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3588 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_25
timestamp 1606821651
transform 1 0 3404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_36
timestamp 1606821651
transform 1 0 4416 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4968 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606821651
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 5980 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_51
timestamp 1606821651
transform 1 0 5796 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_56
timestamp 1606821651
transform 1 0 6256 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1606821651
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_62
timestamp 1606821651
transform 1 0 6808 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8740 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1606821651
transform 1 0 7452 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 8464 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_68
timestamp 1606821651
transform 1 0 7360 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_78
timestamp 1606821651
transform 1 0 8280 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10396 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1606821651
transform 1 0 10212 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1606821651
transform 1 0 12420 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606821651
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1606821651
transform 1 0 11868 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606821651
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 13892 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1606821651
transform 1 0 13432 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1606821651
transform 1 0 13248 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1606821651
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 15548 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_155
timestamp 1606821651
transform 1 0 15364 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1606821651
transform 1 0 18032 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 17204 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606821651
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_173
timestamp 1606821651
transform 1 0 17020 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606821651
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 19044 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1606821651
transform 1 0 18860 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _081_
timestamp 1606821651
transform 1 0 20700 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606821651
transform -1 0 21620 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_211
timestamp 1606821651
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 1606821651
transform 1 0 21068 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1606821651
transform 1 0 1380 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1606821651
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606821651
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_12
timestamp 1606821651
transform 1 0 2208 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _076_
timestamp 1606821651
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606821651
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1606821651
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1606821651
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 6256 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_18_48
timestamp 1606821651
transform 1 0 5520 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1606821651
transform 1 0 7912 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1606821651
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_83
timestamp 1606821651
transform 1 0 8740 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1606821651
transform 1 0 9752 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606821651
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1606821651
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1606821651
transform 1 0 9660 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_103
timestamp 1606821651
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 10764 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1606821651
transform 1 0 12420 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1606821651
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1606821651
transform 1 0 13432 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1606821651
transform 1 0 14076 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_132
timestamp 1606821651
transform 1 0 13248 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_137
timestamp 1606821651
transform 1 0 13708 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1606821651
transform 1 0 15916 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606821651
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_150
timestamp 1606821651
transform 1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_154
timestamp 1606821651
transform 1 0 15272 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_160
timestamp 1606821651
transform 1 0 15824 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1606821651
transform 1 0 17940 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1606821651
transform 1 0 16928 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1606821651
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1606821651
transform 1 0 17756 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _095_
timestamp 1606821651
transform 1 0 20240 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1606821651
transform 1 0 19136 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1606821651
transform 1 0 18952 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_192
timestamp 1606821651
transform 1 0 18768 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_205
timestamp 1606821651
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1606821651
transform 1 0 20884 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606821651
transform -1 0 21620 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606821651
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606821651
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_218
timestamp 1606821651
transform 1 0 21160 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1606821651
transform 1 0 1748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1606821651
transform 1 0 1380 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606821651
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606821651
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1606821651
transform 1 0 1932 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1748 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _074_
timestamp 1606821651
transform 1 0 1380 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_18
timestamp 1606821651
transform 1 0 2760 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1606821651
transform 1 0 2300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1606821651
transform 1 0 2484 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1606821651
transform 1 0 2944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 1606821651
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_28
timestamp 1606821651
transform 1 0 3680 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_24
timestamp 1606821651
transform 1 0 3312 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606821651
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1606821651
transform 1 0 3772 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1606821651
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1606821651
transform 1 0 4600 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1606821651
transform 1 0 4692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _075_
timestamp 1606821651
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 4784 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1606821651
transform 1 0 6256 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606821651
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_56
timestamp 1606821651
transform 1 0 6256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_60
timestamp 1606821651
transform 1 0 6624 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_48
timestamp 1606821651
transform 1 0 5520 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 7268 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1606821651
transform 1 0 7820 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1606821651
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_82
timestamp 1606821651
transform 1 0 8648 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1606821651
transform 1 0 7084 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1606821651
transform 1 0 8740 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1606821651
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1606821651
transform 1 0 10028 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1606821651
transform 1 0 9016 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1606821651
transform 1 0 10120 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606821651
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_95
timestamp 1606821651
transform 1 0 9844 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606821651
transform 1 0 9476 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_96
timestamp 1606821651
transform 1 0 9936 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_107
timestamp 1606821651
transform 1 0 10948 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1606821651
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1606821651
transform 1 0 11040 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1606821651
transform 1 0 11132 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_118
timestamp 1606821651
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1606821651
transform 1 0 12236 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1606821651
transform 1 0 11868 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606821651
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1606821651
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1606821651
transform 1 0 12512 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 13064 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1606821651
transform 1 0 13800 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_19_132
timestamp 1606821651
transform 1 0 13248 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_127
timestamp 1606821651
transform 1 0 12788 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_154
timestamp 1606821651
transform 1 0 15272 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1606821651
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_146
timestamp 1606821651
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1606821651
transform 1 0 15364 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_147
timestamp 1606821651
transform 1 0 14628 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606821651
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1606821651
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1606821651
transform 1 0 16376 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1606821651
transform 1 0 15548 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 15548 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 17756 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 18216 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1606821651
transform 1 0 16560 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606821651
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1606821651
transform 1 0 17388 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_184
timestamp 1606821651
transform 1 0 18032 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_173
timestamp 1606821651
transform 1 0 17020 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1606821651
transform 1 0 19412 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19964 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_19_202
timestamp 1606821651
transform 1 0 19688 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_197
timestamp 1606821651
transform 1 0 19228 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_208
timestamp 1606821651
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _077_
timestamp 1606821651
transform 1 0 20700 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606821651
transform -1 0 21620 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606821651
transform -1 0 21620 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606821651
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_211
timestamp 1606821651
transform 1 0 20516 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 1606821651
transform 1 0 21068 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_215
timestamp 1606821651
transform 1 0 20884 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_219
timestamp 1606821651
transform 1 0 21252 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 2392 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_4  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 1656 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606821651
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1606821651
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1606821651
transform 1 0 2208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 4048 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_30
timestamp 1606821651
transform 1 0 3864 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1606821651
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606821651
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_48
timestamp 1606821651
transform 1 0 5520 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp 1606821651
transform 1 0 6624 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1606821651
transform 1 0 7820 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1606821651
transform 1 0 8372 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1606821651
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_76
timestamp 1606821651
transform 1 0 8096 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 10672 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_21_95
timestamp 1606821651
transform 1 0 9844 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_103
timestamp 1606821651
transform 1 0 10580 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606821651
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_120
timestamp 1606821651
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_123
timestamp 1606821651
transform 1 0 12420 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1606821651
transform 1 0 13156 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 14812 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1606821651
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_165
timestamp 1606821651
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1606821651
transform 1 0 17480 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1606821651
transform 1 0 16468 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18032 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606821651
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1606821651
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606821651
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _093_
timestamp 1606821651
transform 1 0 19320 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _094_
timestamp 1606821651
transform 1 0 18768 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19872 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_190
timestamp 1606821651
transform 1 0 18584 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1606821651
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1606821651
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_4  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 20608 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606821651
transform -1 0 21620 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1606821651
transform 1 0 20424 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_218
timestamp 1606821651
transform 1 0 21160 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _073_
timestamp 1606821651
transform 1 0 1472 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1606821651
transform 1 0 2760 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2024 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606821651
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 1606821651
transform 1 0 1380 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_8
timestamp 1606821651
transform 1 0 1840 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_16
timestamp 1606821651
transform 1 0 2576 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _058_
timestamp 1606821651
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606821651
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606821651
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_36
timestamp 1606821651
transform 1 0 4416 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_48
timestamp 1606821651
transform 1 0 5520 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_60
timestamp 1606821651
transform 1 0 6624 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_72
timestamp 1606821651
transform 1 0 7728 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606821651
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1606821651
transform 1 0 8832 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 11776 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_22_109
timestamp 1606821651
transform 1 0 11132 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_115
timestamp 1606821651
transform 1 0 11684 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1606821651
transform 1 0 13432 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_132
timestamp 1606821651
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_143
timestamp 1606821651
transform 1 0 14260 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1606821651
transform 1 0 15732 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606821651
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606821651
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1606821651
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1606821651
transform 1 0 15640 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1606821651
transform 1 0 16744 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1606821651
transform 1 0 16560 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_186
timestamp 1606821651
transform 1 0 18216 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _096_
timestamp 1606821651
transform 1 0 19136 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19688 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1606821651
transform 1 0 18952 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_200
timestamp 1606821651
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_208
timestamp 1606821651
transform 1 0 20240 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606821651
transform -1 0 21620 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606821651
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1606821651
transform 1 0 20884 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_219
timestamp 1606821651
transform 1 0 21252 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _071_
timestamp 1606821651
transform 1 0 2300 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _072_
timestamp 1606821651
transform 1 0 1748 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1606821651
transform 1 0 2944 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606821651
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1606821651
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1606821651
transform 1 0 2116 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_17
timestamp 1606821651
transform 1 0 2668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_36
timestamp 1606821651
transform 1 0 4416 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606821651
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_48
timestamp 1606821651
transform 1 0 5520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1606821651
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1606821651
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1606821651
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1606821651
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1606821651
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606821651
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1606821651
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1606821651
transform 1 0 12420 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1606821651
transform 1 0 13708 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_135
timestamp 1606821651
transform 1 0 13524 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_146
timestamp 1606821651
transform 1 0 14536 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_158
timestamp 1606821651
transform 1 0 15640 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606821651
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_170
timestamp 1606821651
transform 1 0 16744 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1606821651
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606821651
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _079_
timestamp 1606821651
transform 1 0 19964 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _092_
timestamp 1606821651
transform 1 0 19412 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_196
timestamp 1606821651
transform 1 0 19136 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_203
timestamp 1606821651
transform 1 0 19780 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1606821651
transform 1 0 20516 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606821651
transform -1 0 21620 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1606821651
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_215
timestamp 1606821651
transform 1 0 20884 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_219
timestamp 1606821651
transform 1 0 21252 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _059_
timestamp 1606821651
transform 1 0 2300 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _070_
timestamp 1606821651
transform 1 0 1748 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606821651
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1606821651
transform 1 0 1380 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_11
timestamp 1606821651
transform 1 0 2116 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_17
timestamp 1606821651
transform 1 0 2668 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 4048 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606821651
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1606821651
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_38
timestamp 1606821651
transform 1 0 4600 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_50
timestamp 1606821651
transform 1 0 5704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_62
timestamp 1606821651
transform 1 0 6808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_74
timestamp 1606821651
transform 1 0 7912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606821651
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_86
timestamp 1606821651
transform 1 0 9016 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606821651
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 12512 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606821651
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_117
timestamp 1606821651
transform 1 0 11868 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_123
timestamp 1606821651
transform 1 0 12420 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_130
timestamp 1606821651
transform 1 0 13064 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_142
timestamp 1606821651
transform 1 0 14168 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606821651
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_150
timestamp 1606821651
transform 1 0 14904 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1606821651
transform 1 0 15272 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1606821651
transform 1 0 16376 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1606821651
transform 1 0 17480 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _090_
timestamp 1606821651
transform 1 0 20240 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606821651
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_202
timestamp 1606821651
transform 1 0 19688 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606821651
transform -1 0 21620 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606821651
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1606821651
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_215
timestamp 1606821651
transform 1 0 20884 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_219
timestamp 1606821651
transform 1 0 21252 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _057_
timestamp 1606821651
transform 1 0 2300 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _069_
timestamp 1606821651
transform 1 0 1748 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606821651
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1606821651
transform 1 0 1380 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_11
timestamp 1606821651
transform 1 0 2116 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_17
timestamp 1606821651
transform 1 0 2668 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _068_
timestamp 1606821651
transform 1 0 3220 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1606821651
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1606821651
transform 1 0 4692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606821651
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1606821651
transform 1 0 5796 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1606821651
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606821651
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606821651
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1606821651
transform 1 0 9016 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1606821651
transform 1 0 10120 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606821651
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1606821651
transform 1 0 11224 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1606821651
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _088_
timestamp 1606821651
transform 1 0 13340 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1606821651
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1606821651
transform 1 0 13708 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1606821651
transform 1 0 14812 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_161
timestamp 1606821651
transform 1 0 15916 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606821651
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_173
timestamp 1606821651
transform 1 0 17020 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1606821651
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606821651
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _089_
timestamp 1606821651
transform 1 0 19964 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_196
timestamp 1606821651
transform 1 0 19136 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1606821651
transform 1 0 19872 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _087_
timestamp 1606821651
transform 1 0 20516 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606821651
transform -1 0 21620 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1606821651
transform 1 0 20332 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_215
timestamp 1606821651
transform 1 0 20884 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_219
timestamp 1606821651
transform 1 0 21252 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _066_
timestamp 1606821651
transform 1 0 1748 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _067_
timestamp 1606821651
transform 1 0 1748 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606821651
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606821651
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1606821651
transform 1 0 1380 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1606821651
transform 1 0 2116 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606821651
transform 1 0 1380 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_11
timestamp 1606821651
transform 1 0 2116 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606821651
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1606821651
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606821651
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_23
timestamp 1606821651
transform 1 0 3220 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_35
timestamp 1606821651
transform 1 0 4324 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606821651
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606821651
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606821651
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_47
timestamp 1606821651
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606821651
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606821651
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606821651
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606821651
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_74
timestamp 1606821651
transform 1 0 7912 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606821651
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606821651
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1606821651
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1606821651
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606821651
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606821651
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1606821651
transform 1 0 11868 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_110
timestamp 1606821651
transform 1 0 11224 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1606821651
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1606821651
transform 1 0 12972 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1606821651
transform 1 0 14076 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1606821651
transform 1 0 13524 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606821651
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1606821651
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1606821651
transform 1 0 16376 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1606821651
transform 1 0 14628 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1606821651
transform 1 0 15732 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606821651
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606821651
transform 1 0 17480 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1606821651
transform 1 0 16836 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606821651
transform 1 0 18032 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _083_
timestamp 1606821651
transform 1 0 20240 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606821651
transform 1 0 18584 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_202
timestamp 1606821651
transform 1 0 19688 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606821651
transform 1 0 19136 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_208
timestamp 1606821651
transform 1 0 20240 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _086_
timestamp 1606821651
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606821651
transform -1 0 21620 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606821651
transform -1 0 21620 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606821651
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1606821651
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_215
timestamp 1606821651
transform 1 0 20884 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_219
timestamp 1606821651
transform 1 0 21252 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1606821651
transform 1 0 20884 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_219
timestamp 1606821651
transform 1 0 21252 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _065_
timestamp 1606821651
transform 1 0 1656 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 2208 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606821651
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1606821651
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_10
timestamp 1606821651
transform 1 0 2024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_18
timestamp 1606821651
transform 1 0 2760 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606821651
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1606821651
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606821651
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606821651
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606821651
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1606821651
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606821651
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606821651
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1606821651
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1606821651
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1606821651
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1606821651
transform 1 0 12972 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1606821651
transform 1 0 14076 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606821651
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1606821651
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1606821651
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1606821651
transform 1 0 17480 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 19688 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1606821651
transform 1 0 18584 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_208
timestamp 1606821651
transform 1 0 20240 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606821651
transform -1 0 21620 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606821651
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_215
timestamp 1606821651
transform 1 0 20884 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_219
timestamp 1606821651
transform 1 0 21252 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _064_
timestamp 1606821651
transform 1 0 1748 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606821651
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1606821651
transform 1 0 1380 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_11
timestamp 1606821651
transform 1 0 2116 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_23
timestamp 1606821651
transform 1 0 3220 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_35
timestamp 1606821651
transform 1 0 4324 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606821651
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_47
timestamp 1606821651
transform 1 0 5428 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606821651
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606821651
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1606821651
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_86
timestamp 1606821651
transform 1 0 9016 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_98
timestamp 1606821651
transform 1 0 10120 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606821651
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_110
timestamp 1606821651
transform 1 0 11224 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1606821651
transform 1 0 12420 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1606821651
transform 1 0 13524 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1606821651
transform 1 0 14628 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1606821651
transform 1 0 15732 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606821651
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1606821651
transform 1 0 16836 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606821651
transform 1 0 18032 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606821651
transform 1 0 19136 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_208
timestamp 1606821651
transform 1 0 20240 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _084_
timestamp 1606821651
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606821651
transform -1 0 21620 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_215
timestamp 1606821651
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_219
timestamp 1606821651
transform 1 0 21252 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _063_
timestamp 1606821651
transform 1 0 1748 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606821651
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_3
timestamp 1606821651
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_11
timestamp 1606821651
transform 1 0 2116 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606821651
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_23
timestamp 1606821651
transform 1 0 3220 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606821651
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 6072 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_44
timestamp 1606821651
transform 1 0 5152 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1606821651
transform 1 0 5888 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_60
timestamp 1606821651
transform 1 0 6624 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_72
timestamp 1606821651
transform 1 0 7728 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606821651
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_84
timestamp 1606821651
transform 1 0 8832 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1606821651
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1606821651
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1606821651
transform 1 0 11868 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1606821651
transform 1 0 12972 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1606821651
transform 1 0 14076 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606821651
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1606821651
transform 1 0 15272 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_166
timestamp 1606821651
transform 1 0 16376 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1606821651
transform 1 0 18124 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_178
timestamp 1606821651
transform 1 0 17480 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_184
timestamp 1606821651
transform 1 0 18032 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_191
timestamp 1606821651
transform 1 0 18676 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_203
timestamp 1606821651
transform 1 0 19780 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606821651
transform -1 0 21620 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606821651
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1606821651
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_215
timestamp 1606821651
transform 1 0 20884 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_219
timestamp 1606821651
transform 1 0 21252 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _061_
timestamp 1606821651
transform 1 0 2300 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _062_
timestamp 1606821651
transform 1 0 1748 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606821651
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1606821651
transform 1 0 1380 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 1606821651
transform 1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_17
timestamp 1606821651
transform 1 0 2668 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1606821651
transform 1 0 3772 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_41
timestamp 1606821651
transform 1 0 4876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _060_
timestamp 1606821651
transform 1 0 5796 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606821651
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1606821651
transform 1 0 5612 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_55
timestamp 1606821651
transform 1 0 6164 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606821651
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1606821651
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1606821651
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1606821651
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606821651
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_110
timestamp 1606821651
transform 1 0 11224 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_123
timestamp 1606821651
transform 1 0 12420 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_135
timestamp 1606821651
transform 1 0 13524 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1606821651
transform 1 0 14628 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_159
timestamp 1606821651
transform 1 0 15732 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606821651
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_171
timestamp 1606821651
transform 1 0 16836 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_184
timestamp 1606821651
transform 1 0 18032 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _080_
timestamp 1606821651
transform 1 0 18952 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1606821651
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_198
timestamp 1606821651
transform 1 0 19320 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _082_
timestamp 1606821651
transform 1 0 20516 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606821651
transform -1 0 21620 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_210
timestamp 1606821651
transform 1 0 20424 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_215
timestamp 1606821651
transform 1 0 20884 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_219
timestamp 1606821651
transform 1 0 21252 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606821651
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606821651
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606821651
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1606821651
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606821651
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606821651
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1606821651
transform 1 0 6808 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606821651
transform 1 0 5152 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1606821651
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_63
timestamp 1606821651
transform 1 0 6900 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_75
timestamp 1606821651
transform 1 0 8004 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1606821651
transform 1 0 9660 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_87
timestamp 1606821651
transform 1 0 9108 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_94
timestamp 1606821651
transform 1 0 9752 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1606821651
transform 1 0 12512 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_106
timestamp 1606821651
transform 1 0 10856 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_118
timestamp 1606821651
transform 1 0 11960 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606821651
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_137
timestamp 1606821651
transform 1 0 13708 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1606821651
transform 1 0 15364 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_149
timestamp 1606821651
transform 1 0 14812 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_156
timestamp 1606821651
transform 1 0 15456 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1606821651
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_168
timestamp 1606821651
transform 1 0 16560 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_180
timestamp 1606821651
transform 1 0 17664 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_187
timestamp 1606821651
transform 1 0 18308 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_199
timestamp 1606821651
transform 1 0 19412 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606821651
transform -1 0 21620 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1606821651
transform 1 0 21068 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_211
timestamp 1606821651
transform 1 0 20516 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606821651
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 21638 0 21694 480 6 SC_IN_BOT
port 0 nsew default input
rlabel metal2 s 22098 0 22154 480 6 SC_OUT_BOT
port 1 nsew default tristate
rlabel metal2 s 202 0 258 480 6 bottom_left_grid_pin_42_
port 2 nsew default input
rlabel metal2 s 570 0 626 480 6 bottom_left_grid_pin_43_
port 3 nsew default input
rlabel metal2 s 1030 0 1086 480 6 bottom_left_grid_pin_44_
port 4 nsew default input
rlabel metal2 s 1490 0 1546 480 6 bottom_left_grid_pin_45_
port 5 nsew default input
rlabel metal2 s 1950 0 2006 480 6 bottom_left_grid_pin_46_
port 6 nsew default input
rlabel metal2 s 2410 0 2466 480 6 bottom_left_grid_pin_47_
port 7 nsew default input
rlabel metal2 s 2870 0 2926 480 6 bottom_left_grid_pin_48_
port 8 nsew default input
rlabel metal2 s 3330 0 3386 480 6 bottom_left_grid_pin_49_
port 9 nsew default input
rlabel metal2 s 5722 22320 5778 22800 6 ccff_head
port 10 nsew default input
rlabel metal2 s 17130 22320 17186 22800 6 ccff_tail
port 11 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_in[0]
port 12 nsew default input
rlabel metal3 s 0 8440 480 8560 6 chanx_left_in[10]
port 13 nsew default input
rlabel metal3 s 0 8984 480 9104 6 chanx_left_in[11]
port 14 nsew default input
rlabel metal3 s 0 9392 480 9512 6 chanx_left_in[12]
port 15 nsew default input
rlabel metal3 s 0 9936 480 10056 6 chanx_left_in[13]
port 16 nsew default input
rlabel metal3 s 0 10344 480 10464 6 chanx_left_in[14]
port 17 nsew default input
rlabel metal3 s 0 10752 480 10872 6 chanx_left_in[15]
port 18 nsew default input
rlabel metal3 s 0 11296 480 11416 6 chanx_left_in[16]
port 19 nsew default input
rlabel metal3 s 0 11704 480 11824 6 chanx_left_in[17]
port 20 nsew default input
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[18]
port 21 nsew default input
rlabel metal3 s 0 12656 480 12776 6 chanx_left_in[19]
port 22 nsew default input
rlabel metal3 s 0 4224 480 4344 6 chanx_left_in[1]
port 23 nsew default input
rlabel metal3 s 0 4768 480 4888 6 chanx_left_in[2]
port 24 nsew default input
rlabel metal3 s 0 5176 480 5296 6 chanx_left_in[3]
port 25 nsew default input
rlabel metal3 s 0 5720 480 5840 6 chanx_left_in[4]
port 26 nsew default input
rlabel metal3 s 0 6128 480 6248 6 chanx_left_in[5]
port 27 nsew default input
rlabel metal3 s 0 6672 480 6792 6 chanx_left_in[6]
port 28 nsew default input
rlabel metal3 s 0 7080 480 7200 6 chanx_left_in[7]
port 29 nsew default input
rlabel metal3 s 0 7488 480 7608 6 chanx_left_in[8]
port 30 nsew default input
rlabel metal3 s 0 8032 480 8152 6 chanx_left_in[9]
port 31 nsew default input
rlabel metal3 s 0 13200 480 13320 6 chanx_left_out[0]
port 32 nsew default tristate
rlabel metal3 s 0 17824 480 17944 6 chanx_left_out[10]
port 33 nsew default tristate
rlabel metal3 s 0 18232 480 18352 6 chanx_left_out[11]
port 34 nsew default tristate
rlabel metal3 s 0 18776 480 18896 6 chanx_left_out[12]
port 35 nsew default tristate
rlabel metal3 s 0 19184 480 19304 6 chanx_left_out[13]
port 36 nsew default tristate
rlabel metal3 s 0 19728 480 19848 6 chanx_left_out[14]
port 37 nsew default tristate
rlabel metal3 s 0 20136 480 20256 6 chanx_left_out[15]
port 38 nsew default tristate
rlabel metal3 s 0 20544 480 20664 6 chanx_left_out[16]
port 39 nsew default tristate
rlabel metal3 s 0 21088 480 21208 6 chanx_left_out[17]
port 40 nsew default tristate
rlabel metal3 s 0 21496 480 21616 6 chanx_left_out[18]
port 41 nsew default tristate
rlabel metal3 s 0 22040 480 22160 6 chanx_left_out[19]
port 42 nsew default tristate
rlabel metal3 s 0 13608 480 13728 6 chanx_left_out[1]
port 43 nsew default tristate
rlabel metal3 s 0 14016 480 14136 6 chanx_left_out[2]
port 44 nsew default tristate
rlabel metal3 s 0 14560 480 14680 6 chanx_left_out[3]
port 45 nsew default tristate
rlabel metal3 s 0 14968 480 15088 6 chanx_left_out[4]
port 46 nsew default tristate
rlabel metal3 s 0 15512 480 15632 6 chanx_left_out[5]
port 47 nsew default tristate
rlabel metal3 s 0 15920 480 16040 6 chanx_left_out[6]
port 48 nsew default tristate
rlabel metal3 s 0 16464 480 16584 6 chanx_left_out[7]
port 49 nsew default tristate
rlabel metal3 s 0 16872 480 16992 6 chanx_left_out[8]
port 50 nsew default tristate
rlabel metal3 s 0 17280 480 17400 6 chanx_left_out[9]
port 51 nsew default tristate
rlabel metal3 s 22320 3816 22800 3936 6 chanx_right_in[0]
port 52 nsew default input
rlabel metal3 s 22320 8440 22800 8560 6 chanx_right_in[10]
port 53 nsew default input
rlabel metal3 s 22320 8984 22800 9104 6 chanx_right_in[11]
port 54 nsew default input
rlabel metal3 s 22320 9392 22800 9512 6 chanx_right_in[12]
port 55 nsew default input
rlabel metal3 s 22320 9936 22800 10056 6 chanx_right_in[13]
port 56 nsew default input
rlabel metal3 s 22320 10344 22800 10464 6 chanx_right_in[14]
port 57 nsew default input
rlabel metal3 s 22320 10752 22800 10872 6 chanx_right_in[15]
port 58 nsew default input
rlabel metal3 s 22320 11296 22800 11416 6 chanx_right_in[16]
port 59 nsew default input
rlabel metal3 s 22320 11704 22800 11824 6 chanx_right_in[17]
port 60 nsew default input
rlabel metal3 s 22320 12248 22800 12368 6 chanx_right_in[18]
port 61 nsew default input
rlabel metal3 s 22320 12656 22800 12776 6 chanx_right_in[19]
port 62 nsew default input
rlabel metal3 s 22320 4224 22800 4344 6 chanx_right_in[1]
port 63 nsew default input
rlabel metal3 s 22320 4768 22800 4888 6 chanx_right_in[2]
port 64 nsew default input
rlabel metal3 s 22320 5176 22800 5296 6 chanx_right_in[3]
port 65 nsew default input
rlabel metal3 s 22320 5720 22800 5840 6 chanx_right_in[4]
port 66 nsew default input
rlabel metal3 s 22320 6128 22800 6248 6 chanx_right_in[5]
port 67 nsew default input
rlabel metal3 s 22320 6672 22800 6792 6 chanx_right_in[6]
port 68 nsew default input
rlabel metal3 s 22320 7080 22800 7200 6 chanx_right_in[7]
port 69 nsew default input
rlabel metal3 s 22320 7488 22800 7608 6 chanx_right_in[8]
port 70 nsew default input
rlabel metal3 s 22320 8032 22800 8152 6 chanx_right_in[9]
port 71 nsew default input
rlabel metal3 s 22320 13200 22800 13320 6 chanx_right_out[0]
port 72 nsew default tristate
rlabel metal3 s 22320 17824 22800 17944 6 chanx_right_out[10]
port 73 nsew default tristate
rlabel metal3 s 22320 18232 22800 18352 6 chanx_right_out[11]
port 74 nsew default tristate
rlabel metal3 s 22320 18776 22800 18896 6 chanx_right_out[12]
port 75 nsew default tristate
rlabel metal3 s 22320 19184 22800 19304 6 chanx_right_out[13]
port 76 nsew default tristate
rlabel metal3 s 22320 19728 22800 19848 6 chanx_right_out[14]
port 77 nsew default tristate
rlabel metal3 s 22320 20136 22800 20256 6 chanx_right_out[15]
port 78 nsew default tristate
rlabel metal3 s 22320 20544 22800 20664 6 chanx_right_out[16]
port 79 nsew default tristate
rlabel metal3 s 22320 21088 22800 21208 6 chanx_right_out[17]
port 80 nsew default tristate
rlabel metal3 s 22320 21496 22800 21616 6 chanx_right_out[18]
port 81 nsew default tristate
rlabel metal3 s 22320 22040 22800 22160 6 chanx_right_out[19]
port 82 nsew default tristate
rlabel metal3 s 22320 13608 22800 13728 6 chanx_right_out[1]
port 83 nsew default tristate
rlabel metal3 s 22320 14016 22800 14136 6 chanx_right_out[2]
port 84 nsew default tristate
rlabel metal3 s 22320 14560 22800 14680 6 chanx_right_out[3]
port 85 nsew default tristate
rlabel metal3 s 22320 14968 22800 15088 6 chanx_right_out[4]
port 86 nsew default tristate
rlabel metal3 s 22320 15512 22800 15632 6 chanx_right_out[5]
port 87 nsew default tristate
rlabel metal3 s 22320 15920 22800 16040 6 chanx_right_out[6]
port 88 nsew default tristate
rlabel metal3 s 22320 16464 22800 16584 6 chanx_right_out[7]
port 89 nsew default tristate
rlabel metal3 s 22320 16872 22800 16992 6 chanx_right_out[8]
port 90 nsew default tristate
rlabel metal3 s 22320 17280 22800 17400 6 chanx_right_out[9]
port 91 nsew default tristate
rlabel metal2 s 3698 0 3754 480 6 chany_bottom_in[0]
port 92 nsew default input
rlabel metal2 s 8206 0 8262 480 6 chany_bottom_in[10]
port 93 nsew default input
rlabel metal2 s 8666 0 8722 480 6 chany_bottom_in[11]
port 94 nsew default input
rlabel metal2 s 9126 0 9182 480 6 chany_bottom_in[12]
port 95 nsew default input
rlabel metal2 s 9586 0 9642 480 6 chany_bottom_in[13]
port 96 nsew default input
rlabel metal2 s 9954 0 10010 480 6 chany_bottom_in[14]
port 97 nsew default input
rlabel metal2 s 10414 0 10470 480 6 chany_bottom_in[15]
port 98 nsew default input
rlabel metal2 s 10874 0 10930 480 6 chany_bottom_in[16]
port 99 nsew default input
rlabel metal2 s 11334 0 11390 480 6 chany_bottom_in[17]
port 100 nsew default input
rlabel metal2 s 11794 0 11850 480 6 chany_bottom_in[18]
port 101 nsew default input
rlabel metal2 s 12254 0 12310 480 6 chany_bottom_in[19]
port 102 nsew default input
rlabel metal2 s 4158 0 4214 480 6 chany_bottom_in[1]
port 103 nsew default input
rlabel metal2 s 4618 0 4674 480 6 chany_bottom_in[2]
port 104 nsew default input
rlabel metal2 s 5078 0 5134 480 6 chany_bottom_in[3]
port 105 nsew default input
rlabel metal2 s 5538 0 5594 480 6 chany_bottom_in[4]
port 106 nsew default input
rlabel metal2 s 5998 0 6054 480 6 chany_bottom_in[5]
port 107 nsew default input
rlabel metal2 s 6458 0 6514 480 6 chany_bottom_in[6]
port 108 nsew default input
rlabel metal2 s 6826 0 6882 480 6 chany_bottom_in[7]
port 109 nsew default input
rlabel metal2 s 7286 0 7342 480 6 chany_bottom_in[8]
port 110 nsew default input
rlabel metal2 s 7746 0 7802 480 6 chany_bottom_in[9]
port 111 nsew default input
rlabel metal2 s 12714 0 12770 480 6 chany_bottom_out[0]
port 112 nsew default tristate
rlabel metal2 s 17130 0 17186 480 6 chany_bottom_out[10]
port 113 nsew default tristate
rlabel metal2 s 17590 0 17646 480 6 chany_bottom_out[11]
port 114 nsew default tristate
rlabel metal2 s 18050 0 18106 480 6 chany_bottom_out[12]
port 115 nsew default tristate
rlabel metal2 s 18510 0 18566 480 6 chany_bottom_out[13]
port 116 nsew default tristate
rlabel metal2 s 18970 0 19026 480 6 chany_bottom_out[14]
port 117 nsew default tristate
rlabel metal2 s 19430 0 19486 480 6 chany_bottom_out[15]
port 118 nsew default tristate
rlabel metal2 s 19798 0 19854 480 6 chany_bottom_out[16]
port 119 nsew default tristate
rlabel metal2 s 20258 0 20314 480 6 chany_bottom_out[17]
port 120 nsew default tristate
rlabel metal2 s 20718 0 20774 480 6 chany_bottom_out[18]
port 121 nsew default tristate
rlabel metal2 s 21178 0 21234 480 6 chany_bottom_out[19]
port 122 nsew default tristate
rlabel metal2 s 13174 0 13230 480 6 chany_bottom_out[1]
port 123 nsew default tristate
rlabel metal2 s 13542 0 13598 480 6 chany_bottom_out[2]
port 124 nsew default tristate
rlabel metal2 s 14002 0 14058 480 6 chany_bottom_out[3]
port 125 nsew default tristate
rlabel metal2 s 14462 0 14518 480 6 chany_bottom_out[4]
port 126 nsew default tristate
rlabel metal2 s 14922 0 14978 480 6 chany_bottom_out[5]
port 127 nsew default tristate
rlabel metal2 s 15382 0 15438 480 6 chany_bottom_out[6]
port 128 nsew default tristate
rlabel metal2 s 15842 0 15898 480 6 chany_bottom_out[7]
port 129 nsew default tristate
rlabel metal2 s 16302 0 16358 480 6 chany_bottom_out[8]
port 130 nsew default tristate
rlabel metal2 s 16670 0 16726 480 6 chany_bottom_out[9]
port 131 nsew default tristate
rlabel metal3 s 0 144 480 264 6 left_bottom_grid_pin_34_
port 132 nsew default input
rlabel metal3 s 0 552 480 672 6 left_bottom_grid_pin_35_
port 133 nsew default input
rlabel metal3 s 0 960 480 1080 6 left_bottom_grid_pin_36_
port 134 nsew default input
rlabel metal3 s 0 1504 480 1624 6 left_bottom_grid_pin_37_
port 135 nsew default input
rlabel metal3 s 0 1912 480 2032 6 left_bottom_grid_pin_38_
port 136 nsew default input
rlabel metal3 s 0 2456 480 2576 6 left_bottom_grid_pin_39_
port 137 nsew default input
rlabel metal3 s 0 2864 480 2984 6 left_bottom_grid_pin_40_
port 138 nsew default input
rlabel metal3 s 0 3408 480 3528 6 left_bottom_grid_pin_41_
port 139 nsew default input
rlabel metal3 s 0 22448 480 22568 6 left_top_grid_pin_1_
port 140 nsew default input
rlabel metal2 s 22558 0 22614 480 6 prog_clk_0_S_in
port 141 nsew default input
rlabel metal3 s 22320 144 22800 264 6 right_bottom_grid_pin_34_
port 142 nsew default input
rlabel metal3 s 22320 552 22800 672 6 right_bottom_grid_pin_35_
port 143 nsew default input
rlabel metal3 s 22320 960 22800 1080 6 right_bottom_grid_pin_36_
port 144 nsew default input
rlabel metal3 s 22320 1504 22800 1624 6 right_bottom_grid_pin_37_
port 145 nsew default input
rlabel metal3 s 22320 1912 22800 2032 6 right_bottom_grid_pin_38_
port 146 nsew default input
rlabel metal3 s 22320 2456 22800 2576 6 right_bottom_grid_pin_39_
port 147 nsew default input
rlabel metal3 s 22320 2864 22800 2984 6 right_bottom_grid_pin_40_
port 148 nsew default input
rlabel metal3 s 22320 3408 22800 3528 6 right_bottom_grid_pin_41_
port 149 nsew default input
rlabel metal3 s 22320 22448 22800 22568 6 right_top_grid_pin_1_
port 150 nsew default input
rlabel metal4 s 4376 2128 4696 20176 6 VPWR
port 151 nsew default input
rlabel metal4 s 7808 2128 8128 20176 6 VGND
port 152 nsew default input
<< properties >>
string FIXED_BBOX 0 0 22800 22800
<< end >>
