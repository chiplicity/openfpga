magic
tech sky130A
magscale 1 2
timestamp 1606228978
<< locali >>
rect 16497 22049 16681 22083
rect 16497 22015 16531 22049
rect 4905 21335 4939 21641
rect 8401 21335 8435 21437
rect 6469 20791 6503 21029
rect 20729 20927 20763 21029
rect 15669 19363 15703 19465
rect 8677 17527 8711 17629
rect 12265 17119 12299 17221
rect 14013 17119 14047 17221
rect 12265 17085 12357 17119
rect 13955 17085 14047 17119
rect 7665 15895 7699 16201
rect 7021 15555 7055 15657
rect 17877 14467 17911 14569
rect 20453 13855 20487 14025
rect 11621 13379 11655 13481
rect 9781 12087 9815 12189
rect 4445 10455 4479 10761
rect 8953 10455 8987 10557
rect 12909 10455 12943 10557
rect 5733 10115 5767 10217
rect 5825 10047 5859 10217
rect 8125 9367 8159 9469
rect 9413 9027 9447 9129
rect 10241 8279 10275 8381
rect 12265 8279 12299 8585
rect 11713 7803 11747 8041
rect 13369 7803 13403 7973
rect 15301 7735 15335 7905
rect 16037 7327 16071 7429
rect 16129 7327 16163 7497
rect 20637 6647 20671 6817
rect 13093 4675 13127 4777
rect 11989 4471 12023 4641
rect 19533 4471 19567 4573
rect 20085 3043 20119 3145
rect 20177 2975 20211 3077
rect 15209 2295 15243 2601
<< viali >>
rect 16681 22049 16715 22083
rect 16497 21981 16531 22015
rect 1593 21641 1627 21675
rect 4905 21641 4939 21675
rect 2605 21505 2639 21539
rect 3433 21505 3467 21539
rect 3525 21505 3559 21539
rect 4629 21505 4663 21539
rect 1409 21437 1443 21471
rect 4537 21437 4571 21471
rect 2329 21369 2363 21403
rect 6285 21573 6319 21607
rect 14841 21573 14875 21607
rect 17877 21573 17911 21607
rect 5641 21505 5675 21539
rect 6929 21505 6963 21539
rect 9137 21505 9171 21539
rect 11897 21505 11931 21539
rect 11989 21505 12023 21539
rect 13461 21505 13495 21539
rect 16037 21505 16071 21539
rect 16957 21505 16991 21539
rect 17049 21505 17083 21539
rect 18797 21505 18831 21539
rect 18981 21505 19015 21539
rect 20269 21505 20303 21539
rect 21741 21505 21775 21539
rect 6101 21437 6135 21471
rect 8401 21437 8435 21471
rect 8953 21437 8987 21471
rect 9781 21437 9815 21471
rect 12633 21437 12667 21471
rect 15853 21437 15887 21471
rect 17693 21437 17727 21471
rect 21649 21437 21683 21471
rect 5457 21369 5491 21403
rect 7196 21369 7230 21403
rect 10026 21369 10060 21403
rect 13728 21369 13762 21403
rect 18705 21369 18739 21403
rect 20085 21369 20119 21403
rect 21557 21369 21591 21403
rect 22017 21369 22051 21403
rect 1961 21301 1995 21335
rect 2421 21301 2455 21335
rect 2973 21301 3007 21335
rect 3341 21301 3375 21335
rect 4077 21301 4111 21335
rect 4445 21301 4479 21335
rect 4905 21301 4939 21335
rect 5089 21301 5123 21335
rect 5549 21301 5583 21335
rect 8309 21301 8343 21335
rect 8401 21301 8435 21335
rect 8585 21301 8619 21335
rect 9045 21301 9079 21335
rect 11161 21301 11195 21335
rect 11437 21301 11471 21335
rect 11805 21301 11839 21335
rect 12817 21301 12851 21335
rect 15485 21301 15519 21335
rect 15945 21301 15979 21335
rect 16497 21301 16531 21335
rect 16865 21301 16899 21335
rect 18337 21301 18371 21335
rect 19717 21301 19751 21335
rect 20177 21301 20211 21335
rect 21189 21301 21223 21335
rect 3525 21097 3559 21131
rect 7113 21097 7147 21131
rect 14841 21097 14875 21131
rect 15485 21097 15519 21131
rect 17233 21097 17267 21131
rect 2412 21029 2446 21063
rect 6469 21029 6503 21063
rect 13176 21029 13210 21063
rect 20729 21029 20763 21063
rect 1593 20961 1627 20995
rect 4077 20961 4111 20995
rect 5264 20961 5298 20995
rect 2145 20893 2179 20927
rect 4997 20893 5031 20927
rect 7021 20961 7055 20995
rect 8197 20961 8231 20995
rect 10425 20961 10459 20995
rect 11336 20961 11370 20995
rect 14657 20961 14691 20995
rect 15301 20961 15335 20995
rect 16120 20961 16154 20995
rect 17776 20961 17810 20995
rect 19432 20961 19466 20995
rect 21281 20961 21315 20995
rect 21925 20961 21959 20995
rect 7205 20893 7239 20927
rect 7941 20893 7975 20927
rect 10517 20893 10551 20927
rect 10701 20893 10735 20927
rect 11069 20893 11103 20927
rect 12909 20893 12943 20927
rect 15853 20893 15887 20927
rect 17509 20893 17543 20927
rect 19165 20893 19199 20927
rect 20729 20893 20763 20927
rect 21373 20893 21407 20927
rect 21465 20893 21499 20927
rect 1777 20757 1811 20791
rect 4261 20757 4295 20791
rect 6377 20757 6411 20791
rect 6469 20757 6503 20791
rect 6653 20757 6687 20791
rect 9321 20757 9355 20791
rect 10057 20757 10091 20791
rect 12449 20757 12483 20791
rect 14289 20757 14323 20791
rect 18889 20757 18923 20791
rect 20545 20757 20579 20791
rect 20913 20757 20947 20791
rect 22109 20757 22143 20791
rect 2789 20553 2823 20587
rect 8217 20553 8251 20587
rect 12081 20553 12115 20587
rect 13829 20553 13863 20587
rect 20913 20553 20947 20587
rect 16313 20485 16347 20519
rect 6837 20417 6871 20451
rect 10241 20417 10275 20451
rect 17049 20417 17083 20451
rect 17233 20417 17267 20451
rect 19073 20417 19107 20451
rect 19533 20417 19567 20451
rect 21741 20417 21775 20451
rect 1409 20349 1443 20383
rect 3157 20349 3191 20383
rect 4813 20349 4847 20383
rect 5080 20349 5114 20383
rect 7104 20349 7138 20383
rect 8585 20349 8619 20383
rect 10701 20349 10735 20383
rect 12449 20349 12483 20383
rect 14381 20349 14415 20383
rect 14933 20349 14967 20383
rect 15200 20349 15234 20383
rect 16957 20349 16991 20383
rect 18061 20349 18095 20383
rect 18889 20349 18923 20383
rect 19800 20349 19834 20383
rect 1676 20281 1710 20315
rect 3424 20281 3458 20315
rect 8852 20281 8886 20315
rect 10968 20281 11002 20315
rect 12716 20281 12750 20315
rect 4537 20213 4571 20247
rect 6193 20213 6227 20247
rect 9965 20213 9999 20247
rect 14565 20213 14599 20247
rect 16589 20213 16623 20247
rect 18521 20213 18555 20247
rect 18981 20213 19015 20247
rect 21189 20213 21223 20247
rect 21557 20213 21591 20247
rect 21649 20213 21683 20247
rect 2421 20009 2455 20043
rect 3617 20009 3651 20043
rect 4077 20009 4111 20043
rect 5549 20009 5583 20043
rect 8493 20009 8527 20043
rect 10149 20009 10183 20043
rect 13001 20009 13035 20043
rect 14933 20009 14967 20043
rect 15301 20009 15335 20043
rect 15761 20009 15795 20043
rect 16681 20009 16715 20043
rect 18337 20009 18371 20043
rect 18797 20009 18831 20043
rect 20545 20009 20579 20043
rect 2789 19941 2823 19975
rect 16313 19941 16347 19975
rect 17224 19941 17258 19975
rect 21158 19941 21192 19975
rect 1777 19873 1811 19907
rect 2881 19873 2915 19907
rect 3433 19873 3467 19907
rect 4445 19873 4479 19907
rect 5457 19873 5491 19907
rect 8861 19873 8895 19907
rect 10057 19873 10091 19907
rect 12817 19873 12851 19907
rect 13820 19873 13854 19907
rect 15669 19873 15703 19907
rect 16129 19873 16163 19907
rect 16497 19873 16531 19907
rect 18613 19873 18647 19907
rect 19165 19873 19199 19907
rect 19432 19873 19466 19907
rect 1869 19805 1903 19839
rect 1961 19805 1995 19839
rect 2973 19805 3007 19839
rect 4537 19805 4571 19839
rect 4629 19805 4663 19839
rect 5641 19805 5675 19839
rect 6377 19805 6411 19839
rect 6700 19805 6734 19839
rect 6883 19805 6917 19839
rect 7113 19805 7147 19839
rect 8953 19805 8987 19839
rect 9045 19805 9079 19839
rect 10333 19805 10367 19839
rect 10701 19805 10735 19839
rect 11024 19805 11058 19839
rect 11207 19805 11241 19839
rect 11437 19805 11471 19839
rect 13553 19805 13587 19839
rect 15853 19805 15887 19839
rect 16957 19805 16991 19839
rect 20913 19805 20947 19839
rect 1409 19737 1443 19771
rect 5089 19669 5123 19703
rect 8217 19669 8251 19703
rect 9689 19669 9723 19703
rect 12541 19669 12575 19703
rect 22293 19669 22327 19703
rect 2789 19465 2823 19499
rect 6285 19465 6319 19499
rect 15669 19465 15703 19499
rect 20821 19465 20855 19499
rect 12081 19397 12115 19431
rect 18061 19397 18095 19431
rect 3709 19329 3743 19363
rect 4951 19329 4985 19363
rect 7481 19329 7515 19363
rect 8723 19329 8757 19363
rect 13093 19329 13127 19363
rect 15669 19329 15703 19363
rect 16405 19329 16439 19363
rect 17601 19329 17635 19363
rect 18521 19329 18555 19363
rect 18613 19329 18647 19363
rect 21465 19329 21499 19363
rect 1409 19261 1443 19295
rect 3525 19261 3559 19295
rect 4445 19261 4479 19295
rect 5181 19261 5215 19295
rect 8217 19261 8251 19295
rect 8953 19261 8987 19295
rect 10517 19261 10551 19295
rect 10701 19261 10735 19295
rect 10968 19261 11002 19295
rect 13461 19261 13495 19295
rect 14197 19261 14231 19295
rect 16221 19261 16255 19295
rect 17325 19261 17359 19295
rect 18429 19261 18463 19295
rect 19441 19261 19475 19295
rect 1676 19193 1710 19227
rect 7205 19193 7239 19227
rect 13645 19193 13679 19227
rect 14464 19193 14498 19227
rect 17417 19193 17451 19227
rect 19708 19193 19742 19227
rect 21281 19193 21315 19227
rect 3065 19125 3099 19159
rect 3433 19125 3467 19159
rect 4911 19125 4945 19159
rect 6837 19125 6871 19159
rect 7297 19125 7331 19159
rect 8683 19125 8717 19159
rect 10057 19125 10091 19159
rect 10333 19125 10367 19159
rect 12449 19125 12483 19159
rect 12817 19125 12851 19159
rect 12909 19125 12943 19159
rect 13829 19125 13863 19159
rect 15577 19125 15611 19159
rect 15853 19125 15887 19159
rect 16313 19125 16347 19159
rect 16957 19125 16991 19159
rect 20913 19125 20947 19159
rect 21373 19125 21407 19159
rect 21925 19125 21959 19159
rect 22109 19125 22143 19159
rect 1593 18921 1627 18955
rect 3341 18921 3375 18955
rect 4261 18921 4295 18955
rect 5917 18921 5951 18955
rect 7849 18921 7883 18955
rect 8309 18921 8343 18955
rect 9045 18921 9079 18955
rect 10057 18921 10091 18955
rect 17141 18921 17175 18955
rect 18889 18921 18923 18955
rect 20545 18921 20579 18955
rect 2206 18853 2240 18887
rect 5273 18853 5307 18887
rect 6460 18853 6494 18887
rect 15568 18853 15602 18887
rect 17776 18853 17810 18887
rect 19432 18853 19466 18887
rect 1409 18785 1443 18819
rect 4077 18785 4111 18819
rect 6101 18785 6135 18819
rect 6193 18785 6227 18819
rect 8217 18785 8251 18819
rect 8861 18785 8895 18819
rect 10425 18785 10459 18819
rect 11069 18785 11103 18819
rect 11989 18785 12023 18819
rect 12081 18785 12115 18819
rect 12633 18785 12667 18819
rect 12900 18785 12934 18819
rect 14289 18785 14323 18819
rect 16957 18785 16991 18819
rect 21281 18785 21315 18819
rect 1961 18717 1995 18751
rect 5365 18717 5399 18751
rect 5457 18717 5491 18751
rect 8401 18717 8435 18751
rect 10517 18717 10551 18751
rect 10609 18717 10643 18751
rect 12173 18717 12207 18751
rect 15301 18717 15335 18751
rect 17509 18717 17543 18751
rect 19165 18717 19199 18751
rect 21373 18717 21407 18751
rect 21465 18717 21499 18751
rect 22109 18717 22143 18751
rect 4905 18649 4939 18683
rect 11621 18649 11655 18683
rect 14473 18649 14507 18683
rect 7573 18581 7607 18615
rect 11253 18581 11287 18615
rect 14013 18581 14047 18615
rect 16681 18581 16715 18615
rect 20913 18581 20947 18615
rect 21925 18581 21959 18615
rect 2973 18377 3007 18411
rect 3617 18377 3651 18411
rect 6469 18377 6503 18411
rect 10149 18377 10183 18411
rect 13829 18377 13863 18411
rect 14289 18377 14323 18411
rect 18337 18377 18371 18411
rect 20085 18377 20119 18411
rect 4721 18241 4755 18275
rect 6837 18241 6871 18275
rect 10793 18241 10827 18275
rect 11989 18241 12023 18275
rect 12449 18241 12483 18275
rect 17141 18241 17175 18275
rect 17233 18241 17267 18275
rect 21005 18241 21039 18275
rect 21925 18241 21959 18275
rect 1593 18173 1627 18207
rect 1860 18173 1894 18207
rect 3433 18173 3467 18207
rect 4537 18173 4571 18207
rect 5089 18173 5123 18207
rect 7104 18173 7138 18207
rect 8493 18173 8527 18207
rect 11713 18173 11747 18207
rect 14105 18173 14139 18207
rect 14841 18173 14875 18207
rect 14933 18173 14967 18207
rect 17049 18173 17083 18207
rect 18153 18173 18187 18207
rect 18705 18173 18739 18207
rect 3249 18105 3283 18139
rect 5356 18105 5390 18139
rect 8760 18105 8794 18139
rect 10517 18105 10551 18139
rect 12716 18105 12750 18139
rect 15200 18105 15234 18139
rect 18950 18105 18984 18139
rect 21833 18105 21867 18139
rect 4077 18037 4111 18071
rect 4445 18037 4479 18071
rect 8217 18037 8251 18071
rect 9873 18037 9907 18071
rect 10609 18037 10643 18071
rect 11345 18037 11379 18071
rect 11805 18037 11839 18071
rect 14657 18037 14691 18071
rect 16313 18037 16347 18071
rect 16681 18037 16715 18071
rect 20361 18037 20395 18071
rect 20729 18037 20763 18071
rect 20821 18037 20855 18071
rect 21373 18037 21407 18071
rect 21741 18037 21775 18071
rect 2973 17833 3007 17867
rect 3433 17833 3467 17867
rect 5733 17833 5767 17867
rect 6193 17833 6227 17867
rect 9045 17833 9079 17867
rect 9689 17833 9723 17867
rect 11805 17833 11839 17867
rect 13829 17833 13863 17867
rect 14105 17833 14139 17867
rect 15761 17833 15795 17867
rect 16497 17833 16531 17867
rect 19901 17833 19935 17867
rect 21281 17833 21315 17867
rect 22109 17833 22143 17867
rect 15669 17765 15703 17799
rect 17110 17765 17144 17799
rect 18788 17765 18822 17799
rect 1860 17697 1894 17731
rect 3249 17697 3283 17731
rect 4353 17697 4387 17731
rect 4620 17697 4654 17731
rect 6009 17697 6043 17731
rect 6745 17697 6779 17731
rect 7068 17697 7102 17731
rect 8861 17697 8895 17731
rect 10057 17697 10091 17731
rect 10701 17697 10735 17731
rect 11897 17697 11931 17731
rect 12716 17697 12750 17731
rect 14473 17697 14507 17731
rect 16313 17697 16347 17731
rect 20177 17697 20211 17731
rect 21373 17697 21407 17731
rect 21925 17697 21959 17731
rect 1593 17629 1627 17663
rect 7208 17629 7242 17663
rect 7481 17629 7515 17663
rect 8677 17629 8711 17663
rect 10149 17629 10183 17663
rect 10333 17629 10367 17663
rect 11989 17629 12023 17663
rect 12449 17629 12483 17663
rect 14565 17629 14599 17663
rect 14749 17629 14783 17663
rect 15853 17629 15887 17663
rect 16865 17629 16899 17663
rect 18521 17629 18555 17663
rect 21465 17629 21499 17663
rect 10885 17561 10919 17595
rect 11437 17561 11471 17595
rect 20913 17561 20947 17595
rect 8585 17493 8619 17527
rect 8677 17493 8711 17527
rect 15301 17493 15335 17527
rect 18245 17493 18279 17527
rect 20361 17493 20395 17527
rect 1869 17289 1903 17323
rect 3617 17289 3651 17323
rect 10517 17289 10551 17323
rect 11345 17289 11379 17323
rect 13829 17289 13863 17323
rect 21465 17289 21499 17323
rect 6469 17221 6503 17255
rect 10977 17221 11011 17255
rect 12265 17221 12299 17255
rect 5092 17153 5126 17187
rect 9144 17153 9178 17187
rect 11897 17153 11931 17187
rect 14013 17221 14047 17255
rect 14105 17221 14139 17255
rect 18797 17221 18831 17255
rect 19257 17153 19291 17187
rect 19441 17153 19475 17187
rect 22017 17153 22051 17187
rect 1685 17085 1719 17119
rect 2237 17085 2271 17119
rect 2504 17085 2538 17119
rect 4077 17085 4111 17119
rect 4629 17085 4663 17119
rect 5365 17085 5399 17119
rect 6837 17085 6871 17119
rect 7481 17085 7515 17119
rect 7737 17085 7771 17119
rect 9404 17085 9438 17119
rect 10793 17085 10827 17119
rect 12357 17085 12391 17119
rect 12449 17085 12483 17119
rect 13921 17085 13955 17119
rect 14289 17085 14323 17119
rect 14381 17085 14415 17119
rect 16037 17085 16071 17119
rect 17877 17085 17911 17119
rect 18245 17085 18279 17119
rect 19809 17085 19843 17119
rect 21925 17085 21959 17119
rect 11713 17017 11747 17051
rect 12716 17017 12750 17051
rect 14648 17017 14682 17051
rect 16304 17017 16338 17051
rect 19165 17017 19199 17051
rect 20076 17017 20110 17051
rect 4261 16949 4295 16983
rect 5095 16949 5129 16983
rect 7021 16949 7055 16983
rect 8861 16949 8895 16983
rect 11805 16949 11839 16983
rect 15761 16949 15795 16983
rect 17417 16949 17451 16983
rect 17693 16949 17727 16983
rect 18429 16949 18463 16983
rect 21189 16949 21223 16983
rect 21833 16949 21867 16983
rect 1777 16745 1811 16779
rect 4261 16745 4295 16779
rect 4629 16745 4663 16779
rect 4997 16745 5031 16779
rect 5641 16745 5675 16779
rect 8769 16745 8803 16779
rect 9321 16745 9355 16779
rect 11069 16745 11103 16779
rect 11805 16745 11839 16779
rect 18797 16745 18831 16779
rect 20545 16745 20579 16779
rect 2412 16677 2446 16711
rect 5089 16677 5123 16711
rect 6101 16677 6135 16711
rect 8677 16677 8711 16711
rect 9956 16677 9990 16711
rect 1593 16609 1627 16643
rect 2145 16609 2179 16643
rect 4077 16609 4111 16643
rect 6009 16609 6043 16643
rect 6653 16609 6687 16643
rect 6920 16609 6954 16643
rect 9505 16609 9539 16643
rect 9689 16609 9723 16643
rect 11713 16609 11747 16643
rect 12449 16609 12483 16643
rect 12716 16609 12750 16643
rect 14473 16609 14507 16643
rect 15301 16609 15335 16643
rect 16037 16609 16071 16643
rect 16865 16609 16899 16643
rect 18613 16609 18647 16643
rect 19432 16609 19466 16643
rect 20913 16609 20947 16643
rect 21180 16609 21214 16643
rect 5181 16541 5215 16575
rect 6193 16541 6227 16575
rect 8861 16541 8895 16575
rect 11897 16541 11931 16575
rect 14565 16541 14599 16575
rect 14749 16541 14783 16575
rect 16129 16541 16163 16575
rect 16452 16541 16486 16575
rect 16592 16541 16626 16575
rect 19165 16541 19199 16575
rect 3525 16473 3559 16507
rect 8033 16473 8067 16507
rect 8309 16473 8343 16507
rect 11345 16473 11379 16507
rect 13829 16473 13863 16507
rect 17969 16473 18003 16507
rect 14105 16405 14139 16439
rect 15485 16405 15519 16439
rect 15853 16405 15887 16439
rect 22293 16405 22327 16439
rect 3249 16201 3283 16235
rect 6009 16201 6043 16235
rect 7665 16201 7699 16235
rect 7849 16201 7883 16235
rect 10701 16201 10735 16235
rect 12081 16201 12115 16235
rect 13921 16201 13955 16235
rect 16129 16201 16163 16235
rect 16957 16201 16991 16235
rect 19993 16201 20027 16235
rect 1409 16065 1443 16099
rect 4169 16065 4203 16099
rect 6285 16065 6319 16099
rect 7389 16065 7423 16099
rect 1869 15997 1903 16031
rect 4629 15997 4663 16031
rect 7297 15997 7331 16031
rect 2136 15929 2170 15963
rect 3985 15929 4019 15963
rect 4896 15929 4930 15963
rect 10977 16133 11011 16167
rect 8493 16065 8527 16099
rect 11621 16065 11655 16099
rect 14752 16065 14786 16099
rect 17509 16065 17543 16099
rect 20821 16065 20855 16099
rect 8217 15997 8251 16031
rect 9321 15997 9355 16031
rect 9588 15997 9622 16031
rect 12265 15997 12299 16031
rect 12541 15997 12575 16031
rect 12808 15997 12842 16031
rect 14289 15997 14323 16031
rect 15025 15997 15059 16031
rect 16405 15997 16439 16031
rect 18061 15997 18095 16031
rect 18613 15997 18647 16031
rect 20269 15997 20303 16031
rect 21088 15997 21122 16031
rect 8309 15929 8343 15963
rect 18880 15929 18914 15963
rect 3617 15861 3651 15895
rect 4077 15861 4111 15895
rect 6837 15861 6871 15895
rect 7205 15861 7239 15895
rect 7665 15861 7699 15895
rect 8861 15861 8895 15895
rect 11345 15861 11379 15895
rect 11437 15861 11471 15895
rect 14755 15861 14789 15895
rect 16589 15861 16623 15895
rect 17325 15861 17359 15895
rect 17417 15861 17451 15895
rect 18245 15861 18279 15895
rect 20453 15861 20487 15895
rect 22201 15861 22235 15895
rect 3065 15657 3099 15691
rect 4261 15657 4295 15691
rect 6193 15657 6227 15691
rect 6837 15657 6871 15691
rect 7021 15657 7055 15691
rect 9229 15657 9263 15691
rect 11345 15657 11379 15691
rect 13921 15657 13955 15691
rect 18521 15657 18555 15691
rect 19257 15657 19291 15691
rect 20913 15657 20947 15691
rect 21373 15657 21407 15691
rect 9045 15589 9079 15623
rect 9956 15589 9990 15623
rect 12808 15589 12842 15623
rect 14565 15589 14599 15623
rect 21281 15589 21315 15623
rect 1685 15521 1719 15555
rect 1952 15521 1986 15555
rect 3433 15521 3467 15555
rect 4077 15521 4111 15555
rect 4813 15521 4847 15555
rect 5080 15521 5114 15555
rect 6653 15521 6687 15555
rect 7021 15521 7055 15555
rect 7472 15521 7506 15555
rect 8861 15521 8895 15555
rect 11713 15521 11747 15555
rect 14657 15521 14691 15555
rect 15568 15521 15602 15555
rect 17141 15521 17175 15555
rect 17408 15521 17442 15555
rect 19165 15521 19199 15555
rect 20177 15521 20211 15555
rect 21925 15521 21959 15555
rect 7205 15453 7239 15487
rect 9689 15453 9723 15487
rect 11805 15453 11839 15487
rect 11897 15453 11931 15487
rect 12541 15453 12575 15487
rect 14841 15453 14875 15487
rect 15301 15453 15335 15487
rect 19349 15453 19383 15487
rect 20269 15453 20303 15487
rect 20361 15453 20395 15487
rect 21465 15453 21499 15487
rect 22109 15385 22143 15419
rect 3617 15317 3651 15351
rect 8585 15317 8619 15351
rect 11069 15317 11103 15351
rect 14197 15317 14231 15351
rect 16681 15317 16715 15351
rect 18797 15317 18831 15351
rect 19809 15317 19843 15351
rect 5733 15113 5767 15147
rect 6377 15113 6411 15147
rect 8493 15113 8527 15147
rect 10701 15113 10735 15147
rect 11989 15113 12023 15147
rect 13829 15113 13863 15147
rect 14197 15113 14231 15147
rect 17693 15113 17727 15147
rect 19441 15113 19475 15147
rect 22293 15113 22327 15147
rect 3341 15045 3375 15079
rect 3893 14977 3927 15011
rect 7113 14977 7147 15011
rect 9321 14977 9355 15011
rect 11529 14977 11563 15011
rect 14473 14977 14507 15011
rect 16313 14977 16347 15011
rect 18061 14977 18095 15011
rect 20361 14977 20395 15011
rect 20545 14977 20579 15011
rect 1501 14909 1535 14943
rect 4353 14909 4387 14943
rect 6193 14909 6227 14943
rect 8769 14909 8803 14943
rect 9588 14909 9622 14943
rect 12173 14909 12207 14943
rect 12449 14909 12483 14943
rect 12716 14909 12750 14943
rect 14381 14909 14415 14943
rect 18328 14909 18362 14943
rect 20269 14909 20303 14943
rect 20913 14909 20947 14943
rect 21180 14909 21214 14943
rect 1768 14841 1802 14875
rect 4598 14841 4632 14875
rect 7358 14841 7392 14875
rect 11345 14841 11379 14875
rect 14740 14841 14774 14875
rect 16580 14841 16614 14875
rect 2881 14773 2915 14807
rect 3709 14773 3743 14807
rect 3801 14773 3835 14807
rect 8953 14773 8987 14807
rect 10977 14773 11011 14807
rect 11437 14773 11471 14807
rect 15853 14773 15887 14807
rect 19901 14773 19935 14807
rect 1961 14569 1995 14603
rect 5457 14569 5491 14603
rect 5825 14569 5859 14603
rect 6653 14569 6687 14603
rect 8125 14569 8159 14603
rect 12725 14569 12759 14603
rect 14381 14569 14415 14603
rect 15761 14569 15795 14603
rect 17785 14569 17819 14603
rect 17877 14569 17911 14603
rect 18061 14569 18095 14603
rect 19073 14569 19107 14603
rect 22293 14569 22327 14603
rect 4322 14501 4356 14535
rect 9956 14501 9990 14535
rect 11590 14501 11624 14535
rect 13246 14501 13280 14535
rect 18429 14501 18463 14535
rect 21158 14501 21192 14535
rect 2973 14433 3007 14467
rect 3893 14433 3927 14467
rect 6009 14433 6043 14467
rect 6101 14433 6135 14467
rect 7021 14433 7055 14467
rect 8033 14433 8067 14467
rect 8677 14433 8711 14467
rect 9413 14433 9447 14467
rect 9689 14433 9723 14467
rect 14657 14433 14691 14467
rect 15853 14433 15887 14467
rect 16405 14433 16439 14467
rect 16672 14433 16706 14467
rect 17877 14433 17911 14467
rect 18521 14433 18555 14467
rect 19441 14433 19475 14467
rect 20269 14433 20303 14467
rect 20913 14433 20947 14467
rect 2053 14365 2087 14399
rect 2237 14365 2271 14399
rect 3065 14365 3099 14399
rect 3249 14365 3283 14399
rect 4077 14365 4111 14399
rect 7113 14365 7147 14399
rect 7297 14365 7331 14399
rect 8217 14365 8251 14399
rect 11345 14365 11379 14399
rect 13001 14365 13035 14399
rect 16037 14365 16071 14399
rect 18705 14365 18739 14399
rect 19533 14365 19567 14399
rect 19625 14365 19659 14399
rect 9229 14297 9263 14331
rect 14841 14297 14875 14331
rect 20453 14297 20487 14331
rect 1593 14229 1627 14263
rect 2605 14229 2639 14263
rect 3709 14229 3743 14263
rect 6285 14229 6319 14263
rect 7665 14229 7699 14263
rect 8861 14229 8895 14263
rect 11069 14229 11103 14263
rect 15393 14229 15427 14263
rect 1869 14025 1903 14059
rect 4629 14025 4663 14059
rect 6285 14025 6319 14059
rect 9229 14025 9263 14059
rect 9505 14025 9539 14059
rect 11253 14025 11287 14059
rect 12633 14025 12667 14059
rect 16957 14025 16991 14059
rect 19441 14025 19475 14059
rect 20269 14025 20303 14059
rect 20453 14025 20487 14059
rect 21925 14025 21959 14059
rect 2237 13957 2271 13991
rect 11897 13957 11931 13991
rect 14565 13957 14599 13991
rect 2789 13889 2823 13923
rect 4905 13889 4939 13923
rect 7297 13889 7331 13923
rect 7481 13889 7515 13923
rect 7849 13889 7883 13923
rect 9873 13889 9907 13923
rect 17601 13889 17635 13923
rect 1685 13821 1719 13855
rect 3249 13821 3283 13855
rect 3516 13821 3550 13855
rect 5161 13821 5195 13855
rect 8105 13821 8139 13855
rect 9689 13821 9723 13855
rect 10140 13821 10174 13855
rect 11713 13821 11747 13855
rect 12449 13821 12483 13855
rect 13185 13821 13219 13855
rect 13441 13821 13475 13855
rect 14841 13821 14875 13855
rect 15108 13821 15142 13855
rect 18061 13821 18095 13855
rect 18328 13821 18362 13855
rect 19901 13821 19935 13855
rect 20085 13821 20119 13855
rect 20453 13821 20487 13855
rect 20545 13821 20579 13855
rect 2697 13753 2731 13787
rect 17325 13753 17359 13787
rect 20812 13753 20846 13787
rect 2605 13685 2639 13719
rect 6837 13685 6871 13719
rect 7205 13685 7239 13719
rect 16221 13685 16255 13719
rect 16497 13685 16531 13719
rect 17417 13685 17451 13719
rect 3525 13481 3559 13515
rect 4353 13481 4387 13515
rect 4813 13481 4847 13515
rect 7481 13481 7515 13515
rect 9229 13481 9263 13515
rect 10149 13481 10183 13515
rect 11161 13481 11195 13515
rect 11621 13481 11655 13515
rect 15025 13481 15059 13515
rect 15761 13481 15795 13515
rect 17693 13481 17727 13515
rect 19349 13481 19383 13515
rect 20269 13481 20303 13515
rect 2412 13413 2446 13447
rect 5632 13413 5666 13447
rect 13890 13413 13924 13447
rect 20177 13413 20211 13447
rect 21180 13413 21214 13447
rect 1593 13345 1627 13379
rect 4721 13345 4755 13379
rect 7297 13345 7331 13379
rect 8105 13345 8139 13379
rect 10241 13345 10275 13379
rect 11621 13345 11655 13379
rect 11805 13345 11839 13379
rect 15669 13345 15703 13379
rect 16313 13345 16347 13379
rect 16580 13345 16614 13379
rect 18236 13345 18270 13379
rect 20913 13345 20947 13379
rect 2145 13277 2179 13311
rect 4905 13277 4939 13311
rect 5365 13277 5399 13311
rect 7849 13277 7883 13311
rect 10333 13277 10367 13311
rect 11253 13277 11287 13311
rect 11437 13277 11471 13311
rect 13645 13277 13679 13311
rect 15945 13277 15979 13311
rect 17969 13277 18003 13311
rect 20453 13277 20487 13311
rect 1777 13141 1811 13175
rect 6745 13141 6779 13175
rect 9781 13141 9815 13175
rect 10793 13141 10827 13175
rect 13093 13141 13127 13175
rect 15301 13141 15335 13175
rect 19809 13141 19843 13175
rect 22293 13141 22327 13175
rect 3065 12937 3099 12971
rect 4721 12937 4755 12971
rect 7021 12937 7055 12971
rect 9137 12937 9171 12971
rect 9229 12937 9263 12971
rect 13829 12937 13863 12971
rect 17601 12937 17635 12971
rect 19441 12937 19475 12971
rect 22293 12937 22327 12971
rect 7481 12869 7515 12903
rect 11437 12869 11471 12903
rect 16773 12869 16807 12903
rect 1685 12801 1719 12835
rect 7757 12801 7791 12835
rect 9689 12801 9723 12835
rect 9781 12801 9815 12835
rect 11989 12801 12023 12835
rect 12173 12801 12207 12835
rect 14565 12801 14599 12835
rect 20545 12801 20579 12835
rect 20913 12801 20947 12835
rect 3341 12733 3375 12767
rect 3608 12733 3642 12767
rect 5089 12733 5123 12767
rect 5356 12733 5390 12767
rect 6837 12733 6871 12767
rect 7665 12733 7699 12767
rect 10057 12733 10091 12767
rect 12449 12733 12483 12767
rect 14381 12733 14415 12767
rect 14749 12733 14783 12767
rect 15393 12733 15427 12767
rect 15660 12733 15694 12767
rect 17325 12733 17359 12767
rect 17417 12733 17451 12767
rect 18061 12733 18095 12767
rect 21180 12733 21214 12767
rect 1952 12665 1986 12699
rect 8024 12665 8058 12699
rect 9597 12665 9631 12699
rect 10324 12665 10358 12699
rect 11897 12665 11931 12699
rect 12694 12665 12728 12699
rect 15117 12665 15151 12699
rect 18306 12665 18340 12699
rect 20269 12665 20303 12699
rect 6469 12597 6503 12631
rect 11529 12597 11563 12631
rect 13921 12597 13955 12631
rect 14289 12597 14323 12631
rect 14933 12597 14967 12631
rect 17141 12597 17175 12631
rect 19901 12597 19935 12631
rect 20361 12597 20395 12631
rect 2789 12393 2823 12427
rect 3617 12393 3651 12427
rect 4353 12393 4387 12427
rect 6377 12393 6411 12427
rect 8585 12393 8619 12427
rect 10701 12393 10735 12427
rect 12449 12393 12483 12427
rect 14381 12393 14415 12427
rect 15301 12393 15335 12427
rect 20269 12393 20303 12427
rect 22293 12393 22327 12427
rect 13246 12325 13280 12359
rect 14933 12325 14967 12359
rect 21158 12325 21192 12359
rect 1665 12257 1699 12291
rect 3341 12257 3375 12291
rect 3433 12257 3467 12291
rect 4169 12257 4203 12291
rect 4988 12257 5022 12291
rect 6745 12257 6779 12291
rect 7941 12257 7975 12291
rect 8953 12257 8987 12291
rect 10057 12257 10091 12291
rect 10885 12257 10919 12291
rect 11161 12257 11195 12291
rect 14749 12257 14783 12291
rect 15669 12257 15703 12291
rect 16221 12257 16255 12291
rect 16488 12257 16522 12291
rect 17969 12257 18003 12291
rect 18225 12257 18259 12291
rect 20177 12257 20211 12291
rect 20913 12257 20947 12291
rect 1409 12189 1443 12223
rect 4721 12189 4755 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 8033 12189 8067 12223
rect 8125 12189 8159 12223
rect 9045 12189 9079 12223
rect 9137 12189 9171 12223
rect 9781 12189 9815 12223
rect 13001 12189 13035 12223
rect 15117 12189 15151 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 20453 12189 20487 12223
rect 19349 12121 19383 12155
rect 3157 12053 3191 12087
rect 6101 12053 6135 12087
rect 7573 12053 7607 12087
rect 9781 12053 9815 12087
rect 9873 12053 9907 12087
rect 17601 12053 17635 12087
rect 19809 12053 19843 12087
rect 2789 11849 2823 11883
rect 3065 11849 3099 11883
rect 6377 11849 6411 11883
rect 7297 11849 7331 11883
rect 9045 11849 9079 11883
rect 9505 11849 9539 11883
rect 11253 11849 11287 11883
rect 13829 11849 13863 11883
rect 14105 11849 14139 11883
rect 19993 11849 20027 11883
rect 21741 11849 21775 11883
rect 11989 11781 12023 11815
rect 15117 11781 15151 11815
rect 22201 11781 22235 11815
rect 1409 11713 1443 11747
rect 3525 11713 3559 11747
rect 3709 11713 3743 11747
rect 4721 11713 4755 11747
rect 7665 11713 7699 11747
rect 9873 11713 9907 11747
rect 14933 11713 14967 11747
rect 15577 11713 15611 11747
rect 15761 11713 15795 11747
rect 16589 11713 16623 11747
rect 17601 11713 17635 11747
rect 1676 11645 1710 11679
rect 3433 11645 3467 11679
rect 4169 11645 4203 11679
rect 6561 11645 6595 11679
rect 7113 11645 7147 11679
rect 9321 11645 9355 11679
rect 11713 11645 11747 11679
rect 11805 11645 11839 11679
rect 12449 11645 12483 11679
rect 12716 11645 12750 11679
rect 13921 11645 13955 11679
rect 16405 11645 16439 11679
rect 17325 11645 17359 11679
rect 18061 11645 18095 11679
rect 18317 11645 18351 11679
rect 19809 11645 19843 11679
rect 20361 11645 20395 11679
rect 20617 11645 20651 11679
rect 22017 11645 22051 11679
rect 4988 11577 5022 11611
rect 7910 11577 7944 11611
rect 10140 11577 10174 11611
rect 14657 11577 14691 11611
rect 14749 11577 14783 11611
rect 4353 11509 4387 11543
rect 6101 11509 6135 11543
rect 11529 11509 11563 11543
rect 14289 11509 14323 11543
rect 15485 11509 15519 11543
rect 15945 11509 15979 11543
rect 16313 11509 16347 11543
rect 16957 11509 16991 11543
rect 17417 11509 17451 11543
rect 19441 11509 19475 11543
rect 1409 11305 1443 11339
rect 1869 11305 1903 11339
rect 2421 11305 2455 11339
rect 2789 11305 2823 11339
rect 6285 11305 6319 11339
rect 6561 11305 6595 11339
rect 11069 11305 11103 11339
rect 12725 11305 12759 11339
rect 15025 11305 15059 11339
rect 16773 11305 16807 11339
rect 17693 11305 17727 11339
rect 19901 11305 19935 11339
rect 22293 11305 22327 11339
rect 1777 11237 1811 11271
rect 8002 11237 8036 11271
rect 9956 11237 9990 11271
rect 21158 11237 21192 11271
rect 2881 11169 2915 11203
rect 3433 11169 3467 11203
rect 4353 11169 4387 11203
rect 4905 11169 4939 11203
rect 5172 11169 5206 11203
rect 6929 11169 6963 11203
rect 7021 11169 7055 11203
rect 7757 11169 7791 11203
rect 9689 11169 9723 11203
rect 11345 11169 11379 11203
rect 11612 11169 11646 11203
rect 13268 11169 13302 11203
rect 14473 11169 14507 11203
rect 14841 11169 14875 11203
rect 15660 11169 15694 11203
rect 17601 11169 17635 11203
rect 18512 11169 18546 11203
rect 20085 11169 20119 11203
rect 20177 11169 20211 11203
rect 20913 11169 20947 11203
rect 2053 11101 2087 11135
rect 3065 11101 3099 11135
rect 7205 11101 7239 11135
rect 13001 11101 13035 11135
rect 15393 11101 15427 11135
rect 17877 11101 17911 11135
rect 18245 11101 18279 11135
rect 3617 11033 3651 11067
rect 4537 11033 4571 11067
rect 14657 11033 14691 11067
rect 9137 10965 9171 10999
rect 14381 10965 14415 10999
rect 17233 10965 17267 10999
rect 19625 10965 19659 10999
rect 20361 10965 20395 10999
rect 2605 10761 2639 10795
rect 3617 10761 3651 10795
rect 4445 10761 4479 10795
rect 7113 10761 7147 10795
rect 8861 10761 8895 10795
rect 10977 10761 11011 10795
rect 14841 10761 14875 10795
rect 20361 10761 20395 10795
rect 2237 10625 2271 10659
rect 3157 10625 3191 10659
rect 4077 10625 4111 10659
rect 4261 10625 4295 10659
rect 1961 10557 1995 10591
rect 2053 10557 2087 10591
rect 3065 10557 3099 10591
rect 3985 10557 4019 10591
rect 10517 10693 10551 10727
rect 11989 10693 12023 10727
rect 17417 10693 17451 10727
rect 11621 10625 11655 10659
rect 15577 10625 15611 10659
rect 16040 10625 16074 10659
rect 18567 10625 18601 10659
rect 20913 10625 20947 10659
rect 5089 10557 5123 10591
rect 6929 10557 6963 10591
rect 7481 10557 7515 10591
rect 8953 10557 8987 10591
rect 9137 10557 9171 10591
rect 12173 10557 12207 10591
rect 12449 10557 12483 10591
rect 12909 10557 12943 10591
rect 13001 10557 13035 10591
rect 14657 10557 14691 10591
rect 15393 10557 15427 10591
rect 16313 10557 16347 10591
rect 17877 10557 17911 10591
rect 18061 10557 18095 10591
rect 18797 10557 18831 10591
rect 20177 10557 20211 10591
rect 4629 10489 4663 10523
rect 5334 10489 5368 10523
rect 7748 10489 7782 10523
rect 9382 10489 9416 10523
rect 13268 10489 13302 10523
rect 21158 10489 21192 10523
rect 1593 10421 1627 10455
rect 2973 10421 3007 10455
rect 4445 10421 4479 10455
rect 6469 10421 6503 10455
rect 8953 10421 8987 10455
rect 11345 10421 11379 10455
rect 11437 10421 11471 10455
rect 12633 10421 12667 10455
rect 12909 10421 12943 10455
rect 14381 10421 14415 10455
rect 15209 10421 15243 10455
rect 16043 10421 16077 10455
rect 17693 10421 17727 10455
rect 18527 10421 18561 10455
rect 19901 10421 19935 10455
rect 22293 10421 22327 10455
rect 1961 10217 1995 10251
rect 5365 10217 5399 10251
rect 5733 10217 5767 10251
rect 3433 10149 3467 10183
rect 5273 10149 5307 10183
rect 2329 10081 2363 10115
rect 3341 10081 3375 10115
rect 4353 10081 4387 10115
rect 5733 10081 5767 10115
rect 5825 10217 5859 10251
rect 13369 10217 13403 10251
rect 14105 10217 14139 10251
rect 16681 10217 16715 10251
rect 17141 10217 17175 10251
rect 18061 10217 18095 10251
rect 18613 10217 18647 10251
rect 19073 10217 19107 10251
rect 20085 10217 20119 10251
rect 14013 10149 14047 10183
rect 21158 10149 21192 10183
rect 5917 10081 5951 10115
rect 6184 10081 6218 10115
rect 7573 10081 7607 10115
rect 7829 10081 7863 10115
rect 9413 10081 9447 10115
rect 9781 10081 9815 10115
rect 10333 10081 10367 10115
rect 10600 10081 10634 10115
rect 12245 10081 12279 10115
rect 14657 10081 14691 10115
rect 15301 10081 15335 10115
rect 15568 10081 15602 10115
rect 16957 10081 16991 10115
rect 17969 10081 18003 10115
rect 18981 10081 19015 10115
rect 19993 10081 20027 10115
rect 20913 10081 20947 10115
rect 1501 10013 1535 10047
rect 2421 10013 2455 10047
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 5549 10013 5583 10047
rect 5825 10013 5859 10047
rect 11989 10013 12023 10047
rect 14197 10013 14231 10047
rect 18245 10013 18279 10047
rect 19165 10013 19199 10047
rect 20177 10013 20211 10047
rect 1869 9945 1903 9979
rect 2973 9945 3007 9979
rect 4905 9945 4939 9979
rect 8953 9945 8987 9979
rect 14841 9945 14875 9979
rect 4537 9877 4571 9911
rect 7297 9877 7331 9911
rect 9229 9877 9263 9911
rect 9965 9877 9999 9911
rect 11713 9877 11747 9911
rect 13645 9877 13679 9911
rect 17601 9877 17635 9911
rect 19625 9877 19659 9911
rect 22293 9877 22327 9911
rect 2053 9605 2087 9639
rect 7205 9605 7239 9639
rect 9229 9605 9263 9639
rect 14841 9605 14875 9639
rect 16037 9605 16071 9639
rect 17233 9605 17267 9639
rect 2513 9537 2547 9571
rect 2697 9537 2731 9571
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 5089 9537 5123 9571
rect 7849 9537 7883 9571
rect 8861 9537 8895 9571
rect 9873 9537 9907 9571
rect 12817 9537 12851 9571
rect 15393 9537 15427 9571
rect 16589 9537 16623 9571
rect 18521 9537 18555 9571
rect 18705 9537 18739 9571
rect 19579 9537 19613 9571
rect 21649 9537 21683 9571
rect 21833 9537 21867 9571
rect 1593 9469 1627 9503
rect 2421 9469 2455 9503
rect 3433 9469 3467 9503
rect 3525 9469 3559 9503
rect 5356 9469 5390 9503
rect 8125 9469 8159 9503
rect 8585 9469 8619 9503
rect 9597 9469 9631 9503
rect 10241 9469 10275 9503
rect 10508 9469 10542 9503
rect 12449 9469 12483 9503
rect 13185 9469 13219 9503
rect 15209 9469 15243 9503
rect 17049 9469 17083 9503
rect 17785 9469 17819 9503
rect 18429 9469 18463 9503
rect 18889 9469 18923 9503
rect 19073 9469 19107 9503
rect 19809 9469 19843 9503
rect 4445 9401 4479 9435
rect 7665 9401 7699 9435
rect 8677 9401 8711 9435
rect 12633 9401 12667 9435
rect 13430 9401 13464 9435
rect 15301 9401 15335 9435
rect 16497 9401 16531 9435
rect 21557 9401 21591 9435
rect 3065 9333 3099 9367
rect 4077 9333 4111 9367
rect 4537 9333 4571 9367
rect 6469 9333 6503 9367
rect 7573 9333 7607 9367
rect 8125 9333 8159 9367
rect 8217 9333 8251 9367
rect 9689 9333 9723 9367
rect 11621 9333 11655 9367
rect 11897 9333 11931 9367
rect 14565 9333 14599 9367
rect 16405 9333 16439 9367
rect 17601 9333 17635 9367
rect 18061 9333 18095 9367
rect 19539 9333 19573 9367
rect 20913 9333 20947 9367
rect 21189 9333 21223 9367
rect 2513 9129 2547 9163
rect 4537 9129 4571 9163
rect 4905 9129 4939 9163
rect 5549 9129 5583 9163
rect 5917 9129 5951 9163
rect 6009 9129 6043 9163
rect 6561 9129 6595 9163
rect 9413 9129 9447 9163
rect 14749 9129 14783 9163
rect 18245 9129 18279 9163
rect 20453 9129 20487 9163
rect 3433 9061 3467 9095
rect 8033 9061 8067 9095
rect 8953 9061 8987 9095
rect 9956 9061 9990 9095
rect 13338 9061 13372 9095
rect 16650 9061 16684 9095
rect 21180 9061 21214 9095
rect 3341 8993 3375 9027
rect 4997 8993 5031 9027
rect 6929 8993 6963 9027
rect 7941 8993 7975 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 11437 8993 11471 9027
rect 11704 8993 11738 9027
rect 15669 8993 15703 9027
rect 16405 8993 16439 9027
rect 18061 8993 18095 9027
rect 18936 8993 18970 9027
rect 20913 8993 20947 9027
rect 2053 8925 2087 8959
rect 3617 8925 3651 8959
rect 4077 8925 4111 8959
rect 5181 8925 5215 8959
rect 6101 8925 6135 8959
rect 7021 8925 7055 8959
rect 7205 8925 7239 8959
rect 8217 8925 8251 8959
rect 9045 8925 9079 8959
rect 9229 8925 9263 8959
rect 13093 8925 13127 8959
rect 15761 8925 15795 8959
rect 15853 8925 15887 8959
rect 18613 8925 18647 8959
rect 19119 8925 19153 8959
rect 19349 8925 19383 8959
rect 4445 8857 4479 8891
rect 7573 8857 7607 8891
rect 22293 8857 22327 8891
rect 2973 8789 3007 8823
rect 8585 8789 8619 8823
rect 11069 8789 11103 8823
rect 12817 8789 12851 8823
rect 14473 8789 14507 8823
rect 15301 8789 15335 8823
rect 17785 8789 17819 8823
rect 2697 8585 2731 8619
rect 5733 8585 5767 8619
rect 7297 8585 7331 8619
rect 11713 8585 11747 8619
rect 12265 8585 12299 8619
rect 17417 8585 17451 8619
rect 19717 8585 19751 8619
rect 4721 8517 4755 8551
rect 7665 8517 7699 8551
rect 11989 8517 12023 8551
rect 2789 8449 2823 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 8309 8449 8343 8483
rect 10333 8449 10367 8483
rect 3893 8381 3927 8415
rect 4629 8381 4663 8415
rect 5089 8381 5123 8415
rect 6101 8381 6135 8415
rect 7113 8381 7147 8415
rect 8677 8381 8711 8415
rect 10241 8381 10275 8415
rect 12173 8381 12207 8415
rect 3249 8313 3283 8347
rect 5181 8313 5215 8347
rect 6193 8313 6227 8347
rect 8033 8313 8067 8347
rect 8922 8313 8956 8347
rect 10600 8313 10634 8347
rect 3525 8245 3559 8279
rect 8125 8245 8159 8279
rect 10057 8245 10091 8279
rect 10241 8245 10275 8279
rect 14841 8517 14875 8551
rect 16957 8517 16991 8551
rect 20729 8517 20763 8551
rect 22293 8517 22327 8551
rect 13001 8449 13035 8483
rect 15117 8449 15151 8483
rect 15440 8449 15474 8483
rect 15580 8449 15614 8483
rect 20177 8449 20211 8483
rect 20361 8449 20395 8483
rect 20913 8449 20947 8483
rect 12817 8381 12851 8415
rect 13461 8381 13495 8415
rect 13728 8381 13762 8415
rect 15853 8381 15887 8415
rect 17233 8381 17267 8415
rect 18889 8381 18923 8415
rect 20545 8381 20579 8415
rect 21180 8381 21214 8415
rect 19533 8313 19567 8347
rect 20085 8313 20119 8347
rect 12265 8245 12299 8279
rect 12449 8245 12483 8279
rect 12909 8245 12943 8279
rect 18705 8245 18739 8279
rect 5273 8041 5307 8075
rect 5917 8041 5951 8075
rect 6377 8041 6411 8075
rect 6929 8041 6963 8075
rect 9321 8041 9355 8075
rect 11713 8041 11747 8075
rect 16773 8041 16807 8075
rect 18429 8041 18463 8075
rect 19901 8041 19935 8075
rect 3525 7973 3559 8007
rect 7297 7973 7331 8007
rect 9956 7973 9990 8007
rect 5365 7905 5399 7939
rect 6285 7905 6319 7939
rect 8208 7905 8242 7939
rect 9689 7905 9723 7939
rect 11345 7905 11379 7939
rect 4353 7837 4387 7871
rect 4445 7837 4479 7871
rect 5457 7837 5491 7871
rect 6469 7837 6503 7871
rect 7389 7837 7423 7871
rect 7573 7837 7607 7871
rect 7941 7837 7975 7871
rect 12164 7973 12198 8007
rect 13369 7973 13403 8007
rect 13820 7973 13854 8007
rect 18766 7973 18800 8007
rect 21281 7973 21315 8007
rect 11897 7837 11931 7871
rect 15301 7905 15335 7939
rect 15649 7905 15683 7939
rect 17305 7905 17339 7939
rect 20361 7905 20395 7939
rect 21925 7905 21959 7939
rect 13553 7837 13587 7871
rect 11713 7769 11747 7803
rect 13277 7769 13311 7803
rect 13369 7769 13403 7803
rect 15393 7837 15427 7871
rect 17049 7837 17083 7871
rect 18521 7837 18555 7871
rect 20453 7837 20487 7871
rect 20545 7837 20579 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 4905 7701 4939 7735
rect 11069 7701 11103 7735
rect 11529 7701 11563 7735
rect 14933 7701 14967 7735
rect 15301 7701 15335 7735
rect 19993 7701 20027 7735
rect 20913 7701 20947 7735
rect 22109 7701 22143 7735
rect 5733 7497 5767 7531
rect 7205 7497 7239 7531
rect 9597 7497 9631 7531
rect 12449 7497 12483 7531
rect 16129 7497 16163 7531
rect 16405 7497 16439 7531
rect 21189 7497 21223 7531
rect 10977 7429 11011 7463
rect 15945 7429 15979 7463
rect 16037 7429 16071 7463
rect 5365 7361 5399 7395
rect 6193 7361 6227 7395
rect 6377 7361 6411 7395
rect 7665 7361 7699 7395
rect 7849 7361 7883 7395
rect 10333 7361 10367 7395
rect 10425 7361 10459 7395
rect 11529 7361 11563 7395
rect 13001 7361 13035 7395
rect 14568 7361 14602 7395
rect 5089 7293 5123 7327
rect 7573 7293 7607 7327
rect 8217 7293 8251 7327
rect 12265 7293 12299 7327
rect 13461 7293 13495 7327
rect 14105 7293 14139 7327
rect 14841 7293 14875 7327
rect 16037 7293 16071 7327
rect 20545 7429 20579 7463
rect 17509 7361 17543 7395
rect 19211 7361 19245 7395
rect 19441 7361 19475 7395
rect 21741 7361 21775 7395
rect 16129 7293 16163 7327
rect 16221 7293 16255 7327
rect 17325 7293 17359 7327
rect 18153 7293 18187 7327
rect 18705 7293 18739 7327
rect 19028 7293 19062 7327
rect 21649 7293 21683 7327
rect 4261 7225 4295 7259
rect 5181 7225 5215 7259
rect 6101 7225 6135 7259
rect 8484 7225 8518 7259
rect 10241 7225 10275 7259
rect 11437 7225 11471 7259
rect 17417 7225 17451 7259
rect 4721 7157 4755 7191
rect 9873 7157 9907 7191
rect 11345 7157 11379 7191
rect 12081 7157 12115 7191
rect 12817 7157 12851 7191
rect 12909 7157 12943 7191
rect 13645 7157 13679 7191
rect 14571 7157 14605 7191
rect 16957 7157 16991 7191
rect 18337 7157 18371 7191
rect 21557 7157 21591 7191
rect 6837 6953 6871 6987
rect 7297 6953 7331 6987
rect 10057 6953 10091 6987
rect 12357 6953 12391 6987
rect 13093 6953 13127 6987
rect 17515 6953 17549 6987
rect 11253 6885 11287 6919
rect 15546 6885 15580 6919
rect 19432 6885 19466 6919
rect 5457 6817 5491 6851
rect 6101 6817 6135 6851
rect 8208 6817 8242 6851
rect 10149 6817 10183 6851
rect 12265 6817 12299 6851
rect 12909 6817 12943 6851
rect 13553 6817 13587 6851
rect 13820 6817 13854 6851
rect 17785 6817 17819 6851
rect 19165 6817 19199 6851
rect 20637 6817 20671 6851
rect 21169 6817 21203 6851
rect 6193 6749 6227 6783
rect 6377 6749 6411 6783
rect 7389 6749 7423 6783
rect 7573 6749 7607 6783
rect 7941 6749 7975 6783
rect 10333 6749 10367 6783
rect 11345 6749 11379 6783
rect 11529 6749 11563 6783
rect 12449 6749 12483 6783
rect 15301 6749 15335 6783
rect 17049 6749 17083 6783
rect 17512 6749 17546 6783
rect 5733 6681 5767 6715
rect 11897 6681 11931 6715
rect 20913 6749 20947 6783
rect 6929 6613 6963 6647
rect 9321 6613 9355 6647
rect 9689 6613 9723 6647
rect 10885 6613 10919 6647
rect 14933 6613 14967 6647
rect 16681 6613 16715 6647
rect 18889 6613 18923 6647
rect 20545 6613 20579 6647
rect 20637 6613 20671 6647
rect 22293 6613 22327 6647
rect 9689 6409 9723 6443
rect 12633 6409 12667 6443
rect 14749 6409 14783 6443
rect 15945 6409 15979 6443
rect 19809 6409 19843 6443
rect 20269 6409 20303 6443
rect 6285 6273 6319 6307
rect 7941 6273 7975 6307
rect 15301 6273 15335 6307
rect 7665 6205 7699 6239
rect 8309 6205 8343 6239
rect 8576 6205 8610 6239
rect 10057 6205 10091 6239
rect 10609 6205 10643 6239
rect 12449 6205 12483 6239
rect 13093 6205 13127 6239
rect 15761 6205 15795 6239
rect 16313 6205 16347 6239
rect 18429 6205 18463 6239
rect 20085 6205 20119 6239
rect 20637 6205 20671 6239
rect 20904 6205 20938 6239
rect 7757 6137 7791 6171
rect 10876 6137 10910 6171
rect 13360 6137 13394 6171
rect 15209 6137 15243 6171
rect 16580 6137 16614 6171
rect 18696 6137 18730 6171
rect 6837 6069 6871 6103
rect 7297 6069 7331 6103
rect 10241 6069 10275 6103
rect 11989 6069 12023 6103
rect 14473 6069 14507 6103
rect 15117 6069 15151 6103
rect 17693 6069 17727 6103
rect 22017 6069 22051 6103
rect 6929 5865 6963 5899
rect 10057 5865 10091 5899
rect 14841 5865 14875 5899
rect 17509 5865 17543 5899
rect 20269 5865 20303 5899
rect 18797 5797 18831 5831
rect 7297 5729 7331 5763
rect 7389 5729 7423 5763
rect 8208 5729 8242 5763
rect 11244 5729 11278 5763
rect 12909 5729 12943 5763
rect 13001 5729 13035 5763
rect 13268 5729 13302 5763
rect 14657 5729 14691 5763
rect 15577 5729 15611 5763
rect 16385 5729 16419 5763
rect 17877 5729 17911 5763
rect 20177 5729 20211 5763
rect 21180 5729 21214 5763
rect 7573 5661 7607 5695
rect 7941 5661 7975 5695
rect 10149 5661 10183 5695
rect 10241 5661 10275 5695
rect 10977 5661 11011 5695
rect 16129 5661 16163 5695
rect 18889 5661 18923 5695
rect 19073 5661 19107 5695
rect 20453 5661 20487 5695
rect 20913 5661 20947 5695
rect 19809 5593 19843 5627
rect 9321 5525 9355 5559
rect 9689 5525 9723 5559
rect 12357 5525 12391 5559
rect 12725 5525 12759 5559
rect 14381 5525 14415 5559
rect 15761 5525 15795 5559
rect 18061 5525 18095 5559
rect 18429 5525 18463 5559
rect 22293 5525 22327 5559
rect 9597 5321 9631 5355
rect 12081 5321 12115 5355
rect 19441 5321 19475 5355
rect 19717 5321 19751 5355
rect 10241 5185 10275 5219
rect 12909 5185 12943 5219
rect 17601 5185 17635 5219
rect 20269 5185 20303 5219
rect 8217 5117 8251 5151
rect 10057 5117 10091 5151
rect 10701 5117 10735 5151
rect 10968 5117 11002 5151
rect 14749 5117 14783 5151
rect 15301 5117 15335 5151
rect 17417 5117 17451 5151
rect 18061 5117 18095 5151
rect 20913 5117 20947 5151
rect 8484 5049 8518 5083
rect 13176 5049 13210 5083
rect 15568 5049 15602 5083
rect 18328 5049 18362 5083
rect 20085 5049 20119 5083
rect 21158 5049 21192 5083
rect 9873 4981 9907 5015
rect 12449 4981 12483 5015
rect 14289 4981 14323 5015
rect 14933 4981 14967 5015
rect 16681 4981 16715 5015
rect 16957 4981 16991 5015
rect 17325 4981 17359 5015
rect 20177 4981 20211 5015
rect 22293 4981 22327 5015
rect 10057 4777 10091 4811
rect 12633 4777 12667 4811
rect 13093 4777 13127 4811
rect 13185 4777 13219 4811
rect 13553 4777 13587 4811
rect 13645 4777 13679 4811
rect 14565 4777 14599 4811
rect 14657 4777 14691 4811
rect 15853 4777 15887 4811
rect 17877 4777 17911 4811
rect 18705 4777 18739 4811
rect 19165 4777 19199 4811
rect 19717 4777 19751 4811
rect 20085 4777 20119 4811
rect 10784 4709 10818 4743
rect 19073 4709 19107 4743
rect 21180 4709 21214 4743
rect 9137 4641 9171 4675
rect 11989 4641 12023 4675
rect 12541 4641 12575 4675
rect 13093 4641 13127 4675
rect 15669 4641 15703 4675
rect 16589 4641 16623 4675
rect 17785 4641 17819 4675
rect 10517 4573 10551 4607
rect 12817 4573 12851 4607
rect 13829 4573 13863 4607
rect 14749 4573 14783 4607
rect 16681 4573 16715 4607
rect 16865 4573 16899 4607
rect 17969 4573 18003 4607
rect 19257 4573 19291 4607
rect 19533 4573 19567 4607
rect 20177 4573 20211 4607
rect 20269 4573 20303 4607
rect 20913 4573 20947 4607
rect 11897 4437 11931 4471
rect 11989 4437 12023 4471
rect 12173 4437 12207 4471
rect 14197 4437 14231 4471
rect 16221 4437 16255 4471
rect 17417 4437 17451 4471
rect 19533 4437 19567 4471
rect 22293 4437 22327 4471
rect 13277 4233 13311 4267
rect 20269 4233 20303 4267
rect 9597 4097 9631 4131
rect 9781 4097 9815 4131
rect 10701 4097 10735 4131
rect 10885 4097 10919 4131
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 13829 4097 13863 4131
rect 15945 4097 15979 4131
rect 18705 4097 18739 4131
rect 19717 4097 19751 4131
rect 9505 4029 9539 4063
rect 10609 4029 10643 4063
rect 11621 4029 11655 4063
rect 12725 4029 12759 4063
rect 13645 4029 13679 4063
rect 14289 4029 14323 4063
rect 18521 4029 18555 4063
rect 20085 4029 20119 4063
rect 20729 4029 20763 4063
rect 14556 3961 14590 3995
rect 16190 3961 16224 3995
rect 18429 3961 18463 3995
rect 19441 3961 19475 3995
rect 20974 3961 21008 3995
rect 9137 3893 9171 3927
rect 10241 3893 10275 3927
rect 11253 3893 11287 3927
rect 12909 3893 12943 3927
rect 13737 3893 13771 3927
rect 15669 3893 15703 3927
rect 17325 3893 17359 3927
rect 18061 3893 18095 3927
rect 19073 3893 19107 3927
rect 19533 3893 19567 3927
rect 22109 3893 22143 3927
rect 11161 3689 11195 3723
rect 13185 3689 13219 3723
rect 13553 3689 13587 3723
rect 20453 3689 20487 3723
rect 22293 3689 22327 3723
rect 11529 3621 11563 3655
rect 12541 3621 12575 3655
rect 13645 3621 13679 3655
rect 14565 3621 14599 3655
rect 17202 3621 17236 3655
rect 10701 3553 10735 3587
rect 12633 3553 12667 3587
rect 14657 3553 14691 3587
rect 15557 3553 15591 3587
rect 18613 3553 18647 3587
rect 18869 3553 18903 3587
rect 20269 3553 20303 3587
rect 21180 3553 21214 3587
rect 11621 3485 11655 3519
rect 11805 3485 11839 3519
rect 12817 3485 12851 3519
rect 13737 3485 13771 3519
rect 14841 3485 14875 3519
rect 15301 3485 15335 3519
rect 16957 3485 16991 3519
rect 20913 3485 20947 3519
rect 14197 3417 14231 3451
rect 12173 3349 12207 3383
rect 16681 3349 16715 3383
rect 18337 3349 18371 3383
rect 19993 3349 20027 3383
rect 17417 3145 17451 3179
rect 18245 3145 18279 3179
rect 19993 3145 20027 3179
rect 20085 3145 20119 3179
rect 13185 3077 13219 3111
rect 15577 3077 15611 3111
rect 12725 3009 12759 3043
rect 13737 3009 13771 3043
rect 20085 3009 20119 3043
rect 20177 3077 20211 3111
rect 11713 2941 11747 2975
rect 14197 2941 14231 2975
rect 16037 2941 16071 2975
rect 16304 2941 16338 2975
rect 18061 2941 18095 2975
rect 18613 2941 18647 2975
rect 18880 2941 18914 2975
rect 20177 2941 20211 2975
rect 20269 2941 20303 2975
rect 20525 2941 20559 2975
rect 21925 2941 21959 2975
rect 22109 2941 22143 2975
rect 13645 2873 13679 2907
rect 14464 2873 14498 2907
rect 22293 2873 22327 2907
rect 11897 2805 11931 2839
rect 13553 2805 13587 2839
rect 21649 2805 21683 2839
rect 14381 2601 14415 2635
rect 14841 2601 14875 2635
rect 15209 2601 15243 2635
rect 16865 2601 16899 2635
rect 17601 2601 17635 2635
rect 19717 2601 19751 2635
rect 20085 2601 20119 2635
rect 20453 2601 20487 2635
rect 12909 2533 12943 2567
rect 14749 2533 14783 2567
rect 13737 2465 13771 2499
rect 13829 2397 13863 2431
rect 13921 2397 13955 2431
rect 14933 2397 14967 2431
rect 15752 2533 15786 2567
rect 18582 2533 18616 2567
rect 21557 2533 21591 2567
rect 15485 2465 15519 2499
rect 17693 2465 17727 2499
rect 20545 2465 20579 2499
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 20637 2397 20671 2431
rect 21649 2397 21683 2431
rect 21833 2397 21867 2431
rect 21189 2329 21223 2363
rect 13369 2261 13403 2295
rect 15209 2261 15243 2295
rect 17233 2261 17267 2295
<< metal1 >>
rect 14274 22788 14280 22840
rect 14332 22828 14338 22840
rect 19426 22828 19432 22840
rect 14332 22800 19432 22828
rect 14332 22788 14338 22800
rect 19426 22788 19432 22800
rect 19484 22788 19490 22840
rect 10502 22312 10508 22364
rect 10560 22352 10566 22364
rect 17862 22352 17868 22364
rect 10560 22324 17868 22352
rect 10560 22312 10566 22324
rect 17862 22312 17868 22324
rect 17920 22312 17926 22364
rect 12158 22244 12164 22296
rect 12216 22284 12222 22296
rect 17218 22284 17224 22296
rect 12216 22256 17224 22284
rect 12216 22244 12222 22256
rect 17218 22244 17224 22256
rect 17276 22244 17282 22296
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 19334 22216 19340 22228
rect 16632 22188 19340 22216
rect 16632 22176 16638 22188
rect 19334 22176 19340 22188
rect 19392 22176 19398 22228
rect 16669 22083 16727 22089
rect 16669 22049 16681 22083
rect 16715 22080 16727 22083
rect 19610 22080 19616 22092
rect 16715 22052 19616 22080
rect 16715 22049 16727 22052
rect 16669 22043 16727 22049
rect 19610 22040 19616 22052
rect 19668 22040 19674 22092
rect 14918 21972 14924 22024
rect 14976 22012 14982 22024
rect 16485 22015 16543 22021
rect 16485 22012 16497 22015
rect 14976 21984 16497 22012
rect 14976 21972 14982 21984
rect 16485 21981 16497 21984
rect 16531 21981 16543 22015
rect 16485 21975 16543 21981
rect 8662 21904 8668 21956
rect 8720 21944 8726 21956
rect 18598 21944 18604 21956
rect 8720 21916 18604 21944
rect 8720 21904 8726 21916
rect 18598 21904 18604 21916
rect 18656 21904 18662 21956
rect 12710 21836 12716 21888
rect 12768 21876 12774 21888
rect 21726 21876 21732 21888
rect 12768 21848 21732 21876
rect 12768 21836 12774 21848
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 1104 21786 22816 21808
rect 1104 21734 4614 21786
rect 4666 21734 4678 21786
rect 4730 21734 4742 21786
rect 4794 21734 4806 21786
rect 4858 21734 11878 21786
rect 11930 21734 11942 21786
rect 11994 21734 12006 21786
rect 12058 21734 12070 21786
rect 12122 21734 19142 21786
rect 19194 21734 19206 21786
rect 19258 21734 19270 21786
rect 19322 21734 19334 21786
rect 19386 21734 22816 21786
rect 1104 21712 22816 21734
rect 290 21632 296 21684
rect 348 21672 354 21684
rect 1581 21675 1639 21681
rect 1581 21672 1593 21675
rect 348 21644 1593 21672
rect 348 21632 354 21644
rect 1581 21641 1593 21644
rect 1627 21641 1639 21675
rect 4338 21672 4344 21684
rect 1581 21635 1639 21641
rect 3436 21644 4344 21672
rect 2593 21539 2651 21545
rect 2593 21505 2605 21539
rect 2639 21536 2651 21539
rect 3234 21536 3240 21548
rect 2639 21508 3240 21536
rect 2639 21505 2651 21508
rect 2593 21499 2651 21505
rect 3234 21496 3240 21508
rect 3292 21496 3298 21548
rect 3436 21545 3464 21644
rect 4338 21632 4344 21644
rect 4396 21632 4402 21684
rect 4893 21675 4951 21681
rect 4893 21641 4905 21675
rect 4939 21672 4951 21675
rect 4939 21644 8064 21672
rect 4939 21641 4951 21644
rect 4893 21635 4951 21641
rect 3602 21564 3608 21616
rect 3660 21604 3666 21616
rect 3660 21576 4752 21604
rect 3660 21564 3666 21576
rect 3421 21539 3479 21545
rect 3421 21505 3433 21539
rect 3467 21505 3479 21539
rect 3421 21499 3479 21505
rect 3513 21539 3571 21545
rect 3513 21505 3525 21539
rect 3559 21505 3571 21539
rect 3513 21499 3571 21505
rect 1394 21468 1400 21480
rect 1355 21440 1400 21468
rect 1394 21428 1400 21440
rect 1452 21428 1458 21480
rect 3528 21468 3556 21499
rect 3694 21496 3700 21548
rect 3752 21536 3758 21548
rect 4617 21539 4675 21545
rect 4617 21536 4629 21539
rect 3752 21508 4629 21536
rect 3752 21496 3758 21508
rect 4617 21505 4629 21508
rect 4663 21505 4675 21539
rect 4724 21536 4752 21576
rect 4982 21564 4988 21616
rect 5040 21604 5046 21616
rect 6273 21607 6331 21613
rect 6273 21604 6285 21607
rect 5040 21576 6285 21604
rect 5040 21564 5046 21576
rect 6273 21573 6285 21576
rect 6319 21573 6331 21607
rect 8036 21604 8064 21644
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 17310 21672 17316 21684
rect 8168 21644 10732 21672
rect 8168 21632 8174 21644
rect 9674 21604 9680 21616
rect 8036 21576 9680 21604
rect 6273 21567 6331 21573
rect 9674 21564 9680 21576
rect 9732 21564 9738 21616
rect 10704 21604 10732 21644
rect 17052 21644 17316 21672
rect 14826 21604 14832 21616
rect 10704 21576 12020 21604
rect 14739 21576 14832 21604
rect 5629 21539 5687 21545
rect 5629 21536 5641 21539
rect 4724 21508 5641 21536
rect 4617 21499 4675 21505
rect 5629 21505 5641 21508
rect 5675 21505 5687 21539
rect 6822 21536 6828 21548
rect 5629 21499 5687 21505
rect 6012 21508 6828 21536
rect 3878 21468 3884 21480
rect 3528 21440 3884 21468
rect 3878 21428 3884 21440
rect 3936 21428 3942 21480
rect 4154 21428 4160 21480
rect 4212 21468 4218 21480
rect 4525 21471 4583 21477
rect 4525 21468 4537 21471
rect 4212 21440 4537 21468
rect 4212 21428 4218 21440
rect 4525 21437 4537 21440
rect 4571 21437 4583 21471
rect 4525 21431 4583 21437
rect 4890 21428 4896 21480
rect 4948 21468 4954 21480
rect 6012 21468 6040 21508
rect 6822 21496 6828 21508
rect 6880 21536 6886 21548
rect 6917 21539 6975 21545
rect 6917 21536 6929 21539
rect 6880 21508 6929 21536
rect 6880 21496 6886 21508
rect 6917 21505 6929 21508
rect 6963 21505 6975 21539
rect 6917 21499 6975 21505
rect 7926 21496 7932 21548
rect 7984 21536 7990 21548
rect 11992 21545 12020 21576
rect 14826 21564 14832 21576
rect 14884 21604 14890 21616
rect 14884 21576 16988 21604
rect 14884 21564 14890 21576
rect 9125 21539 9183 21545
rect 9125 21536 9137 21539
rect 7984 21508 9137 21536
rect 7984 21496 7990 21508
rect 9125 21505 9137 21508
rect 9171 21505 9183 21539
rect 11885 21539 11943 21545
rect 11885 21536 11897 21539
rect 9125 21499 9183 21505
rect 10796 21508 11897 21536
rect 4948 21440 6040 21468
rect 6089 21471 6147 21477
rect 4948 21428 4954 21440
rect 6089 21437 6101 21471
rect 6135 21468 6147 21471
rect 6638 21468 6644 21480
rect 6135 21440 6644 21468
rect 6135 21437 6147 21440
rect 6089 21431 6147 21437
rect 6638 21428 6644 21440
rect 6696 21428 6702 21480
rect 8389 21471 8447 21477
rect 7116 21440 7328 21468
rect 2317 21403 2375 21409
rect 2317 21369 2329 21403
rect 2363 21400 2375 21403
rect 5445 21403 5503 21409
rect 5445 21400 5457 21403
rect 2363 21372 2728 21400
rect 2363 21369 2375 21372
rect 2317 21363 2375 21369
rect 1394 21292 1400 21344
rect 1452 21332 1458 21344
rect 1949 21335 2007 21341
rect 1949 21332 1961 21335
rect 1452 21304 1961 21332
rect 1452 21292 1458 21304
rect 1949 21301 1961 21304
rect 1995 21301 2007 21335
rect 1949 21295 2007 21301
rect 2409 21335 2467 21341
rect 2409 21301 2421 21335
rect 2455 21332 2467 21335
rect 2590 21332 2596 21344
rect 2455 21304 2596 21332
rect 2455 21301 2467 21304
rect 2409 21295 2467 21301
rect 2590 21292 2596 21304
rect 2648 21292 2654 21344
rect 2700 21332 2728 21372
rect 4080 21372 5457 21400
rect 2958 21332 2964 21344
rect 2700 21304 2964 21332
rect 2958 21292 2964 21304
rect 3016 21292 3022 21344
rect 3326 21332 3332 21344
rect 3287 21304 3332 21332
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 4080 21341 4108 21372
rect 5445 21369 5457 21372
rect 5491 21400 5503 21403
rect 7116 21400 7144 21440
rect 5491 21372 7144 21400
rect 7184 21403 7242 21409
rect 5491 21369 5503 21372
rect 5445 21363 5503 21369
rect 7184 21369 7196 21403
rect 7230 21369 7242 21403
rect 7300 21400 7328 21440
rect 8389 21437 8401 21471
rect 8435 21468 8447 21471
rect 8570 21468 8576 21480
rect 8435 21440 8576 21468
rect 8435 21437 8447 21440
rect 8389 21431 8447 21437
rect 8570 21428 8576 21440
rect 8628 21428 8634 21480
rect 8938 21468 8944 21480
rect 8899 21440 8944 21468
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9582 21428 9588 21480
rect 9640 21468 9646 21480
rect 9769 21471 9827 21477
rect 9769 21468 9781 21471
rect 9640 21440 9781 21468
rect 9640 21428 9646 21440
rect 9769 21437 9781 21440
rect 9815 21437 9827 21471
rect 10796 21468 10824 21508
rect 11885 21505 11897 21508
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 11977 21539 12035 21545
rect 11977 21505 11989 21539
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12526 21496 12532 21548
rect 12584 21536 12590 21548
rect 13449 21539 13507 21545
rect 13449 21536 13461 21539
rect 12584 21508 13461 21536
rect 12584 21496 12590 21508
rect 13449 21505 13461 21508
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 14458 21496 14464 21548
rect 14516 21536 14522 21548
rect 16960 21545 16988 21576
rect 17052 21545 17080 21644
rect 17310 21632 17316 21644
rect 17368 21672 17374 21684
rect 17368 21644 19012 21672
rect 17368 21632 17374 21644
rect 17865 21607 17923 21613
rect 17865 21573 17877 21607
rect 17911 21604 17923 21607
rect 17911 21576 18920 21604
rect 17911 21573 17923 21576
rect 17865 21567 17923 21573
rect 16025 21539 16083 21545
rect 16025 21536 16037 21539
rect 14516 21508 16037 21536
rect 14516 21496 14522 21508
rect 16025 21505 16037 21508
rect 16071 21505 16083 21539
rect 16025 21499 16083 21505
rect 16945 21539 17003 21545
rect 16945 21505 16957 21539
rect 16991 21505 17003 21539
rect 16945 21499 17003 21505
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21505 17095 21539
rect 18785 21539 18843 21545
rect 18785 21536 18797 21539
rect 17037 21499 17095 21505
rect 17144 21508 18797 21536
rect 12618 21468 12624 21480
rect 9769 21431 9827 21437
rect 9876 21440 10824 21468
rect 12579 21440 12624 21468
rect 9876 21400 9904 21440
rect 12618 21428 12624 21440
rect 12676 21428 12682 21480
rect 15841 21471 15899 21477
rect 15841 21437 15853 21471
rect 15887 21468 15899 21471
rect 16206 21468 16212 21480
rect 15887 21440 16212 21468
rect 15887 21437 15899 21440
rect 15841 21431 15899 21437
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 16390 21428 16396 21480
rect 16448 21468 16454 21480
rect 17144 21468 17172 21508
rect 18785 21505 18797 21508
rect 18831 21505 18843 21539
rect 18785 21499 18843 21505
rect 17678 21468 17684 21480
rect 16448 21440 17172 21468
rect 17639 21440 17684 21468
rect 16448 21428 16454 21440
rect 17678 21428 17684 21440
rect 17736 21428 17742 21480
rect 7300 21372 9904 21400
rect 7184 21363 7242 21369
rect 4065 21335 4123 21341
rect 4065 21301 4077 21335
rect 4111 21301 4123 21335
rect 4065 21295 4123 21301
rect 4433 21335 4491 21341
rect 4433 21301 4445 21335
rect 4479 21332 4491 21335
rect 4893 21335 4951 21341
rect 4893 21332 4905 21335
rect 4479 21304 4905 21332
rect 4479 21301 4491 21304
rect 4433 21295 4491 21301
rect 4893 21301 4905 21304
rect 4939 21301 4951 21335
rect 5074 21332 5080 21344
rect 5035 21304 5080 21332
rect 4893 21295 4951 21301
rect 5074 21292 5080 21304
rect 5132 21292 5138 21344
rect 5258 21292 5264 21344
rect 5316 21332 5322 21344
rect 5537 21335 5595 21341
rect 5537 21332 5549 21335
rect 5316 21304 5549 21332
rect 5316 21292 5322 21304
rect 5537 21301 5549 21304
rect 5583 21301 5595 21335
rect 7208 21332 7236 21363
rect 9950 21360 9956 21412
rect 10008 21409 10014 21412
rect 10008 21403 10072 21409
rect 10008 21369 10026 21403
rect 10060 21369 10072 21403
rect 13716 21403 13774 21409
rect 10008 21363 10072 21369
rect 11440 21372 13676 21400
rect 10008 21360 10014 21363
rect 8110 21332 8116 21344
rect 7208 21304 8116 21332
rect 5537 21295 5595 21301
rect 8110 21292 8116 21304
rect 8168 21292 8174 21344
rect 8297 21335 8355 21341
rect 8297 21301 8309 21335
rect 8343 21332 8355 21335
rect 8389 21335 8447 21341
rect 8389 21332 8401 21335
rect 8343 21304 8401 21332
rect 8343 21301 8355 21304
rect 8297 21295 8355 21301
rect 8389 21301 8401 21304
rect 8435 21301 8447 21335
rect 8389 21295 8447 21301
rect 8573 21335 8631 21341
rect 8573 21301 8585 21335
rect 8619 21332 8631 21335
rect 8662 21332 8668 21344
rect 8619 21304 8668 21332
rect 8619 21301 8631 21304
rect 8573 21295 8631 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 9030 21332 9036 21344
rect 8991 21304 9036 21332
rect 9030 21292 9036 21304
rect 9088 21292 9094 21344
rect 11054 21292 11060 21344
rect 11112 21332 11118 21344
rect 11440 21341 11468 21372
rect 11149 21335 11207 21341
rect 11149 21332 11161 21335
rect 11112 21304 11161 21332
rect 11112 21292 11118 21304
rect 11149 21301 11161 21304
rect 11195 21301 11207 21335
rect 11149 21295 11207 21301
rect 11425 21335 11483 21341
rect 11425 21301 11437 21335
rect 11471 21301 11483 21335
rect 11425 21295 11483 21301
rect 11793 21335 11851 21341
rect 11793 21301 11805 21335
rect 11839 21332 11851 21335
rect 12158 21332 12164 21344
rect 11839 21304 12164 21332
rect 11839 21301 11851 21304
rect 11793 21295 11851 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12802 21332 12808 21344
rect 12763 21304 12808 21332
rect 12802 21292 12808 21304
rect 12860 21292 12866 21344
rect 13648 21332 13676 21372
rect 13716 21369 13728 21403
rect 13762 21400 13774 21403
rect 13906 21400 13912 21412
rect 13762 21372 13912 21400
rect 13762 21369 13774 21372
rect 13716 21363 13774 21369
rect 13906 21360 13912 21372
rect 13964 21360 13970 21412
rect 14642 21360 14648 21412
rect 14700 21400 14706 21412
rect 14700 21372 15516 21400
rect 14700 21360 14706 21372
rect 15378 21332 15384 21344
rect 13648 21304 15384 21332
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15488 21341 15516 21372
rect 17218 21360 17224 21412
rect 17276 21400 17282 21412
rect 18693 21403 18751 21409
rect 18693 21400 18705 21403
rect 17276 21372 18705 21400
rect 17276 21360 17282 21372
rect 18693 21369 18705 21372
rect 18739 21369 18751 21403
rect 18892 21400 18920 21576
rect 18984 21545 19012 21644
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 20257 21539 20315 21545
rect 20257 21536 20269 21539
rect 19015 21508 20269 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 20257 21505 20269 21508
rect 20303 21536 20315 21539
rect 20530 21536 20536 21548
rect 20303 21508 20536 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 21726 21536 21732 21548
rect 21687 21508 21732 21536
rect 21726 21496 21732 21508
rect 21784 21496 21790 21548
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 21637 21471 21695 21477
rect 21637 21468 21649 21471
rect 19116 21440 21649 21468
rect 19116 21428 19122 21440
rect 21637 21437 21649 21440
rect 21683 21437 21695 21471
rect 21637 21431 21695 21437
rect 19978 21400 19984 21412
rect 18892 21372 19984 21400
rect 18693 21363 18751 21369
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 20073 21403 20131 21409
rect 20073 21369 20085 21403
rect 20119 21400 20131 21403
rect 20714 21400 20720 21412
rect 20119 21372 20720 21400
rect 20119 21369 20131 21372
rect 20073 21363 20131 21369
rect 20714 21360 20720 21372
rect 20772 21360 20778 21412
rect 21545 21403 21603 21409
rect 21545 21369 21557 21403
rect 21591 21400 21603 21403
rect 21726 21400 21732 21412
rect 21591 21372 21732 21400
rect 21591 21369 21603 21372
rect 21545 21363 21603 21369
rect 21726 21360 21732 21372
rect 21784 21400 21790 21412
rect 22005 21403 22063 21409
rect 22005 21400 22017 21403
rect 21784 21372 22017 21400
rect 21784 21360 21790 21372
rect 22005 21369 22017 21372
rect 22051 21369 22063 21403
rect 22005 21363 22063 21369
rect 15473 21335 15531 21341
rect 15473 21301 15485 21335
rect 15519 21301 15531 21335
rect 15930 21332 15936 21344
rect 15891 21304 15936 21332
rect 15473 21295 15531 21301
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 16022 21292 16028 21344
rect 16080 21332 16086 21344
rect 16485 21335 16543 21341
rect 16485 21332 16497 21335
rect 16080 21304 16497 21332
rect 16080 21292 16086 21304
rect 16485 21301 16497 21304
rect 16531 21301 16543 21335
rect 16850 21332 16856 21344
rect 16811 21304 16856 21332
rect 16485 21295 16543 21301
rect 16850 21292 16856 21304
rect 16908 21292 16914 21344
rect 17126 21292 17132 21344
rect 17184 21332 17190 21344
rect 18325 21335 18383 21341
rect 18325 21332 18337 21335
rect 17184 21304 18337 21332
rect 17184 21292 17190 21304
rect 18325 21301 18337 21304
rect 18371 21301 18383 21335
rect 18325 21295 18383 21301
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19705 21335 19763 21341
rect 19705 21332 19717 21335
rect 19484 21304 19717 21332
rect 19484 21292 19490 21304
rect 19705 21301 19717 21304
rect 19751 21301 19763 21335
rect 19705 21295 19763 21301
rect 20165 21335 20223 21341
rect 20165 21301 20177 21335
rect 20211 21332 20223 21335
rect 20806 21332 20812 21344
rect 20211 21304 20812 21332
rect 20211 21301 20223 21304
rect 20165 21295 20223 21301
rect 20806 21292 20812 21304
rect 20864 21292 20870 21344
rect 21174 21332 21180 21344
rect 21135 21304 21180 21332
rect 21174 21292 21180 21304
rect 21232 21292 21238 21344
rect 1104 21242 22816 21264
rect 1104 21190 8246 21242
rect 8298 21190 8310 21242
rect 8362 21190 8374 21242
rect 8426 21190 8438 21242
rect 8490 21190 15510 21242
rect 15562 21190 15574 21242
rect 15626 21190 15638 21242
rect 15690 21190 15702 21242
rect 15754 21190 22816 21242
rect 1104 21168 22816 21190
rect 3513 21131 3571 21137
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 3602 21128 3608 21140
rect 3559 21100 3608 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 3602 21088 3608 21100
rect 3660 21088 3666 21140
rect 5074 21088 5080 21140
rect 5132 21128 5138 21140
rect 7101 21131 7159 21137
rect 7101 21128 7113 21131
rect 5132 21100 7113 21128
rect 5132 21088 5138 21100
rect 7101 21097 7113 21100
rect 7147 21097 7159 21131
rect 7101 21091 7159 21097
rect 8570 21088 8576 21140
rect 8628 21128 8634 21140
rect 9306 21128 9312 21140
rect 8628 21100 9312 21128
rect 8628 21088 8634 21100
rect 9306 21088 9312 21100
rect 9364 21088 9370 21140
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 14458 21128 14464 21140
rect 12308 21100 14464 21128
rect 12308 21088 12314 21100
rect 14458 21088 14464 21100
rect 14516 21088 14522 21140
rect 14829 21131 14887 21137
rect 14829 21097 14841 21131
rect 14875 21128 14887 21131
rect 14918 21128 14924 21140
rect 14875 21100 14924 21128
rect 14875 21097 14887 21100
rect 14829 21091 14887 21097
rect 14918 21088 14924 21100
rect 14976 21088 14982 21140
rect 15473 21131 15531 21137
rect 15473 21097 15485 21131
rect 15519 21128 15531 21131
rect 16574 21128 16580 21140
rect 15519 21100 16580 21128
rect 15519 21097 15531 21100
rect 15473 21091 15531 21097
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 17218 21128 17224 21140
rect 17179 21100 17224 21128
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 17678 21088 17684 21140
rect 17736 21128 17742 21140
rect 19702 21128 19708 21140
rect 17736 21100 19708 21128
rect 17736 21088 17742 21100
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 2400 21063 2458 21069
rect 2400 21029 2412 21063
rect 2446 21060 2458 21063
rect 2774 21060 2780 21072
rect 2446 21032 2780 21060
rect 2446 21029 2458 21032
rect 2400 21023 2458 21029
rect 2774 21020 2780 21032
rect 2832 21060 2838 21072
rect 3694 21060 3700 21072
rect 2832 21032 3700 21060
rect 2832 21020 2838 21032
rect 3694 21020 3700 21032
rect 3752 21020 3758 21072
rect 6457 21063 6515 21069
rect 4080 21032 6408 21060
rect 4080 21001 4108 21032
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20992 1639 20995
rect 4065 20995 4123 21001
rect 1627 20964 4016 20992
rect 1627 20961 1639 20964
rect 1581 20955 1639 20961
rect 2130 20924 2136 20936
rect 2091 20896 2136 20924
rect 2130 20884 2136 20896
rect 2188 20884 2194 20936
rect 3988 20924 4016 20964
rect 4065 20961 4077 20995
rect 4111 20961 4123 20995
rect 4065 20955 4123 20961
rect 5252 20995 5310 21001
rect 5252 20961 5264 20995
rect 5298 20992 5310 20995
rect 6178 20992 6184 21004
rect 5298 20964 6184 20992
rect 5298 20961 5310 20964
rect 5252 20955 5310 20961
rect 6178 20952 6184 20964
rect 6236 20952 6242 21004
rect 6380 20992 6408 21032
rect 6457 21029 6469 21063
rect 6503 21060 6515 21063
rect 7926 21060 7932 21072
rect 6503 21032 7932 21060
rect 6503 21029 6515 21032
rect 6457 21023 6515 21029
rect 7116 21004 7144 21032
rect 7926 21020 7932 21032
rect 7984 21020 7990 21072
rect 13164 21063 13222 21069
rect 13164 21029 13176 21063
rect 13210 21060 13222 21063
rect 13814 21060 13820 21072
rect 13210 21032 13820 21060
rect 13210 21029 13222 21032
rect 13164 21023 13222 21029
rect 13814 21020 13820 21032
rect 13872 21020 13878 21072
rect 16758 21060 16764 21072
rect 15304 21032 16764 21060
rect 6914 20992 6920 21004
rect 6380 20964 6920 20992
rect 6914 20952 6920 20964
rect 6972 20952 6978 21004
rect 7009 20995 7067 21001
rect 7009 20961 7021 20995
rect 7055 20961 7067 20995
rect 7009 20955 7067 20961
rect 4246 20924 4252 20936
rect 3988 20896 4252 20924
rect 4246 20884 4252 20896
rect 4304 20884 4310 20936
rect 4982 20924 4988 20936
rect 4943 20896 4988 20924
rect 4982 20884 4988 20896
rect 5040 20884 5046 20936
rect 6270 20884 6276 20936
rect 6328 20924 6334 20936
rect 7024 20924 7052 20955
rect 7098 20952 7104 21004
rect 7156 20952 7162 21004
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 8185 20995 8243 21001
rect 8185 20992 8197 20995
rect 7800 20964 8197 20992
rect 7800 20952 7806 20964
rect 8185 20961 8197 20964
rect 8231 20961 8243 20995
rect 10410 20992 10416 21004
rect 10371 20964 10416 20992
rect 8185 20955 8243 20961
rect 10410 20952 10416 20964
rect 10468 20952 10474 21004
rect 11324 20995 11382 21001
rect 11324 20961 11336 20995
rect 11370 20992 11382 20995
rect 12250 20992 12256 21004
rect 11370 20964 12256 20992
rect 11370 20961 11382 20964
rect 11324 20955 11382 20961
rect 12250 20952 12256 20964
rect 12308 20952 12314 21004
rect 14550 20952 14556 21004
rect 14608 20992 14614 21004
rect 15304 21001 15332 21032
rect 16758 21020 16764 21032
rect 16816 21020 16822 21072
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 19058 21060 19064 21072
rect 17920 21032 19064 21060
rect 17920 21020 17926 21032
rect 19058 21020 19064 21032
rect 19116 21020 19122 21072
rect 20717 21063 20775 21069
rect 20717 21029 20729 21063
rect 20763 21060 20775 21063
rect 20763 21032 21404 21060
rect 20763 21029 20775 21032
rect 20717 21023 20775 21029
rect 16114 21001 16120 21004
rect 14645 20995 14703 21001
rect 14645 20992 14657 20995
rect 14608 20964 14657 20992
rect 14608 20952 14614 20964
rect 14645 20961 14657 20964
rect 14691 20961 14703 20995
rect 14645 20955 14703 20961
rect 15289 20995 15347 21001
rect 15289 20961 15301 20995
rect 15335 20961 15347 20995
rect 15289 20955 15347 20961
rect 16108 20955 16120 21001
rect 16172 20992 16178 21004
rect 17764 20995 17822 21001
rect 16172 20964 16208 20992
rect 16114 20952 16120 20955
rect 16172 20952 16178 20964
rect 17764 20961 17776 20995
rect 17810 20992 17822 20995
rect 18322 20992 18328 21004
rect 17810 20964 18328 20992
rect 17810 20961 17822 20964
rect 17764 20955 17822 20961
rect 18322 20952 18328 20964
rect 18380 20952 18386 21004
rect 19420 20995 19478 21001
rect 19420 20961 19432 20995
rect 19466 20992 19478 20995
rect 20806 20992 20812 21004
rect 19466 20964 20812 20992
rect 19466 20961 19478 20964
rect 19420 20955 19478 20961
rect 20806 20952 20812 20964
rect 20864 20952 20870 21004
rect 20898 20952 20904 21004
rect 20956 20992 20962 21004
rect 21269 20995 21327 21001
rect 21269 20992 21281 20995
rect 20956 20964 21281 20992
rect 20956 20952 20962 20964
rect 21269 20961 21281 20964
rect 21315 20961 21327 20995
rect 21376 20992 21404 21032
rect 21913 20995 21971 21001
rect 21376 20964 21496 20992
rect 21269 20955 21327 20961
rect 6328 20896 7052 20924
rect 7193 20927 7251 20933
rect 6328 20884 6334 20896
rect 7193 20893 7205 20927
rect 7239 20893 7251 20927
rect 7193 20887 7251 20893
rect 7929 20927 7987 20933
rect 7929 20893 7941 20927
rect 7975 20893 7987 20927
rect 7929 20887 7987 20893
rect 7208 20856 7236 20887
rect 5920 20828 7236 20856
rect 1765 20791 1823 20797
rect 1765 20757 1777 20791
rect 1811 20788 1823 20791
rect 1946 20788 1952 20800
rect 1811 20760 1952 20788
rect 1811 20757 1823 20760
rect 1765 20751 1823 20757
rect 1946 20748 1952 20760
rect 2004 20748 2010 20800
rect 3878 20748 3884 20800
rect 3936 20788 3942 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 3936 20760 4261 20788
rect 3936 20748 3942 20760
rect 4249 20757 4261 20760
rect 4295 20757 4307 20791
rect 4249 20751 4307 20757
rect 5350 20748 5356 20800
rect 5408 20788 5414 20800
rect 5920 20788 5948 20828
rect 5408 20760 5948 20788
rect 6365 20791 6423 20797
rect 5408 20748 5414 20760
rect 6365 20757 6377 20791
rect 6411 20788 6423 20791
rect 6457 20791 6515 20797
rect 6457 20788 6469 20791
rect 6411 20760 6469 20788
rect 6411 20757 6423 20760
rect 6365 20751 6423 20757
rect 6457 20757 6469 20760
rect 6503 20757 6515 20791
rect 6638 20788 6644 20800
rect 6599 20760 6644 20788
rect 6457 20751 6515 20757
rect 6638 20748 6644 20760
rect 6696 20748 6702 20800
rect 7944 20788 7972 20887
rect 9766 20884 9772 20936
rect 9824 20924 9830 20936
rect 10505 20927 10563 20933
rect 10505 20924 10517 20927
rect 9824 20896 10517 20924
rect 9824 20884 9830 20896
rect 10505 20893 10517 20896
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10962 20924 10968 20936
rect 10735 20896 10968 20924
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 10962 20884 10968 20896
rect 11020 20884 11026 20936
rect 11057 20927 11115 20933
rect 11057 20893 11069 20927
rect 11103 20893 11115 20927
rect 11057 20887 11115 20893
rect 10594 20816 10600 20868
rect 10652 20856 10658 20868
rect 11072 20856 11100 20887
rect 12526 20884 12532 20936
rect 12584 20924 12590 20936
rect 12897 20927 12955 20933
rect 12897 20924 12909 20927
rect 12584 20896 12909 20924
rect 12584 20884 12590 20896
rect 12897 20893 12909 20896
rect 12943 20893 12955 20927
rect 12897 20887 12955 20893
rect 15841 20927 15899 20933
rect 15841 20893 15853 20927
rect 15887 20893 15899 20927
rect 17497 20927 17555 20933
rect 17497 20924 17509 20927
rect 15841 20887 15899 20893
rect 17420 20896 17509 20924
rect 10652 20828 11100 20856
rect 10652 20816 10658 20828
rect 8570 20788 8576 20800
rect 7944 20760 8576 20788
rect 8570 20748 8576 20760
rect 8628 20748 8634 20800
rect 9309 20791 9367 20797
rect 9309 20757 9321 20791
rect 9355 20788 9367 20791
rect 9490 20788 9496 20800
rect 9355 20760 9496 20788
rect 9355 20757 9367 20760
rect 9309 20751 9367 20757
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 10045 20791 10103 20797
rect 10045 20757 10057 20791
rect 10091 20788 10103 20791
rect 10778 20788 10784 20800
rect 10091 20760 10784 20788
rect 10091 20757 10103 20760
rect 10045 20751 10103 20757
rect 10778 20748 10784 20760
rect 10836 20748 10842 20800
rect 12434 20748 12440 20800
rect 12492 20788 12498 20800
rect 12492 20760 12537 20788
rect 12492 20748 12498 20760
rect 13906 20748 13912 20800
rect 13964 20788 13970 20800
rect 14277 20791 14335 20797
rect 14277 20788 14289 20791
rect 13964 20760 14289 20788
rect 13964 20748 13970 20760
rect 14277 20757 14289 20760
rect 14323 20788 14335 20791
rect 15470 20788 15476 20800
rect 14323 20760 15476 20788
rect 14323 20757 14335 20760
rect 14277 20751 14335 20757
rect 15470 20748 15476 20760
rect 15528 20748 15534 20800
rect 15856 20788 15884 20887
rect 16942 20788 16948 20800
rect 15856 20760 16948 20788
rect 16942 20748 16948 20760
rect 17000 20788 17006 20800
rect 17420 20788 17448 20896
rect 17497 20893 17509 20896
rect 17543 20893 17555 20927
rect 17497 20887 17555 20893
rect 18966 20884 18972 20936
rect 19024 20924 19030 20936
rect 19153 20927 19211 20933
rect 19153 20924 19165 20927
rect 19024 20896 19165 20924
rect 19024 20884 19030 20896
rect 19153 20893 19165 20896
rect 19199 20893 19211 20927
rect 20717 20927 20775 20933
rect 20717 20924 20729 20927
rect 19153 20887 19211 20893
rect 20180 20896 20729 20924
rect 18690 20816 18696 20868
rect 18748 20856 18754 20868
rect 18748 20828 19196 20856
rect 18748 20816 18754 20828
rect 17000 20760 17448 20788
rect 17000 20748 17006 20760
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 18877 20791 18935 20797
rect 18877 20788 18889 20791
rect 18472 20760 18889 20788
rect 18472 20748 18478 20760
rect 18877 20757 18889 20760
rect 18923 20757 18935 20791
rect 19168 20788 19196 20828
rect 20180 20788 20208 20896
rect 20717 20893 20729 20896
rect 20763 20893 20775 20927
rect 21358 20924 21364 20936
rect 21319 20896 21364 20924
rect 20717 20887 20775 20893
rect 21358 20884 21364 20896
rect 21416 20884 21422 20936
rect 21468 20933 21496 20964
rect 21913 20961 21925 20995
rect 21959 20961 21971 20995
rect 21913 20955 21971 20961
rect 21453 20927 21511 20933
rect 21453 20893 21465 20927
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 21928 20856 21956 20955
rect 21324 20828 21956 20856
rect 21324 20816 21330 20828
rect 19168 20760 20208 20788
rect 20533 20791 20591 20797
rect 18877 20751 18935 20757
rect 20533 20757 20545 20791
rect 20579 20788 20591 20791
rect 20714 20788 20720 20800
rect 20579 20760 20720 20788
rect 20579 20757 20591 20760
rect 20533 20751 20591 20757
rect 20714 20748 20720 20760
rect 20772 20748 20778 20800
rect 20901 20791 20959 20797
rect 20901 20757 20913 20791
rect 20947 20788 20959 20791
rect 20990 20788 20996 20800
rect 20947 20760 20996 20788
rect 20947 20757 20959 20760
rect 20901 20751 20959 20757
rect 20990 20748 20996 20760
rect 21048 20748 21054 20800
rect 22094 20748 22100 20800
rect 22152 20788 22158 20800
rect 22152 20760 22197 20788
rect 22152 20748 22158 20760
rect 1104 20698 22816 20720
rect 1104 20646 4614 20698
rect 4666 20646 4678 20698
rect 4730 20646 4742 20698
rect 4794 20646 4806 20698
rect 4858 20646 11878 20698
rect 11930 20646 11942 20698
rect 11994 20646 12006 20698
rect 12058 20646 12070 20698
rect 12122 20646 19142 20698
rect 19194 20646 19206 20698
rect 19258 20646 19270 20698
rect 19322 20646 19334 20698
rect 19386 20646 22816 20698
rect 1104 20624 22816 20646
rect 2774 20544 2780 20596
rect 2832 20584 2838 20596
rect 2832 20556 2877 20584
rect 2832 20544 2838 20556
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 3786 20584 3792 20596
rect 3016 20556 3792 20584
rect 3016 20544 3022 20556
rect 3786 20544 3792 20556
rect 3844 20544 3850 20596
rect 4062 20544 4068 20596
rect 4120 20544 4126 20596
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 5902 20584 5908 20596
rect 4304 20556 5908 20584
rect 4304 20544 4310 20556
rect 5902 20544 5908 20556
rect 5960 20544 5966 20596
rect 8018 20584 8024 20596
rect 6012 20556 8024 20584
rect 4080 20516 4108 20544
rect 4798 20516 4804 20528
rect 4080 20488 4804 20516
rect 4798 20476 4804 20488
rect 4856 20476 4862 20528
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1486 20380 1492 20392
rect 1443 20352 1492 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1486 20340 1492 20352
rect 1544 20380 1550 20392
rect 2130 20380 2136 20392
rect 1544 20352 2136 20380
rect 1544 20340 1550 20352
rect 2130 20340 2136 20352
rect 2188 20380 2194 20392
rect 3145 20383 3203 20389
rect 3145 20380 3157 20383
rect 2188 20352 3157 20380
rect 2188 20340 2194 20352
rect 3145 20349 3157 20352
rect 3191 20380 3203 20383
rect 4801 20383 4859 20389
rect 4801 20380 4813 20383
rect 3191 20352 4813 20380
rect 3191 20349 3203 20352
rect 3145 20343 3203 20349
rect 4801 20349 4813 20352
rect 4847 20380 4859 20383
rect 4890 20380 4896 20392
rect 4847 20352 4896 20380
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 4890 20340 4896 20352
rect 4948 20340 4954 20392
rect 5068 20383 5126 20389
rect 5068 20349 5080 20383
rect 5114 20380 5126 20383
rect 5350 20380 5356 20392
rect 5114 20352 5356 20380
rect 5114 20349 5126 20352
rect 5068 20343 5126 20349
rect 5350 20340 5356 20352
rect 5408 20340 5414 20392
rect 5442 20340 5448 20392
rect 5500 20380 5506 20392
rect 6012 20380 6040 20556
rect 8018 20544 8024 20556
rect 8076 20544 8082 20596
rect 8110 20544 8116 20596
rect 8168 20584 8174 20596
rect 8205 20587 8263 20593
rect 8205 20584 8217 20587
rect 8168 20556 8217 20584
rect 8168 20544 8174 20556
rect 8205 20553 8217 20556
rect 8251 20553 8263 20587
rect 11330 20584 11336 20596
rect 8205 20547 8263 20553
rect 8312 20556 11336 20584
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7098 20389 7104 20392
rect 7092 20380 7104 20389
rect 5500 20352 6040 20380
rect 7059 20352 7104 20380
rect 5500 20340 5506 20352
rect 7092 20343 7104 20352
rect 7098 20340 7104 20343
rect 7156 20340 7162 20392
rect 1664 20315 1722 20321
rect 1664 20281 1676 20315
rect 1710 20312 1722 20315
rect 2958 20312 2964 20324
rect 1710 20284 2964 20312
rect 1710 20281 1722 20284
rect 1664 20275 1722 20281
rect 2958 20272 2964 20284
rect 3016 20272 3022 20324
rect 3412 20315 3470 20321
rect 3412 20281 3424 20315
rect 3458 20312 3470 20315
rect 3602 20312 3608 20324
rect 3458 20284 3608 20312
rect 3458 20281 3470 20284
rect 3412 20275 3470 20281
rect 3602 20272 3608 20284
rect 3660 20272 3666 20324
rect 4430 20272 4436 20324
rect 4488 20312 4494 20324
rect 8312 20312 8340 20556
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 11606 20544 11612 20596
rect 11664 20544 11670 20596
rect 12069 20587 12127 20593
rect 12069 20553 12081 20587
rect 12115 20584 12127 20587
rect 12250 20584 12256 20596
rect 12115 20556 12256 20584
rect 12115 20553 12127 20556
rect 12069 20547 12127 20553
rect 12250 20544 12256 20556
rect 12308 20544 12314 20596
rect 13814 20584 13820 20596
rect 12452 20556 13400 20584
rect 13727 20556 13820 20584
rect 11624 20516 11652 20544
rect 12452 20516 12480 20556
rect 11624 20488 12480 20516
rect 13372 20516 13400 20556
rect 13814 20544 13820 20556
rect 13872 20584 13878 20596
rect 13872 20556 17080 20584
rect 13872 20544 13878 20556
rect 14734 20516 14740 20528
rect 13372 20488 14740 20516
rect 14734 20476 14740 20488
rect 14792 20476 14798 20528
rect 16114 20476 16120 20528
rect 16172 20516 16178 20528
rect 16301 20519 16359 20525
rect 16301 20516 16313 20519
rect 16172 20488 16313 20516
rect 16172 20476 16178 20488
rect 16301 20485 16313 20488
rect 16347 20516 16359 20519
rect 16390 20516 16396 20528
rect 16347 20488 16396 20516
rect 16347 20485 16359 20488
rect 16301 20479 16359 20485
rect 16390 20476 16396 20488
rect 16448 20476 16454 20528
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 17052 20457 17080 20556
rect 20806 20544 20812 20596
rect 20864 20584 20870 20596
rect 20901 20587 20959 20593
rect 20901 20584 20913 20587
rect 20864 20556 20913 20584
rect 20864 20544 20870 20556
rect 20901 20553 20913 20556
rect 20947 20553 20959 20587
rect 20901 20547 20959 20553
rect 18966 20476 18972 20528
rect 19024 20516 19030 20528
rect 19024 20488 19380 20516
rect 19024 20476 19030 20488
rect 19352 20460 19380 20488
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 9732 20420 10241 20448
rect 9732 20408 9738 20420
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 17037 20451 17095 20457
rect 10229 20411 10287 20417
rect 14384 20420 15056 20448
rect 8570 20380 8576 20392
rect 8483 20352 8576 20380
rect 8570 20340 8576 20352
rect 8628 20380 8634 20392
rect 9122 20380 9128 20392
rect 8628 20352 9128 20380
rect 8628 20340 8634 20352
rect 9122 20340 9128 20352
rect 9180 20380 9186 20392
rect 9582 20380 9588 20392
rect 9180 20352 9588 20380
rect 9180 20340 9186 20352
rect 9582 20340 9588 20352
rect 9640 20380 9646 20392
rect 10594 20380 10600 20392
rect 9640 20352 10600 20380
rect 9640 20340 9646 20352
rect 10594 20340 10600 20352
rect 10652 20380 10658 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10652 20352 10701 20380
rect 10652 20340 10658 20352
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 12158 20380 12164 20392
rect 10689 20343 10747 20349
rect 10796 20352 12164 20380
rect 4488 20284 8340 20312
rect 8840 20315 8898 20321
rect 4488 20272 4494 20284
rect 8840 20281 8852 20315
rect 8886 20312 8898 20315
rect 9490 20312 9496 20324
rect 8886 20284 9496 20312
rect 8886 20281 8898 20284
rect 8840 20275 8898 20281
rect 9490 20272 9496 20284
rect 9548 20272 9554 20324
rect 10796 20312 10824 20352
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 12526 20380 12532 20392
rect 12483 20352 12532 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 12526 20340 12532 20352
rect 12584 20340 12590 20392
rect 14384 20389 14412 20420
rect 15028 20392 15056 20420
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17221 20451 17279 20457
rect 17221 20417 17233 20451
rect 17267 20448 17279 20451
rect 17310 20448 17316 20460
rect 17267 20420 17316 20448
rect 17267 20417 17279 20420
rect 17221 20411 17279 20417
rect 17310 20408 17316 20420
rect 17368 20448 17374 20460
rect 17494 20448 17500 20460
rect 17368 20420 17500 20448
rect 17368 20408 17374 20420
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19061 20451 19119 20457
rect 19061 20448 19073 20451
rect 18748 20420 19073 20448
rect 18748 20408 18754 20420
rect 19061 20417 19073 20420
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 19334 20408 19340 20460
rect 19392 20448 19398 20460
rect 19521 20451 19579 20457
rect 19521 20448 19533 20451
rect 19392 20420 19533 20448
rect 19392 20408 19398 20420
rect 19521 20417 19533 20420
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 21450 20448 21456 20460
rect 20588 20420 21456 20448
rect 20588 20408 20594 20420
rect 21450 20408 21456 20420
rect 21508 20448 21514 20460
rect 21729 20451 21787 20457
rect 21729 20448 21741 20451
rect 21508 20420 21741 20448
rect 21508 20408 21514 20420
rect 21729 20417 21741 20420
rect 21775 20417 21787 20451
rect 21729 20411 21787 20417
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20349 14427 20383
rect 14918 20380 14924 20392
rect 14879 20352 14924 20380
rect 14369 20343 14427 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 15010 20340 15016 20392
rect 15068 20340 15074 20392
rect 15194 20389 15200 20392
rect 15188 20380 15200 20389
rect 15155 20352 15200 20380
rect 15188 20343 15200 20352
rect 15194 20340 15200 20343
rect 15252 20340 15258 20392
rect 15470 20340 15476 20392
rect 15528 20380 15534 20392
rect 16945 20383 17003 20389
rect 16945 20380 16957 20383
rect 15528 20352 16957 20380
rect 15528 20340 15534 20352
rect 16945 20349 16957 20352
rect 16991 20349 17003 20383
rect 16945 20343 17003 20349
rect 18049 20383 18107 20389
rect 18049 20349 18061 20383
rect 18095 20380 18107 20383
rect 18506 20380 18512 20392
rect 18095 20352 18512 20380
rect 18095 20349 18107 20352
rect 18049 20343 18107 20349
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20380 18935 20383
rect 19426 20380 19432 20392
rect 18923 20352 19432 20380
rect 18923 20349 18935 20352
rect 18877 20343 18935 20349
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 19788 20383 19846 20389
rect 19788 20349 19800 20383
rect 19834 20380 19846 20383
rect 19834 20352 21588 20380
rect 19834 20349 19846 20352
rect 19788 20343 19846 20349
rect 10962 20321 10968 20324
rect 10956 20312 10968 20321
rect 9784 20284 10824 20312
rect 10923 20284 10968 20312
rect 2406 20204 2412 20256
rect 2464 20244 2470 20256
rect 4154 20244 4160 20256
rect 2464 20216 4160 20244
rect 2464 20204 2470 20216
rect 4154 20204 4160 20216
rect 4212 20204 4218 20256
rect 4525 20247 4583 20253
rect 4525 20213 4537 20247
rect 4571 20244 4583 20247
rect 5350 20244 5356 20256
rect 4571 20216 5356 20244
rect 4571 20213 4583 20216
rect 4525 20207 4583 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 6178 20244 6184 20256
rect 6139 20216 6184 20244
rect 6178 20204 6184 20216
rect 6236 20204 6242 20256
rect 8662 20204 8668 20256
rect 8720 20244 8726 20256
rect 9784 20244 9812 20284
rect 10956 20275 10968 20284
rect 10962 20272 10968 20275
rect 11020 20272 11026 20324
rect 12710 20321 12716 20324
rect 12704 20275 12716 20321
rect 12768 20312 12774 20324
rect 12768 20284 12804 20312
rect 12710 20272 12716 20275
rect 12768 20272 12774 20284
rect 16850 20272 16856 20324
rect 16908 20312 16914 20324
rect 19978 20312 19984 20324
rect 16908 20284 19984 20312
rect 16908 20272 16914 20284
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 20088 20284 21220 20312
rect 9950 20244 9956 20256
rect 8720 20216 9812 20244
rect 9911 20216 9956 20244
rect 8720 20204 8726 20216
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 11330 20204 11336 20256
rect 11388 20244 11394 20256
rect 12802 20244 12808 20256
rect 11388 20216 12808 20244
rect 11388 20204 11394 20216
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14553 20247 14611 20253
rect 14553 20244 14565 20247
rect 14332 20216 14565 20244
rect 14332 20204 14338 20216
rect 14553 20213 14565 20216
rect 14599 20213 14611 20247
rect 14553 20207 14611 20213
rect 16390 20204 16396 20256
rect 16448 20244 16454 20256
rect 16577 20247 16635 20253
rect 16577 20244 16589 20247
rect 16448 20216 16589 20244
rect 16448 20204 16454 20216
rect 16577 20213 16589 20216
rect 16623 20213 16635 20247
rect 16577 20207 16635 20213
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 18782 20244 18788 20256
rect 18555 20216 18788 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 18782 20204 18788 20216
rect 18840 20204 18846 20256
rect 18969 20247 19027 20253
rect 18969 20213 18981 20247
rect 19015 20244 19027 20247
rect 20088 20244 20116 20284
rect 21192 20253 21220 20284
rect 21560 20256 21588 20352
rect 19015 20216 20116 20244
rect 21177 20247 21235 20253
rect 19015 20213 19027 20216
rect 18969 20207 19027 20213
rect 21177 20213 21189 20247
rect 21223 20213 21235 20247
rect 21542 20244 21548 20256
rect 21503 20216 21548 20244
rect 21177 20207 21235 20213
rect 21542 20204 21548 20216
rect 21600 20204 21606 20256
rect 21634 20204 21640 20256
rect 21692 20244 21698 20256
rect 21692 20216 21737 20244
rect 21692 20204 21698 20216
rect 1104 20154 22816 20176
rect 1104 20102 8246 20154
rect 8298 20102 8310 20154
rect 8362 20102 8374 20154
rect 8426 20102 8438 20154
rect 8490 20102 15510 20154
rect 15562 20102 15574 20154
rect 15626 20102 15638 20154
rect 15690 20102 15702 20154
rect 15754 20102 22816 20154
rect 1104 20080 22816 20102
rect 2406 20040 2412 20052
rect 2367 20012 2412 20040
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 3234 20000 3240 20052
rect 3292 20040 3298 20052
rect 3605 20043 3663 20049
rect 3605 20040 3617 20043
rect 3292 20012 3617 20040
rect 3292 20000 3298 20012
rect 3605 20009 3617 20012
rect 3651 20009 3663 20043
rect 3605 20003 3663 20009
rect 4065 20043 4123 20049
rect 4065 20009 4077 20043
rect 4111 20040 4123 20043
rect 5537 20043 5595 20049
rect 5537 20040 5549 20043
rect 4111 20012 5549 20040
rect 4111 20009 4123 20012
rect 4065 20003 4123 20009
rect 5537 20009 5549 20012
rect 5583 20009 5595 20043
rect 5537 20003 5595 20009
rect 6178 20000 6184 20052
rect 6236 20040 6242 20052
rect 8481 20043 8539 20049
rect 6236 20012 7788 20040
rect 6236 20000 6242 20012
rect 2777 19975 2835 19981
rect 2777 19941 2789 19975
rect 2823 19972 2835 19975
rect 4246 19972 4252 19984
rect 2823 19944 4252 19972
rect 2823 19941 2835 19944
rect 2777 19935 2835 19941
rect 4246 19932 4252 19944
rect 4304 19932 4310 19984
rect 4798 19932 4804 19984
rect 4856 19972 4862 19984
rect 6086 19972 6092 19984
rect 4856 19944 6092 19972
rect 4856 19932 4862 19944
rect 6086 19932 6092 19944
rect 6144 19932 6150 19984
rect 7760 19972 7788 20012
rect 8481 20009 8493 20043
rect 8527 20040 8539 20043
rect 9030 20040 9036 20052
rect 8527 20012 9036 20040
rect 8527 20009 8539 20012
rect 8481 20003 8539 20009
rect 9030 20000 9036 20012
rect 9088 20000 9094 20052
rect 10137 20043 10195 20049
rect 10137 20009 10149 20043
rect 10183 20040 10195 20043
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 10183 20012 13001 20040
rect 10183 20009 10195 20012
rect 10137 20003 10195 20009
rect 12989 20009 13001 20012
rect 13035 20009 13047 20043
rect 12989 20003 13047 20009
rect 14921 20043 14979 20049
rect 14921 20009 14933 20043
rect 14967 20040 14979 20043
rect 15194 20040 15200 20052
rect 14967 20012 15200 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15194 20000 15200 20012
rect 15252 20000 15258 20052
rect 15289 20043 15347 20049
rect 15289 20009 15301 20043
rect 15335 20009 15347 20043
rect 15289 20003 15347 20009
rect 7760 19944 9076 19972
rect 1762 19904 1768 19916
rect 1723 19876 1768 19904
rect 1762 19864 1768 19876
rect 1820 19864 1826 19916
rect 2866 19904 2872 19916
rect 2827 19876 2872 19904
rect 2866 19864 2872 19876
rect 2924 19864 2930 19916
rect 3418 19904 3424 19916
rect 3379 19876 3424 19904
rect 3418 19864 3424 19876
rect 3476 19864 3482 19916
rect 3602 19864 3608 19916
rect 3660 19904 3666 19916
rect 4433 19907 4491 19913
rect 4433 19904 4445 19907
rect 3660 19876 4445 19904
rect 3660 19864 3666 19876
rect 4433 19873 4445 19876
rect 4479 19873 4491 19907
rect 5445 19907 5503 19913
rect 5445 19904 5457 19907
rect 4433 19867 4491 19873
rect 4816 19876 5457 19904
rect 1854 19836 1860 19848
rect 1815 19808 1860 19836
rect 1854 19796 1860 19808
rect 1912 19796 1918 19848
rect 1946 19796 1952 19848
rect 2004 19836 2010 19848
rect 2406 19836 2412 19848
rect 2004 19808 2412 19836
rect 2004 19796 2010 19808
rect 2406 19796 2412 19808
rect 2464 19796 2470 19848
rect 2958 19836 2964 19848
rect 2919 19808 2964 19836
rect 2958 19796 2964 19808
rect 3016 19796 3022 19848
rect 3694 19796 3700 19848
rect 3752 19836 3758 19848
rect 4525 19839 4583 19845
rect 4525 19836 4537 19839
rect 3752 19808 4537 19836
rect 3752 19796 3758 19808
rect 4525 19805 4537 19808
rect 4571 19805 4583 19839
rect 4525 19799 4583 19805
rect 4614 19796 4620 19848
rect 4672 19836 4678 19848
rect 4672 19808 4717 19836
rect 4672 19796 4678 19808
rect 1397 19771 1455 19777
rect 1397 19737 1409 19771
rect 1443 19768 1455 19771
rect 4816 19768 4844 19876
rect 5445 19873 5457 19876
rect 5491 19873 5503 19907
rect 8662 19904 8668 19916
rect 5445 19867 5503 19873
rect 7024 19876 8668 19904
rect 5074 19796 5080 19848
rect 5132 19836 5138 19848
rect 5350 19836 5356 19848
rect 5132 19808 5356 19836
rect 5132 19796 5138 19808
rect 5350 19796 5356 19808
rect 5408 19836 5414 19848
rect 5629 19839 5687 19845
rect 5629 19836 5641 19839
rect 5408 19808 5641 19836
rect 5408 19796 5414 19808
rect 5629 19805 5641 19808
rect 5675 19805 5687 19839
rect 5629 19799 5687 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 6546 19836 6552 19848
rect 6411 19808 6552 19836
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 6546 19796 6552 19808
rect 6604 19796 6610 19848
rect 6730 19845 6736 19848
rect 6688 19839 6736 19845
rect 6688 19805 6700 19839
rect 6734 19805 6736 19839
rect 6688 19799 6736 19805
rect 6730 19796 6736 19799
rect 6788 19796 6794 19848
rect 6871 19839 6929 19845
rect 6871 19805 6883 19839
rect 6917 19836 6929 19839
rect 7024 19836 7052 19876
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 8846 19904 8852 19916
rect 8807 19876 8852 19904
rect 8846 19864 8852 19876
rect 8904 19864 8910 19916
rect 6917 19808 7052 19836
rect 6917 19805 6929 19808
rect 6871 19799 6929 19805
rect 7098 19796 7104 19848
rect 7156 19836 7162 19848
rect 9048 19845 9076 19944
rect 12158 19932 12164 19984
rect 12216 19972 12222 19984
rect 15304 19972 15332 20003
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15749 20043 15807 20049
rect 15749 20040 15761 20043
rect 15436 20012 15761 20040
rect 15436 20000 15442 20012
rect 15749 20009 15761 20012
rect 15795 20009 15807 20043
rect 15749 20003 15807 20009
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 15988 20012 16252 20040
rect 15988 20000 15994 20012
rect 12216 19944 15332 19972
rect 12216 19932 12222 19944
rect 15838 19932 15844 19984
rect 15896 19932 15902 19984
rect 10045 19907 10103 19913
rect 10045 19873 10057 19907
rect 10091 19904 10103 19907
rect 12066 19904 12072 19916
rect 10091 19876 12072 19904
rect 10091 19873 10103 19876
rect 10045 19867 10103 19873
rect 12066 19864 12072 19876
rect 12124 19864 12130 19916
rect 12805 19907 12863 19913
rect 12805 19904 12817 19907
rect 12176 19876 12817 19904
rect 8941 19839 8999 19845
rect 8941 19836 8953 19839
rect 7156 19808 7201 19836
rect 8855 19808 8953 19836
rect 7156 19796 7162 19808
rect 1443 19740 4844 19768
rect 1443 19737 1455 19740
rect 1397 19731 1455 19737
rect 3510 19660 3516 19712
rect 3568 19700 3574 19712
rect 5077 19703 5135 19709
rect 5077 19700 5089 19703
rect 3568 19672 5089 19700
rect 3568 19660 3574 19672
rect 5077 19669 5089 19672
rect 5123 19669 5135 19703
rect 5077 19663 5135 19669
rect 5258 19660 5264 19712
rect 5316 19700 5322 19712
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 5316 19672 8217 19700
rect 5316 19660 5322 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 8205 19663 8263 19669
rect 8662 19660 8668 19712
rect 8720 19700 8726 19712
rect 8855 19700 8883 19808
rect 8941 19805 8953 19808
rect 8987 19805 8999 19839
rect 8941 19799 8999 19805
rect 9033 19839 9091 19845
rect 9033 19805 9045 19839
rect 9079 19805 9091 19839
rect 10318 19836 10324 19848
rect 10279 19808 10324 19836
rect 9033 19799 9091 19805
rect 10318 19796 10324 19808
rect 10376 19796 10382 19848
rect 10594 19796 10600 19848
rect 10652 19836 10658 19848
rect 11054 19845 11060 19848
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 10652 19808 10701 19836
rect 10652 19796 10658 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 11012 19839 11060 19845
rect 11012 19805 11024 19839
rect 11058 19805 11060 19839
rect 11012 19799 11060 19805
rect 11054 19796 11060 19799
rect 11112 19796 11118 19848
rect 11238 19845 11244 19848
rect 11195 19839 11244 19845
rect 11195 19805 11207 19839
rect 11241 19805 11244 19839
rect 11195 19799 11244 19805
rect 11238 19796 11244 19799
rect 11296 19796 11302 19848
rect 11422 19836 11428 19848
rect 11383 19808 11428 19836
rect 11422 19796 11428 19808
rect 11480 19796 11486 19848
rect 11606 19796 11612 19848
rect 11664 19836 11670 19848
rect 12176 19836 12204 19876
rect 12805 19873 12817 19876
rect 12851 19873 12863 19907
rect 12805 19867 12863 19873
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 13808 19907 13866 19913
rect 12952 19876 13584 19904
rect 12952 19864 12958 19876
rect 13556 19848 13584 19876
rect 13808 19873 13820 19907
rect 13854 19904 13866 19907
rect 14826 19904 14832 19916
rect 13854 19876 14832 19904
rect 13854 19873 13866 19876
rect 13808 19867 13866 19873
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 15657 19907 15715 19913
rect 15657 19873 15669 19907
rect 15703 19904 15715 19907
rect 15856 19904 15884 19932
rect 16117 19907 16175 19913
rect 16117 19904 16129 19907
rect 15703 19876 16129 19904
rect 15703 19873 15715 19876
rect 15657 19867 15715 19873
rect 16117 19873 16129 19876
rect 16163 19873 16175 19907
rect 16224 19904 16252 20012
rect 16482 20000 16488 20052
rect 16540 20000 16546 20052
rect 16669 20043 16727 20049
rect 16669 20009 16681 20043
rect 16715 20040 16727 20043
rect 18322 20040 18328 20052
rect 16715 20012 18184 20040
rect 18283 20012 18328 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 16301 19975 16359 19981
rect 16301 19941 16313 19975
rect 16347 19972 16359 19975
rect 16500 19972 16528 20000
rect 17218 19981 17224 19984
rect 17212 19972 17224 19981
rect 16347 19944 16528 19972
rect 17179 19944 17224 19972
rect 16347 19941 16359 19944
rect 16301 19935 16359 19941
rect 17212 19935 17224 19944
rect 17218 19932 17224 19935
rect 17276 19932 17282 19984
rect 18156 19972 18184 20012
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18785 20043 18843 20049
rect 18785 20009 18797 20043
rect 18831 20040 18843 20043
rect 19518 20040 19524 20052
rect 18831 20012 19524 20040
rect 18831 20009 18843 20012
rect 18785 20003 18843 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 20533 20043 20591 20049
rect 20533 20009 20545 20043
rect 20579 20040 20591 20043
rect 21542 20040 21548 20052
rect 20579 20012 21548 20040
rect 20579 20009 20591 20012
rect 20533 20003 20591 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 20254 19972 20260 19984
rect 18156 19944 20260 19972
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 20714 19932 20720 19984
rect 20772 19972 20778 19984
rect 21146 19975 21204 19981
rect 21146 19972 21158 19975
rect 20772 19944 21158 19972
rect 20772 19932 20778 19944
rect 21146 19941 21158 19944
rect 21192 19941 21204 19975
rect 21146 19935 21204 19941
rect 16485 19907 16543 19913
rect 16485 19904 16497 19907
rect 16224 19876 16497 19904
rect 16117 19867 16175 19873
rect 16485 19873 16497 19876
rect 16531 19904 16543 19907
rect 18598 19904 18604 19916
rect 16531 19876 18092 19904
rect 18559 19876 18604 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 11664 19808 12204 19836
rect 11664 19796 11670 19808
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 13446 19836 13452 19848
rect 12584 19808 13452 19836
rect 12584 19796 12590 19808
rect 13446 19796 13452 19808
rect 13504 19796 13510 19848
rect 13538 19796 13544 19848
rect 13596 19836 13602 19848
rect 13596 19808 13641 19836
rect 13596 19796 13602 19808
rect 14642 19796 14648 19848
rect 14700 19836 14706 19848
rect 15562 19836 15568 19848
rect 14700 19808 15568 19836
rect 14700 19796 14706 19808
rect 15562 19796 15568 19808
rect 15620 19796 15626 19848
rect 15841 19839 15899 19845
rect 15841 19805 15853 19839
rect 15887 19805 15899 19839
rect 16942 19836 16948 19848
rect 16903 19808 16948 19836
rect 15841 19799 15899 19805
rect 9214 19728 9220 19780
rect 9272 19768 9278 19780
rect 10502 19768 10508 19780
rect 9272 19740 10508 19768
rect 9272 19728 9278 19740
rect 10502 19728 10508 19740
rect 10560 19728 10566 19780
rect 15856 19768 15884 19799
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 14476 19740 15884 19768
rect 8720 19672 8883 19700
rect 9677 19703 9735 19709
rect 8720 19660 8726 19672
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 9766 19700 9772 19712
rect 9723 19672 9772 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 12526 19700 12532 19712
rect 12487 19672 12532 19700
rect 12526 19660 12532 19672
rect 12584 19660 12590 19712
rect 12618 19660 12624 19712
rect 12676 19700 12682 19712
rect 14476 19700 14504 19740
rect 12676 19672 14504 19700
rect 12676 19660 12682 19672
rect 14734 19660 14740 19712
rect 14792 19700 14798 19712
rect 16574 19700 16580 19712
rect 14792 19672 16580 19700
rect 14792 19660 14798 19672
rect 16574 19660 16580 19672
rect 16632 19660 16638 19712
rect 18064 19700 18092 19876
rect 18598 19864 18604 19876
rect 18656 19864 18662 19916
rect 19153 19907 19211 19913
rect 19153 19873 19165 19907
rect 19199 19904 19211 19907
rect 19242 19904 19248 19916
rect 19199 19876 19248 19904
rect 19199 19873 19211 19876
rect 19153 19867 19211 19873
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 19420 19907 19478 19913
rect 19420 19873 19432 19907
rect 19466 19904 19478 19907
rect 20806 19904 20812 19916
rect 19466 19876 20812 19904
rect 19466 19873 19478 19876
rect 19420 19867 19478 19873
rect 20806 19864 20812 19876
rect 20864 19864 20870 19916
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 20901 19839 20959 19845
rect 20901 19836 20913 19839
rect 20404 19808 20913 19836
rect 20404 19796 20410 19808
rect 20901 19805 20913 19808
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 22281 19703 22339 19709
rect 22281 19700 22293 19703
rect 18064 19672 22293 19700
rect 22281 19669 22293 19672
rect 22327 19669 22339 19703
rect 22281 19663 22339 19669
rect 1104 19610 22816 19632
rect 1104 19558 4614 19610
rect 4666 19558 4678 19610
rect 4730 19558 4742 19610
rect 4794 19558 4806 19610
rect 4858 19558 11878 19610
rect 11930 19558 11942 19610
rect 11994 19558 12006 19610
rect 12058 19558 12070 19610
rect 12122 19558 19142 19610
rect 19194 19558 19206 19610
rect 19258 19558 19270 19610
rect 19322 19558 19334 19610
rect 19386 19558 22816 19610
rect 1104 19536 22816 19558
rect 2314 19456 2320 19508
rect 2372 19456 2378 19508
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19496 2835 19499
rect 2958 19496 2964 19508
rect 2823 19468 2964 19496
rect 2823 19465 2835 19468
rect 2777 19459 2835 19465
rect 2958 19456 2964 19468
rect 3016 19456 3022 19508
rect 3050 19456 3056 19508
rect 3108 19496 3114 19508
rect 4154 19496 4160 19508
rect 3108 19468 4160 19496
rect 3108 19456 3114 19468
rect 4154 19456 4160 19468
rect 4212 19456 4218 19508
rect 4430 19456 4436 19508
rect 4488 19496 4494 19508
rect 4982 19496 4988 19508
rect 4488 19468 4988 19496
rect 4488 19456 4494 19468
rect 4982 19456 4988 19468
rect 5040 19456 5046 19508
rect 5166 19456 5172 19508
rect 5224 19496 5230 19508
rect 6178 19496 6184 19508
rect 5224 19468 6184 19496
rect 5224 19456 5230 19468
rect 6178 19456 6184 19468
rect 6236 19456 6242 19508
rect 6273 19499 6331 19505
rect 6273 19465 6285 19499
rect 6319 19496 6331 19499
rect 6362 19496 6368 19508
rect 6319 19468 6368 19496
rect 6319 19465 6331 19468
rect 6273 19459 6331 19465
rect 6362 19456 6368 19468
rect 6420 19496 6426 19508
rect 8662 19496 8668 19508
rect 6420 19468 8668 19496
rect 6420 19456 6426 19468
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 8846 19456 8852 19508
rect 8904 19496 8910 19508
rect 10134 19496 10140 19508
rect 8904 19468 10140 19496
rect 8904 19456 8910 19468
rect 10134 19456 10140 19468
rect 10192 19456 10198 19508
rect 13170 19496 13176 19508
rect 10520 19468 13176 19496
rect 2332 19428 2360 19456
rect 2332 19400 4476 19428
rect 2406 19320 2412 19372
rect 2464 19360 2470 19372
rect 3697 19363 3755 19369
rect 3697 19360 3709 19363
rect 2464 19332 3709 19360
rect 2464 19320 2470 19332
rect 3697 19329 3709 19332
rect 3743 19360 3755 19363
rect 4062 19360 4068 19372
rect 3743 19332 4068 19360
rect 3743 19329 3755 19332
rect 3697 19323 3755 19329
rect 4062 19320 4068 19332
rect 4120 19320 4126 19372
rect 4448 19360 4476 19400
rect 5828 19400 7696 19428
rect 4982 19369 4988 19372
rect 4939 19363 4988 19369
rect 4448 19332 4844 19360
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19292 1455 19295
rect 1486 19292 1492 19304
rect 1443 19264 1492 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1486 19252 1492 19264
rect 1544 19252 1550 19304
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3513 19295 3571 19301
rect 3513 19292 3525 19295
rect 3108 19264 3525 19292
rect 3108 19252 3114 19264
rect 3513 19261 3525 19264
rect 3559 19261 3571 19295
rect 3513 19255 3571 19261
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4522 19292 4528 19304
rect 4479 19264 4528 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4522 19252 4528 19264
rect 4580 19252 4586 19304
rect 4816 19292 4844 19332
rect 4939 19329 4951 19363
rect 4985 19329 4988 19363
rect 4939 19323 4988 19329
rect 4982 19320 4988 19323
rect 5040 19320 5046 19372
rect 5828 19360 5856 19400
rect 5092 19332 5856 19360
rect 5092 19292 5120 19332
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6914 19360 6920 19372
rect 6144 19332 6920 19360
rect 6144 19320 6150 19332
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7558 19360 7564 19372
rect 7515 19332 7564 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 7668 19360 7696 19400
rect 8570 19360 8576 19372
rect 7668 19332 8576 19360
rect 8570 19320 8576 19332
rect 8628 19320 8634 19372
rect 8711 19363 8769 19369
rect 8711 19329 8723 19363
rect 8757 19360 8769 19363
rect 10520 19360 10548 19468
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 15657 19499 15715 19505
rect 15657 19496 15669 19499
rect 13372 19468 15669 19496
rect 12069 19431 12127 19437
rect 12069 19397 12081 19431
rect 12115 19397 12127 19431
rect 12069 19391 12127 19397
rect 8757 19332 10548 19360
rect 12084 19360 12112 19391
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 13262 19428 13268 19440
rect 12400 19400 13268 19428
rect 12400 19388 12406 19400
rect 13262 19388 13268 19400
rect 13320 19388 13326 19440
rect 12802 19360 12808 19372
rect 12084 19332 12808 19360
rect 8757 19329 8769 19332
rect 8711 19323 8769 19329
rect 12802 19320 12808 19332
rect 12860 19320 12866 19372
rect 13078 19360 13084 19372
rect 13039 19332 13084 19360
rect 13078 19320 13084 19332
rect 13136 19320 13142 19372
rect 4816 19264 5120 19292
rect 5169 19295 5227 19301
rect 5169 19261 5181 19295
rect 5215 19292 5227 19295
rect 5258 19292 5264 19304
rect 5215 19264 5264 19292
rect 5215 19261 5227 19264
rect 5169 19255 5227 19261
rect 5258 19252 5264 19264
rect 5316 19252 5322 19304
rect 6822 19292 6828 19304
rect 5828 19264 6828 19292
rect 1664 19227 1722 19233
rect 1664 19193 1676 19227
rect 1710 19224 1722 19227
rect 3234 19224 3240 19236
rect 1710 19196 3240 19224
rect 1710 19193 1722 19196
rect 1664 19187 1722 19193
rect 3234 19184 3240 19196
rect 3292 19184 3298 19236
rect 2958 19116 2964 19168
rect 3016 19156 3022 19168
rect 3053 19159 3111 19165
rect 3053 19156 3065 19159
rect 3016 19128 3065 19156
rect 3016 19116 3022 19128
rect 3053 19125 3065 19128
rect 3099 19125 3111 19159
rect 3053 19119 3111 19125
rect 3142 19116 3148 19168
rect 3200 19156 3206 19168
rect 3421 19159 3479 19165
rect 3421 19156 3433 19159
rect 3200 19128 3433 19156
rect 3200 19116 3206 19128
rect 3421 19125 3433 19128
rect 3467 19125 3479 19159
rect 3421 19119 3479 19125
rect 4899 19159 4957 19165
rect 4899 19125 4911 19159
rect 4945 19156 4957 19159
rect 5828 19156 5856 19264
rect 6822 19252 6828 19264
rect 6880 19292 6886 19304
rect 8202 19292 8208 19304
rect 6880 19264 7972 19292
rect 8163 19264 8208 19292
rect 6880 19252 6886 19264
rect 7193 19227 7251 19233
rect 7193 19193 7205 19227
rect 7239 19224 7251 19227
rect 7374 19224 7380 19236
rect 7239 19196 7380 19224
rect 7239 19193 7251 19196
rect 7193 19187 7251 19193
rect 7374 19184 7380 19196
rect 7432 19184 7438 19236
rect 4945 19128 5856 19156
rect 4945 19125 4957 19128
rect 4899 19119 4957 19125
rect 6638 19116 6644 19168
rect 6696 19156 6702 19168
rect 6825 19159 6883 19165
rect 6825 19156 6837 19159
rect 6696 19128 6837 19156
rect 6696 19116 6702 19128
rect 6825 19125 6837 19128
rect 6871 19125 6883 19159
rect 6825 19119 6883 19125
rect 7285 19159 7343 19165
rect 7285 19125 7297 19159
rect 7331 19156 7343 19159
rect 7834 19156 7840 19168
rect 7331 19128 7840 19156
rect 7331 19125 7343 19128
rect 7285 19119 7343 19125
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 7944 19156 7972 19264
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8941 19295 8999 19301
rect 8941 19292 8953 19295
rect 8312 19264 8953 19292
rect 8110 19184 8116 19236
rect 8168 19224 8174 19236
rect 8312 19224 8340 19264
rect 8941 19261 8953 19264
rect 8987 19292 8999 19295
rect 8987 19264 9628 19292
rect 8987 19261 8999 19264
rect 8941 19255 8999 19261
rect 8168 19196 8340 19224
rect 9600 19224 9628 19264
rect 9674 19252 9680 19304
rect 9732 19292 9738 19304
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 9732 19264 10517 19292
rect 9732 19252 9738 19264
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10594 19252 10600 19304
rect 10652 19292 10658 19304
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 10652 19264 10701 19292
rect 10652 19252 10658 19264
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 10689 19255 10747 19261
rect 10956 19295 11014 19301
rect 10956 19261 10968 19295
rect 11002 19292 11014 19295
rect 12434 19292 12440 19304
rect 11002 19264 12440 19292
rect 11002 19261 11014 19264
rect 10956 19255 11014 19261
rect 12434 19252 12440 19264
rect 12492 19292 12498 19304
rect 13372 19292 13400 19468
rect 15657 19465 15669 19468
rect 15703 19465 15715 19499
rect 20806 19496 20812 19508
rect 15657 19459 15715 19465
rect 16480 19468 20392 19496
rect 20719 19468 20812 19496
rect 13538 19388 13544 19440
rect 13596 19428 13602 19440
rect 13596 19400 14228 19428
rect 13596 19388 13602 19400
rect 13630 19320 13636 19372
rect 13688 19320 13694 19372
rect 12492 19264 13400 19292
rect 13449 19295 13507 19301
rect 12492 19252 12498 19264
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 13648 19292 13676 19320
rect 14200 19304 14228 19400
rect 15194 19388 15200 19440
rect 15252 19428 15258 19440
rect 16480 19428 16508 19468
rect 17862 19428 17868 19440
rect 15252 19400 16508 19428
rect 17236 19400 17868 19428
rect 15252 19388 15258 19400
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 16393 19363 16451 19369
rect 16393 19360 16405 19363
rect 15703 19332 16405 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 16393 19329 16405 19332
rect 16439 19329 16451 19363
rect 16393 19323 16451 19329
rect 14182 19292 14188 19304
rect 13495 19264 13676 19292
rect 14143 19264 14188 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 14182 19252 14188 19264
rect 14240 19252 14246 19304
rect 16209 19295 16267 19301
rect 16209 19292 16221 19295
rect 14292 19264 16221 19292
rect 12250 19224 12256 19236
rect 9600 19196 12256 19224
rect 8168 19184 8174 19196
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 12526 19184 12532 19236
rect 12584 19224 12590 19236
rect 13630 19224 13636 19236
rect 12584 19196 13124 19224
rect 13591 19196 13636 19224
rect 12584 19184 12590 19196
rect 8671 19159 8729 19165
rect 8671 19156 8683 19159
rect 7944 19128 8683 19156
rect 8671 19125 8683 19128
rect 8717 19156 8729 19159
rect 9582 19156 9588 19168
rect 8717 19128 9588 19156
rect 8717 19125 8729 19128
rect 8671 19119 8729 19125
rect 9582 19116 9588 19128
rect 9640 19116 9646 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10318 19156 10324 19168
rect 10279 19128 10324 19156
rect 10318 19116 10324 19128
rect 10376 19116 10382 19168
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10962 19156 10968 19168
rect 10468 19128 10968 19156
rect 10468 19116 10474 19128
rect 10962 19116 10968 19128
rect 11020 19156 11026 19168
rect 12437 19159 12495 19165
rect 12437 19156 12449 19159
rect 11020 19128 12449 19156
rect 11020 19116 11026 19128
rect 12437 19125 12449 19128
rect 12483 19125 12495 19159
rect 12802 19156 12808 19168
rect 12763 19128 12808 19156
rect 12437 19119 12495 19125
rect 12802 19116 12808 19128
rect 12860 19116 12866 19168
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 13096 19156 13124 19196
rect 13630 19184 13636 19196
rect 13688 19184 13694 19236
rect 14292 19224 14320 19264
rect 16209 19261 16221 19264
rect 16255 19261 16267 19295
rect 16209 19255 16267 19261
rect 13740 19196 14320 19224
rect 14452 19227 14510 19233
rect 13740 19156 13768 19196
rect 14452 19193 14464 19227
rect 14498 19224 14510 19227
rect 14642 19224 14648 19236
rect 14498 19196 14648 19224
rect 14498 19193 14510 19196
rect 14452 19187 14510 19193
rect 14642 19184 14648 19196
rect 14700 19184 14706 19236
rect 17236 19224 17264 19400
rect 17862 19388 17868 19400
rect 17920 19388 17926 19440
rect 18046 19428 18052 19440
rect 18007 19400 18052 19428
rect 18046 19388 18052 19400
rect 18104 19388 18110 19440
rect 20364 19428 20392 19468
rect 20806 19456 20812 19468
rect 20864 19496 20870 19508
rect 21634 19496 21640 19508
rect 20864 19468 21640 19496
rect 20864 19456 20870 19468
rect 21634 19456 21640 19468
rect 21692 19456 21698 19508
rect 21174 19428 21180 19440
rect 18248 19400 18644 19428
rect 20364 19400 21180 19428
rect 17494 19320 17500 19372
rect 17552 19360 17558 19372
rect 17586 19360 17592 19372
rect 17552 19332 17592 19360
rect 17552 19320 17558 19332
rect 17586 19320 17592 19332
rect 17644 19360 17650 19372
rect 18248 19360 18276 19400
rect 17644 19332 18276 19360
rect 17644 19320 17650 19332
rect 18322 19320 18328 19372
rect 18380 19360 18386 19372
rect 18616 19369 18644 19400
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 18509 19363 18567 19369
rect 18509 19360 18521 19363
rect 18380 19332 18521 19360
rect 18380 19320 18386 19332
rect 18509 19329 18521 19332
rect 18555 19329 18567 19363
rect 18509 19323 18567 19329
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19329 18659 19363
rect 21450 19360 21456 19372
rect 21411 19332 21456 19360
rect 18601 19323 18659 19329
rect 21450 19320 21456 19332
rect 21508 19320 21514 19372
rect 17313 19295 17371 19301
rect 17313 19261 17325 19295
rect 17359 19292 17371 19295
rect 18230 19292 18236 19304
rect 17359 19264 18236 19292
rect 17359 19261 17371 19264
rect 17313 19255 17371 19261
rect 18230 19252 18236 19264
rect 18288 19252 18294 19304
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19429 19295 19487 19301
rect 19429 19292 19441 19295
rect 19392 19264 19441 19292
rect 19392 19252 19398 19264
rect 19429 19261 19441 19264
rect 19475 19261 19487 19295
rect 21358 19292 21364 19304
rect 19429 19255 19487 19261
rect 19536 19264 21364 19292
rect 15856 19196 17264 19224
rect 17405 19227 17463 19233
rect 12952 19128 12997 19156
rect 13096 19128 13768 19156
rect 13817 19159 13875 19165
rect 12952 19116 12958 19128
rect 13817 19125 13829 19159
rect 13863 19156 13875 19159
rect 14274 19156 14280 19168
rect 13863 19128 14280 19156
rect 13863 19125 13875 19128
rect 13817 19119 13875 19125
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 15378 19116 15384 19168
rect 15436 19156 15442 19168
rect 15856 19165 15884 19196
rect 17405 19193 17417 19227
rect 17451 19224 17463 19227
rect 18874 19224 18880 19236
rect 17451 19196 18880 19224
rect 17451 19193 17463 19196
rect 17405 19187 17463 19193
rect 18874 19184 18880 19196
rect 18932 19184 18938 19236
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15436 19128 15577 19156
rect 15436 19116 15442 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15565 19119 15623 19125
rect 15841 19159 15899 19165
rect 15841 19125 15853 19159
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16301 19159 16359 19165
rect 16301 19156 16313 19159
rect 16172 19128 16313 19156
rect 16172 19116 16178 19128
rect 16301 19125 16313 19128
rect 16347 19125 16359 19159
rect 16301 19119 16359 19125
rect 16945 19159 17003 19165
rect 16945 19125 16957 19159
rect 16991 19156 17003 19159
rect 19536 19156 19564 19264
rect 21358 19252 21364 19264
rect 21416 19252 21422 19304
rect 19696 19227 19754 19233
rect 19696 19193 19708 19227
rect 19742 19224 19754 19227
rect 20530 19224 20536 19236
rect 19742 19196 20536 19224
rect 19742 19193 19754 19196
rect 19696 19187 19754 19193
rect 20530 19184 20536 19196
rect 20588 19224 20594 19236
rect 21269 19227 21327 19233
rect 21269 19224 21281 19227
rect 20588 19196 21281 19224
rect 20588 19184 20594 19196
rect 21269 19193 21281 19196
rect 21315 19193 21327 19227
rect 21269 19187 21327 19193
rect 16991 19128 19564 19156
rect 16991 19125 17003 19128
rect 16945 19119 17003 19125
rect 20898 19116 20904 19168
rect 20956 19156 20962 19168
rect 21358 19156 21364 19168
rect 20956 19128 21001 19156
rect 21319 19128 21364 19156
rect 20956 19116 20962 19128
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 21910 19156 21916 19168
rect 21871 19128 21916 19156
rect 21910 19116 21916 19128
rect 21968 19156 21974 19168
rect 22097 19159 22155 19165
rect 22097 19156 22109 19159
rect 21968 19128 22109 19156
rect 21968 19116 21974 19128
rect 22097 19125 22109 19128
rect 22143 19125 22155 19159
rect 22097 19119 22155 19125
rect 1104 19066 22816 19088
rect 1104 19014 8246 19066
rect 8298 19014 8310 19066
rect 8362 19014 8374 19066
rect 8426 19014 8438 19066
rect 8490 19014 15510 19066
rect 15562 19014 15574 19066
rect 15626 19014 15638 19066
rect 15690 19014 15702 19066
rect 15754 19014 22816 19066
rect 1104 18992 22816 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 2866 18952 2872 18964
rect 1627 18924 2872 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 2866 18912 2872 18924
rect 2924 18912 2930 18964
rect 3234 18912 3240 18964
rect 3292 18952 3298 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 3292 18924 3341 18952
rect 3292 18912 3298 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 4246 18952 4252 18964
rect 4207 18924 4252 18952
rect 3329 18915 3387 18921
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 5905 18955 5963 18961
rect 5905 18952 5917 18955
rect 5224 18924 5917 18952
rect 5224 18912 5230 18924
rect 5905 18921 5917 18924
rect 5951 18921 5963 18955
rect 6546 18952 6552 18964
rect 5905 18915 5963 18921
rect 6196 18924 6552 18952
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 2222 18893 2228 18896
rect 2194 18887 2228 18893
rect 2194 18884 2206 18887
rect 1820 18856 2206 18884
rect 1820 18844 1826 18856
rect 2194 18853 2206 18856
rect 2280 18884 2286 18896
rect 5261 18887 5319 18893
rect 2280 18856 2342 18884
rect 2194 18847 2228 18853
rect 2222 18844 2228 18847
rect 2280 18844 2286 18856
rect 5261 18853 5273 18887
rect 5307 18884 5319 18887
rect 5442 18884 5448 18896
rect 5307 18856 5448 18884
rect 5307 18853 5319 18856
rect 5261 18847 5319 18853
rect 5442 18844 5448 18856
rect 5500 18844 5506 18896
rect 5920 18884 5948 18915
rect 6196 18884 6224 18924
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7834 18952 7840 18964
rect 7795 18924 7840 18952
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8110 18912 8116 18964
rect 8168 18952 8174 18964
rect 8297 18955 8355 18961
rect 8297 18952 8309 18955
rect 8168 18924 8309 18952
rect 8168 18912 8174 18924
rect 8297 18921 8309 18924
rect 8343 18952 8355 18955
rect 8343 18924 8524 18952
rect 8343 18921 8355 18924
rect 8297 18915 8355 18921
rect 6454 18893 6460 18896
rect 6448 18884 6460 18893
rect 5920 18856 6224 18884
rect 6367 18856 6460 18884
rect 1394 18816 1400 18828
rect 1355 18788 1400 18816
rect 1394 18776 1400 18788
rect 1452 18776 1458 18828
rect 2498 18776 2504 18828
rect 2556 18816 2562 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 2556 18788 4077 18816
rect 2556 18776 2562 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 6086 18816 6092 18828
rect 6047 18788 6092 18816
rect 4065 18779 4123 18785
rect 6086 18776 6092 18788
rect 6144 18776 6150 18828
rect 6196 18825 6224 18856
rect 6448 18847 6460 18856
rect 6512 18884 6518 18896
rect 6512 18856 8432 18884
rect 6454 18844 6460 18847
rect 6512 18844 6518 18856
rect 6181 18819 6239 18825
rect 6181 18785 6193 18819
rect 6227 18785 6239 18819
rect 6181 18779 6239 18785
rect 6730 18776 6736 18828
rect 6788 18816 6794 18828
rect 7006 18816 7012 18828
rect 6788 18788 7012 18816
rect 6788 18776 6794 18788
rect 7006 18776 7012 18788
rect 7064 18776 7070 18828
rect 7190 18776 7196 18828
rect 7248 18816 7254 18828
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 7248 18788 8217 18816
rect 7248 18776 7254 18788
rect 8205 18785 8217 18788
rect 8251 18785 8263 18819
rect 8205 18779 8263 18785
rect 1486 18708 1492 18760
rect 1544 18748 1550 18760
rect 1949 18751 2007 18757
rect 1949 18748 1961 18751
rect 1544 18720 1961 18748
rect 1544 18708 1550 18720
rect 1949 18717 1961 18720
rect 1995 18717 2007 18751
rect 1949 18711 2007 18717
rect 4982 18708 4988 18760
rect 5040 18748 5046 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5040 18720 5365 18748
rect 5040 18708 5046 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5445 18751 5503 18757
rect 5445 18717 5457 18751
rect 5491 18748 5503 18751
rect 5718 18748 5724 18760
rect 5491 18720 5724 18748
rect 5491 18717 5503 18720
rect 5445 18711 5503 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 8404 18757 8432 18856
rect 8496 18816 8524 18924
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 9033 18955 9091 18961
rect 9033 18952 9045 18955
rect 8628 18924 9045 18952
rect 8628 18912 8634 18924
rect 9033 18921 9045 18924
rect 9079 18921 9091 18955
rect 9033 18915 9091 18921
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10091 18924 12756 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 12158 18884 12164 18896
rect 8864 18856 12164 18884
rect 8570 18816 8576 18828
rect 8496 18788 8576 18816
rect 8570 18776 8576 18788
rect 8628 18776 8634 18828
rect 8864 18825 8892 18856
rect 12158 18844 12164 18856
rect 12216 18844 12222 18896
rect 12728 18884 12756 18924
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 16482 18952 16488 18964
rect 12860 18924 16488 18952
rect 12860 18912 12866 18924
rect 16482 18912 16488 18924
rect 16540 18912 16546 18964
rect 17129 18955 17187 18961
rect 17129 18921 17141 18955
rect 17175 18921 17187 18955
rect 18874 18952 18880 18964
rect 18835 18924 18880 18952
rect 17129 18915 17187 18921
rect 15556 18887 15614 18893
rect 12728 18856 14136 18884
rect 8849 18819 8907 18825
rect 8849 18785 8861 18819
rect 8895 18785 8907 18819
rect 10410 18816 10416 18828
rect 10371 18788 10416 18816
rect 8849 18779 8907 18785
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18717 8447 18751
rect 8389 18711 8447 18717
rect 4893 18683 4951 18689
rect 4893 18649 4905 18683
rect 4939 18680 4951 18683
rect 8864 18680 8892 18779
rect 10410 18776 10416 18788
rect 10468 18776 10474 18828
rect 11054 18816 11060 18828
rect 11015 18788 11060 18816
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11572 18788 11989 18816
rect 11572 18776 11578 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12069 18819 12127 18825
rect 12069 18785 12081 18819
rect 12115 18816 12127 18819
rect 12434 18816 12440 18828
rect 12115 18788 12440 18816
rect 12115 18785 12127 18788
rect 12069 18779 12127 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 12621 18819 12679 18825
rect 12621 18785 12633 18819
rect 12667 18816 12679 18819
rect 12710 18816 12716 18828
rect 12667 18788 12716 18816
rect 12667 18785 12679 18788
rect 12621 18779 12679 18785
rect 12710 18776 12716 18788
rect 12768 18776 12774 18828
rect 12888 18819 12946 18825
rect 12888 18785 12900 18819
rect 12934 18816 12946 18819
rect 13630 18816 13636 18828
rect 12934 18788 13636 18816
rect 12934 18785 12946 18788
rect 12888 18779 12946 18785
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 10505 18751 10563 18757
rect 10505 18717 10517 18751
rect 10551 18717 10563 18751
rect 10505 18711 10563 18717
rect 4939 18652 6224 18680
rect 4939 18649 4951 18652
rect 4893 18643 4951 18649
rect 4338 18572 4344 18624
rect 4396 18612 4402 18624
rect 5350 18612 5356 18624
rect 4396 18584 5356 18612
rect 4396 18572 4402 18584
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 6196 18612 6224 18652
rect 7392 18652 8892 18680
rect 10520 18680 10548 18711
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 12158 18748 12164 18760
rect 10652 18720 10697 18748
rect 12119 18720 12164 18748
rect 10652 18708 10658 18720
rect 12158 18708 12164 18720
rect 12216 18708 12222 18760
rect 11054 18680 11060 18692
rect 10520 18652 11060 18680
rect 7392 18612 7420 18652
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 11609 18683 11667 18689
rect 11164 18652 11560 18680
rect 7558 18612 7564 18624
rect 6196 18584 7420 18612
rect 7519 18584 7564 18612
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 8938 18572 8944 18624
rect 8996 18612 9002 18624
rect 11164 18612 11192 18652
rect 8996 18584 11192 18612
rect 8996 18572 9002 18584
rect 11238 18572 11244 18624
rect 11296 18612 11302 18624
rect 11532 18612 11560 18652
rect 11609 18649 11621 18683
rect 11655 18680 11667 18683
rect 12618 18680 12624 18692
rect 11655 18652 12624 18680
rect 11655 18649 11667 18652
rect 11609 18643 11667 18649
rect 12618 18640 12624 18652
rect 12676 18640 12682 18692
rect 12342 18612 12348 18624
rect 11296 18584 11341 18612
rect 11532 18584 12348 18612
rect 11296 18572 11302 18584
rect 12342 18572 12348 18584
rect 12400 18572 12406 18624
rect 12526 18572 12532 18624
rect 12584 18612 12590 18624
rect 14001 18615 14059 18621
rect 14001 18612 14013 18615
rect 12584 18584 14013 18612
rect 12584 18572 12590 18584
rect 14001 18581 14013 18584
rect 14047 18581 14059 18615
rect 14108 18612 14136 18856
rect 15556 18853 15568 18887
rect 15602 18884 15614 18887
rect 15930 18884 15936 18896
rect 15602 18856 15936 18884
rect 15602 18853 15614 18856
rect 15556 18847 15614 18853
rect 15930 18844 15936 18856
rect 15988 18844 15994 18896
rect 17144 18884 17172 18915
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 19150 18912 19156 18964
rect 19208 18952 19214 18964
rect 19334 18952 19340 18964
rect 19208 18924 19340 18952
rect 19208 18912 19214 18924
rect 19334 18912 19340 18924
rect 19392 18952 19398 18964
rect 20346 18952 20352 18964
rect 19392 18924 20352 18952
rect 19392 18912 19398 18924
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 20530 18952 20536 18964
rect 20491 18924 20536 18952
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 16040 18856 17172 18884
rect 17764 18887 17822 18893
rect 14274 18816 14280 18828
rect 14235 18788 14280 18816
rect 14274 18776 14280 18788
rect 14332 18776 14338 18828
rect 14734 18776 14740 18828
rect 14792 18816 14798 18828
rect 16040 18816 16068 18856
rect 17764 18853 17776 18887
rect 17810 18884 17822 18887
rect 18414 18884 18420 18896
rect 17810 18856 18420 18884
rect 17810 18853 17822 18856
rect 17764 18847 17822 18853
rect 18414 18844 18420 18856
rect 18472 18844 18478 18896
rect 19420 18887 19478 18893
rect 19420 18853 19432 18887
rect 19466 18884 19478 18887
rect 21358 18884 21364 18896
rect 19466 18856 21364 18884
rect 19466 18853 19478 18856
rect 19420 18847 19478 18853
rect 21358 18844 21364 18856
rect 21416 18844 21422 18896
rect 14792 18788 16068 18816
rect 14792 18776 14798 18788
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16632 18788 16957 18816
rect 16632 18776 16638 18788
rect 16945 18785 16957 18788
rect 16991 18785 17003 18819
rect 16945 18779 17003 18785
rect 21082 18776 21088 18828
rect 21140 18816 21146 18828
rect 21269 18819 21327 18825
rect 21269 18816 21281 18819
rect 21140 18788 21281 18816
rect 21140 18776 21146 18788
rect 21269 18785 21281 18788
rect 21315 18785 21327 18819
rect 21269 18779 21327 18785
rect 14182 18708 14188 18760
rect 14240 18748 14246 18760
rect 14918 18748 14924 18760
rect 14240 18720 14924 18748
rect 14240 18708 14246 18720
rect 14918 18708 14924 18720
rect 14976 18748 14982 18760
rect 15289 18751 15347 18757
rect 15289 18748 15301 18751
rect 14976 18720 15301 18748
rect 14976 18708 14982 18720
rect 15289 18717 15301 18720
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 17497 18751 17555 18757
rect 17497 18717 17509 18751
rect 17543 18717 17555 18751
rect 19150 18748 19156 18760
rect 19111 18720 19156 18748
rect 17497 18711 17555 18717
rect 14458 18680 14464 18692
rect 14419 18652 14464 18680
rect 14458 18640 14464 18652
rect 14516 18640 14522 18692
rect 16942 18640 16948 18692
rect 17000 18680 17006 18692
rect 17512 18680 17540 18711
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 21361 18751 21419 18757
rect 21361 18717 21373 18751
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 21453 18751 21511 18757
rect 21453 18717 21465 18751
rect 21499 18748 21511 18751
rect 21818 18748 21824 18760
rect 21499 18720 21824 18748
rect 21499 18717 21511 18720
rect 21453 18711 21511 18717
rect 17000 18652 17540 18680
rect 21376 18680 21404 18711
rect 21818 18708 21824 18720
rect 21876 18708 21882 18760
rect 22097 18751 22155 18757
rect 22097 18717 22109 18751
rect 22143 18717 22155 18751
rect 22097 18711 22155 18717
rect 21542 18680 21548 18692
rect 21376 18652 21548 18680
rect 17000 18640 17006 18652
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 15930 18612 15936 18624
rect 14108 18584 15936 18612
rect 14001 18575 14059 18581
rect 15930 18572 15936 18584
rect 15988 18572 15994 18624
rect 16666 18612 16672 18624
rect 16627 18584 16672 18612
rect 16666 18572 16672 18584
rect 16724 18572 16730 18624
rect 16850 18572 16856 18624
rect 16908 18612 16914 18624
rect 20622 18612 20628 18624
rect 16908 18584 20628 18612
rect 16908 18572 16914 18584
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 20898 18612 20904 18624
rect 20859 18584 20904 18612
rect 20898 18572 20904 18584
rect 20956 18572 20962 18624
rect 20990 18572 20996 18624
rect 21048 18612 21054 18624
rect 21913 18615 21971 18621
rect 21913 18612 21925 18615
rect 21048 18584 21925 18612
rect 21048 18572 21054 18584
rect 21913 18581 21925 18584
rect 21959 18612 21971 18615
rect 22112 18612 22140 18711
rect 21959 18584 22140 18612
rect 21959 18581 21971 18584
rect 21913 18575 21971 18581
rect 1104 18522 22816 18544
rect 1104 18470 4614 18522
rect 4666 18470 4678 18522
rect 4730 18470 4742 18522
rect 4794 18470 4806 18522
rect 4858 18470 11878 18522
rect 11930 18470 11942 18522
rect 11994 18470 12006 18522
rect 12058 18470 12070 18522
rect 12122 18470 19142 18522
rect 19194 18470 19206 18522
rect 19258 18470 19270 18522
rect 19322 18470 19334 18522
rect 19386 18470 22816 18522
rect 1104 18448 22816 18470
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 2961 18411 3019 18417
rect 2961 18408 2973 18411
rect 2280 18380 2973 18408
rect 2280 18368 2286 18380
rect 2961 18377 2973 18380
rect 3007 18377 3019 18411
rect 2961 18371 3019 18377
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3476 18380 3617 18408
rect 3476 18368 3482 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 6454 18408 6460 18420
rect 3605 18371 3663 18377
rect 4724 18380 6316 18408
rect 6415 18380 6460 18408
rect 3234 18232 3240 18284
rect 3292 18232 3298 18284
rect 4724 18281 4752 18380
rect 6288 18340 6316 18380
rect 6454 18368 6460 18380
rect 6512 18368 6518 18420
rect 6730 18368 6736 18420
rect 6788 18408 6794 18420
rect 9858 18408 9864 18420
rect 6788 18380 9864 18408
rect 6788 18368 6794 18380
rect 9858 18368 9864 18380
rect 9916 18368 9922 18420
rect 10137 18411 10195 18417
rect 10137 18377 10149 18411
rect 10183 18408 10195 18411
rect 11606 18408 11612 18420
rect 10183 18380 11612 18408
rect 10183 18377 10195 18380
rect 10137 18371 10195 18377
rect 11606 18368 11612 18380
rect 11664 18368 11670 18420
rect 12710 18408 12716 18420
rect 12452 18380 12716 18408
rect 6638 18340 6644 18352
rect 6288 18312 6644 18340
rect 6638 18300 6644 18312
rect 6696 18300 6702 18352
rect 10042 18300 10048 18352
rect 10100 18340 10106 18352
rect 11422 18340 11428 18352
rect 10100 18312 11428 18340
rect 10100 18300 10106 18312
rect 11422 18300 11428 18312
rect 11480 18300 11486 18352
rect 11514 18300 11520 18352
rect 11572 18340 11578 18352
rect 11790 18340 11796 18352
rect 11572 18312 11796 18340
rect 11572 18300 11578 18312
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 4709 18275 4767 18281
rect 4709 18241 4721 18275
rect 4755 18241 4767 18275
rect 4709 18235 4767 18241
rect 5000 18244 5212 18272
rect 1486 18164 1492 18216
rect 1544 18204 1550 18216
rect 1854 18213 1860 18216
rect 1581 18207 1639 18213
rect 1581 18204 1593 18207
rect 1544 18176 1593 18204
rect 1544 18164 1550 18176
rect 1581 18173 1593 18176
rect 1627 18173 1639 18207
rect 1848 18204 1860 18213
rect 1815 18176 1860 18204
rect 1581 18167 1639 18173
rect 1848 18167 1860 18176
rect 1854 18164 1860 18167
rect 1912 18164 1918 18216
rect 3252 18204 3280 18232
rect 3421 18207 3479 18213
rect 3421 18204 3433 18207
rect 3252 18176 3433 18204
rect 3421 18173 3433 18176
rect 3467 18173 3479 18207
rect 3421 18167 3479 18173
rect 4338 18164 4344 18216
rect 4396 18164 4402 18216
rect 4525 18207 4583 18213
rect 4525 18173 4537 18207
rect 4571 18204 4583 18207
rect 5000 18204 5028 18244
rect 4571 18176 5028 18204
rect 5077 18207 5135 18213
rect 4571 18173 4583 18176
rect 4525 18167 4583 18173
rect 5077 18173 5089 18207
rect 5123 18173 5135 18207
rect 5184 18204 5212 18244
rect 6546 18232 6552 18284
rect 6604 18272 6610 18284
rect 6825 18275 6883 18281
rect 6825 18272 6837 18275
rect 6604 18244 6837 18272
rect 6604 18232 6610 18244
rect 6825 18241 6837 18244
rect 6871 18241 6883 18275
rect 6825 18235 6883 18241
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10652 18244 10793 18272
rect 10652 18232 10658 18244
rect 10781 18241 10793 18244
rect 10827 18272 10839 18275
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 10827 18244 11989 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 11977 18241 11989 18244
rect 12023 18272 12035 18275
rect 12158 18272 12164 18284
rect 12023 18244 12164 18272
rect 12023 18241 12035 18244
rect 11977 18235 12035 18241
rect 12158 18232 12164 18244
rect 12216 18232 12222 18284
rect 12250 18232 12256 18284
rect 12308 18272 12314 18284
rect 12452 18281 12480 18380
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 13817 18411 13875 18417
rect 13817 18408 13829 18411
rect 13688 18380 13829 18408
rect 13688 18368 13694 18380
rect 13817 18377 13829 18380
rect 13863 18377 13875 18411
rect 14274 18408 14280 18420
rect 14235 18380 14280 18408
rect 13817 18371 13875 18377
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 14642 18408 14648 18420
rect 14516 18380 14648 18408
rect 14516 18368 14522 18380
rect 14642 18368 14648 18380
rect 14700 18408 14706 18420
rect 16666 18408 16672 18420
rect 14700 18380 16672 18408
rect 14700 18368 14706 18380
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 18325 18411 18383 18417
rect 18325 18377 18337 18411
rect 18371 18408 18383 18411
rect 19610 18408 19616 18420
rect 18371 18380 19616 18408
rect 18371 18377 18383 18380
rect 18325 18371 18383 18377
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 20073 18411 20131 18417
rect 20073 18377 20085 18411
rect 20119 18408 20131 18411
rect 21358 18408 21364 18420
rect 20119 18380 21364 18408
rect 20119 18377 20131 18380
rect 20073 18371 20131 18377
rect 21358 18368 21364 18380
rect 21416 18368 21422 18420
rect 18690 18340 18696 18352
rect 17236 18312 18696 18340
rect 17236 18284 17264 18312
rect 18690 18300 18696 18312
rect 18748 18300 18754 18352
rect 12437 18275 12495 18281
rect 12437 18272 12449 18275
rect 12308 18244 12449 18272
rect 12308 18232 12314 18244
rect 12437 18241 12449 18244
rect 12483 18241 12495 18275
rect 17126 18272 17132 18284
rect 17087 18244 17132 18272
rect 12437 18235 12495 18241
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17218 18232 17224 18284
rect 17276 18272 17282 18284
rect 20993 18275 21051 18281
rect 17276 18244 17321 18272
rect 18156 18244 18828 18272
rect 17276 18232 17282 18244
rect 6730 18204 6736 18216
rect 5184 18176 6736 18204
rect 5077 18167 5135 18173
rect 3237 18139 3295 18145
rect 3237 18105 3249 18139
rect 3283 18136 3295 18139
rect 4356 18136 4384 18164
rect 3283 18108 4384 18136
rect 5092 18136 5120 18167
rect 6730 18164 6736 18176
rect 6788 18164 6794 18216
rect 7092 18207 7150 18213
rect 7092 18173 7104 18207
rect 7138 18204 7150 18207
rect 7558 18204 7564 18216
rect 7138 18176 7564 18204
rect 7138 18173 7150 18176
rect 7092 18167 7150 18173
rect 7558 18164 7564 18176
rect 7616 18164 7622 18216
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 9122 18204 9128 18216
rect 8527 18176 9128 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 9122 18164 9128 18176
rect 9180 18204 9186 18216
rect 10318 18204 10324 18216
rect 9180 18176 10324 18204
rect 9180 18164 9186 18176
rect 10318 18164 10324 18176
rect 10376 18164 10382 18216
rect 11701 18207 11759 18213
rect 11701 18173 11713 18207
rect 11747 18204 11759 18207
rect 13170 18204 13176 18216
rect 11747 18176 13176 18204
rect 11747 18173 11759 18176
rect 11701 18167 11759 18173
rect 13170 18164 13176 18176
rect 13228 18164 13234 18216
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 13320 18176 14105 18204
rect 13320 18164 13326 18176
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14182 18164 14188 18216
rect 14240 18204 14246 18216
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 14240 18176 14841 18204
rect 14240 18164 14246 18176
rect 14829 18173 14841 18176
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 14921 18207 14979 18213
rect 14921 18173 14933 18207
rect 14967 18173 14979 18207
rect 14921 18167 14979 18173
rect 17037 18207 17095 18213
rect 17037 18173 17049 18207
rect 17083 18204 17095 18207
rect 18046 18204 18052 18216
rect 17083 18176 18052 18204
rect 17083 18173 17095 18176
rect 17037 18167 17095 18173
rect 5166 18136 5172 18148
rect 5092 18108 5172 18136
rect 3283 18105 3295 18108
rect 3237 18099 3295 18105
rect 5166 18096 5172 18108
rect 5224 18096 5230 18148
rect 5344 18139 5402 18145
rect 5344 18105 5356 18139
rect 5390 18136 5402 18139
rect 5718 18136 5724 18148
rect 5390 18108 5724 18136
rect 5390 18105 5402 18108
rect 5344 18099 5402 18105
rect 5718 18096 5724 18108
rect 5776 18096 5782 18148
rect 7742 18096 7748 18148
rect 7800 18136 7806 18148
rect 8748 18139 8806 18145
rect 7800 18108 8432 18136
rect 7800 18096 7806 18108
rect 4065 18071 4123 18077
rect 4065 18037 4077 18071
rect 4111 18068 4123 18071
rect 4338 18068 4344 18080
rect 4111 18040 4344 18068
rect 4111 18037 4123 18040
rect 4065 18031 4123 18037
rect 4338 18028 4344 18040
rect 4396 18028 4402 18080
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 5074 18068 5080 18080
rect 4479 18040 5080 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 8110 18028 8116 18080
rect 8168 18068 8174 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 8168 18040 8217 18068
rect 8168 18028 8174 18040
rect 8205 18037 8217 18040
rect 8251 18037 8263 18071
rect 8404 18068 8432 18108
rect 8748 18105 8760 18139
rect 8794 18136 8806 18139
rect 8938 18136 8944 18148
rect 8794 18108 8944 18136
rect 8794 18105 8806 18108
rect 8748 18099 8806 18105
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 10505 18139 10563 18145
rect 10505 18105 10517 18139
rect 10551 18136 10563 18139
rect 11146 18136 11152 18148
rect 10551 18108 11152 18136
rect 10551 18105 10563 18108
rect 10505 18099 10563 18105
rect 11146 18096 11152 18108
rect 11204 18096 11210 18148
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 12526 18136 12532 18148
rect 12400 18108 12532 18136
rect 12400 18096 12406 18108
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 12710 18145 12716 18148
rect 12704 18099 12716 18145
rect 12768 18136 12774 18148
rect 12768 18108 12804 18136
rect 12710 18096 12716 18099
rect 12768 18096 12774 18108
rect 14936 18080 14964 18167
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 18156 18213 18184 18244
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18173 18199 18207
rect 18141 18167 18199 18173
rect 18414 18164 18420 18216
rect 18472 18204 18478 18216
rect 18693 18207 18751 18213
rect 18693 18204 18705 18207
rect 18472 18176 18705 18204
rect 18472 18164 18478 18176
rect 18693 18173 18705 18176
rect 18739 18173 18751 18207
rect 18800 18204 18828 18244
rect 20993 18241 21005 18275
rect 21039 18272 21051 18275
rect 21174 18272 21180 18284
rect 21039 18244 21180 18272
rect 21039 18241 21051 18244
rect 20993 18235 21051 18241
rect 21174 18232 21180 18244
rect 21232 18232 21238 18284
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 21913 18275 21971 18281
rect 21913 18272 21925 18275
rect 21876 18244 21925 18272
rect 21876 18232 21882 18244
rect 21913 18241 21925 18244
rect 21959 18241 21971 18275
rect 21913 18235 21971 18241
rect 20622 18204 20628 18216
rect 18800 18176 20628 18204
rect 18693 18167 18751 18173
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 15194 18145 15200 18148
rect 15188 18136 15200 18145
rect 15155 18108 15200 18136
rect 15188 18099 15200 18108
rect 15194 18096 15200 18099
rect 15252 18096 15258 18148
rect 15304 18108 16804 18136
rect 9861 18071 9919 18077
rect 9861 18068 9873 18071
rect 8404 18040 9873 18068
rect 8205 18031 8263 18037
rect 9861 18037 9873 18040
rect 9907 18037 9919 18071
rect 9861 18031 9919 18037
rect 10594 18028 10600 18080
rect 10652 18068 10658 18080
rect 11330 18068 11336 18080
rect 10652 18040 10697 18068
rect 11291 18040 11336 18068
rect 10652 18028 10658 18040
rect 11330 18028 11336 18040
rect 11388 18028 11394 18080
rect 11422 18028 11428 18080
rect 11480 18068 11486 18080
rect 11793 18071 11851 18077
rect 11793 18068 11805 18071
rect 11480 18040 11805 18068
rect 11480 18028 11486 18040
rect 11793 18037 11805 18040
rect 11839 18037 11851 18071
rect 11793 18031 11851 18037
rect 13262 18028 13268 18080
rect 13320 18068 13326 18080
rect 13722 18068 13728 18080
rect 13320 18040 13728 18068
rect 13320 18028 13326 18040
rect 13722 18028 13728 18040
rect 13780 18028 13786 18080
rect 14645 18071 14703 18077
rect 14645 18037 14657 18071
rect 14691 18068 14703 18071
rect 14918 18068 14924 18080
rect 14691 18040 14924 18068
rect 14691 18037 14703 18040
rect 14645 18031 14703 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15010 18028 15016 18080
rect 15068 18068 15074 18080
rect 15304 18068 15332 18108
rect 15068 18040 15332 18068
rect 15068 18028 15074 18040
rect 16114 18028 16120 18080
rect 16172 18068 16178 18080
rect 16301 18071 16359 18077
rect 16301 18068 16313 18071
rect 16172 18040 16313 18068
rect 16172 18028 16178 18040
rect 16301 18037 16313 18040
rect 16347 18037 16359 18071
rect 16666 18068 16672 18080
rect 16627 18040 16672 18068
rect 16301 18031 16359 18037
rect 16666 18028 16672 18040
rect 16724 18028 16730 18080
rect 16776 18068 16804 18108
rect 18230 18096 18236 18148
rect 18288 18136 18294 18148
rect 18938 18139 18996 18145
rect 18938 18136 18950 18139
rect 18288 18108 18950 18136
rect 18288 18096 18294 18108
rect 18938 18105 18950 18108
rect 18984 18136 18996 18139
rect 19242 18136 19248 18148
rect 18984 18108 19248 18136
rect 18984 18105 18996 18108
rect 18938 18099 18996 18105
rect 19242 18096 19248 18108
rect 19300 18096 19306 18148
rect 21450 18096 21456 18148
rect 21508 18136 21514 18148
rect 21821 18139 21879 18145
rect 21821 18136 21833 18139
rect 21508 18108 21833 18136
rect 21508 18096 21514 18108
rect 21821 18105 21833 18108
rect 21867 18105 21879 18139
rect 21821 18099 21879 18105
rect 19886 18068 19892 18080
rect 16776 18040 19892 18068
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 20162 18028 20168 18080
rect 20220 18068 20226 18080
rect 20349 18071 20407 18077
rect 20349 18068 20361 18071
rect 20220 18040 20361 18068
rect 20220 18028 20226 18040
rect 20349 18037 20361 18040
rect 20395 18037 20407 18071
rect 20714 18068 20720 18080
rect 20675 18040 20720 18068
rect 20349 18031 20407 18037
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 20806 18028 20812 18080
rect 20864 18068 20870 18080
rect 21358 18068 21364 18080
rect 20864 18040 20909 18068
rect 21319 18040 21364 18068
rect 20864 18028 20870 18040
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 21726 18068 21732 18080
rect 21687 18040 21732 18068
rect 21726 18028 21732 18040
rect 21784 18028 21790 18080
rect 1104 17978 22816 18000
rect 1104 17926 8246 17978
rect 8298 17926 8310 17978
rect 8362 17926 8374 17978
rect 8426 17926 8438 17978
rect 8490 17926 15510 17978
rect 15562 17926 15574 17978
rect 15626 17926 15638 17978
rect 15690 17926 15702 17978
rect 15754 17926 22816 17978
rect 1104 17904 22816 17926
rect 1854 17824 1860 17876
rect 1912 17864 1918 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 1912 17836 2973 17864
rect 1912 17824 1918 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 2961 17827 3019 17833
rect 3326 17824 3332 17876
rect 3384 17864 3390 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3384 17836 3433 17864
rect 3384 17824 3390 17836
rect 3421 17833 3433 17836
rect 3467 17833 3479 17867
rect 3421 17827 3479 17833
rect 5166 17824 5172 17876
rect 5224 17824 5230 17876
rect 5718 17864 5724 17876
rect 5679 17836 5724 17864
rect 5718 17824 5724 17836
rect 5776 17824 5782 17876
rect 6178 17864 6184 17876
rect 6139 17836 6184 17864
rect 6178 17824 6184 17836
rect 6236 17824 6242 17876
rect 7006 17864 7012 17876
rect 6748 17836 7012 17864
rect 2130 17756 2136 17808
rect 2188 17796 2194 17808
rect 3970 17796 3976 17808
rect 2188 17768 3976 17796
rect 2188 17756 2194 17768
rect 3970 17756 3976 17768
rect 4028 17756 4034 17808
rect 5184 17796 5212 17824
rect 5350 17796 5356 17808
rect 4356 17768 5356 17796
rect 1848 17731 1906 17737
rect 1848 17697 1860 17731
rect 1894 17728 1906 17731
rect 2222 17728 2228 17740
rect 1894 17700 2228 17728
rect 1894 17697 1906 17700
rect 1848 17691 1906 17697
rect 2222 17688 2228 17700
rect 2280 17688 2286 17740
rect 3237 17731 3295 17737
rect 3237 17697 3249 17731
rect 3283 17728 3295 17731
rect 3510 17728 3516 17740
rect 3283 17700 3516 17728
rect 3283 17697 3295 17700
rect 3237 17691 3295 17697
rect 3510 17688 3516 17700
rect 3568 17688 3574 17740
rect 4356 17737 4384 17768
rect 5350 17756 5356 17768
rect 5408 17756 5414 17808
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17697 4399 17731
rect 4341 17691 4399 17697
rect 4608 17731 4666 17737
rect 4608 17697 4620 17731
rect 4654 17728 4666 17731
rect 5166 17728 5172 17740
rect 4654 17700 5172 17728
rect 4654 17697 4666 17700
rect 4608 17691 4666 17697
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5902 17688 5908 17740
rect 5960 17728 5966 17740
rect 5997 17731 6055 17737
rect 5997 17728 6009 17731
rect 5960 17700 6009 17728
rect 5960 17688 5966 17700
rect 5997 17697 6009 17700
rect 6043 17728 6055 17731
rect 6454 17728 6460 17740
rect 6043 17700 6460 17728
rect 6043 17697 6055 17700
rect 5997 17691 6055 17697
rect 6454 17688 6460 17700
rect 6512 17688 6518 17740
rect 6546 17688 6552 17740
rect 6604 17728 6610 17740
rect 6748 17737 6776 17836
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 7282 17824 7288 17876
rect 7340 17864 7346 17876
rect 9033 17867 9091 17873
rect 9033 17864 9045 17867
rect 7340 17836 9045 17864
rect 7340 17824 7346 17836
rect 9033 17833 9045 17836
rect 9079 17833 9091 17867
rect 9033 17827 9091 17833
rect 9677 17867 9735 17873
rect 9677 17833 9689 17867
rect 9723 17864 9735 17867
rect 10594 17864 10600 17876
rect 9723 17836 10600 17864
rect 9723 17833 9735 17836
rect 9677 17827 9735 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11793 17867 11851 17873
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 12710 17864 12716 17876
rect 11839 17836 12716 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 12710 17824 12716 17836
rect 12768 17864 12774 17876
rect 13817 17867 13875 17873
rect 13817 17864 13829 17867
rect 12768 17836 13829 17864
rect 12768 17824 12774 17836
rect 13817 17833 13829 17836
rect 13863 17833 13875 17867
rect 13817 17827 13875 17833
rect 14093 17867 14151 17873
rect 14093 17833 14105 17867
rect 14139 17833 14151 17867
rect 14093 17827 14151 17833
rect 15749 17867 15807 17873
rect 15749 17833 15761 17867
rect 15795 17864 15807 17867
rect 16390 17864 16396 17876
rect 15795 17836 16396 17864
rect 15795 17833 15807 17836
rect 15749 17827 15807 17833
rect 9766 17756 9772 17808
rect 9824 17796 9830 17808
rect 9824 17768 10732 17796
rect 9824 17756 9830 17768
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 6604 17700 6745 17728
rect 6604 17688 6610 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 7056 17731 7114 17737
rect 7056 17728 7068 17731
rect 6880 17700 7068 17728
rect 6880 17688 6886 17700
rect 7056 17697 7068 17700
rect 7102 17697 7114 17731
rect 8846 17728 8852 17740
rect 8807 17700 8852 17728
rect 7056 17691 7114 17697
rect 8846 17688 8852 17700
rect 8904 17688 8910 17740
rect 10045 17731 10103 17737
rect 10045 17697 10057 17731
rect 10091 17728 10103 17731
rect 10502 17728 10508 17740
rect 10091 17700 10508 17728
rect 10091 17697 10103 17700
rect 10045 17691 10103 17697
rect 10502 17688 10508 17700
rect 10560 17688 10566 17740
rect 10704 17737 10732 17768
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 12250 17796 12256 17808
rect 11756 17768 12256 17796
rect 11756 17756 11762 17768
rect 12250 17756 12256 17768
rect 12308 17756 12314 17808
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 14108 17796 14136 17827
rect 16390 17824 16396 17836
rect 16448 17824 16454 17876
rect 16482 17824 16488 17876
rect 16540 17864 16546 17876
rect 17218 17864 17224 17876
rect 16540 17836 16585 17864
rect 16960 17836 17224 17864
rect 16540 17824 16546 17836
rect 12492 17768 14136 17796
rect 15657 17799 15715 17805
rect 12492 17756 12498 17768
rect 15657 17765 15669 17799
rect 15703 17796 15715 17799
rect 16022 17796 16028 17808
rect 15703 17768 16028 17796
rect 15703 17765 15715 17768
rect 15657 17759 15715 17765
rect 16022 17756 16028 17768
rect 16080 17756 16086 17808
rect 16960 17796 16988 17836
rect 17218 17824 17224 17836
rect 17276 17824 17282 17876
rect 19242 17824 19248 17876
rect 19300 17864 19306 17876
rect 19889 17867 19947 17873
rect 19889 17864 19901 17867
rect 19300 17836 19901 17864
rect 19300 17824 19306 17836
rect 19889 17833 19901 17836
rect 19935 17833 19947 17867
rect 19889 17827 19947 17833
rect 21269 17867 21327 17873
rect 21269 17833 21281 17867
rect 21315 17864 21327 17867
rect 21358 17864 21364 17876
rect 21315 17836 21364 17864
rect 21315 17833 21327 17836
rect 21269 17827 21327 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22152 17836 22197 17864
rect 22152 17824 22158 17836
rect 16224 17768 16988 17796
rect 10689 17731 10747 17737
rect 10689 17697 10701 17731
rect 10735 17697 10747 17731
rect 10689 17691 10747 17697
rect 11885 17731 11943 17737
rect 11885 17697 11897 17731
rect 11931 17728 11943 17731
rect 12704 17731 12762 17737
rect 12704 17728 12716 17731
rect 11931 17700 12716 17728
rect 11931 17697 11943 17700
rect 11885 17691 11943 17697
rect 12704 17697 12716 17700
rect 12750 17728 12762 17731
rect 13814 17728 13820 17740
rect 12750 17700 13820 17728
rect 12750 17697 12762 17700
rect 12704 17691 12762 17697
rect 13814 17688 13820 17700
rect 13872 17688 13878 17740
rect 13998 17688 14004 17740
rect 14056 17728 14062 17740
rect 14461 17731 14519 17737
rect 14461 17728 14473 17731
rect 14056 17700 14473 17728
rect 14056 17688 14062 17700
rect 14461 17697 14473 17700
rect 14507 17697 14519 17731
rect 14461 17691 14519 17697
rect 1486 17620 1492 17672
rect 1544 17660 1550 17672
rect 1581 17663 1639 17669
rect 1581 17660 1593 17663
rect 1544 17632 1593 17660
rect 1544 17620 1550 17632
rect 1581 17629 1593 17632
rect 1627 17629 1639 17663
rect 1581 17623 1639 17629
rect 1596 17524 1624 17623
rect 7190 17620 7196 17672
rect 7248 17660 7254 17672
rect 7466 17660 7472 17672
rect 7248 17632 7293 17660
rect 7427 17632 7472 17660
rect 7248 17620 7254 17632
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 7834 17620 7840 17672
rect 7892 17660 7898 17672
rect 8665 17663 8723 17669
rect 8665 17660 8677 17663
rect 7892 17632 8677 17660
rect 7892 17620 7898 17632
rect 8665 17629 8677 17632
rect 8711 17629 8723 17663
rect 10134 17660 10140 17672
rect 10095 17632 10140 17660
rect 8665 17623 8723 17629
rect 10134 17620 10140 17632
rect 10192 17620 10198 17672
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17660 10379 17663
rect 11698 17660 11704 17672
rect 10367 17632 11704 17660
rect 10367 17629 10379 17632
rect 10321 17623 10379 17629
rect 11698 17620 11704 17632
rect 11756 17660 11762 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 11756 17632 11989 17660
rect 11756 17620 11762 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 12158 17620 12164 17672
rect 12216 17660 12222 17672
rect 12437 17663 12495 17669
rect 12437 17660 12449 17663
rect 12216 17632 12449 17660
rect 12216 17620 12222 17632
rect 12437 17629 12449 17632
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 14553 17663 14611 17669
rect 14553 17660 14565 17663
rect 14148 17632 14565 17660
rect 14148 17620 14154 17632
rect 14553 17629 14565 17632
rect 14599 17629 14611 17663
rect 14734 17660 14740 17672
rect 14695 17632 14740 17660
rect 14553 17623 14611 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 15010 17620 15016 17672
rect 15068 17660 15074 17672
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15068 17632 15853 17660
rect 15068 17620 15074 17632
rect 15841 17629 15853 17632
rect 15887 17660 15899 17663
rect 16224 17660 16252 17768
rect 17034 17756 17040 17808
rect 17092 17805 17098 17808
rect 17092 17799 17156 17805
rect 17092 17765 17110 17799
rect 17144 17765 17156 17799
rect 17092 17759 17156 17765
rect 18776 17799 18834 17805
rect 18776 17765 18788 17799
rect 18822 17796 18834 17799
rect 18874 17796 18880 17808
rect 18822 17768 18880 17796
rect 18822 17765 18834 17768
rect 18776 17759 18834 17765
rect 17092 17756 17098 17759
rect 18874 17756 18880 17768
rect 18932 17756 18938 17808
rect 18966 17756 18972 17808
rect 19024 17796 19030 17808
rect 23566 17796 23572 17808
rect 19024 17768 23572 17796
rect 19024 17756 19030 17768
rect 23566 17756 23572 17768
rect 23624 17756 23630 17808
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17697 16359 17731
rect 20162 17728 20168 17740
rect 20123 17700 20168 17728
rect 16301 17691 16359 17697
rect 15887 17632 16252 17660
rect 15887 17629 15899 17632
rect 15841 17623 15899 17629
rect 10873 17595 10931 17601
rect 10873 17592 10885 17595
rect 8128 17564 10885 17592
rect 2314 17524 2320 17536
rect 1596 17496 2320 17524
rect 2314 17484 2320 17496
rect 2372 17484 2378 17536
rect 4062 17484 4068 17536
rect 4120 17524 4126 17536
rect 8128 17524 8156 17564
rect 10873 17561 10885 17564
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 11425 17595 11483 17601
rect 11425 17561 11437 17595
rect 11471 17592 11483 17595
rect 11790 17592 11796 17604
rect 11471 17564 11796 17592
rect 11471 17561 11483 17564
rect 11425 17555 11483 17561
rect 11790 17552 11796 17564
rect 11848 17552 11854 17604
rect 16316 17592 16344 17691
rect 20162 17688 20168 17700
rect 20220 17688 20226 17740
rect 20898 17688 20904 17740
rect 20956 17728 20962 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 20956 17700 21373 17728
rect 20956 17688 20962 17700
rect 21361 17697 21373 17700
rect 21407 17697 21419 17731
rect 21361 17691 21419 17697
rect 21913 17731 21971 17737
rect 21913 17697 21925 17731
rect 21959 17697 21971 17731
rect 21913 17691 21971 17697
rect 16850 17660 16856 17672
rect 16811 17632 16856 17660
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 18138 17620 18144 17672
rect 18196 17660 18202 17672
rect 18414 17660 18420 17672
rect 18196 17632 18420 17660
rect 18196 17620 18202 17632
rect 18414 17620 18420 17632
rect 18472 17660 18478 17672
rect 18509 17663 18567 17669
rect 18509 17660 18521 17663
rect 18472 17632 18521 17660
rect 18472 17620 18478 17632
rect 18509 17629 18521 17632
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 21453 17663 21511 17669
rect 21453 17629 21465 17663
rect 21499 17629 21511 17663
rect 21453 17623 21511 17629
rect 20901 17595 20959 17601
rect 20901 17592 20913 17595
rect 13372 17564 16344 17592
rect 19444 17564 20913 17592
rect 8570 17524 8576 17536
rect 4120 17496 8156 17524
rect 8531 17496 8576 17524
rect 4120 17484 4126 17496
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 8665 17527 8723 17533
rect 8665 17493 8677 17527
rect 8711 17524 8723 17527
rect 12342 17524 12348 17536
rect 8711 17496 12348 17524
rect 8711 17493 8723 17496
rect 8665 17487 8723 17493
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 13372 17524 13400 17564
rect 12676 17496 13400 17524
rect 12676 17484 12682 17496
rect 14642 17484 14648 17536
rect 14700 17524 14706 17536
rect 15289 17527 15347 17533
rect 15289 17524 15301 17527
rect 14700 17496 15301 17524
rect 14700 17484 14706 17496
rect 15289 17493 15301 17496
rect 15335 17493 15347 17527
rect 15289 17487 15347 17493
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 18233 17527 18291 17533
rect 18233 17524 18245 17527
rect 17184 17496 18245 17524
rect 17184 17484 17190 17496
rect 18233 17493 18245 17496
rect 18279 17493 18291 17527
rect 18233 17487 18291 17493
rect 18690 17484 18696 17536
rect 18748 17524 18754 17536
rect 19444 17524 19472 17564
rect 20901 17561 20913 17564
rect 20947 17561 20959 17595
rect 20901 17555 20959 17561
rect 21174 17552 21180 17604
rect 21232 17592 21238 17604
rect 21358 17592 21364 17604
rect 21232 17564 21364 17592
rect 21232 17552 21238 17564
rect 21358 17552 21364 17564
rect 21416 17592 21422 17604
rect 21468 17592 21496 17623
rect 21416 17564 21496 17592
rect 21416 17552 21422 17564
rect 20346 17524 20352 17536
rect 18748 17496 19472 17524
rect 20307 17496 20352 17524
rect 18748 17484 18754 17496
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 20530 17484 20536 17536
rect 20588 17524 20594 17536
rect 21928 17524 21956 17691
rect 20588 17496 21956 17524
rect 20588 17484 20594 17496
rect 1104 17434 22816 17456
rect 1104 17382 4614 17434
rect 4666 17382 4678 17434
rect 4730 17382 4742 17434
rect 4794 17382 4806 17434
rect 4858 17382 11878 17434
rect 11930 17382 11942 17434
rect 11994 17382 12006 17434
rect 12058 17382 12070 17434
rect 12122 17382 19142 17434
rect 19194 17382 19206 17434
rect 19258 17382 19270 17434
rect 19322 17382 19334 17434
rect 19386 17382 22816 17434
rect 1104 17360 22816 17382
rect 934 17280 940 17332
rect 992 17320 998 17332
rect 1857 17323 1915 17329
rect 1857 17320 1869 17323
rect 992 17292 1869 17320
rect 992 17280 998 17292
rect 1857 17289 1869 17292
rect 1903 17289 1915 17323
rect 1857 17283 1915 17289
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 3602 17320 3608 17332
rect 2280 17292 3608 17320
rect 2280 17280 2286 17292
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 10502 17320 10508 17332
rect 4264 17292 10088 17320
rect 10463 17292 10508 17320
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17116 1731 17119
rect 2130 17116 2136 17128
rect 1719 17088 2136 17116
rect 1719 17085 1731 17088
rect 1673 17079 1731 17085
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 2222 17076 2228 17128
rect 2280 17116 2286 17128
rect 2492 17119 2550 17125
rect 2280 17088 2325 17116
rect 2280 17076 2286 17088
rect 2492 17085 2504 17119
rect 2538 17116 2550 17119
rect 3694 17116 3700 17128
rect 2538 17088 3700 17116
rect 2538 17085 2550 17088
rect 2492 17079 2550 17085
rect 3694 17076 3700 17088
rect 3752 17076 3758 17128
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 4065 17119 4123 17125
rect 4065 17116 4077 17119
rect 3844 17088 4077 17116
rect 3844 17076 3850 17088
rect 4065 17085 4077 17088
rect 4111 17085 4123 17119
rect 4065 17079 4123 17085
rect 4264 17048 4292 17292
rect 6457 17255 6515 17261
rect 6457 17221 6469 17255
rect 6503 17252 6515 17255
rect 7466 17252 7472 17264
rect 6503 17224 7472 17252
rect 6503 17221 6515 17224
rect 6457 17215 6515 17221
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 5080 17187 5138 17193
rect 5080 17184 5092 17187
rect 4396 17156 5092 17184
rect 4396 17144 4402 17156
rect 5080 17153 5092 17156
rect 5126 17153 5138 17187
rect 5080 17147 5138 17153
rect 5258 17144 5264 17196
rect 5316 17184 5322 17196
rect 6472 17184 6500 17215
rect 7466 17212 7472 17224
rect 7524 17212 7530 17264
rect 10060 17252 10088 17292
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 11333 17323 11391 17329
rect 11333 17289 11345 17323
rect 11379 17320 11391 17323
rect 11422 17320 11428 17332
rect 11379 17292 11428 17320
rect 11379 17289 11391 17292
rect 11333 17283 11391 17289
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 12434 17320 12440 17332
rect 11900 17292 12440 17320
rect 10965 17255 11023 17261
rect 10965 17252 10977 17255
rect 10060 17224 10977 17252
rect 10965 17221 10977 17224
rect 11011 17221 11023 17255
rect 10965 17215 11023 17221
rect 11900 17196 11928 17292
rect 12434 17280 12440 17292
rect 12492 17280 12498 17332
rect 13814 17320 13820 17332
rect 13775 17292 13820 17320
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 20806 17280 20812 17332
rect 20864 17320 20870 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 20864 17292 21465 17320
rect 20864 17280 20870 17292
rect 21453 17289 21465 17292
rect 21499 17289 21511 17323
rect 21453 17283 21511 17289
rect 12158 17212 12164 17264
rect 12216 17252 12222 17264
rect 12253 17255 12311 17261
rect 12253 17252 12265 17255
rect 12216 17224 12265 17252
rect 12216 17212 12222 17224
rect 12253 17221 12265 17224
rect 12299 17221 12311 17255
rect 12253 17215 12311 17221
rect 14001 17255 14059 17261
rect 14001 17221 14013 17255
rect 14047 17252 14059 17255
rect 14093 17255 14151 17261
rect 14093 17252 14105 17255
rect 14047 17224 14105 17252
rect 14047 17221 14059 17224
rect 14001 17215 14059 17221
rect 14093 17221 14105 17224
rect 14139 17252 14151 17255
rect 14182 17252 14188 17264
rect 14139 17224 14188 17252
rect 14139 17221 14151 17224
rect 14093 17215 14151 17221
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 14274 17212 14280 17264
rect 14332 17212 14338 17264
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18785 17255 18843 17261
rect 18785 17252 18797 17255
rect 18012 17224 18797 17252
rect 18012 17212 18018 17224
rect 18785 17221 18797 17224
rect 18831 17221 18843 17255
rect 18785 17215 18843 17221
rect 5316 17156 6500 17184
rect 5316 17144 5322 17156
rect 6638 17144 6644 17196
rect 6696 17184 6702 17196
rect 9132 17187 9190 17193
rect 6696 17156 7604 17184
rect 6696 17144 6702 17156
rect 4614 17116 4620 17128
rect 4575 17088 4620 17116
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17116 5411 17119
rect 6362 17116 6368 17128
rect 5399 17088 6368 17116
rect 5399 17085 5411 17088
rect 5353 17079 5411 17085
rect 6362 17076 6368 17088
rect 6420 17076 6426 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6604 17088 6837 17116
rect 6604 17076 6610 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7064 17088 7481 17116
rect 7064 17076 7070 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 7576 17116 7604 17156
rect 9132 17153 9144 17187
rect 9178 17184 9190 17187
rect 9178 17156 9260 17184
rect 9178 17153 9190 17156
rect 9132 17147 9190 17153
rect 7725 17119 7783 17125
rect 7725 17116 7737 17119
rect 7576 17088 7737 17116
rect 7469 17079 7527 17085
rect 7725 17085 7737 17088
rect 7771 17116 7783 17119
rect 8018 17116 8024 17128
rect 7771 17088 8024 17116
rect 7771 17085 7783 17088
rect 7725 17079 7783 17085
rect 2516 17020 4292 17048
rect 2516 16992 2544 17020
rect 6730 17008 6736 17060
rect 6788 17048 6794 17060
rect 7484 17048 7512 17079
rect 8018 17076 8024 17088
rect 8076 17076 8082 17128
rect 9122 17048 9128 17060
rect 6788 17020 7420 17048
rect 7484 17020 9128 17048
rect 6788 17008 6794 17020
rect 2498 16940 2504 16992
rect 2556 16940 2562 16992
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4430 16980 4436 16992
rect 4295 16952 4436 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 5083 16983 5141 16989
rect 5083 16949 5095 16983
rect 5129 16980 5141 16983
rect 6822 16980 6828 16992
rect 5129 16952 6828 16980
rect 5129 16949 5141 16952
rect 5083 16943 5141 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 6914 16940 6920 16992
rect 6972 16980 6978 16992
rect 7009 16983 7067 16989
rect 7009 16980 7021 16983
rect 6972 16952 7021 16980
rect 6972 16940 6978 16952
rect 7009 16949 7021 16952
rect 7055 16949 7067 16983
rect 7392 16980 7420 17020
rect 9122 17008 9128 17020
rect 9180 17048 9186 17060
rect 9232 17048 9260 17156
rect 11698 17144 11704 17196
rect 11756 17184 11762 17196
rect 11882 17184 11888 17196
rect 11756 17156 11888 17184
rect 11756 17144 11762 17156
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 14292 17184 14320 17212
rect 12268 17156 12572 17184
rect 9392 17119 9450 17125
rect 9392 17116 9404 17119
rect 9180 17020 9260 17048
rect 9324 17088 9404 17116
rect 9180 17008 9186 17020
rect 8570 16980 8576 16992
rect 7392 16952 8576 16980
rect 7009 16943 7067 16949
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 8849 16983 8907 16989
rect 8849 16949 8861 16983
rect 8895 16980 8907 16983
rect 9324 16980 9352 17088
rect 9392 17085 9404 17088
rect 9438 17116 9450 17119
rect 10134 17116 10140 17128
rect 9438 17088 10140 17116
rect 9438 17085 9450 17088
rect 9392 17079 9450 17085
rect 10134 17076 10140 17088
rect 10192 17076 10198 17128
rect 10778 17116 10784 17128
rect 10739 17088 10784 17116
rect 10778 17076 10784 17088
rect 10836 17076 10842 17128
rect 12268 17116 12296 17156
rect 11624 17088 12296 17116
rect 12345 17119 12403 17125
rect 9582 17008 9588 17060
rect 9640 17048 9646 17060
rect 11624 17048 11652 17088
rect 12345 17085 12357 17119
rect 12391 17116 12403 17119
rect 12434 17116 12440 17128
rect 12391 17088 12440 17116
rect 12391 17085 12403 17088
rect 12345 17079 12403 17085
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12544 17116 12572 17156
rect 13464 17156 14320 17184
rect 12544 17088 13124 17116
rect 9640 17020 11652 17048
rect 11701 17051 11759 17057
rect 9640 17008 9646 17020
rect 11701 17017 11713 17051
rect 11747 17048 11759 17051
rect 12526 17048 12532 17060
rect 11747 17020 12532 17048
rect 11747 17017 11759 17020
rect 11701 17011 11759 17017
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 12704 17051 12762 17057
rect 12704 17017 12716 17051
rect 12750 17048 12762 17051
rect 12802 17048 12808 17060
rect 12750 17020 12808 17048
rect 12750 17017 12762 17020
rect 12704 17011 12762 17017
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 8895 16952 9352 16980
rect 11793 16983 11851 16989
rect 8895 16949 8907 16952
rect 8849 16943 8907 16949
rect 11793 16949 11805 16983
rect 11839 16980 11851 16983
rect 12618 16980 12624 16992
rect 11839 16952 12624 16980
rect 11839 16949 11851 16952
rect 11793 16943 11851 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13096 16980 13124 17088
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 13464 17116 13492 17156
rect 17494 17144 17500 17196
rect 17552 17184 17558 17196
rect 19245 17187 19303 17193
rect 19245 17184 19257 17187
rect 17552 17156 19257 17184
rect 17552 17144 17558 17156
rect 19245 17153 19257 17156
rect 19291 17153 19303 17187
rect 19245 17147 19303 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19702 17184 19708 17196
rect 19475 17156 19708 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 21818 17184 21824 17196
rect 20864 17156 21824 17184
rect 20864 17144 20870 17156
rect 21818 17144 21824 17156
rect 21876 17184 21882 17196
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 21876 17156 22017 17184
rect 21876 17144 21882 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 13228 17088 13492 17116
rect 13228 17076 13234 17088
rect 13538 17076 13544 17128
rect 13596 17116 13602 17128
rect 13909 17119 13967 17125
rect 13909 17116 13921 17119
rect 13596 17088 13921 17116
rect 13596 17076 13602 17088
rect 13909 17085 13921 17088
rect 13955 17085 13967 17119
rect 13909 17079 13967 17085
rect 14182 17076 14188 17128
rect 14240 17116 14246 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 14240 17088 14289 17116
rect 14240 17076 14246 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 14369 17119 14427 17125
rect 14369 17085 14381 17119
rect 14415 17116 14427 17119
rect 14918 17116 14924 17128
rect 14415 17088 14924 17116
rect 14415 17085 14427 17088
rect 14369 17079 14427 17085
rect 14918 17076 14924 17088
rect 14976 17076 14982 17128
rect 16025 17119 16083 17125
rect 16025 17085 16037 17119
rect 16071 17116 16083 17119
rect 16850 17116 16856 17128
rect 16071 17088 16856 17116
rect 16071 17085 16083 17088
rect 16025 17079 16083 17085
rect 16850 17076 16856 17088
rect 16908 17116 16914 17128
rect 17862 17116 17868 17128
rect 16908 17088 17724 17116
rect 17823 17088 17868 17116
rect 16908 17076 16914 17088
rect 14636 17051 14694 17057
rect 14636 17017 14648 17051
rect 14682 17048 14694 17051
rect 14734 17048 14740 17060
rect 14682 17020 14740 17048
rect 14682 17017 14694 17020
rect 14636 17011 14694 17017
rect 14734 17008 14740 17020
rect 14792 17048 14798 17060
rect 15378 17048 15384 17060
rect 14792 17020 15384 17048
rect 14792 17008 14798 17020
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 16114 17008 16120 17060
rect 16172 17048 16178 17060
rect 16292 17051 16350 17057
rect 16292 17048 16304 17051
rect 16172 17020 16304 17048
rect 16172 17008 16178 17020
rect 16292 17017 16304 17020
rect 16338 17048 16350 17051
rect 16482 17048 16488 17060
rect 16338 17020 16488 17048
rect 16338 17017 16350 17020
rect 16292 17011 16350 17017
rect 16482 17008 16488 17020
rect 16540 17008 16546 17060
rect 15194 16980 15200 16992
rect 13096 16952 15200 16980
rect 15194 16940 15200 16952
rect 15252 16980 15258 16992
rect 15749 16983 15807 16989
rect 15749 16980 15761 16983
rect 15252 16952 15761 16980
rect 15252 16940 15258 16952
rect 15749 16949 15761 16952
rect 15795 16949 15807 16983
rect 15749 16943 15807 16949
rect 17034 16940 17040 16992
rect 17092 16980 17098 16992
rect 17696 16989 17724 17088
rect 17862 17076 17868 17088
rect 17920 17076 17926 17128
rect 18230 17116 18236 17128
rect 18191 17088 18236 17116
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 19797 17119 19855 17125
rect 19797 17116 19809 17119
rect 19116 17088 19809 17116
rect 19116 17076 19122 17088
rect 19797 17085 19809 17088
rect 19843 17085 19855 17119
rect 19797 17079 19855 17085
rect 19153 17051 19211 17057
rect 19153 17048 19165 17051
rect 18432 17020 19165 17048
rect 17405 16983 17463 16989
rect 17405 16980 17417 16983
rect 17092 16952 17417 16980
rect 17092 16940 17098 16952
rect 17405 16949 17417 16952
rect 17451 16949 17463 16983
rect 17405 16943 17463 16949
rect 17681 16983 17739 16989
rect 17681 16949 17693 16983
rect 17727 16980 17739 16983
rect 18138 16980 18144 16992
rect 17727 16952 18144 16980
rect 17727 16949 17739 16952
rect 17681 16943 17739 16949
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 18432 16989 18460 17020
rect 19153 17017 19165 17020
rect 19199 17017 19211 17051
rect 19153 17011 19211 17017
rect 18417 16983 18475 16989
rect 18417 16949 18429 16983
rect 18463 16949 18475 16983
rect 19812 16980 19840 17079
rect 20438 17076 20444 17128
rect 20496 17116 20502 17128
rect 21913 17119 21971 17125
rect 21913 17116 21925 17119
rect 20496 17088 21925 17116
rect 20496 17076 20502 17088
rect 21913 17085 21925 17088
rect 21959 17085 21971 17119
rect 21913 17079 21971 17085
rect 20064 17051 20122 17057
rect 20064 17017 20076 17051
rect 20110 17048 20122 17051
rect 20110 17020 21864 17048
rect 20110 17017 20122 17020
rect 20064 17011 20122 17017
rect 21836 16992 21864 17020
rect 20990 16980 20996 16992
rect 19812 16952 20996 16980
rect 18417 16943 18475 16949
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 21174 16980 21180 16992
rect 21135 16952 21180 16980
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21818 16980 21824 16992
rect 21779 16952 21824 16980
rect 21818 16940 21824 16952
rect 21876 16940 21882 16992
rect 1104 16890 22816 16912
rect 1104 16838 8246 16890
rect 8298 16838 8310 16890
rect 8362 16838 8374 16890
rect 8426 16838 8438 16890
rect 8490 16838 15510 16890
rect 15562 16838 15574 16890
rect 15626 16838 15638 16890
rect 15690 16838 15702 16890
rect 15754 16838 22816 16890
rect 1104 16816 22816 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1765 16779 1823 16785
rect 1765 16776 1777 16779
rect 1728 16748 1777 16776
rect 1728 16736 1734 16748
rect 1765 16745 1777 16748
rect 1811 16745 1823 16779
rect 1765 16739 1823 16745
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 4062 16776 4068 16788
rect 2188 16748 4068 16776
rect 2188 16736 2194 16748
rect 4062 16736 4068 16748
rect 4120 16736 4126 16788
rect 4246 16776 4252 16788
rect 4207 16748 4252 16776
rect 4246 16736 4252 16748
rect 4304 16736 4310 16788
rect 4617 16779 4675 16785
rect 4617 16745 4629 16779
rect 4663 16776 4675 16779
rect 4890 16776 4896 16788
rect 4663 16748 4896 16776
rect 4663 16745 4675 16748
rect 4617 16739 4675 16745
rect 4890 16736 4896 16748
rect 4948 16736 4954 16788
rect 4985 16779 5043 16785
rect 4985 16745 4997 16779
rect 5031 16776 5043 16779
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5031 16748 5641 16776
rect 5031 16745 5043 16748
rect 4985 16739 5043 16745
rect 5629 16745 5641 16748
rect 5675 16776 5687 16779
rect 8757 16779 8815 16785
rect 8757 16776 8769 16779
rect 5675 16748 8769 16776
rect 5675 16745 5687 16748
rect 5629 16739 5687 16745
rect 8757 16745 8769 16748
rect 8803 16745 8815 16779
rect 8757 16739 8815 16745
rect 9309 16779 9367 16785
rect 9309 16745 9321 16779
rect 9355 16776 9367 16779
rect 9674 16776 9680 16788
rect 9355 16748 9680 16776
rect 9355 16745 9367 16748
rect 9309 16739 9367 16745
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 10778 16736 10784 16788
rect 10836 16776 10842 16788
rect 11057 16779 11115 16785
rect 11057 16776 11069 16779
rect 10836 16748 11069 16776
rect 10836 16736 10842 16748
rect 11057 16745 11069 16748
rect 11103 16776 11115 16779
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11103 16748 11805 16776
rect 11103 16745 11115 16748
rect 11057 16739 11115 16745
rect 11793 16745 11805 16748
rect 11839 16745 11851 16779
rect 18785 16779 18843 16785
rect 11793 16739 11851 16745
rect 11900 16748 17540 16776
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 2400 16711 2458 16717
rect 1912 16680 2360 16708
rect 1912 16668 1918 16680
rect 1578 16640 1584 16652
rect 1539 16612 1584 16640
rect 1578 16600 1584 16612
rect 1636 16600 1642 16652
rect 2133 16643 2191 16649
rect 2133 16609 2145 16643
rect 2179 16640 2191 16643
rect 2222 16640 2228 16652
rect 2179 16612 2228 16640
rect 2179 16609 2191 16612
rect 2133 16603 2191 16609
rect 2222 16600 2228 16612
rect 2280 16600 2286 16652
rect 2332 16640 2360 16680
rect 2400 16677 2412 16711
rect 2446 16708 2458 16711
rect 3142 16708 3148 16720
rect 2446 16680 3148 16708
rect 2446 16677 2458 16680
rect 2400 16671 2458 16677
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 5077 16711 5135 16717
rect 5077 16677 5089 16711
rect 5123 16708 5135 16711
rect 5258 16708 5264 16720
rect 5123 16680 5264 16708
rect 5123 16677 5135 16680
rect 5077 16671 5135 16677
rect 5258 16668 5264 16680
rect 5316 16668 5322 16720
rect 6089 16711 6147 16717
rect 6089 16677 6101 16711
rect 6135 16708 6147 16711
rect 7834 16708 7840 16720
rect 6135 16680 7840 16708
rect 6135 16677 6147 16680
rect 6089 16671 6147 16677
rect 7834 16668 7840 16680
rect 7892 16668 7898 16720
rect 8662 16708 8668 16720
rect 8623 16680 8668 16708
rect 8662 16668 8668 16680
rect 8720 16668 8726 16720
rect 9122 16668 9128 16720
rect 9180 16708 9186 16720
rect 9944 16711 10002 16717
rect 9180 16680 9720 16708
rect 9180 16668 9186 16680
rect 4065 16643 4123 16649
rect 4065 16640 4077 16643
rect 2332 16612 4077 16640
rect 4065 16609 4077 16612
rect 4111 16609 4123 16643
rect 5994 16640 6000 16652
rect 5955 16612 6000 16640
rect 4065 16603 4123 16609
rect 5994 16600 6000 16612
rect 6052 16600 6058 16652
rect 6362 16600 6368 16652
rect 6420 16640 6426 16652
rect 6546 16640 6552 16652
rect 6420 16612 6552 16640
rect 6420 16600 6426 16612
rect 6546 16600 6552 16612
rect 6604 16600 6610 16652
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16640 6699 16643
rect 6730 16640 6736 16652
rect 6687 16612 6736 16640
rect 6687 16609 6699 16612
rect 6641 16603 6699 16609
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 6908 16643 6966 16649
rect 6908 16609 6920 16643
rect 6954 16640 6966 16643
rect 6954 16612 8033 16640
rect 6954 16609 6966 16612
rect 6908 16603 6966 16609
rect 5166 16532 5172 16584
rect 5224 16572 5230 16584
rect 6178 16572 6184 16584
rect 5224 16544 5269 16572
rect 6139 16544 6184 16572
rect 5224 16532 5230 16544
rect 6178 16532 6184 16544
rect 6236 16532 6242 16584
rect 8005 16572 8033 16612
rect 9214 16600 9220 16652
rect 9272 16640 9278 16652
rect 9692 16649 9720 16680
rect 9944 16677 9956 16711
rect 9990 16708 10002 16711
rect 10502 16708 10508 16720
rect 9990 16680 10508 16708
rect 9990 16677 10002 16680
rect 9944 16671 10002 16677
rect 10502 16668 10508 16680
rect 10560 16668 10566 16720
rect 11900 16708 11928 16748
rect 11072 16680 11928 16708
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9272 16612 9505 16640
rect 9272 16600 9278 16612
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 9493 16603 9551 16609
rect 9677 16643 9735 16649
rect 9677 16609 9689 16643
rect 9723 16609 9735 16643
rect 11072 16640 11100 16680
rect 12802 16668 12808 16720
rect 12860 16708 12866 16720
rect 13998 16708 14004 16720
rect 12860 16680 14004 16708
rect 12860 16668 12866 16680
rect 9677 16603 9735 16609
rect 9784 16612 11100 16640
rect 8110 16572 8116 16584
rect 8005 16544 8116 16572
rect 8110 16532 8116 16544
rect 8168 16572 8174 16584
rect 8849 16575 8907 16581
rect 8849 16572 8861 16575
rect 8168 16544 8861 16572
rect 8168 16532 8174 16544
rect 8849 16541 8861 16544
rect 8895 16541 8907 16575
rect 8849 16535 8907 16541
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 9784 16572 9812 16612
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11698 16640 11704 16652
rect 11204 16612 11376 16640
rect 11659 16612 11704 16640
rect 11204 16600 11210 16612
rect 9640 16544 9812 16572
rect 9640 16532 9646 16544
rect 3513 16507 3571 16513
rect 3513 16473 3525 16507
rect 3559 16504 3571 16507
rect 3694 16504 3700 16516
rect 3559 16476 3700 16504
rect 3559 16473 3571 16476
rect 3513 16467 3571 16473
rect 3694 16464 3700 16476
rect 3752 16464 3758 16516
rect 8018 16504 8024 16516
rect 7979 16476 8024 16504
rect 8018 16464 8024 16476
rect 8076 16464 8082 16516
rect 8297 16507 8355 16513
rect 8297 16473 8309 16507
rect 8343 16504 8355 16507
rect 8570 16504 8576 16516
rect 8343 16476 8576 16504
rect 8343 16473 8355 16476
rect 8297 16467 8355 16473
rect 8570 16464 8576 16476
rect 8628 16464 8634 16516
rect 11348 16513 11376 16612
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 12434 16640 12440 16652
rect 12395 16612 12440 16640
rect 12434 16600 12440 16612
rect 12492 16600 12498 16652
rect 12704 16643 12762 16649
rect 12704 16609 12716 16643
rect 12750 16640 12762 16643
rect 13722 16640 13728 16652
rect 12750 16612 13728 16640
rect 12750 16609 12762 16612
rect 12704 16603 12762 16609
rect 13722 16600 13728 16612
rect 13780 16600 13786 16652
rect 11606 16532 11612 16584
rect 11664 16572 11670 16584
rect 11882 16572 11888 16584
rect 11664 16544 11888 16572
rect 11664 16532 11670 16544
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 13832 16513 13860 16680
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 14182 16668 14188 16720
rect 14240 16708 14246 16720
rect 17512 16708 17540 16748
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 18874 16776 18880 16788
rect 18831 16748 18880 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 18874 16736 18880 16748
rect 18932 16736 18938 16788
rect 20533 16779 20591 16785
rect 20533 16745 20545 16779
rect 20579 16776 20591 16779
rect 21818 16776 21824 16788
rect 20579 16748 21824 16776
rect 20579 16745 20591 16748
rect 20533 16739 20591 16745
rect 21818 16736 21824 16748
rect 21876 16736 21882 16788
rect 22278 16708 22284 16720
rect 14240 16680 16068 16708
rect 17512 16680 22284 16708
rect 14240 16668 14246 16680
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 13964 16612 14473 16640
rect 13964 16600 13970 16612
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 15289 16643 15347 16649
rect 15289 16609 15301 16643
rect 15335 16640 15347 16643
rect 15930 16640 15936 16652
rect 15335 16612 15936 16640
rect 15335 16609 15347 16612
rect 15289 16603 15347 16609
rect 15930 16600 15936 16612
rect 15988 16600 15994 16652
rect 16040 16649 16068 16680
rect 22278 16668 22284 16680
rect 22336 16668 22342 16720
rect 16025 16643 16083 16649
rect 16025 16609 16037 16643
rect 16071 16609 16083 16643
rect 16025 16603 16083 16609
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 16850 16640 16856 16652
rect 16264 16612 16623 16640
rect 16811 16612 16856 16640
rect 16264 16600 16270 16612
rect 13998 16532 14004 16584
rect 14056 16572 14062 16584
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14056 16544 14565 16572
rect 14056 16532 14062 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 14737 16575 14795 16581
rect 14737 16541 14749 16575
rect 14783 16572 14795 16575
rect 14826 16572 14832 16584
rect 14783 16544 14832 16572
rect 14783 16541 14795 16544
rect 14737 16535 14795 16541
rect 14826 16532 14832 16544
rect 14884 16532 14890 16584
rect 16114 16572 16120 16584
rect 16075 16544 16120 16572
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 16390 16532 16396 16584
rect 16448 16581 16454 16584
rect 16595 16581 16623 16612
rect 16850 16600 16856 16612
rect 16908 16600 16914 16652
rect 18601 16643 18659 16649
rect 18601 16609 18613 16643
rect 18647 16640 18659 16643
rect 18690 16640 18696 16652
rect 18647 16612 18696 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 19420 16643 19478 16649
rect 19420 16609 19432 16643
rect 19466 16640 19478 16643
rect 20438 16640 20444 16652
rect 19466 16612 20444 16640
rect 19466 16609 19478 16612
rect 19420 16603 19478 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20901 16643 20959 16649
rect 20901 16609 20913 16643
rect 20947 16640 20959 16643
rect 20990 16640 20996 16652
rect 20947 16612 20996 16640
rect 20947 16609 20959 16612
rect 20901 16603 20959 16609
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 21174 16649 21180 16652
rect 21168 16640 21180 16649
rect 21135 16612 21180 16640
rect 21168 16603 21180 16612
rect 21174 16600 21180 16603
rect 21232 16600 21238 16652
rect 16448 16575 16498 16581
rect 16448 16541 16452 16575
rect 16486 16541 16498 16575
rect 16448 16535 16498 16541
rect 16580 16575 16638 16581
rect 16580 16541 16592 16575
rect 16626 16541 16638 16575
rect 16580 16535 16638 16541
rect 16448 16532 16454 16535
rect 18138 16532 18144 16584
rect 18196 16572 18202 16584
rect 19058 16572 19064 16584
rect 18196 16544 19064 16572
rect 18196 16532 18202 16544
rect 19058 16532 19064 16544
rect 19116 16572 19122 16584
rect 19153 16575 19211 16581
rect 19153 16572 19165 16575
rect 19116 16544 19165 16572
rect 19116 16532 19122 16544
rect 19153 16541 19165 16544
rect 19199 16541 19211 16575
rect 19153 16535 19211 16541
rect 11333 16507 11391 16513
rect 11333 16473 11345 16507
rect 11379 16473 11391 16507
rect 11333 16467 11391 16473
rect 13817 16507 13875 16513
rect 13817 16473 13829 16507
rect 13863 16473 13875 16507
rect 16132 16504 16160 16532
rect 13817 16467 13875 16473
rect 14016 16476 16160 16504
rect 1394 16396 1400 16448
rect 1452 16436 1458 16448
rect 6546 16436 6552 16448
rect 1452 16408 6552 16436
rect 1452 16396 1458 16408
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 7926 16436 7932 16448
rect 6696 16408 7932 16436
rect 6696 16396 6702 16408
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 11514 16396 11520 16448
rect 11572 16436 11578 16448
rect 12342 16436 12348 16448
rect 11572 16408 12348 16436
rect 11572 16396 11578 16408
rect 12342 16396 12348 16408
rect 12400 16436 12406 16448
rect 14016 16436 14044 16476
rect 17770 16464 17776 16516
rect 17828 16504 17834 16516
rect 17957 16507 18015 16513
rect 17957 16504 17969 16507
rect 17828 16476 17969 16504
rect 17828 16464 17834 16476
rect 17957 16473 17969 16476
rect 18003 16473 18015 16507
rect 17957 16467 18015 16473
rect 12400 16408 14044 16436
rect 14093 16439 14151 16445
rect 12400 16396 12406 16408
rect 14093 16405 14105 16439
rect 14139 16436 14151 16439
rect 14274 16436 14280 16448
rect 14139 16408 14280 16436
rect 14139 16405 14151 16408
rect 14093 16399 14151 16405
rect 14274 16396 14280 16408
rect 14332 16396 14338 16448
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 15841 16439 15899 16445
rect 15841 16405 15853 16439
rect 15887 16436 15899 16439
rect 17862 16436 17868 16448
rect 15887 16408 17868 16436
rect 15887 16405 15899 16408
rect 15841 16399 15899 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 22278 16436 22284 16448
rect 22239 16408 22284 16436
rect 22278 16396 22284 16408
rect 22336 16396 22342 16448
rect 1104 16346 22816 16368
rect 1104 16294 4614 16346
rect 4666 16294 4678 16346
rect 4730 16294 4742 16346
rect 4794 16294 4806 16346
rect 4858 16294 11878 16346
rect 11930 16294 11942 16346
rect 11994 16294 12006 16346
rect 12058 16294 12070 16346
rect 12122 16294 19142 16346
rect 19194 16294 19206 16346
rect 19258 16294 19270 16346
rect 19322 16294 19334 16346
rect 19386 16294 22816 16346
rect 1104 16272 22816 16294
rect 3142 16192 3148 16244
rect 3200 16232 3206 16244
rect 3237 16235 3295 16241
rect 3237 16232 3249 16235
rect 3200 16204 3249 16232
rect 3200 16192 3206 16204
rect 3237 16201 3249 16204
rect 3283 16201 3295 16235
rect 3237 16195 3295 16201
rect 5258 16192 5264 16244
rect 5316 16232 5322 16244
rect 5997 16235 6055 16241
rect 5997 16232 6009 16235
rect 5316 16204 6009 16232
rect 5316 16192 5322 16204
rect 5997 16201 6009 16204
rect 6043 16201 6055 16235
rect 5997 16195 6055 16201
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7653 16235 7711 16241
rect 7653 16232 7665 16235
rect 6788 16204 7665 16232
rect 6788 16192 6794 16204
rect 7653 16201 7665 16204
rect 7699 16201 7711 16235
rect 7834 16232 7840 16244
rect 7795 16204 7840 16232
rect 7653 16195 7711 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 10689 16235 10747 16241
rect 7984 16204 10364 16232
rect 7984 16192 7990 16204
rect 5718 16124 5724 16176
rect 5776 16164 5782 16176
rect 5776 16136 8248 16164
rect 5776 16124 5782 16136
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 3970 16056 3976 16108
rect 4028 16096 4034 16108
rect 4157 16099 4215 16105
rect 4157 16096 4169 16099
rect 4028 16068 4169 16096
rect 4028 16056 4034 16068
rect 4157 16065 4169 16068
rect 4203 16065 4215 16099
rect 6270 16096 6276 16108
rect 6231 16068 6276 16096
rect 4157 16059 4215 16065
rect 6270 16056 6276 16068
rect 6328 16056 6334 16108
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 6880 16068 7389 16096
rect 6880 16056 6886 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 1670 15988 1676 16040
rect 1728 16028 1734 16040
rect 1857 16031 1915 16037
rect 1857 16028 1869 16031
rect 1728 16000 1869 16028
rect 1728 15988 1734 16000
rect 1857 15997 1869 16000
rect 1903 15997 1915 16031
rect 1857 15991 1915 15997
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 3988 16028 4016 16056
rect 3660 16000 4016 16028
rect 3660 15988 3666 16000
rect 4430 15988 4436 16040
rect 4488 16028 4494 16040
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4488 16000 4629 16028
rect 4488 15988 4494 16000
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 5350 15988 5356 16040
rect 5408 16028 5414 16040
rect 8220 16037 8248 16136
rect 8481 16099 8539 16105
rect 8481 16065 8493 16099
rect 8527 16096 8539 16099
rect 8662 16096 8668 16108
rect 8527 16068 8668 16096
rect 8527 16065 8539 16068
rect 8481 16059 8539 16065
rect 8662 16056 8668 16068
rect 8720 16056 8726 16108
rect 10336 16096 10364 16204
rect 10689 16201 10701 16235
rect 10735 16232 10747 16235
rect 11054 16232 11060 16244
rect 10735 16204 11060 16232
rect 10735 16201 10747 16204
rect 10689 16195 10747 16201
rect 11054 16192 11060 16204
rect 11112 16232 11118 16244
rect 11698 16232 11704 16244
rect 11112 16204 11704 16232
rect 11112 16192 11118 16204
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12069 16235 12127 16241
rect 12069 16201 12081 16235
rect 12115 16232 12127 16235
rect 12434 16232 12440 16244
rect 12115 16204 12440 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 12434 16192 12440 16204
rect 12492 16192 12498 16244
rect 12544 16204 13768 16232
rect 10410 16124 10416 16176
rect 10468 16164 10474 16176
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 10468 16136 10977 16164
rect 10468 16124 10474 16136
rect 10965 16133 10977 16136
rect 11011 16133 11023 16167
rect 12544 16164 12572 16204
rect 10965 16127 11023 16133
rect 11072 16136 12572 16164
rect 13740 16164 13768 16204
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 13909 16235 13967 16241
rect 13909 16232 13921 16235
rect 13872 16204 13921 16232
rect 13872 16192 13878 16204
rect 13909 16201 13921 16204
rect 13955 16232 13967 16235
rect 14090 16232 14096 16244
rect 13955 16204 14096 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 14292 16204 16129 16232
rect 14292 16164 14320 16204
rect 16117 16201 16129 16204
rect 16163 16232 16175 16235
rect 16850 16232 16856 16244
rect 16163 16204 16856 16232
rect 16163 16201 16175 16204
rect 16117 16195 16175 16201
rect 16850 16192 16856 16204
rect 16908 16192 16914 16244
rect 16945 16235 17003 16241
rect 16945 16201 16957 16235
rect 16991 16232 17003 16235
rect 18230 16232 18236 16244
rect 16991 16204 18236 16232
rect 16991 16201 17003 16204
rect 16945 16195 17003 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19981 16235 20039 16241
rect 19981 16201 19993 16235
rect 20027 16232 20039 16235
rect 20438 16232 20444 16244
rect 20027 16204 20444 16232
rect 20027 16201 20039 16204
rect 19981 16195 20039 16201
rect 20438 16192 20444 16204
rect 20496 16192 20502 16244
rect 20990 16232 20996 16244
rect 20824 16204 20996 16232
rect 13740 16136 14320 16164
rect 11072 16096 11100 16136
rect 11606 16096 11612 16108
rect 10336 16068 11100 16096
rect 11567 16068 11612 16096
rect 11606 16056 11612 16068
rect 11664 16056 11670 16108
rect 14740 16099 14798 16105
rect 14740 16096 14752 16099
rect 14016 16068 14752 16096
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 5408 16000 7297 16028
rect 5408 15988 5414 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 8205 16031 8263 16037
rect 8205 15997 8217 16031
rect 8251 15997 8263 16031
rect 8205 15991 8263 15997
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9576 16031 9634 16037
rect 9576 15997 9588 16031
rect 9622 16028 9634 16031
rect 10778 16028 10784 16040
rect 9622 16000 10784 16028
rect 9622 15997 9634 16000
rect 9576 15991 9634 15997
rect 2124 15963 2182 15969
rect 2124 15929 2136 15963
rect 2170 15960 2182 15963
rect 3050 15960 3056 15972
rect 2170 15932 3056 15960
rect 2170 15929 2182 15932
rect 2124 15923 2182 15929
rect 3050 15920 3056 15932
rect 3108 15920 3114 15972
rect 3694 15920 3700 15972
rect 3752 15960 3758 15972
rect 3973 15963 4031 15969
rect 3973 15960 3985 15963
rect 3752 15932 3985 15960
rect 3752 15920 3758 15932
rect 3973 15929 3985 15932
rect 4019 15929 4031 15963
rect 3973 15923 4031 15929
rect 4884 15963 4942 15969
rect 4884 15929 4896 15963
rect 4930 15960 4942 15963
rect 6178 15960 6184 15972
rect 4930 15932 6184 15960
rect 4930 15929 4942 15932
rect 4884 15923 4942 15929
rect 6178 15920 6184 15932
rect 6236 15920 6242 15972
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 8297 15963 8355 15969
rect 8297 15960 8309 15963
rect 6972 15932 8309 15960
rect 6972 15920 6978 15932
rect 8297 15929 8309 15932
rect 8343 15929 8355 15963
rect 9324 15960 9352 15991
rect 10778 15988 10784 16000
rect 10836 15988 10842 16040
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 15997 12311 16031
rect 12253 15991 12311 15997
rect 9766 15960 9772 15972
rect 8297 15923 8355 15929
rect 8404 15932 8984 15960
rect 9324 15932 9772 15960
rect 3605 15895 3663 15901
rect 3605 15861 3617 15895
rect 3651 15892 3663 15895
rect 3878 15892 3884 15904
rect 3651 15864 3884 15892
rect 3651 15861 3663 15864
rect 3605 15855 3663 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4062 15892 4068 15904
rect 4023 15864 4068 15892
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4798 15852 4804 15904
rect 4856 15892 4862 15904
rect 5258 15892 5264 15904
rect 4856 15864 5264 15892
rect 4856 15852 4862 15864
rect 5258 15852 5264 15864
rect 5316 15852 5322 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6825 15895 6883 15901
rect 6825 15892 6837 15895
rect 6420 15864 6837 15892
rect 6420 15852 6426 15864
rect 6825 15861 6837 15864
rect 6871 15861 6883 15895
rect 7190 15892 7196 15904
rect 7151 15864 7196 15892
rect 6825 15855 6883 15861
rect 7190 15852 7196 15864
rect 7248 15852 7254 15904
rect 7653 15895 7711 15901
rect 7653 15861 7665 15895
rect 7699 15892 7711 15895
rect 8404 15892 8432 15932
rect 8846 15892 8852 15904
rect 7699 15864 8432 15892
rect 8807 15864 8852 15892
rect 7699 15861 7711 15864
rect 7653 15855 7711 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 8956 15892 8984 15932
rect 9766 15920 9772 15932
rect 9824 15920 9830 15972
rect 12268 15960 12296 15991
rect 12434 15988 12440 16040
rect 12492 16028 12498 16040
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 12492 16000 12541 16028
rect 12492 15988 12498 16000
rect 12529 15997 12541 16000
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 12796 16031 12854 16037
rect 12796 15997 12808 16031
rect 12842 16028 12854 16031
rect 13906 16028 13912 16040
rect 12842 16000 13912 16028
rect 12842 15997 12854 16000
rect 12796 15991 12854 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 13538 15960 13544 15972
rect 9876 15932 11652 15960
rect 12268 15932 13544 15960
rect 9876 15892 9904 15932
rect 11330 15892 11336 15904
rect 8956 15864 9904 15892
rect 11291 15864 11336 15892
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11425 15895 11483 15901
rect 11425 15861 11437 15895
rect 11471 15892 11483 15895
rect 11514 15892 11520 15904
rect 11471 15864 11520 15892
rect 11471 15861 11483 15864
rect 11425 15855 11483 15861
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 11624 15892 11652 15932
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 14016 15892 14044 16068
rect 14740 16065 14752 16068
rect 14786 16065 14798 16099
rect 16114 16096 16120 16108
rect 14740 16059 14798 16065
rect 14844 16068 16120 16096
rect 14277 16031 14335 16037
rect 14277 15997 14289 16031
rect 14323 16028 14335 16031
rect 14844 16028 14872 16068
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 20824 16105 20852 16204
rect 20990 16192 20996 16204
rect 21048 16192 21054 16244
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 16224 16068 17509 16096
rect 15010 16028 15016 16040
rect 14323 16000 14872 16028
rect 14971 16000 15016 16028
rect 14323 15997 14335 16000
rect 14277 15991 14335 15997
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 16224 16028 16252 16068
rect 17497 16065 17509 16068
rect 17543 16096 17555 16099
rect 20809 16099 20867 16105
rect 17543 16068 18736 16096
rect 17543 16065 17555 16068
rect 17497 16059 17555 16065
rect 16040 16000 16252 16028
rect 11624 15864 14044 15892
rect 14274 15852 14280 15904
rect 14332 15892 14338 15904
rect 14743 15895 14801 15901
rect 14743 15892 14755 15895
rect 14332 15864 14755 15892
rect 14332 15852 14338 15864
rect 14743 15861 14755 15864
rect 14789 15861 14801 15895
rect 14743 15855 14801 15861
rect 15010 15852 15016 15904
rect 15068 15892 15074 15904
rect 16040 15892 16068 16000
rect 16298 15988 16304 16040
rect 16356 16028 16362 16040
rect 16393 16031 16451 16037
rect 16393 16028 16405 16031
rect 16356 16000 16405 16028
rect 16356 15988 16362 16000
rect 16393 15997 16405 16000
rect 16439 15997 16451 16031
rect 16393 15991 16451 15997
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 15997 18107 16031
rect 18049 15991 18107 15997
rect 16114 15920 16120 15972
rect 16172 15960 16178 15972
rect 16482 15960 16488 15972
rect 16172 15932 16488 15960
rect 16172 15920 16178 15932
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 18064 15960 18092 15991
rect 18230 15988 18236 16040
rect 18288 16028 18294 16040
rect 18601 16031 18659 16037
rect 18601 16028 18613 16031
rect 18288 16000 18613 16028
rect 18288 15988 18294 16000
rect 18601 15997 18613 16000
rect 18647 15997 18659 16031
rect 18708 16028 18736 16068
rect 20809 16065 20821 16099
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20254 16028 20260 16040
rect 18708 16000 19564 16028
rect 20215 16000 20260 16028
rect 18601 15991 18659 15997
rect 18868 15963 18926 15969
rect 18064 15932 18828 15960
rect 16574 15892 16580 15904
rect 15068 15864 16068 15892
rect 16535 15864 16580 15892
rect 15068 15852 15074 15864
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 17310 15892 17316 15904
rect 17271 15864 17316 15892
rect 17310 15852 17316 15864
rect 17368 15852 17374 15904
rect 17405 15895 17463 15901
rect 17405 15861 17417 15895
rect 17451 15892 17463 15895
rect 18046 15892 18052 15904
rect 17451 15864 18052 15892
rect 17451 15861 17463 15864
rect 17405 15855 17463 15861
rect 18046 15852 18052 15864
rect 18104 15852 18110 15904
rect 18233 15895 18291 15901
rect 18233 15861 18245 15895
rect 18279 15892 18291 15895
rect 18506 15892 18512 15904
rect 18279 15864 18512 15892
rect 18279 15861 18291 15864
rect 18233 15855 18291 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18800 15892 18828 15932
rect 18868 15929 18880 15963
rect 18914 15960 18926 15963
rect 19426 15960 19432 15972
rect 18914 15932 19432 15960
rect 18914 15929 18926 15932
rect 18868 15923 18926 15929
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 19536 15960 19564 16000
rect 20254 15988 20260 16000
rect 20312 15988 20318 16040
rect 21076 16031 21134 16037
rect 21076 15997 21088 16031
rect 21122 16028 21134 16031
rect 22278 16028 22284 16040
rect 21122 16000 22284 16028
rect 21122 15997 21134 16000
rect 21076 15991 21134 15997
rect 22278 15988 22284 16000
rect 22336 15988 22342 16040
rect 21358 15960 21364 15972
rect 19536 15932 21364 15960
rect 19886 15892 19892 15904
rect 18800 15864 19892 15892
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 19978 15852 19984 15904
rect 20036 15892 20042 15904
rect 20254 15892 20260 15904
rect 20036 15864 20260 15892
rect 20036 15852 20042 15864
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 20456 15901 20484 15932
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 20441 15895 20499 15901
rect 20441 15861 20453 15895
rect 20487 15861 20499 15895
rect 20441 15855 20499 15861
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 22189 15895 22247 15901
rect 22189 15892 22201 15895
rect 21600 15864 22201 15892
rect 21600 15852 21606 15864
rect 22189 15861 22201 15864
rect 22235 15861 22247 15895
rect 22189 15855 22247 15861
rect 1104 15802 22816 15824
rect 1104 15750 8246 15802
rect 8298 15750 8310 15802
rect 8362 15750 8374 15802
rect 8426 15750 8438 15802
rect 8490 15750 15510 15802
rect 15562 15750 15574 15802
rect 15626 15750 15638 15802
rect 15690 15750 15702 15802
rect 15754 15750 22816 15802
rect 1104 15728 22816 15750
rect 3050 15688 3056 15700
rect 3011 15660 3056 15688
rect 3050 15648 3056 15660
rect 3108 15648 3114 15700
rect 4154 15648 4160 15700
rect 4212 15688 4218 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 4212 15660 4261 15688
rect 4212 15648 4218 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 6178 15688 6184 15700
rect 6139 15660 6184 15688
rect 4249 15651 4307 15657
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 6822 15688 6828 15700
rect 6783 15660 6828 15688
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7009 15691 7067 15697
rect 7009 15657 7021 15691
rect 7055 15688 7067 15691
rect 9217 15691 9275 15697
rect 9217 15688 9229 15691
rect 7055 15660 9229 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 9217 15657 9229 15660
rect 9263 15657 9275 15691
rect 10410 15688 10416 15700
rect 9217 15651 9275 15657
rect 9876 15660 10416 15688
rect 4080 15592 8432 15620
rect 1670 15552 1676 15564
rect 1631 15524 1676 15552
rect 1670 15512 1676 15524
rect 1728 15512 1734 15564
rect 1946 15561 1952 15564
rect 1940 15515 1952 15561
rect 2004 15552 2010 15564
rect 3421 15555 3479 15561
rect 2004 15524 2040 15552
rect 1946 15512 1952 15515
rect 2004 15512 2010 15524
rect 3421 15521 3433 15555
rect 3467 15552 3479 15555
rect 3510 15552 3516 15564
rect 3467 15524 3516 15552
rect 3467 15521 3479 15524
rect 3421 15515 3479 15521
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4080 15561 4108 15592
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15521 4123 15555
rect 4798 15552 4804 15564
rect 4759 15524 4804 15552
rect 4065 15515 4123 15521
rect 4798 15512 4804 15524
rect 4856 15512 4862 15564
rect 5068 15555 5126 15561
rect 5068 15521 5080 15555
rect 5114 15552 5126 15555
rect 6641 15555 6699 15561
rect 5114 15524 6592 15552
rect 5114 15521 5126 15524
rect 5068 15515 5126 15521
rect 3605 15351 3663 15357
rect 3605 15317 3617 15351
rect 3651 15348 3663 15351
rect 3970 15348 3976 15360
rect 3651 15320 3976 15348
rect 3651 15317 3663 15320
rect 3605 15311 3663 15317
rect 3970 15308 3976 15320
rect 4028 15308 4034 15360
rect 6564 15348 6592 15524
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 7009 15555 7067 15561
rect 7009 15552 7021 15555
rect 6687 15524 7021 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 7009 15521 7021 15524
rect 7055 15521 7067 15555
rect 7009 15515 7067 15521
rect 7460 15555 7518 15561
rect 7460 15521 7472 15555
rect 7506 15552 7518 15555
rect 8294 15552 8300 15564
rect 7506 15524 8300 15552
rect 7506 15521 7518 15524
rect 7460 15515 7518 15521
rect 8294 15512 8300 15524
rect 8352 15512 8358 15564
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7193 15487 7251 15493
rect 7193 15484 7205 15487
rect 7156 15456 7205 15484
rect 7156 15444 7162 15456
rect 7193 15453 7205 15456
rect 7239 15453 7251 15487
rect 8404 15484 8432 15592
rect 8478 15580 8484 15632
rect 8536 15620 8542 15632
rect 9033 15623 9091 15629
rect 9033 15620 9045 15623
rect 8536 15592 9045 15620
rect 8536 15580 8542 15592
rect 9033 15589 9045 15592
rect 9079 15589 9091 15623
rect 9876 15620 9904 15660
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 11146 15648 11152 15700
rect 11204 15688 11210 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11204 15660 11345 15688
rect 11204 15648 11210 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 13906 15688 13912 15700
rect 13867 15660 13912 15688
rect 11333 15651 11391 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 18322 15648 18328 15700
rect 18380 15688 18386 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 18380 15660 18521 15688
rect 18380 15648 18386 15660
rect 18509 15657 18521 15660
rect 18555 15688 18567 15691
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 18555 15660 19257 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 20901 15691 20959 15697
rect 20901 15688 20913 15691
rect 20772 15660 20913 15688
rect 20772 15648 20778 15660
rect 20901 15657 20913 15660
rect 20947 15657 20959 15691
rect 20901 15651 20959 15657
rect 21174 15648 21180 15700
rect 21232 15688 21238 15700
rect 21361 15691 21419 15697
rect 21361 15688 21373 15691
rect 21232 15660 21373 15688
rect 21232 15648 21238 15660
rect 21361 15657 21373 15660
rect 21407 15657 21419 15691
rect 21361 15651 21419 15657
rect 9033 15583 9091 15589
rect 9508 15592 9904 15620
rect 9944 15623 10002 15629
rect 8849 15555 8907 15561
rect 8849 15521 8861 15555
rect 8895 15552 8907 15555
rect 9508 15552 9536 15592
rect 9944 15589 9956 15623
rect 9990 15620 10002 15623
rect 11054 15620 11060 15632
rect 9990 15592 11060 15620
rect 9990 15589 10002 15592
rect 9944 15583 10002 15589
rect 11054 15580 11060 15592
rect 11112 15580 11118 15632
rect 12796 15623 12854 15629
rect 12796 15589 12808 15623
rect 12842 15620 12854 15623
rect 13998 15620 14004 15632
rect 12842 15592 14004 15620
rect 12842 15589 12854 15592
rect 12796 15583 12854 15589
rect 13998 15580 14004 15592
rect 14056 15580 14062 15632
rect 14553 15623 14611 15629
rect 14553 15589 14565 15623
rect 14599 15620 14611 15623
rect 16482 15620 16488 15632
rect 14599 15592 16488 15620
rect 14599 15589 14611 15592
rect 14553 15583 14611 15589
rect 16482 15580 16488 15592
rect 16540 15580 16546 15632
rect 21269 15623 21327 15629
rect 21269 15589 21281 15623
rect 21315 15620 21327 15623
rect 22278 15620 22284 15632
rect 21315 15592 22284 15620
rect 21315 15589 21327 15592
rect 21269 15583 21327 15589
rect 22278 15580 22284 15592
rect 22336 15580 22342 15632
rect 10226 15552 10232 15564
rect 8895 15524 9536 15552
rect 9600 15524 10232 15552
rect 8895 15521 8907 15524
rect 8849 15515 8907 15521
rect 9600 15484 9628 15524
rect 10226 15512 10232 15524
rect 10284 15512 10290 15564
rect 11698 15552 11704 15564
rect 11659 15524 11704 15552
rect 11698 15512 11704 15524
rect 11756 15512 11762 15564
rect 13906 15512 13912 15564
rect 13964 15552 13970 15564
rect 14366 15552 14372 15564
rect 13964 15524 14372 15552
rect 13964 15512 13970 15524
rect 14366 15512 14372 15524
rect 14424 15512 14430 15564
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 15194 15552 15200 15564
rect 14691 15524 15200 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 15194 15512 15200 15524
rect 15252 15512 15258 15564
rect 15562 15561 15568 15564
rect 15556 15552 15568 15561
rect 15523 15524 15568 15552
rect 15556 15515 15568 15524
rect 15562 15512 15568 15515
rect 15620 15512 15626 15564
rect 17129 15555 17187 15561
rect 17129 15521 17141 15555
rect 17175 15552 17187 15555
rect 17218 15552 17224 15564
rect 17175 15524 17224 15552
rect 17175 15521 17187 15524
rect 17129 15515 17187 15521
rect 17218 15512 17224 15524
rect 17276 15512 17282 15564
rect 17396 15555 17454 15561
rect 17396 15521 17408 15555
rect 17442 15552 17454 15555
rect 17678 15552 17684 15564
rect 17442 15524 17684 15552
rect 17442 15521 17454 15524
rect 17396 15515 17454 15521
rect 17678 15512 17684 15524
rect 17736 15512 17742 15564
rect 19153 15555 19211 15561
rect 19153 15521 19165 15555
rect 19199 15552 19211 15555
rect 19426 15552 19432 15564
rect 19199 15524 19432 15552
rect 19199 15521 19211 15524
rect 19153 15515 19211 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15552 20223 15555
rect 21358 15552 21364 15564
rect 20211 15524 21364 15552
rect 20211 15521 20223 15524
rect 20165 15515 20223 15521
rect 21358 15512 21364 15524
rect 21416 15512 21422 15564
rect 21910 15552 21916 15564
rect 21871 15524 21916 15552
rect 21910 15512 21916 15524
rect 21968 15512 21974 15564
rect 8404 15456 9628 15484
rect 9677 15487 9735 15493
rect 7193 15447 7251 15453
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 9677 15447 9735 15453
rect 11072 15456 11805 15484
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 6564 15320 8585 15348
rect 8573 15317 8585 15320
rect 8619 15348 8631 15351
rect 8662 15348 8668 15360
rect 8619 15320 8668 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 9692 15348 9720 15447
rect 9858 15348 9864 15360
rect 9692 15320 9864 15348
rect 9858 15308 9864 15320
rect 9916 15308 9922 15360
rect 10778 15308 10784 15360
rect 10836 15348 10842 15360
rect 11072 15357 11100 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 11606 15376 11612 15428
rect 11664 15416 11670 15428
rect 11900 15416 11928 15447
rect 12434 15444 12440 15496
rect 12492 15484 12498 15496
rect 12529 15487 12587 15493
rect 12529 15484 12541 15487
rect 12492 15456 12541 15484
rect 12492 15444 12498 15456
rect 12529 15453 12541 15456
rect 12575 15453 12587 15487
rect 12529 15447 12587 15453
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15453 14887 15487
rect 14829 15447 14887 15453
rect 11664 15388 11928 15416
rect 14844 15416 14872 15447
rect 14918 15444 14924 15496
rect 14976 15484 14982 15496
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 14976 15456 15301 15484
rect 14976 15444 14982 15456
rect 15289 15453 15301 15456
rect 15335 15453 15347 15487
rect 15289 15447 15347 15453
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 18966 15484 18972 15496
rect 18564 15456 18972 15484
rect 18564 15444 18570 15456
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 19024 15456 19349 15484
rect 19024 15444 19030 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 15010 15416 15016 15428
rect 14844 15388 15016 15416
rect 11664 15376 11670 15388
rect 15010 15376 15016 15388
rect 15068 15376 15074 15428
rect 16942 15416 16948 15428
rect 16595 15388 16948 15416
rect 11057 15351 11115 15357
rect 11057 15348 11069 15351
rect 10836 15320 11069 15348
rect 10836 15308 10842 15320
rect 11057 15317 11069 15320
rect 11103 15317 11115 15351
rect 11057 15311 11115 15317
rect 14185 15351 14243 15357
rect 14185 15317 14197 15351
rect 14231 15348 14243 15351
rect 16595 15348 16623 15388
rect 16942 15376 16948 15388
rect 17000 15376 17006 15428
rect 19352 15416 19380 15447
rect 19978 15444 19984 15496
rect 20036 15484 20042 15496
rect 20257 15487 20315 15493
rect 20257 15484 20269 15487
rect 20036 15456 20269 15484
rect 20036 15444 20042 15456
rect 20257 15453 20269 15456
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15484 20407 15487
rect 20990 15484 20996 15496
rect 20395 15456 20996 15484
rect 20395 15453 20407 15456
rect 20349 15447 20407 15453
rect 20990 15444 20996 15456
rect 21048 15444 21054 15496
rect 21174 15444 21180 15496
rect 21232 15484 21238 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 21232 15456 21465 15484
rect 21232 15444 21238 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 19352 15388 20392 15416
rect 14231 15320 16623 15348
rect 16669 15351 16727 15357
rect 14231 15317 14243 15320
rect 14185 15311 14243 15317
rect 16669 15317 16681 15351
rect 16715 15348 16727 15351
rect 16850 15348 16856 15360
rect 16715 15320 16856 15348
rect 16715 15317 16727 15320
rect 16669 15311 16727 15317
rect 16850 15308 16856 15320
rect 16908 15308 16914 15360
rect 17310 15308 17316 15360
rect 17368 15348 17374 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 17368 15320 18797 15348
rect 17368 15308 17374 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 19794 15348 19800 15360
rect 19755 15320 19800 15348
rect 18785 15311 18843 15317
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 20364 15348 20392 15388
rect 20714 15376 20720 15428
rect 20772 15416 20778 15428
rect 22097 15419 22155 15425
rect 22097 15416 22109 15419
rect 20772 15388 22109 15416
rect 20772 15376 20778 15388
rect 22097 15385 22109 15388
rect 22143 15385 22155 15419
rect 22097 15379 22155 15385
rect 20806 15348 20812 15360
rect 20364 15320 20812 15348
rect 20806 15308 20812 15320
rect 20864 15348 20870 15360
rect 21174 15348 21180 15360
rect 20864 15320 21180 15348
rect 20864 15308 20870 15320
rect 21174 15308 21180 15320
rect 21232 15308 21238 15360
rect 1104 15258 22816 15280
rect 1104 15206 4614 15258
rect 4666 15206 4678 15258
rect 4730 15206 4742 15258
rect 4794 15206 4806 15258
rect 4858 15206 11878 15258
rect 11930 15206 11942 15258
rect 11994 15206 12006 15258
rect 12058 15206 12070 15258
rect 12122 15206 19142 15258
rect 19194 15206 19206 15258
rect 19258 15206 19270 15258
rect 19322 15206 19334 15258
rect 19386 15206 22816 15258
rect 1104 15184 22816 15206
rect 3694 15104 3700 15156
rect 3752 15144 3758 15156
rect 4982 15144 4988 15156
rect 3752 15116 4988 15144
rect 3752 15104 3758 15116
rect 4982 15104 4988 15116
rect 5040 15144 5046 15156
rect 5721 15147 5779 15153
rect 5721 15144 5733 15147
rect 5040 15116 5733 15144
rect 5040 15104 5046 15116
rect 5721 15113 5733 15116
rect 5767 15113 5779 15147
rect 5721 15107 5779 15113
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 6914 15144 6920 15156
rect 6411 15116 6920 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 6914 15104 6920 15116
rect 6972 15104 6978 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 8352 15116 8493 15144
rect 8352 15104 8358 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 11054 15144 11060 15156
rect 10735 15116 11060 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 11054 15104 11060 15116
rect 11112 15144 11118 15156
rect 11698 15144 11704 15156
rect 11112 15116 11704 15144
rect 11112 15104 11118 15116
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15144 12035 15147
rect 12342 15144 12348 15156
rect 12023 15116 12348 15144
rect 12023 15113 12035 15116
rect 11977 15107 12035 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13817 15147 13875 15153
rect 13817 15113 13829 15147
rect 13863 15144 13875 15147
rect 13998 15144 14004 15156
rect 13863 15116 14004 15144
rect 13863 15113 13875 15116
rect 13817 15107 13875 15113
rect 13998 15104 14004 15116
rect 14056 15104 14062 15156
rect 14182 15144 14188 15156
rect 14143 15116 14188 15144
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 15562 15144 15568 15156
rect 15436 15116 15568 15144
rect 15436 15104 15442 15116
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 15930 15104 15936 15156
rect 15988 15144 15994 15156
rect 17678 15144 17684 15156
rect 15988 15116 17264 15144
rect 17639 15116 17684 15144
rect 15988 15104 15994 15116
rect 3329 15079 3387 15085
rect 3329 15045 3341 15079
rect 3375 15076 3387 15079
rect 3786 15076 3792 15088
rect 3375 15048 3792 15076
rect 3375 15045 3387 15048
rect 3329 15039 3387 15045
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 17236 15076 17264 15116
rect 17678 15104 17684 15116
rect 17736 15104 17742 15156
rect 18230 15144 18236 15156
rect 18064 15116 18236 15144
rect 17954 15076 17960 15088
rect 17236 15048 17960 15076
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 3881 15011 3939 15017
rect 3881 15008 3893 15011
rect 3660 14980 3893 15008
rect 3660 14968 3666 14980
rect 3881 14977 3893 14980
rect 3927 14977 3939 15011
rect 7098 15008 7104 15020
rect 7059 14980 7104 15008
rect 3881 14971 3939 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 8680 14980 9321 15008
rect 1489 14943 1547 14949
rect 1489 14909 1501 14943
rect 1535 14940 1547 14943
rect 1578 14940 1584 14952
rect 1535 14912 1584 14940
rect 1535 14909 1547 14912
rect 1489 14903 1547 14909
rect 1578 14900 1584 14912
rect 1636 14900 1642 14952
rect 4154 14900 4160 14952
rect 4212 14940 4218 14952
rect 4341 14943 4399 14949
rect 4341 14940 4353 14943
rect 4212 14912 4353 14940
rect 4212 14900 4218 14912
rect 4341 14909 4353 14912
rect 4387 14940 4399 14943
rect 4430 14940 4436 14952
rect 4387 14912 4436 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 4430 14900 4436 14912
rect 4488 14900 4494 14952
rect 6181 14943 6239 14949
rect 6181 14909 6193 14943
rect 6227 14940 6239 14943
rect 6362 14940 6368 14952
rect 6227 14912 6368 14940
rect 6227 14909 6239 14912
rect 6181 14903 6239 14909
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 7116 14940 7144 14968
rect 8680 14940 8708 14980
rect 9309 14977 9321 14980
rect 9355 14977 9367 15011
rect 9309 14971 9367 14977
rect 7116 14912 8708 14940
rect 8757 14943 8815 14949
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 9324 14940 9352 14971
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 11517 15011 11575 15017
rect 11517 15008 11529 15011
rect 10376 14980 11529 15008
rect 10376 14968 10382 14980
rect 11517 14977 11529 14980
rect 11563 14977 11575 15011
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 11517 14971 11575 14977
rect 13832 14980 14473 15008
rect 9576 14943 9634 14949
rect 9324 14912 9536 14940
rect 8757 14903 8815 14909
rect 1756 14875 1814 14881
rect 1756 14841 1768 14875
rect 1802 14872 1814 14875
rect 2038 14872 2044 14884
rect 1802 14844 2044 14872
rect 1802 14841 1814 14844
rect 1756 14835 1814 14841
rect 2038 14832 2044 14844
rect 2096 14832 2102 14884
rect 4062 14832 4068 14884
rect 4120 14872 4126 14884
rect 4586 14875 4644 14881
rect 4586 14872 4598 14875
rect 4120 14844 4598 14872
rect 4120 14832 4126 14844
rect 4586 14841 4598 14844
rect 4632 14841 4644 14875
rect 4586 14835 4644 14841
rect 6822 14832 6828 14884
rect 6880 14872 6886 14884
rect 7346 14875 7404 14881
rect 7346 14872 7358 14875
rect 6880 14844 7358 14872
rect 6880 14832 6886 14844
rect 7346 14841 7358 14844
rect 7392 14841 7404 14875
rect 8772 14872 8800 14903
rect 9398 14872 9404 14884
rect 8772 14844 9404 14872
rect 7346 14835 7404 14841
rect 9398 14832 9404 14844
rect 9456 14832 9462 14884
rect 9508 14872 9536 14912
rect 9576 14909 9588 14943
rect 9622 14940 9634 14943
rect 10778 14940 10784 14952
rect 9622 14912 10784 14940
rect 9622 14909 9634 14912
rect 9576 14903 9634 14909
rect 10778 14900 10784 14912
rect 10836 14900 10842 14952
rect 11698 14900 11704 14952
rect 11756 14940 11762 14952
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11756 14912 12173 14940
rect 11756 14900 11762 14912
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 12710 14949 12716 14952
rect 12704 14940 12716 14949
rect 12492 14912 12537 14940
rect 12671 14912 12716 14940
rect 12492 14900 12498 14912
rect 12704 14903 12716 14912
rect 12710 14900 12716 14903
rect 12768 14900 12774 14952
rect 9766 14872 9772 14884
rect 9508 14844 9772 14872
rect 9766 14832 9772 14844
rect 9824 14832 9830 14884
rect 11333 14875 11391 14881
rect 11333 14841 11345 14875
rect 11379 14872 11391 14875
rect 12452 14872 12480 14900
rect 13832 14872 13860 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 15746 14968 15752 15020
rect 15804 15008 15810 15020
rect 16301 15011 16359 15017
rect 16301 15008 16313 15011
rect 15804 14980 16313 15008
rect 15804 14968 15810 14980
rect 16301 14977 16313 14980
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 17310 14968 17316 15020
rect 17368 15008 17374 15020
rect 18064 15017 18092 15116
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 19426 15144 19432 15156
rect 19387 15116 19432 15144
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19702 15104 19708 15156
rect 19760 15144 19766 15156
rect 20714 15144 20720 15156
rect 19760 15116 20720 15144
rect 19760 15104 19766 15116
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 17368 14980 18061 15008
rect 17368 14968 17374 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 20346 15008 20352 15020
rect 20307 14980 20352 15008
rect 18049 14971 18107 14977
rect 20346 14968 20352 14980
rect 20404 14968 20410 15020
rect 20548 15017 20576 15116
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 22281 15147 22339 15153
rect 22281 15144 22293 15147
rect 21140 15116 22293 15144
rect 21140 15104 21146 15116
rect 22281 15113 22293 15116
rect 22327 15113 22339 15147
rect 22281 15107 22339 15113
rect 20533 15011 20591 15017
rect 20533 14977 20545 15011
rect 20579 14977 20591 15011
rect 20533 14971 20591 14977
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14940 14427 14943
rect 15010 14940 15016 14952
rect 14415 14912 15016 14940
rect 14415 14909 14427 14912
rect 14369 14903 14427 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 17126 14940 17132 14952
rect 15764 14912 17132 14940
rect 11379 14844 12204 14872
rect 12452 14844 13860 14872
rect 11379 14841 11391 14844
rect 11333 14835 11391 14841
rect 12176 14816 12204 14844
rect 14182 14832 14188 14884
rect 14240 14872 14246 14884
rect 14728 14875 14786 14881
rect 14728 14872 14740 14875
rect 14240 14844 14740 14872
rect 14240 14832 14246 14844
rect 14728 14841 14740 14844
rect 14774 14872 14786 14875
rect 15764 14872 15792 14912
rect 17126 14900 17132 14912
rect 17184 14900 17190 14952
rect 17402 14900 17408 14952
rect 17460 14940 17466 14952
rect 18322 14949 18328 14952
rect 18316 14940 18328 14949
rect 17460 14912 18000 14940
rect 18283 14912 18328 14940
rect 17460 14900 17466 14912
rect 14774 14844 15792 14872
rect 16568 14875 16626 14881
rect 14774 14841 14786 14844
rect 14728 14835 14786 14841
rect 16568 14841 16580 14875
rect 16614 14872 16626 14875
rect 17310 14872 17316 14884
rect 16614 14844 17316 14872
rect 16614 14841 16626 14844
rect 16568 14835 16626 14841
rect 17310 14832 17316 14844
rect 17368 14832 17374 14884
rect 17972 14872 18000 14912
rect 18316 14903 18328 14912
rect 18322 14900 18328 14903
rect 18380 14900 18386 14952
rect 18874 14900 18880 14952
rect 18932 14940 18938 14952
rect 20257 14943 20315 14949
rect 20257 14940 20269 14943
rect 18932 14912 20269 14940
rect 18932 14900 18938 14912
rect 20257 14909 20269 14912
rect 20303 14909 20315 14943
rect 20257 14903 20315 14909
rect 20714 14900 20720 14952
rect 20772 14940 20778 14952
rect 20901 14943 20959 14949
rect 20901 14940 20913 14943
rect 20772 14912 20913 14940
rect 20772 14900 20778 14912
rect 20901 14909 20913 14912
rect 20947 14909 20959 14943
rect 20901 14903 20959 14909
rect 21168 14943 21226 14949
rect 21168 14909 21180 14943
rect 21214 14940 21226 14943
rect 21542 14940 21548 14952
rect 21214 14912 21548 14940
rect 21214 14909 21226 14912
rect 21168 14903 21226 14909
rect 21542 14900 21548 14912
rect 21600 14900 21606 14952
rect 17972 14844 19932 14872
rect 19904 14816 19932 14844
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2869 14807 2927 14813
rect 2869 14804 2881 14807
rect 2004 14776 2881 14804
rect 2004 14764 2010 14776
rect 2869 14773 2881 14776
rect 2915 14773 2927 14807
rect 3694 14804 3700 14816
rect 3655 14776 3700 14804
rect 2869 14767 2927 14773
rect 3694 14764 3700 14776
rect 3752 14764 3758 14816
rect 3789 14807 3847 14813
rect 3789 14773 3801 14807
rect 3835 14804 3847 14807
rect 4246 14804 4252 14816
rect 3835 14776 4252 14804
rect 3835 14773 3847 14776
rect 3789 14767 3847 14773
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 7466 14804 7472 14816
rect 4396 14776 7472 14804
rect 4396 14764 4402 14776
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 8941 14807 8999 14813
rect 8941 14804 8953 14807
rect 8168 14776 8953 14804
rect 8168 14764 8174 14776
rect 8941 14773 8953 14776
rect 8987 14773 8999 14807
rect 8941 14767 8999 14773
rect 10965 14807 11023 14813
rect 10965 14773 10977 14807
rect 11011 14804 11023 14807
rect 11146 14804 11152 14816
rect 11011 14776 11152 14804
rect 11011 14773 11023 14776
rect 10965 14767 11023 14773
rect 11146 14764 11152 14776
rect 11204 14764 11210 14816
rect 11425 14807 11483 14813
rect 11425 14773 11437 14807
rect 11471 14804 11483 14807
rect 11606 14804 11612 14816
rect 11471 14776 11612 14804
rect 11471 14773 11483 14776
rect 11425 14767 11483 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 12158 14764 12164 14816
rect 12216 14764 12222 14816
rect 15378 14764 15384 14816
rect 15436 14804 15442 14816
rect 15841 14807 15899 14813
rect 15841 14804 15853 14807
rect 15436 14776 15853 14804
rect 15436 14764 15442 14776
rect 15841 14773 15853 14776
rect 15887 14773 15899 14807
rect 15841 14767 15899 14773
rect 16482 14764 16488 14816
rect 16540 14804 16546 14816
rect 19058 14804 19064 14816
rect 16540 14776 19064 14804
rect 16540 14764 16546 14776
rect 19058 14764 19064 14776
rect 19116 14764 19122 14816
rect 19886 14804 19892 14816
rect 19799 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 1104 14714 22816 14736
rect 1104 14662 8246 14714
rect 8298 14662 8310 14714
rect 8362 14662 8374 14714
rect 8426 14662 8438 14714
rect 8490 14662 15510 14714
rect 15562 14662 15574 14714
rect 15626 14662 15638 14714
rect 15690 14662 15702 14714
rect 15754 14662 22816 14714
rect 1104 14640 22816 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2682 14560 2688 14612
rect 2740 14600 2746 14612
rect 3234 14600 3240 14612
rect 2740 14572 3240 14600
rect 2740 14560 2746 14572
rect 3234 14560 3240 14572
rect 3292 14600 3298 14612
rect 3602 14600 3608 14612
rect 3292 14572 3608 14600
rect 3292 14560 3298 14572
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 4062 14560 4068 14612
rect 4120 14600 4126 14612
rect 5445 14603 5503 14609
rect 5445 14600 5457 14603
rect 4120 14572 5457 14600
rect 4120 14560 4126 14572
rect 5445 14569 5457 14572
rect 5491 14569 5503 14603
rect 5813 14603 5871 14609
rect 5813 14600 5825 14603
rect 5445 14563 5503 14569
rect 5552 14572 5825 14600
rect 3694 14492 3700 14544
rect 3752 14532 3758 14544
rect 4310 14535 4368 14541
rect 4310 14532 4322 14535
rect 3752 14504 4322 14532
rect 3752 14492 3758 14504
rect 4310 14501 4322 14504
rect 4356 14532 4368 14535
rect 4430 14532 4436 14544
rect 4356 14504 4436 14532
rect 4356 14501 4368 14504
rect 4310 14495 4368 14501
rect 4430 14492 4436 14504
rect 4488 14492 4494 14544
rect 2958 14464 2964 14476
rect 2919 14436 2964 14464
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 3881 14467 3939 14473
rect 3881 14433 3893 14467
rect 3927 14464 3939 14467
rect 5552 14464 5580 14572
rect 5813 14569 5825 14572
rect 5859 14600 5871 14603
rect 6086 14600 6092 14612
rect 5859 14572 6092 14600
rect 5859 14569 5871 14572
rect 5813 14563 5871 14569
rect 6086 14560 6092 14572
rect 6144 14560 6150 14612
rect 6641 14603 6699 14609
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 7190 14600 7196 14612
rect 6687 14572 7196 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7524 14572 8125 14600
rect 7524 14560 7530 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 12618 14560 12624 14612
rect 12676 14600 12682 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12676 14572 12725 14600
rect 12676 14560 12682 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 9944 14535 10002 14541
rect 9944 14501 9956 14535
rect 9990 14532 10002 14535
rect 11054 14532 11060 14544
rect 9990 14504 11060 14532
rect 9990 14501 10002 14504
rect 9944 14495 10002 14501
rect 11054 14492 11060 14504
rect 11112 14492 11118 14544
rect 11330 14492 11336 14544
rect 11388 14532 11394 14544
rect 11578 14535 11636 14541
rect 11578 14532 11590 14535
rect 11388 14504 11590 14532
rect 11388 14492 11394 14504
rect 11578 14501 11590 14504
rect 11624 14501 11636 14535
rect 12728 14532 12756 14563
rect 12802 14560 12808 14612
rect 12860 14600 12866 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 12860 14572 14381 14600
rect 12860 14560 12866 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14369 14563 14427 14569
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 17402 14600 17408 14612
rect 15795 14572 17408 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 17773 14603 17831 14609
rect 17773 14600 17785 14603
rect 17604 14572 17785 14600
rect 13234 14535 13292 14541
rect 13234 14532 13246 14535
rect 12728 14504 13246 14532
rect 11578 14495 11636 14501
rect 13234 14501 13246 14504
rect 13280 14501 13292 14535
rect 13234 14495 13292 14501
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 15102 14532 15108 14544
rect 14056 14504 15108 14532
rect 14056 14492 14062 14504
rect 15102 14492 15108 14504
rect 15160 14492 15166 14544
rect 17310 14492 17316 14544
rect 17368 14532 17374 14544
rect 17604 14532 17632 14572
rect 17773 14569 17785 14572
rect 17819 14600 17831 14603
rect 17865 14603 17923 14609
rect 17865 14600 17877 14603
rect 17819 14572 17877 14600
rect 17819 14569 17831 14572
rect 17773 14563 17831 14569
rect 17865 14569 17877 14572
rect 17911 14569 17923 14603
rect 18046 14600 18052 14612
rect 18007 14572 18052 14600
rect 17865 14563 17923 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 18138 14560 18144 14612
rect 18196 14600 18202 14612
rect 18506 14600 18512 14612
rect 18196 14572 18512 14600
rect 18196 14560 18202 14572
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 19058 14600 19064 14612
rect 19019 14572 19064 14600
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 20806 14560 20812 14612
rect 20864 14600 20870 14612
rect 21450 14600 21456 14612
rect 20864 14572 21456 14600
rect 20864 14560 20870 14572
rect 21450 14560 21456 14572
rect 21508 14600 21514 14612
rect 22281 14603 22339 14609
rect 22281 14600 22293 14603
rect 21508 14572 22293 14600
rect 21508 14560 21514 14572
rect 22281 14569 22293 14572
rect 22327 14569 22339 14603
rect 22281 14563 22339 14569
rect 17368 14504 17632 14532
rect 17368 14492 17374 14504
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 18417 14535 18475 14541
rect 18417 14532 18429 14535
rect 17736 14504 18429 14532
rect 17736 14492 17742 14504
rect 18417 14501 18429 14504
rect 18463 14501 18475 14535
rect 18417 14495 18475 14501
rect 18966 14492 18972 14544
rect 19024 14532 19030 14544
rect 19024 14504 19656 14532
rect 19024 14492 19030 14504
rect 3927 14436 5580 14464
rect 5997 14467 6055 14473
rect 3927 14433 3939 14436
rect 3881 14427 3939 14433
rect 5997 14433 6009 14467
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 2038 14396 2044 14408
rect 1951 14368 2044 14396
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2682 14396 2688 14408
rect 2271 14368 2688 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3050 14396 3056 14408
rect 3011 14368 3056 14396
rect 3050 14356 3056 14368
rect 3108 14356 3114 14408
rect 3234 14396 3240 14408
rect 3195 14368 3240 14396
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3694 14356 3700 14408
rect 3752 14396 3758 14408
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3752 14368 4077 14396
rect 3752 14356 3758 14368
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 2056 14328 2084 14356
rect 6012 14328 6040 14427
rect 6086 14424 6092 14476
rect 6144 14464 6150 14476
rect 7009 14467 7067 14473
rect 6144 14436 6189 14464
rect 6144 14424 6150 14436
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7466 14464 7472 14476
rect 7055 14436 7472 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 7466 14424 7472 14436
rect 7524 14424 7530 14476
rect 8018 14464 8024 14476
rect 7979 14436 8024 14464
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8665 14467 8723 14473
rect 8665 14433 8677 14467
rect 8711 14464 8723 14467
rect 8754 14464 8760 14476
rect 8711 14436 8760 14464
rect 8711 14433 8723 14436
rect 8665 14427 8723 14433
rect 8754 14424 8760 14436
rect 8812 14424 8818 14476
rect 9398 14464 9404 14476
rect 9359 14436 9404 14464
rect 9398 14424 9404 14436
rect 9456 14424 9462 14476
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 9766 14464 9772 14476
rect 9723 14436 9772 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 9766 14424 9772 14436
rect 9824 14464 9830 14476
rect 14642 14464 14648 14476
rect 9824 14436 11376 14464
rect 14603 14436 14648 14464
rect 9824 14424 9830 14436
rect 7098 14396 7104 14408
rect 7059 14368 7104 14396
rect 7098 14356 7104 14368
rect 7156 14356 7162 14408
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14396 7346 14408
rect 7558 14396 7564 14408
rect 7340 14368 7564 14396
rect 7340 14356 7346 14368
rect 7558 14356 7564 14368
rect 7616 14356 7622 14408
rect 8202 14356 8208 14408
rect 8260 14396 8266 14408
rect 11348 14405 11376 14436
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 15841 14467 15899 14473
rect 15841 14433 15853 14467
rect 15887 14464 15899 14467
rect 15930 14464 15936 14476
rect 15887 14436 15936 14464
rect 15887 14433 15899 14436
rect 15841 14427 15899 14433
rect 15930 14424 15936 14436
rect 15988 14424 15994 14476
rect 16393 14467 16451 14473
rect 16393 14433 16405 14467
rect 16439 14464 16451 14467
rect 16482 14464 16488 14476
rect 16439 14436 16488 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 16660 14467 16718 14473
rect 16660 14433 16672 14467
rect 16706 14464 16718 14467
rect 17865 14467 17923 14473
rect 16706 14436 17816 14464
rect 16706 14433 16718 14436
rect 16660 14427 16718 14433
rect 11333 14399 11391 14405
rect 8260 14368 8305 14396
rect 8260 14356 8266 14368
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 12434 14356 12440 14408
rect 12492 14396 12498 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12492 14368 13001 14396
rect 12492 14356 12498 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 16025 14399 16083 14405
rect 16025 14365 16037 14399
rect 16071 14396 16083 14399
rect 17788 14396 17816 14436
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 18509 14467 18567 14473
rect 18509 14464 18521 14467
rect 17911 14436 18521 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18509 14433 18521 14436
rect 18555 14433 18567 14467
rect 19426 14464 19432 14476
rect 18509 14427 18567 14433
rect 18616 14436 19432 14464
rect 18616 14396 18644 14436
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 16071 14368 16436 14396
rect 17788 14368 18644 14396
rect 18693 14399 18751 14405
rect 16071 14365 16083 14368
rect 16025 14359 16083 14365
rect 9214 14328 9220 14340
rect 2056 14300 4108 14328
rect 6012 14300 9220 14328
rect 1581 14263 1639 14269
rect 1581 14229 1593 14263
rect 1627 14260 1639 14263
rect 2314 14260 2320 14272
rect 1627 14232 2320 14260
rect 1627 14229 1639 14232
rect 1581 14223 1639 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 2593 14263 2651 14269
rect 2593 14229 2605 14263
rect 2639 14260 2651 14263
rect 3418 14260 3424 14272
rect 2639 14232 3424 14260
rect 2639 14229 2651 14232
rect 2593 14223 2651 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 3694 14260 3700 14272
rect 3655 14232 3700 14260
rect 3694 14220 3700 14232
rect 3752 14220 3758 14272
rect 4080 14260 4108 14300
rect 9214 14288 9220 14300
rect 9272 14288 9278 14340
rect 5074 14260 5080 14272
rect 4080 14232 5080 14260
rect 5074 14220 5080 14232
rect 5132 14220 5138 14272
rect 6270 14260 6276 14272
rect 6231 14232 6276 14260
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7653 14263 7711 14269
rect 7653 14260 7665 14263
rect 7340 14232 7665 14260
rect 7340 14220 7346 14232
rect 7653 14229 7665 14232
rect 7699 14229 7711 14263
rect 7653 14223 7711 14229
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 8849 14263 8907 14269
rect 8849 14260 8861 14263
rect 7800 14232 8861 14260
rect 7800 14220 7806 14232
rect 8849 14229 8861 14232
rect 8895 14229 8907 14263
rect 11054 14260 11060 14272
rect 10967 14232 11060 14260
rect 8849 14223 8907 14229
rect 11054 14220 11060 14232
rect 11112 14260 11118 14272
rect 11514 14260 11520 14272
rect 11112 14232 11520 14260
rect 11112 14220 11118 14232
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 13004 14260 13032 14359
rect 14829 14331 14887 14337
rect 14829 14297 14841 14331
rect 14875 14328 14887 14331
rect 15930 14328 15936 14340
rect 14875 14300 15936 14328
rect 14875 14297 14887 14300
rect 14829 14291 14887 14297
rect 15930 14288 15936 14300
rect 15988 14288 15994 14340
rect 13170 14260 13176 14272
rect 13004 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 15381 14263 15439 14269
rect 15381 14229 15393 14263
rect 15427 14260 15439 14263
rect 16114 14260 16120 14272
rect 15427 14232 16120 14260
rect 15427 14229 15439 14232
rect 15381 14223 15439 14229
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 16408 14260 16436 14368
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 18966 14396 18972 14408
rect 18739 14368 18972 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 19518 14396 19524 14408
rect 19479 14368 19524 14396
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 19628 14405 19656 14504
rect 20346 14492 20352 14544
rect 20404 14532 20410 14544
rect 20530 14532 20536 14544
rect 20404 14504 20536 14532
rect 20404 14492 20410 14504
rect 20530 14492 20536 14504
rect 20588 14492 20594 14544
rect 21082 14492 21088 14544
rect 21140 14541 21146 14544
rect 21140 14535 21204 14541
rect 21140 14501 21158 14535
rect 21192 14501 21204 14535
rect 21140 14495 21204 14501
rect 21140 14492 21146 14495
rect 20254 14464 20260 14476
rect 20215 14436 20260 14464
rect 20254 14424 20260 14436
rect 20312 14424 20318 14476
rect 20714 14424 20720 14476
rect 20772 14464 20778 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20772 14436 20913 14464
rect 20772 14424 20778 14436
rect 20901 14433 20913 14436
rect 20947 14433 20959 14467
rect 20901 14427 20959 14433
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 20441 14331 20499 14337
rect 20441 14328 20453 14331
rect 17328 14300 20453 14328
rect 17328 14260 17356 14300
rect 20441 14297 20453 14300
rect 20487 14297 20499 14331
rect 20441 14291 20499 14297
rect 16408 14232 17356 14260
rect 17954 14220 17960 14272
rect 18012 14260 18018 14272
rect 19702 14260 19708 14272
rect 18012 14232 19708 14260
rect 18012 14220 18018 14232
rect 19702 14220 19708 14232
rect 19760 14220 19766 14272
rect 1104 14170 22816 14192
rect 1104 14118 4614 14170
rect 4666 14118 4678 14170
rect 4730 14118 4742 14170
rect 4794 14118 4806 14170
rect 4858 14118 11878 14170
rect 11930 14118 11942 14170
rect 11994 14118 12006 14170
rect 12058 14118 12070 14170
rect 12122 14118 19142 14170
rect 19194 14118 19206 14170
rect 19258 14118 19270 14170
rect 19322 14118 19334 14170
rect 19386 14118 22816 14170
rect 1104 14096 22816 14118
rect 1857 14059 1915 14065
rect 1857 14025 1869 14059
rect 1903 14056 1915 14059
rect 3602 14056 3608 14068
rect 1903 14028 3608 14056
rect 1903 14025 1915 14028
rect 1857 14019 1915 14025
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 4154 14016 4160 14068
rect 4212 14016 4218 14068
rect 4430 14016 4436 14068
rect 4488 14056 4494 14068
rect 4617 14059 4675 14065
rect 4617 14056 4629 14059
rect 4488 14028 4629 14056
rect 4488 14016 4494 14028
rect 4617 14025 4629 14028
rect 4663 14025 4675 14059
rect 4617 14019 4675 14025
rect 5074 14016 5080 14068
rect 5132 14056 5138 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 5132 14028 6285 14056
rect 5132 14016 5138 14028
rect 6273 14025 6285 14028
rect 6319 14025 6331 14059
rect 6273 14019 6331 14025
rect 6822 14016 6828 14068
rect 6880 14056 6886 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 6880 14028 9229 14056
rect 6880 14016 6886 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 9493 14059 9551 14065
rect 9493 14025 9505 14059
rect 9539 14056 9551 14059
rect 9766 14056 9772 14068
rect 9539 14028 9772 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 11241 14059 11299 14065
rect 11241 14025 11253 14059
rect 11287 14056 11299 14059
rect 11330 14056 11336 14068
rect 11287 14028 11336 14056
rect 11287 14025 11299 14028
rect 11241 14019 11299 14025
rect 11330 14016 11336 14028
rect 11388 14016 11394 14068
rect 12621 14059 12679 14065
rect 12621 14025 12633 14059
rect 12667 14056 12679 14059
rect 13078 14056 13084 14068
rect 12667 14028 13084 14056
rect 12667 14025 12679 14028
rect 12621 14019 12679 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13228 14028 14228 14056
rect 13228 14016 13234 14028
rect 2225 13991 2283 13997
rect 2225 13957 2237 13991
rect 2271 13988 2283 13991
rect 3234 13988 3240 14000
rect 2271 13960 3240 13988
rect 2271 13957 2283 13960
rect 2225 13951 2283 13957
rect 3234 13948 3240 13960
rect 3292 13948 3298 14000
rect 4172 13988 4200 14016
rect 4172 13960 4936 13988
rect 2682 13880 2688 13932
rect 2740 13920 2746 13932
rect 4908 13929 4936 13960
rect 5902 13948 5908 14000
rect 5960 13988 5966 14000
rect 6362 13988 6368 14000
rect 5960 13960 6368 13988
rect 5960 13948 5966 13960
rect 6362 13948 6368 13960
rect 6420 13948 6426 14000
rect 7006 13948 7012 14000
rect 7064 13988 7070 14000
rect 7064 13960 7880 13988
rect 7064 13948 7070 13960
rect 2777 13923 2835 13929
rect 2777 13920 2789 13923
rect 2740 13892 2789 13920
rect 2740 13880 2746 13892
rect 2777 13889 2789 13892
rect 2823 13889 2835 13923
rect 2777 13883 2835 13889
rect 4893 13923 4951 13929
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 4893 13883 4951 13889
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6328 13892 7297 13920
rect 6328 13880 6334 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 7558 13920 7564 13932
rect 7515 13892 7564 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 7852 13929 7880 13960
rect 7837 13923 7895 13929
rect 7837 13889 7849 13923
rect 7883 13889 7895 13923
rect 9784 13920 9812 14016
rect 11885 13991 11943 13997
rect 11885 13957 11897 13991
rect 11931 13988 11943 13991
rect 12894 13988 12900 14000
rect 11931 13960 12900 13988
rect 11931 13957 11943 13960
rect 11885 13951 11943 13957
rect 12894 13948 12900 13960
rect 12952 13948 12958 14000
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9784 13892 9873 13920
rect 7837 13883 7895 13889
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 10962 13880 10968 13932
rect 11020 13920 11026 13932
rect 11020 13892 13299 13920
rect 11020 13880 11026 13892
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 1719 13824 3188 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 2130 13744 2136 13796
rect 2188 13784 2194 13796
rect 2685 13787 2743 13793
rect 2685 13784 2697 13787
rect 2188 13756 2697 13784
rect 2188 13744 2194 13756
rect 2685 13753 2697 13756
rect 2731 13753 2743 13787
rect 2685 13747 2743 13753
rect 2593 13719 2651 13725
rect 2593 13685 2605 13719
rect 2639 13716 2651 13719
rect 2774 13716 2780 13728
rect 2639 13688 2780 13716
rect 2639 13685 2651 13688
rect 2593 13679 2651 13685
rect 2774 13676 2780 13688
rect 2832 13676 2838 13728
rect 3160 13716 3188 13824
rect 3234 13812 3240 13864
rect 3292 13852 3298 13864
rect 3504 13855 3562 13861
rect 3292 13824 3337 13852
rect 3292 13812 3298 13824
rect 3504 13821 3516 13855
rect 3550 13852 3562 13855
rect 4246 13852 4252 13864
rect 3550 13824 4252 13852
rect 3550 13821 3562 13824
rect 3504 13815 3562 13821
rect 4246 13812 4252 13824
rect 4304 13812 4310 13864
rect 4982 13812 4988 13864
rect 5040 13852 5046 13864
rect 5149 13855 5207 13861
rect 5149 13852 5161 13855
rect 5040 13824 5161 13852
rect 5040 13812 5046 13824
rect 5149 13821 5161 13824
rect 5195 13821 5207 13855
rect 6546 13852 6552 13864
rect 5149 13815 5207 13821
rect 5276 13824 6552 13852
rect 4890 13744 4896 13796
rect 4948 13784 4954 13796
rect 5276 13784 5304 13824
rect 6546 13812 6552 13824
rect 6604 13852 6610 13864
rect 7742 13852 7748 13864
rect 6604 13824 7748 13852
rect 6604 13812 6610 13824
rect 7742 13812 7748 13824
rect 7800 13812 7806 13864
rect 8093 13855 8151 13861
rect 8093 13852 8105 13855
rect 7944 13824 8105 13852
rect 7944 13796 7972 13824
rect 8093 13821 8105 13824
rect 8139 13821 8151 13855
rect 9674 13852 9680 13864
rect 9635 13824 9680 13852
rect 8093 13815 8151 13821
rect 9674 13812 9680 13824
rect 9732 13812 9738 13864
rect 10128 13855 10186 13861
rect 10128 13821 10140 13855
rect 10174 13852 10186 13855
rect 11054 13852 11060 13864
rect 10174 13824 11060 13852
rect 10174 13821 10186 13824
rect 10128 13815 10186 13821
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11422 13812 11428 13864
rect 11480 13852 11486 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11480 13824 11713 13852
rect 11480 13812 11486 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 12437 13855 12495 13861
rect 12437 13821 12449 13855
rect 12483 13852 12495 13855
rect 12986 13852 12992 13864
rect 12483 13824 12992 13852
rect 12483 13821 12495 13824
rect 12437 13815 12495 13821
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13170 13852 13176 13864
rect 13131 13824 13176 13852
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 13271 13852 13299 13892
rect 13429 13855 13487 13861
rect 13429 13852 13441 13855
rect 13271 13824 13441 13852
rect 13429 13821 13441 13824
rect 13475 13852 13487 13855
rect 13722 13852 13728 13864
rect 13475 13824 13728 13852
rect 13475 13821 13487 13824
rect 13429 13815 13487 13821
rect 13722 13812 13728 13824
rect 13780 13812 13786 13864
rect 14200 13852 14228 14028
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 15252 14028 16957 14056
rect 15252 14016 15258 14028
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 18966 14056 18972 14068
rect 16945 14019 17003 14025
rect 17604 14028 18972 14056
rect 14553 13991 14611 13997
rect 14553 13957 14565 13991
rect 14599 13957 14611 13991
rect 14553 13951 14611 13957
rect 14568 13920 14596 13951
rect 17604 13929 17632 14028
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19426 14056 19432 14068
rect 19387 14028 19432 14056
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 20254 14056 20260 14068
rect 20215 14028 20260 14056
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 20441 14059 20499 14065
rect 20441 14025 20453 14059
rect 20487 14056 20499 14059
rect 20714 14056 20720 14068
rect 20487 14028 20720 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 21913 14059 21971 14065
rect 21913 14056 21925 14059
rect 21784 14028 21925 14056
rect 21784 14016 21790 14028
rect 21913 14025 21925 14028
rect 21959 14025 21971 14059
rect 21913 14019 21971 14025
rect 20070 13988 20076 14000
rect 19904 13960 20076 13988
rect 17589 13923 17647 13929
rect 14568 13892 14964 13920
rect 14829 13855 14887 13861
rect 14829 13852 14841 13855
rect 14200 13824 14841 13852
rect 14829 13821 14841 13824
rect 14875 13821 14887 13855
rect 14936 13852 14964 13892
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 15102 13861 15108 13864
rect 15096 13852 15108 13861
rect 14936 13824 15108 13852
rect 14829 13815 14887 13821
rect 15096 13815 15108 13824
rect 15102 13812 15108 13815
rect 15160 13812 15166 13864
rect 16482 13812 16488 13864
rect 16540 13852 16546 13864
rect 17218 13852 17224 13864
rect 16540 13824 17224 13852
rect 16540 13812 16546 13824
rect 17218 13812 17224 13824
rect 17276 13852 17282 13864
rect 17954 13852 17960 13864
rect 17276 13824 17960 13852
rect 17276 13812 17282 13824
rect 17954 13812 17960 13824
rect 18012 13852 18018 13864
rect 18049 13855 18107 13861
rect 18049 13852 18061 13855
rect 18012 13824 18061 13852
rect 18012 13812 18018 13824
rect 18049 13821 18061 13824
rect 18095 13821 18107 13855
rect 18049 13815 18107 13821
rect 18316 13855 18374 13861
rect 18316 13821 18328 13855
rect 18362 13852 18374 13855
rect 19518 13852 19524 13864
rect 18362 13824 19524 13852
rect 18362 13821 18374 13824
rect 18316 13815 18374 13821
rect 19518 13812 19524 13824
rect 19576 13812 19582 13864
rect 19904 13861 19932 13960
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 20088 13892 20668 13920
rect 20088 13861 20116 13892
rect 19889 13855 19947 13861
rect 19889 13821 19901 13855
rect 19935 13821 19947 13855
rect 19889 13815 19947 13821
rect 20073 13855 20131 13861
rect 20073 13821 20085 13855
rect 20119 13821 20131 13855
rect 20073 13815 20131 13821
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13852 20499 13855
rect 20533 13855 20591 13861
rect 20533 13852 20545 13855
rect 20487 13824 20545 13852
rect 20487 13821 20499 13824
rect 20441 13815 20499 13821
rect 20533 13821 20545 13824
rect 20579 13821 20591 13855
rect 20640 13852 20668 13892
rect 21174 13852 21180 13864
rect 20640 13824 21180 13852
rect 20533 13815 20591 13821
rect 21174 13812 21180 13824
rect 21232 13812 21238 13864
rect 4948 13756 5304 13784
rect 4948 13744 4954 13756
rect 6914 13744 6920 13796
rect 6972 13784 6978 13796
rect 7926 13784 7932 13796
rect 6972 13756 7932 13784
rect 6972 13744 6978 13756
rect 7926 13744 7932 13756
rect 7984 13744 7990 13796
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 12526 13784 12532 13796
rect 8904 13756 12532 13784
rect 8904 13744 8910 13756
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 17313 13787 17371 13793
rect 17313 13753 17325 13787
rect 17359 13784 17371 13787
rect 18230 13784 18236 13796
rect 17359 13756 18236 13784
rect 17359 13753 17371 13756
rect 17313 13747 17371 13753
rect 18230 13744 18236 13756
rect 18288 13744 18294 13796
rect 20806 13793 20812 13796
rect 20800 13784 20812 13793
rect 20767 13756 20812 13784
rect 20800 13747 20812 13756
rect 20806 13744 20812 13747
rect 20864 13744 20870 13796
rect 3234 13716 3240 13728
rect 3160 13688 3240 13716
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 5350 13716 5356 13728
rect 4488 13688 5356 13716
rect 4488 13676 4494 13688
rect 5350 13676 5356 13688
rect 5408 13716 5414 13728
rect 6825 13719 6883 13725
rect 6825 13716 6837 13719
rect 5408 13688 6837 13716
rect 5408 13676 5414 13688
rect 6825 13685 6837 13688
rect 6871 13685 6883 13719
rect 6825 13679 6883 13685
rect 7006 13676 7012 13728
rect 7064 13716 7070 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7064 13688 7205 13716
rect 7064 13676 7070 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 7193 13679 7251 13685
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 11790 13716 11796 13728
rect 8812 13688 11796 13716
rect 8812 13676 8818 13688
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 16206 13716 16212 13728
rect 16167 13688 16212 13716
rect 16206 13676 16212 13688
rect 16264 13676 16270 13728
rect 16482 13716 16488 13728
rect 16443 13688 16488 13716
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 17405 13719 17463 13725
rect 17405 13685 17417 13719
rect 17451 13716 17463 13719
rect 17678 13716 17684 13728
rect 17451 13688 17684 13716
rect 17451 13685 17463 13688
rect 17405 13679 17463 13685
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 1104 13626 22816 13648
rect 1104 13574 8246 13626
rect 8298 13574 8310 13626
rect 8362 13574 8374 13626
rect 8426 13574 8438 13626
rect 8490 13574 15510 13626
rect 15562 13574 15574 13626
rect 15626 13574 15638 13626
rect 15690 13574 15702 13626
rect 15754 13574 22816 13626
rect 1104 13552 22816 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2682 13512 2688 13524
rect 1912 13484 2688 13512
rect 1912 13472 1918 13484
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 2958 13472 2964 13524
rect 3016 13512 3022 13524
rect 3513 13515 3571 13521
rect 3513 13512 3525 13515
rect 3016 13484 3525 13512
rect 3016 13472 3022 13484
rect 3513 13481 3525 13484
rect 3559 13512 3571 13515
rect 3602 13512 3608 13524
rect 3559 13484 3608 13512
rect 3559 13481 3571 13484
rect 3513 13475 3571 13481
rect 3602 13472 3608 13484
rect 3660 13472 3666 13524
rect 4246 13472 4252 13524
rect 4304 13472 4310 13524
rect 4341 13515 4399 13521
rect 4341 13481 4353 13515
rect 4387 13512 4399 13515
rect 4522 13512 4528 13524
rect 4387 13484 4528 13512
rect 4387 13481 4399 13484
rect 4341 13475 4399 13481
rect 4522 13472 4528 13484
rect 4580 13472 4586 13524
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 6914 13512 6920 13524
rect 4847 13484 6920 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 6914 13472 6920 13484
rect 6972 13472 6978 13524
rect 7466 13512 7472 13524
rect 7427 13484 7472 13512
rect 7466 13472 7472 13484
rect 7524 13472 7530 13524
rect 7926 13472 7932 13524
rect 7984 13512 7990 13524
rect 9217 13515 9275 13521
rect 9217 13512 9229 13515
rect 7984 13484 9229 13512
rect 7984 13472 7990 13484
rect 9217 13481 9229 13484
rect 9263 13481 9275 13515
rect 9217 13475 9275 13481
rect 10137 13515 10195 13521
rect 10137 13481 10149 13515
rect 10183 13512 10195 13515
rect 10962 13512 10968 13524
rect 10183 13484 10968 13512
rect 10183 13481 10195 13484
rect 10137 13475 10195 13481
rect 10962 13472 10968 13484
rect 11020 13472 11026 13524
rect 11146 13512 11152 13524
rect 11107 13484 11152 13512
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 11609 13515 11667 13521
rect 11609 13481 11621 13515
rect 11655 13512 11667 13515
rect 11655 13484 12848 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 2400 13447 2458 13453
rect 2400 13413 2412 13447
rect 2446 13444 2458 13447
rect 3050 13444 3056 13456
rect 2446 13416 3056 13444
rect 2446 13413 2458 13416
rect 2400 13407 2458 13413
rect 3050 13404 3056 13416
rect 3108 13404 3114 13456
rect 1581 13379 1639 13385
rect 1581 13345 1593 13379
rect 1627 13376 1639 13379
rect 1762 13376 1768 13388
rect 1627 13348 1768 13376
rect 1627 13345 1639 13348
rect 1581 13339 1639 13345
rect 1762 13336 1768 13348
rect 1820 13336 1826 13388
rect 4264 13320 4292 13472
rect 5620 13447 5678 13453
rect 5620 13413 5632 13447
rect 5666 13444 5678 13447
rect 9306 13444 9312 13456
rect 5666 13416 9312 13444
rect 5666 13413 5678 13416
rect 5620 13407 5678 13413
rect 9306 13404 9312 13416
rect 9364 13404 9370 13456
rect 12820 13444 12848 13484
rect 13722 13472 13728 13524
rect 13780 13512 13786 13524
rect 15013 13515 15071 13521
rect 15013 13512 15025 13515
rect 13780 13484 15025 13512
rect 13780 13472 13786 13484
rect 15013 13481 15025 13484
rect 15059 13481 15071 13515
rect 15013 13475 15071 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 16574 13512 16580 13524
rect 15795 13484 16580 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 16574 13472 16580 13484
rect 16632 13472 16638 13524
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 17402 13512 17408 13524
rect 17000 13484 17408 13512
rect 17000 13472 17006 13484
rect 17402 13472 17408 13484
rect 17460 13472 17466 13524
rect 17678 13512 17684 13524
rect 17639 13484 17684 13512
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 18046 13472 18052 13524
rect 18104 13512 18110 13524
rect 19242 13512 19248 13524
rect 18104 13484 19248 13512
rect 18104 13472 18110 13484
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19518 13512 19524 13524
rect 19383 13484 19524 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 19794 13472 19800 13524
rect 19852 13512 19858 13524
rect 20257 13515 20315 13521
rect 20257 13512 20269 13515
rect 19852 13484 20269 13512
rect 19852 13472 19858 13484
rect 20257 13481 20269 13484
rect 20303 13481 20315 13515
rect 20257 13475 20315 13481
rect 13878 13447 13936 13453
rect 13878 13444 13890 13447
rect 12820 13416 13890 13444
rect 13878 13413 13890 13416
rect 13924 13444 13936 13447
rect 14366 13444 14372 13456
rect 13924 13416 14372 13444
rect 13924 13413 13936 13416
rect 13878 13407 13936 13413
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 16482 13404 16488 13456
rect 16540 13444 16546 13456
rect 20165 13447 20223 13453
rect 20165 13444 20177 13447
rect 16540 13416 20177 13444
rect 16540 13404 16546 13416
rect 20165 13413 20177 13416
rect 20211 13413 20223 13447
rect 20165 13407 20223 13413
rect 21168 13447 21226 13453
rect 21168 13413 21180 13447
rect 21214 13444 21226 13447
rect 21726 13444 21732 13456
rect 21214 13416 21732 13444
rect 21214 13413 21226 13416
rect 21168 13407 21226 13413
rect 21726 13404 21732 13416
rect 21784 13404 21790 13456
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 6822 13376 6828 13388
rect 4755 13348 6828 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 6822 13336 6828 13348
rect 6880 13336 6886 13388
rect 7282 13376 7288 13388
rect 7243 13348 7288 13376
rect 7282 13336 7288 13348
rect 7340 13336 7346 13388
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8093 13379 8151 13385
rect 8093 13376 8105 13379
rect 7984 13348 8105 13376
rect 7984 13336 7990 13348
rect 8093 13345 8105 13348
rect 8139 13345 8151 13379
rect 8093 13339 8151 13345
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13376 10287 13379
rect 11609 13379 11667 13385
rect 11609 13376 11621 13379
rect 10275 13348 11621 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 11609 13345 11621 13348
rect 11655 13345 11667 13379
rect 11790 13376 11796 13388
rect 11751 13348 11796 13376
rect 11609 13339 11667 13345
rect 11790 13336 11796 13348
rect 11848 13336 11854 13388
rect 15657 13379 15715 13385
rect 15657 13345 15669 13379
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 1728 13280 2145 13308
rect 1728 13268 1734 13280
rect 2133 13277 2145 13280
rect 2179 13277 2191 13311
rect 2133 13271 2191 13277
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4890 13308 4896 13320
rect 4851 13280 4896 13308
rect 4890 13268 4896 13280
rect 4948 13268 4954 13320
rect 5166 13268 5172 13320
rect 5224 13308 5230 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5224 13280 5365 13308
rect 5224 13268 5230 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 7837 13311 7895 13317
rect 7837 13308 7849 13311
rect 7800 13280 7849 13308
rect 7800 13268 7806 13280
rect 7837 13277 7849 13280
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 9766 13268 9772 13320
rect 9824 13308 9830 13320
rect 10318 13308 10324 13320
rect 9824 13280 10324 13308
rect 9824 13268 9830 13280
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10410 13268 10416 13320
rect 10468 13308 10474 13320
rect 11241 13311 11299 13317
rect 11241 13308 11253 13311
rect 10468 13280 11253 13308
rect 10468 13268 10474 13280
rect 11241 13277 11253 13280
rect 11287 13277 11299 13311
rect 11241 13271 11299 13277
rect 11425 13311 11483 13317
rect 11425 13277 11437 13311
rect 11471 13308 11483 13311
rect 12342 13308 12348 13320
rect 11471 13280 12348 13308
rect 11471 13277 11483 13280
rect 11425 13271 11483 13277
rect 12342 13268 12348 13280
rect 12400 13268 12406 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 13170 13308 13176 13320
rect 12676 13280 13176 13308
rect 12676 13268 12682 13280
rect 13170 13268 13176 13280
rect 13228 13308 13234 13320
rect 13633 13311 13691 13317
rect 13633 13308 13645 13311
rect 13228 13280 13645 13308
rect 13228 13268 13234 13280
rect 13633 13277 13645 13280
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 7098 13200 7104 13252
rect 7156 13240 7162 13252
rect 7282 13240 7288 13252
rect 7156 13212 7288 13240
rect 7156 13200 7162 13212
rect 7282 13200 7288 13212
rect 7340 13200 7346 13252
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 12710 13240 12716 13252
rect 9732 13212 12716 13240
rect 9732 13200 9738 13212
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 1762 13172 1768 13184
rect 1723 13144 1768 13172
rect 1762 13132 1768 13144
rect 1820 13132 1826 13184
rect 5350 13132 5356 13184
rect 5408 13172 5414 13184
rect 6733 13175 6791 13181
rect 6733 13172 6745 13175
rect 5408 13144 6745 13172
rect 5408 13132 5414 13144
rect 6733 13141 6745 13144
rect 6779 13141 6791 13175
rect 6733 13135 6791 13141
rect 9769 13175 9827 13181
rect 9769 13141 9781 13175
rect 9815 13172 9827 13175
rect 10686 13172 10692 13184
rect 9815 13144 10692 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10781 13175 10839 13181
rect 10781 13141 10793 13175
rect 10827 13172 10839 13175
rect 11422 13172 11428 13184
rect 10827 13144 11428 13172
rect 10827 13141 10839 13144
rect 10781 13135 10839 13141
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 13081 13175 13139 13181
rect 13081 13172 13093 13175
rect 11756 13144 13093 13172
rect 11756 13132 11762 13144
rect 13081 13141 13093 13144
rect 13127 13141 13139 13175
rect 15286 13172 15292 13184
rect 15247 13144 15292 13172
rect 13081 13135 13139 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15672 13172 15700 13339
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 16301 13379 16359 13385
rect 16301 13376 16313 13379
rect 15804 13348 16313 13376
rect 15804 13336 15810 13348
rect 16301 13345 16313 13348
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16568 13379 16626 13385
rect 16568 13345 16580 13379
rect 16614 13376 16626 13379
rect 17310 13376 17316 13388
rect 16614 13348 17316 13376
rect 16614 13345 16626 13348
rect 16568 13339 16626 13345
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 18230 13385 18236 13388
rect 18224 13376 18236 13385
rect 18191 13348 18236 13376
rect 18224 13339 18236 13348
rect 18288 13376 18294 13388
rect 19426 13376 19432 13388
rect 18288 13348 19432 13376
rect 18230 13336 18236 13339
rect 18288 13336 18294 13348
rect 19426 13336 19432 13348
rect 19484 13336 19490 13388
rect 20714 13336 20720 13388
rect 20772 13376 20778 13388
rect 20898 13376 20904 13388
rect 20772 13348 20904 13376
rect 20772 13336 20778 13348
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 15933 13311 15991 13317
rect 15933 13277 15945 13311
rect 15979 13308 15991 13311
rect 16206 13308 16212 13320
rect 15979 13280 16212 13308
rect 15979 13277 15991 13280
rect 15933 13271 15991 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 17954 13308 17960 13320
rect 17915 13280 17960 13308
rect 17954 13268 17960 13280
rect 18012 13268 18018 13320
rect 20438 13308 20444 13320
rect 20399 13280 20444 13308
rect 20438 13268 20444 13280
rect 20496 13268 20502 13320
rect 18230 13172 18236 13184
rect 15672 13144 18236 13172
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 19797 13175 19855 13181
rect 19797 13141 19809 13175
rect 19843 13172 19855 13175
rect 20806 13172 20812 13184
rect 19843 13144 20812 13172
rect 19843 13141 19855 13144
rect 19797 13135 19855 13141
rect 20806 13132 20812 13144
rect 20864 13132 20870 13184
rect 21174 13132 21180 13184
rect 21232 13172 21238 13184
rect 22281 13175 22339 13181
rect 22281 13172 22293 13175
rect 21232 13144 22293 13172
rect 21232 13132 21238 13144
rect 22281 13141 22293 13144
rect 22327 13141 22339 13175
rect 22281 13135 22339 13141
rect 1104 13082 22816 13104
rect 1104 13030 4614 13082
rect 4666 13030 4678 13082
rect 4730 13030 4742 13082
rect 4794 13030 4806 13082
rect 4858 13030 11878 13082
rect 11930 13030 11942 13082
rect 11994 13030 12006 13082
rect 12058 13030 12070 13082
rect 12122 13030 19142 13082
rect 19194 13030 19206 13082
rect 19258 13030 19270 13082
rect 19322 13030 19334 13082
rect 19386 13030 22816 13082
rect 1104 13008 22816 13030
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4304 12940 4721 12968
rect 4304 12928 4310 12940
rect 4709 12937 4721 12940
rect 4755 12937 4767 12971
rect 4709 12931 4767 12937
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5718 12968 5724 12980
rect 5316 12940 5724 12968
rect 5316 12928 5322 12940
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7006 12968 7012 12980
rect 6967 12940 7012 12968
rect 7006 12928 7012 12940
rect 7064 12928 7070 12980
rect 7926 12928 7932 12980
rect 7984 12968 7990 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 7984 12940 9137 12968
rect 7984 12928 7990 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 9217 12971 9275 12977
rect 9217 12937 9229 12971
rect 9263 12968 9275 12971
rect 9263 12940 12020 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 7469 12903 7527 12909
rect 7469 12869 7481 12903
rect 7515 12869 7527 12903
rect 7469 12863 7527 12869
rect 11425 12903 11483 12909
rect 11425 12869 11437 12903
rect 11471 12900 11483 12903
rect 11882 12900 11888 12912
rect 11471 12872 11888 12900
rect 11471 12869 11483 12872
rect 11425 12863 11483 12869
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 7484 12832 7512 12863
rect 11882 12860 11888 12872
rect 11940 12860 11946 12912
rect 7742 12832 7748 12844
rect 7484 12804 7748 12832
rect 7742 12792 7748 12804
rect 7800 12792 7806 12844
rect 9674 12832 9680 12844
rect 9635 12804 9680 12832
rect 9674 12792 9680 12804
rect 9732 12792 9738 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9824 12804 9917 12832
rect 9824 12792 9830 12804
rect 11054 12792 11060 12844
rect 11112 12832 11118 12844
rect 11992 12841 12020 12940
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 13817 12971 13875 12977
rect 13817 12968 13829 12971
rect 12768 12940 13829 12968
rect 12768 12928 12774 12940
rect 13817 12937 13829 12940
rect 13863 12937 13875 12971
rect 13817 12931 13875 12937
rect 15304 12940 17448 12968
rect 11977 12835 12035 12841
rect 11112 12804 11928 12832
rect 11112 12792 11118 12804
rect 1688 12764 1716 12792
rect 3602 12773 3608 12776
rect 3329 12767 3387 12773
rect 3329 12764 3341 12767
rect 1688 12736 3341 12764
rect 3329 12733 3341 12736
rect 3375 12733 3387 12767
rect 3596 12764 3608 12773
rect 3563 12736 3608 12764
rect 3329 12727 3387 12733
rect 3596 12727 3608 12736
rect 1940 12699 1998 12705
rect 1940 12665 1952 12699
rect 1986 12696 1998 12699
rect 2774 12696 2780 12708
rect 1986 12668 2780 12696
rect 1986 12665 1998 12668
rect 1940 12659 1998 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 3344 12696 3372 12727
rect 3602 12724 3608 12727
rect 3660 12724 3666 12776
rect 5077 12767 5135 12773
rect 5077 12764 5089 12767
rect 3712 12736 5089 12764
rect 3712 12696 3740 12736
rect 5077 12733 5089 12736
rect 5123 12764 5135 12767
rect 5166 12764 5172 12776
rect 5123 12736 5172 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5166 12724 5172 12736
rect 5224 12724 5230 12776
rect 5350 12773 5356 12776
rect 5344 12764 5356 12773
rect 5311 12736 5356 12764
rect 5344 12727 5356 12736
rect 5350 12724 5356 12727
rect 5408 12724 5414 12776
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 7616 12736 7665 12764
rect 7616 12724 7622 12736
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 8754 12764 8760 12776
rect 7653 12727 7711 12733
rect 7760 12736 8760 12764
rect 3344 12668 3740 12696
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 7760 12696 7788 12736
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9784 12764 9812 12792
rect 9180 12736 9812 12764
rect 9180 12724 9186 12736
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10045 12767 10103 12773
rect 10045 12764 10057 12767
rect 9916 12736 10057 12764
rect 9916 12724 9922 12736
rect 10045 12733 10057 12736
rect 10091 12764 10103 12767
rect 10594 12764 10600 12776
rect 10091 12736 10600 12764
rect 10091 12733 10103 12736
rect 10045 12727 10103 12733
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 10686 12724 10692 12776
rect 10744 12764 10750 12776
rect 11900 12764 11928 12804
rect 11977 12801 11989 12835
rect 12023 12801 12035 12835
rect 11977 12795 12035 12801
rect 12161 12835 12219 12841
rect 12161 12801 12173 12835
rect 12207 12832 12219 12835
rect 12342 12832 12348 12844
rect 12207 12804 12348 12832
rect 12207 12801 12219 12804
rect 12161 12795 12219 12801
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 14918 12832 14924 12844
rect 14599 12804 14924 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 12437 12767 12495 12773
rect 12437 12764 12449 12767
rect 10744 12736 11468 12764
rect 11900 12736 12449 12764
rect 10744 12724 10750 12736
rect 8018 12705 8024 12708
rect 4120 12668 7788 12696
rect 4120 12656 4126 12668
rect 8012 12659 8024 12705
rect 8076 12696 8082 12708
rect 9585 12699 9643 12705
rect 8076 12668 8112 12696
rect 8018 12656 8024 12659
rect 8076 12656 8082 12668
rect 9585 12665 9597 12699
rect 9631 12696 9643 12699
rect 10312 12699 10370 12705
rect 9631 12668 10272 12696
rect 9631 12665 9643 12668
rect 9585 12659 9643 12665
rect 4982 12588 4988 12640
rect 5040 12628 5046 12640
rect 6457 12631 6515 12637
rect 6457 12628 6469 12631
rect 5040 12600 6469 12628
rect 5040 12588 5046 12600
rect 6457 12597 6469 12600
rect 6503 12597 6515 12631
rect 10244 12628 10272 12668
rect 10312 12665 10324 12699
rect 10358 12696 10370 12699
rect 11330 12696 11336 12708
rect 10358 12668 11336 12696
rect 10358 12665 10370 12668
rect 10312 12659 10370 12665
rect 11330 12656 11336 12668
rect 11388 12656 11394 12708
rect 11440 12696 11468 12736
rect 12437 12733 12449 12736
rect 12483 12733 12495 12767
rect 12437 12727 12495 12733
rect 12526 12724 12532 12776
rect 12584 12764 12590 12776
rect 14369 12767 14427 12773
rect 14369 12764 14381 12767
rect 12584 12736 14381 12764
rect 12584 12724 12590 12736
rect 14369 12733 14381 12736
rect 14415 12733 14427 12767
rect 14369 12727 14427 12733
rect 14737 12767 14795 12773
rect 14737 12733 14749 12767
rect 14783 12764 14795 12767
rect 15304 12764 15332 12940
rect 16758 12900 16764 12912
rect 16719 12872 16764 12900
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 17310 12900 17316 12912
rect 16868 12872 17316 12900
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 16868 12832 16896 12872
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 17420 12900 17448 12940
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 17589 12971 17647 12977
rect 17589 12968 17601 12971
rect 17552 12940 17601 12968
rect 17552 12928 17558 12940
rect 17589 12937 17601 12940
rect 17635 12937 17647 12971
rect 19426 12968 19432 12980
rect 19387 12940 19432 12968
rect 17589 12931 17647 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19702 12928 19708 12980
rect 19760 12968 19766 12980
rect 19886 12968 19892 12980
rect 19760 12940 19892 12968
rect 19760 12928 19766 12940
rect 19886 12928 19892 12940
rect 19944 12928 19950 12980
rect 21082 12928 21088 12980
rect 21140 12968 21146 12980
rect 22281 12971 22339 12977
rect 22281 12968 22293 12971
rect 21140 12940 22293 12968
rect 21140 12928 21146 12940
rect 22281 12937 22293 12940
rect 22327 12937 22339 12971
rect 22281 12931 22339 12937
rect 18046 12900 18052 12912
rect 17420 12872 18052 12900
rect 18046 12860 18052 12872
rect 18104 12860 18110 12912
rect 17862 12832 17868 12844
rect 16632 12804 16896 12832
rect 17328 12804 17868 12832
rect 16632 12792 16638 12804
rect 14783 12736 15332 12764
rect 15381 12767 15439 12773
rect 14783 12733 14795 12736
rect 14737 12727 14795 12733
rect 15381 12733 15393 12767
rect 15427 12764 15439 12767
rect 15470 12764 15476 12776
rect 15427 12736 15476 12764
rect 15427 12733 15439 12736
rect 15381 12727 15439 12733
rect 15470 12724 15476 12736
rect 15528 12724 15534 12776
rect 15648 12767 15706 12773
rect 15648 12733 15660 12767
rect 15694 12764 15706 12767
rect 16206 12764 16212 12776
rect 15694 12736 16212 12764
rect 15694 12733 15706 12736
rect 15648 12727 15706 12733
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 17328 12773 17356 12804
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 20533 12835 20591 12841
rect 20533 12801 20545 12835
rect 20579 12832 20591 12835
rect 20714 12832 20720 12844
rect 20579 12804 20720 12832
rect 20579 12801 20591 12804
rect 20533 12795 20591 12801
rect 20714 12792 20720 12804
rect 20772 12792 20778 12844
rect 20898 12832 20904 12844
rect 20859 12804 20904 12832
rect 20898 12792 20904 12804
rect 20956 12792 20962 12844
rect 17313 12767 17371 12773
rect 17313 12733 17325 12767
rect 17359 12733 17371 12767
rect 17313 12727 17371 12733
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 17460 12736 17505 12764
rect 17460 12724 17466 12736
rect 17954 12724 17960 12776
rect 18012 12764 18018 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 18012 12736 18061 12764
rect 18012 12724 18018 12736
rect 18049 12733 18061 12736
rect 18095 12764 18107 12767
rect 20916 12764 20944 12792
rect 21174 12773 21180 12776
rect 21168 12764 21180 12773
rect 18095 12736 20944 12764
rect 21135 12736 21180 12764
rect 18095 12733 18107 12736
rect 18049 12727 18107 12733
rect 21168 12727 21180 12736
rect 21174 12724 21180 12727
rect 21232 12724 21238 12776
rect 11885 12699 11943 12705
rect 11885 12696 11897 12699
rect 11440 12668 11897 12696
rect 11885 12665 11897 12668
rect 11931 12665 11943 12699
rect 11885 12659 11943 12665
rect 12158 12656 12164 12708
rect 12216 12696 12222 12708
rect 12682 12699 12740 12705
rect 12682 12696 12694 12699
rect 12216 12668 12694 12696
rect 12216 12656 12222 12668
rect 12682 12665 12694 12668
rect 12728 12665 12740 12699
rect 15010 12696 15016 12708
rect 12682 12659 12740 12665
rect 13924 12668 15016 12696
rect 11054 12628 11060 12640
rect 10244 12600 11060 12628
rect 6457 12591 6515 12597
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11514 12628 11520 12640
rect 11475 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 13924 12637 13952 12668
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 15105 12699 15163 12705
rect 15105 12665 15117 12699
rect 15151 12696 15163 12699
rect 15151 12668 17632 12696
rect 15151 12665 15163 12668
rect 15105 12659 15163 12665
rect 13909 12631 13967 12637
rect 13909 12597 13921 12631
rect 13955 12597 13967 12631
rect 14274 12628 14280 12640
rect 14235 12600 14280 12628
rect 13909 12591 13967 12597
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 14918 12628 14924 12640
rect 14879 12600 14924 12628
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 15838 12588 15844 12640
rect 15896 12628 15902 12640
rect 16206 12628 16212 12640
rect 15896 12600 16212 12628
rect 15896 12588 15902 12600
rect 16206 12588 16212 12600
rect 16264 12628 16270 12640
rect 17129 12631 17187 12637
rect 17129 12628 17141 12631
rect 16264 12600 17141 12628
rect 16264 12588 16270 12600
rect 17129 12597 17141 12600
rect 17175 12628 17187 12631
rect 17310 12628 17316 12640
rect 17175 12600 17316 12628
rect 17175 12597 17187 12600
rect 17129 12591 17187 12597
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 17604 12628 17632 12668
rect 17678 12656 17684 12708
rect 17736 12696 17742 12708
rect 18294 12699 18352 12705
rect 18294 12696 18306 12699
rect 17736 12668 18306 12696
rect 17736 12656 17742 12668
rect 18294 12665 18306 12668
rect 18340 12665 18352 12699
rect 18294 12659 18352 12665
rect 20257 12699 20315 12705
rect 20257 12665 20269 12699
rect 20303 12696 20315 12699
rect 20806 12696 20812 12708
rect 20303 12668 20812 12696
rect 20303 12665 20315 12668
rect 20257 12659 20315 12665
rect 20806 12656 20812 12668
rect 20864 12696 20870 12708
rect 21634 12696 21640 12708
rect 20864 12668 21640 12696
rect 20864 12656 20870 12668
rect 21634 12656 21640 12668
rect 21692 12656 21698 12708
rect 19334 12628 19340 12640
rect 17604 12600 19340 12628
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 19886 12628 19892 12640
rect 19847 12600 19892 12628
rect 19886 12588 19892 12600
rect 19944 12588 19950 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 20404 12600 20449 12628
rect 20404 12588 20410 12600
rect 1104 12538 22816 12560
rect 1104 12486 8246 12538
rect 8298 12486 8310 12538
rect 8362 12486 8374 12538
rect 8426 12486 8438 12538
rect 8490 12486 15510 12538
rect 15562 12486 15574 12538
rect 15626 12486 15638 12538
rect 15690 12486 15702 12538
rect 15754 12486 22816 12538
rect 1104 12464 22816 12486
rect 1578 12384 1584 12436
rect 1636 12384 1642 12436
rect 2130 12384 2136 12436
rect 2188 12424 2194 12436
rect 2777 12427 2835 12433
rect 2777 12424 2789 12427
rect 2188 12396 2789 12424
rect 2188 12384 2194 12396
rect 2777 12393 2789 12396
rect 2823 12393 2835 12427
rect 2777 12387 2835 12393
rect 2958 12384 2964 12436
rect 3016 12424 3022 12436
rect 3605 12427 3663 12433
rect 3605 12424 3617 12427
rect 3016 12396 3617 12424
rect 3016 12384 3022 12396
rect 3605 12393 3617 12396
rect 3651 12393 3663 12427
rect 3605 12387 3663 12393
rect 4154 12384 4160 12436
rect 4212 12384 4218 12436
rect 4341 12427 4399 12433
rect 4341 12393 4353 12427
rect 4387 12424 4399 12427
rect 5258 12424 5264 12436
rect 4387 12396 5264 12424
rect 4387 12393 4399 12396
rect 4341 12387 4399 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6365 12427 6423 12433
rect 6365 12424 6377 12427
rect 6144 12396 6377 12424
rect 6144 12384 6150 12396
rect 6365 12393 6377 12396
rect 6411 12393 6423 12427
rect 6365 12387 6423 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 10410 12424 10416 12436
rect 8619 12396 10416 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 10410 12384 10416 12396
rect 10468 12384 10474 12436
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 12437 12427 12495 12433
rect 12437 12424 12449 12427
rect 10888 12396 12449 12424
rect 1596 12356 1624 12384
rect 4172 12356 4200 12384
rect 8846 12356 8852 12368
rect 1596 12328 4200 12356
rect 4632 12328 8852 12356
rect 1486 12248 1492 12300
rect 1544 12288 1550 12300
rect 1653 12291 1711 12297
rect 1653 12288 1665 12291
rect 1544 12260 1665 12288
rect 1544 12248 1550 12260
rect 1653 12257 1665 12260
rect 1699 12257 1711 12291
rect 1653 12251 1711 12257
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3329 12291 3387 12297
rect 3329 12288 3341 12291
rect 3108 12260 3341 12288
rect 3108 12248 3114 12260
rect 3329 12257 3341 12260
rect 3375 12257 3387 12291
rect 3329 12251 3387 12257
rect 3421 12291 3479 12297
rect 3421 12257 3433 12291
rect 3467 12257 3479 12291
rect 3421 12251 3479 12257
rect 4157 12291 4215 12297
rect 4157 12257 4169 12291
rect 4203 12288 4215 12291
rect 4338 12288 4344 12300
rect 4203 12260 4344 12288
rect 4203 12257 4215 12260
rect 4157 12251 4215 12257
rect 1394 12220 1400 12232
rect 1355 12192 1400 12220
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 3436 12220 3464 12251
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4632 12220 4660 12328
rect 8846 12316 8852 12328
rect 8904 12316 8910 12368
rect 4982 12297 4988 12300
rect 4976 12288 4988 12297
rect 4943 12260 4988 12288
rect 4976 12251 4988 12260
rect 4982 12248 4988 12251
rect 5040 12248 5046 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 10888 12297 10916 12396
rect 12437 12393 12449 12396
rect 12483 12393 12495 12427
rect 14366 12424 14372 12436
rect 14327 12396 14372 12424
rect 12437 12387 12495 12393
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 15289 12427 15347 12433
rect 15289 12393 15301 12427
rect 15335 12424 15347 12427
rect 16298 12424 16304 12436
rect 15335 12396 16304 12424
rect 15335 12393 15347 12396
rect 15289 12387 15347 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 16390 12384 16396 12436
rect 16448 12424 16454 12436
rect 18782 12424 18788 12436
rect 16448 12396 18788 12424
rect 16448 12384 16454 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 19334 12384 19340 12436
rect 19392 12424 19398 12436
rect 19392 12396 19739 12424
rect 19392 12384 19398 12396
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 13234 12359 13292 12365
rect 13234 12356 13246 12359
rect 11112 12328 13246 12356
rect 11112 12316 11118 12328
rect 13234 12325 13246 12328
rect 13280 12356 13292 12359
rect 13814 12356 13820 12368
rect 13280 12328 13820 12356
rect 13280 12325 13292 12328
rect 13234 12319 13292 12325
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 14921 12359 14979 12365
rect 14921 12325 14933 12359
rect 14967 12356 14979 12359
rect 15102 12356 15108 12368
rect 14967 12328 15108 12356
rect 14967 12325 14979 12328
rect 14921 12319 14979 12325
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 17126 12356 17132 12368
rect 15488 12328 17132 12356
rect 6733 12291 6791 12297
rect 6733 12288 6745 12291
rect 5592 12260 6745 12288
rect 5592 12248 5598 12260
rect 6733 12257 6745 12260
rect 6779 12257 6791 12291
rect 7929 12291 7987 12297
rect 7929 12288 7941 12291
rect 6733 12251 6791 12257
rect 6932 12260 7941 12288
rect 3436 12192 4660 12220
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 4338 12152 4344 12164
rect 3436 12124 4344 12152
rect 1394 12044 1400 12096
rect 1452 12084 1458 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 1452 12056 3157 12084
rect 1452 12044 1458 12056
rect 3145 12053 3157 12056
rect 3191 12084 3203 12087
rect 3436 12084 3464 12124
rect 4338 12112 4344 12124
rect 4396 12152 4402 12164
rect 4724 12152 4752 12183
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6825 12223 6883 12229
rect 6825 12220 6837 12223
rect 5776 12192 6837 12220
rect 5776 12180 5782 12192
rect 6825 12189 6837 12192
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 4396 12124 4752 12152
rect 4396 12112 4402 12124
rect 5810 12112 5816 12164
rect 5868 12152 5874 12164
rect 6932 12152 6960 12260
rect 7929 12257 7941 12260
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 8941 12291 8999 12297
rect 8941 12257 8953 12291
rect 8987 12288 8999 12291
rect 10045 12291 10103 12297
rect 8987 12260 9996 12288
rect 8987 12257 8999 12260
rect 8941 12251 8999 12257
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7190 12220 7196 12232
rect 7055 12192 7196 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 8021 12223 8079 12229
rect 8021 12220 8033 12223
rect 7524 12192 8033 12220
rect 7524 12180 7530 12192
rect 8021 12189 8033 12192
rect 8067 12189 8079 12223
rect 8021 12183 8079 12189
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 9033 12223 9091 12229
rect 8168 12192 8261 12220
rect 8168 12180 8174 12192
rect 9033 12189 9045 12223
rect 9079 12189 9091 12223
rect 9033 12183 9091 12189
rect 5868 12124 6960 12152
rect 7208 12152 7236 12180
rect 8128 12152 8156 12180
rect 7208 12124 8156 12152
rect 9048 12152 9076 12183
rect 9122 12180 9128 12232
rect 9180 12220 9186 12232
rect 9180 12192 9225 12220
rect 9180 12180 9186 12192
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9769 12223 9827 12229
rect 9769 12220 9781 12223
rect 9456 12192 9781 12220
rect 9456 12180 9462 12192
rect 9769 12189 9781 12192
rect 9815 12189 9827 12223
rect 9968 12220 9996 12260
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10873 12291 10931 12297
rect 10873 12288 10885 12291
rect 10091 12260 10885 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10873 12257 10885 12260
rect 10919 12257 10931 12291
rect 10873 12251 10931 12257
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12288 14795 12291
rect 15488 12288 15516 12328
rect 17126 12316 17132 12328
rect 17184 12316 17190 12368
rect 17218 12316 17224 12368
rect 17276 12356 17282 12368
rect 19610 12356 19616 12368
rect 17276 12328 19616 12356
rect 17276 12316 17282 12328
rect 19610 12316 19616 12328
rect 19668 12316 19674 12368
rect 19711 12356 19739 12396
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 19944 12396 20269 12424
rect 19944 12384 19950 12396
rect 20257 12393 20269 12396
rect 20303 12393 20315 12427
rect 20257 12387 20315 12393
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 22281 12427 22339 12433
rect 22281 12424 22293 12427
rect 20496 12396 22293 12424
rect 20496 12384 20502 12396
rect 22281 12393 22293 12396
rect 22327 12393 22339 12427
rect 22281 12387 22339 12393
rect 19711 12328 19932 12356
rect 19904 12300 19932 12328
rect 21082 12316 21088 12368
rect 21140 12365 21146 12368
rect 21140 12359 21204 12365
rect 21140 12325 21158 12359
rect 21192 12325 21204 12359
rect 21140 12319 21204 12325
rect 21140 12316 21146 12319
rect 15654 12288 15660 12300
rect 14783 12260 15516 12288
rect 15615 12260 15660 12288
rect 14783 12257 14795 12260
rect 14737 12251 14795 12257
rect 10134 12220 10140 12232
rect 9968 12192 10140 12220
rect 9769 12183 9827 12189
rect 10134 12180 10140 12192
rect 10192 12180 10198 12232
rect 10226 12180 10232 12232
rect 10284 12220 10290 12232
rect 11164 12220 11192 12251
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 16206 12288 16212 12300
rect 16167 12260 16212 12288
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 16298 12248 16304 12300
rect 16356 12248 16362 12300
rect 16476 12291 16534 12297
rect 16476 12257 16488 12291
rect 16522 12288 16534 12291
rect 16758 12288 16764 12300
rect 16522 12260 16764 12288
rect 16522 12257 16534 12260
rect 16476 12251 16534 12257
rect 16758 12248 16764 12260
rect 16816 12248 16822 12300
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 17954 12288 17960 12300
rect 17368 12260 17960 12288
rect 17368 12248 17374 12260
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18213 12291 18271 12297
rect 18213 12288 18225 12291
rect 18104 12260 18225 12288
rect 18104 12248 18110 12260
rect 18213 12257 18225 12260
rect 18259 12257 18271 12291
rect 18213 12251 18271 12257
rect 18782 12248 18788 12300
rect 18840 12288 18846 12300
rect 18840 12260 19380 12288
rect 18840 12248 18846 12260
rect 10284 12192 11192 12220
rect 10284 12180 10290 12192
rect 12526 12180 12532 12232
rect 12584 12220 12590 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12584 12192 13001 12220
rect 12584 12180 12590 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 12989 12183 13047 12189
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 15105 12223 15163 12229
rect 15105 12220 15117 12223
rect 14700 12192 15117 12220
rect 14700 12180 14706 12192
rect 15105 12189 15117 12192
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 15194 12180 15200 12232
rect 15252 12220 15258 12232
rect 15672 12220 15700 12248
rect 15252 12192 15700 12220
rect 15252 12180 15258 12192
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15930 12220 15936 12232
rect 15804 12192 15849 12220
rect 15891 12192 15936 12220
rect 15804 12180 15810 12192
rect 15930 12180 15936 12192
rect 15988 12180 15994 12232
rect 16316 12220 16344 12248
rect 16040 12192 16344 12220
rect 9306 12152 9312 12164
rect 9048 12124 9312 12152
rect 5868 12112 5874 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 16040 12152 16068 12192
rect 19352 12161 19380 12260
rect 19886 12248 19892 12300
rect 19944 12248 19950 12300
rect 20070 12248 20076 12300
rect 20128 12288 20134 12300
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 20128 12260 20177 12288
rect 20128 12248 20134 12260
rect 20165 12257 20177 12260
rect 20211 12257 20223 12291
rect 20898 12288 20904 12300
rect 20859 12260 20904 12288
rect 20165 12251 20223 12257
rect 20898 12248 20904 12260
rect 20956 12248 20962 12300
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 20806 12220 20812 12232
rect 20487 12192 20812 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 9416 12124 9996 12152
rect 3191 12056 3464 12084
rect 3191 12053 3203 12056
rect 3145 12047 3203 12053
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 6052 12056 6101 12084
rect 6052 12044 6058 12056
rect 6089 12053 6101 12056
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7156 12056 7573 12084
rect 7156 12044 7162 12056
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7561 12047 7619 12053
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9416 12084 9444 12124
rect 8628 12056 9444 12084
rect 9769 12087 9827 12093
rect 8628 12044 8634 12056
rect 9769 12053 9781 12087
rect 9815 12084 9827 12087
rect 9861 12087 9919 12093
rect 9861 12084 9873 12087
rect 9815 12056 9873 12084
rect 9815 12053 9827 12056
rect 9769 12047 9827 12053
rect 9861 12053 9873 12056
rect 9907 12053 9919 12087
rect 9968 12084 9996 12124
rect 15580 12124 16068 12152
rect 19337 12155 19395 12161
rect 15580 12084 15608 12124
rect 19337 12121 19349 12155
rect 19383 12121 19395 12155
rect 19337 12115 19395 12121
rect 9968 12056 15608 12084
rect 9861 12047 9919 12053
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 16850 12084 16856 12096
rect 15712 12056 16856 12084
rect 15712 12044 15718 12056
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17586 12084 17592 12096
rect 17547 12056 17592 12084
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 19797 12087 19855 12093
rect 19797 12053 19809 12087
rect 19843 12084 19855 12087
rect 20530 12084 20536 12096
rect 19843 12056 20536 12084
rect 19843 12053 19855 12056
rect 19797 12047 19855 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 22816 12016
rect 1104 11942 4614 11994
rect 4666 11942 4678 11994
rect 4730 11942 4742 11994
rect 4794 11942 4806 11994
rect 4858 11942 11878 11994
rect 11930 11942 11942 11994
rect 11994 11942 12006 11994
rect 12058 11942 12070 11994
rect 12122 11942 19142 11994
rect 19194 11942 19206 11994
rect 19258 11942 19270 11994
rect 19322 11942 19334 11994
rect 19386 11942 22816 11994
rect 1104 11920 22816 11942
rect 2774 11840 2780 11892
rect 2832 11880 2838 11892
rect 3053 11883 3111 11889
rect 2832 11852 2877 11880
rect 2832 11840 2838 11852
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3234 11880 3240 11892
rect 3099 11852 3240 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3234 11840 3240 11852
rect 3292 11840 3298 11892
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 5810 11880 5816 11892
rect 4212 11852 5816 11880
rect 4212 11840 4218 11852
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6178 11840 6184 11892
rect 6236 11880 6242 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 6236 11852 6377 11880
rect 6236 11840 6242 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 6365 11843 6423 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 8018 11880 8024 11892
rect 7484 11852 8024 11880
rect 4338 11772 4344 11824
rect 4396 11812 4402 11824
rect 4396 11784 4752 11812
rect 4396 11772 4402 11784
rect 4724 11756 4752 11784
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11704 1458 11756
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3513 11747 3571 11753
rect 3513 11744 3525 11747
rect 3384 11716 3525 11744
rect 3384 11704 3390 11716
rect 3513 11713 3525 11716
rect 3559 11713 3571 11747
rect 3513 11707 3571 11713
rect 3697 11747 3755 11753
rect 3697 11713 3709 11747
rect 3743 11744 3755 11747
rect 4062 11744 4068 11756
rect 3743 11716 4068 11744
rect 3743 11713 3755 11716
rect 3697 11707 3755 11713
rect 4062 11704 4068 11716
rect 4120 11744 4126 11756
rect 4430 11744 4436 11756
rect 4120 11716 4436 11744
rect 4120 11704 4126 11716
rect 4430 11704 4436 11716
rect 4488 11704 4494 11756
rect 4706 11744 4712 11756
rect 4619 11716 4712 11744
rect 4706 11704 4712 11716
rect 4764 11704 4770 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 7484 11744 7512 11852
rect 8018 11840 8024 11852
rect 8076 11880 8082 11892
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8076 11852 9045 11880
rect 8076 11840 8082 11852
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 9033 11843 9091 11849
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 11241 11883 11299 11889
rect 9539 11852 11008 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 10980 11812 11008 11852
rect 11241 11849 11253 11883
rect 11287 11880 11299 11883
rect 11330 11880 11336 11892
rect 11287 11852 11336 11880
rect 11287 11849 11299 11852
rect 11241 11843 11299 11849
rect 11330 11840 11336 11852
rect 11388 11840 11394 11892
rect 13814 11880 13820 11892
rect 11440 11852 13584 11880
rect 13775 11852 13820 11880
rect 11440 11812 11468 11852
rect 10980 11784 11468 11812
rect 11977 11815 12035 11821
rect 11977 11781 11989 11815
rect 12023 11812 12035 11815
rect 12434 11812 12440 11824
rect 12023 11784 12440 11812
rect 12023 11781 12035 11784
rect 11977 11775 12035 11781
rect 12434 11772 12440 11784
rect 12492 11772 12498 11824
rect 7650 11744 7656 11756
rect 5868 11716 7512 11744
rect 7611 11716 7656 11744
rect 5868 11704 5874 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 9674 11704 9680 11756
rect 9732 11744 9738 11756
rect 9858 11744 9864 11756
rect 9732 11716 9864 11744
rect 9732 11704 9738 11716
rect 9858 11704 9864 11716
rect 9916 11704 9922 11756
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11480 11716 11836 11744
rect 11480 11704 11486 11716
rect 1664 11679 1722 11685
rect 1664 11645 1676 11679
rect 1710 11676 1722 11679
rect 2130 11676 2136 11688
rect 1710 11648 2136 11676
rect 1710 11645 1722 11648
rect 1664 11639 1722 11645
rect 2130 11636 2136 11648
rect 2188 11636 2194 11688
rect 3418 11676 3424 11688
rect 3379 11648 3424 11676
rect 3418 11636 3424 11648
rect 3476 11636 3482 11688
rect 4157 11679 4215 11685
rect 4157 11645 4169 11679
rect 4203 11676 4215 11679
rect 4246 11676 4252 11688
rect 4203 11648 4252 11676
rect 4203 11645 4215 11648
rect 4157 11639 4215 11645
rect 4246 11636 4252 11648
rect 4304 11636 4310 11688
rect 6549 11679 6607 11685
rect 6549 11645 6561 11679
rect 6595 11645 6607 11679
rect 7098 11676 7104 11688
rect 7059 11648 7104 11676
rect 6549 11639 6607 11645
rect 1854 11568 1860 11620
rect 1912 11608 1918 11620
rect 4798 11608 4804 11620
rect 1912 11580 4804 11608
rect 1912 11568 1918 11580
rect 4798 11568 4804 11580
rect 4856 11568 4862 11620
rect 4976 11611 5034 11617
rect 4976 11577 4988 11611
rect 5022 11608 5034 11611
rect 5626 11608 5632 11620
rect 5022 11580 5632 11608
rect 5022 11577 5034 11580
rect 4976 11571 5034 11577
rect 5626 11568 5632 11580
rect 5684 11568 5690 11620
rect 6564 11608 6592 11639
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 9122 11676 9128 11688
rect 7760 11648 9128 11676
rect 7760 11608 7788 11648
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11676 9367 11679
rect 9766 11676 9772 11688
rect 9355 11648 9772 11676
rect 9355 11645 9367 11648
rect 9309 11639 9367 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 11698 11676 11704 11688
rect 11659 11648 11704 11676
rect 11698 11636 11704 11648
rect 11756 11636 11762 11688
rect 11808 11685 11836 11716
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12710 11685 12716 11688
rect 12492 11648 12537 11676
rect 12492 11636 12498 11648
rect 12704 11639 12716 11685
rect 12768 11676 12774 11688
rect 12768 11648 12804 11676
rect 12710 11636 12716 11639
rect 12768 11636 12774 11648
rect 5736 11580 6224 11608
rect 6564 11580 7788 11608
rect 4341 11543 4399 11549
rect 4341 11509 4353 11543
rect 4387 11540 4399 11543
rect 4890 11540 4896 11552
rect 4387 11512 4896 11540
rect 4387 11509 4399 11512
rect 4341 11503 4399 11509
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5166 11500 5172 11552
rect 5224 11540 5230 11552
rect 5736 11540 5764 11580
rect 5224 11512 5764 11540
rect 5224 11500 5230 11512
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6089 11543 6147 11549
rect 6089 11540 6101 11543
rect 5960 11512 6101 11540
rect 5960 11500 5966 11512
rect 6089 11509 6101 11512
rect 6135 11509 6147 11543
rect 6196 11540 6224 11580
rect 7834 11568 7840 11620
rect 7892 11617 7898 11620
rect 10134 11617 10140 11620
rect 7892 11611 7956 11617
rect 7892 11577 7910 11611
rect 7944 11577 7956 11611
rect 10128 11608 10140 11617
rect 10047 11580 10140 11608
rect 7892 11571 7956 11577
rect 10128 11571 10140 11580
rect 10192 11608 10198 11620
rect 11054 11608 11060 11620
rect 10192 11580 11060 11608
rect 7892 11568 7898 11571
rect 10134 11568 10140 11571
rect 10192 11568 10198 11580
rect 11054 11568 11060 11580
rect 11112 11568 11118 11620
rect 13556 11608 13584 11852
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14274 11880 14280 11892
rect 14139 11852 14280 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14274 11840 14280 11852
rect 14332 11840 14338 11892
rect 15378 11840 15384 11892
rect 15436 11880 15442 11892
rect 18414 11880 18420 11892
rect 15436 11852 18420 11880
rect 15436 11840 15442 11852
rect 18414 11840 18420 11852
rect 18472 11840 18478 11892
rect 19978 11880 19984 11892
rect 19939 11852 19984 11880
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20714 11840 20720 11892
rect 20772 11880 20778 11892
rect 21729 11883 21787 11889
rect 21729 11880 21741 11883
rect 20772 11852 21741 11880
rect 20772 11840 20778 11852
rect 21729 11849 21741 11852
rect 21775 11849 21787 11883
rect 21729 11843 21787 11849
rect 15010 11772 15016 11824
rect 15068 11812 15074 11824
rect 15105 11815 15163 11821
rect 15105 11812 15117 11815
rect 15068 11784 15117 11812
rect 15068 11772 15074 11784
rect 15105 11781 15117 11784
rect 15151 11781 15163 11815
rect 16758 11812 16764 11824
rect 15105 11775 15163 11781
rect 15764 11784 16764 11812
rect 14918 11744 14924 11756
rect 14879 11716 14924 11744
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15764 11753 15792 11784
rect 16758 11772 16764 11784
rect 16816 11772 16822 11824
rect 21358 11772 21364 11824
rect 21416 11812 21422 11824
rect 22189 11815 22247 11821
rect 22189 11812 22201 11815
rect 21416 11784 22201 11812
rect 21416 11772 21422 11784
rect 22189 11781 22201 11784
rect 22235 11781 22247 11815
rect 22189 11775 22247 11781
rect 15565 11747 15623 11753
rect 15565 11744 15577 11747
rect 15528 11716 15577 11744
rect 15528 11704 15534 11716
rect 15565 11713 15577 11716
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 16577 11747 16635 11753
rect 16577 11713 16589 11747
rect 16623 11713 16635 11747
rect 17586 11744 17592 11756
rect 17547 11716 17592 11744
rect 16577 11707 16635 11713
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13780 11648 13921 11676
rect 13780 11636 13786 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 14458 11636 14464 11688
rect 14516 11676 14522 11688
rect 15010 11676 15016 11688
rect 14516 11648 15016 11676
rect 14516 11636 14522 11648
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 16393 11679 16451 11685
rect 16393 11645 16405 11679
rect 16439 11645 16451 11679
rect 16393 11639 16451 11645
rect 14645 11611 14703 11617
rect 14645 11608 14657 11611
rect 11532 11580 12112 11608
rect 13556 11580 14657 11608
rect 8018 11540 8024 11552
rect 6196 11512 8024 11540
rect 6089 11503 6147 11509
rect 8018 11500 8024 11512
rect 8076 11500 8082 11552
rect 11532 11549 11560 11580
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11509 11575 11543
rect 12084 11540 12112 11580
rect 14645 11577 14657 11580
rect 14691 11577 14703 11611
rect 14645 11571 14703 11577
rect 14737 11611 14795 11617
rect 14737 11577 14749 11611
rect 14783 11608 14795 11611
rect 14918 11608 14924 11620
rect 14783 11580 14924 11608
rect 14783 11577 14795 11580
rect 14737 11571 14795 11577
rect 14918 11568 14924 11580
rect 14976 11568 14982 11620
rect 15746 11608 15752 11620
rect 15304 11580 15752 11608
rect 12434 11540 12440 11552
rect 12084 11512 12440 11540
rect 11517 11503 11575 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 14277 11543 14335 11549
rect 14277 11509 14289 11543
rect 14323 11540 14335 11543
rect 15304 11540 15332 11580
rect 15746 11568 15752 11580
rect 15804 11568 15810 11620
rect 14323 11512 15332 11540
rect 14323 11509 14335 11512
rect 14277 11503 14335 11509
rect 15378 11500 15384 11552
rect 15436 11540 15442 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 15436 11512 15485 11540
rect 15436 11500 15442 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 15933 11543 15991 11549
rect 15933 11540 15945 11543
rect 15896 11512 15945 11540
rect 15896 11500 15902 11512
rect 15933 11509 15945 11512
rect 15979 11509 15991 11543
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 15933 11503 15991 11509
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16408 11540 16436 11639
rect 16592 11552 16620 11707
rect 17586 11704 17592 11716
rect 17644 11744 17650 11756
rect 17644 11716 18184 11744
rect 17644 11704 17650 11716
rect 17310 11676 17316 11688
rect 17271 11648 17316 11676
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18156 11676 18184 11716
rect 18305 11679 18363 11685
rect 18305 11676 18317 11679
rect 18156 11648 18317 11676
rect 18049 11639 18107 11645
rect 18305 11645 18317 11648
rect 18351 11645 18363 11679
rect 19794 11676 19800 11688
rect 19755 11648 19800 11676
rect 18305 11639 18363 11645
rect 17770 11608 17776 11620
rect 17328 11580 17776 11608
rect 17328 11552 17356 11580
rect 17770 11568 17776 11580
rect 17828 11608 17834 11620
rect 18064 11608 18092 11639
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19886 11636 19892 11688
rect 19944 11676 19950 11688
rect 20349 11679 20407 11685
rect 20349 11676 20361 11679
rect 19944 11648 20361 11676
rect 19944 11636 19950 11648
rect 20349 11645 20361 11648
rect 20395 11645 20407 11679
rect 20349 11639 20407 11645
rect 20438 11636 20444 11688
rect 20496 11676 20502 11688
rect 20605 11679 20663 11685
rect 20605 11676 20617 11679
rect 20496 11648 20617 11676
rect 20496 11636 20502 11648
rect 20605 11645 20617 11648
rect 20651 11645 20663 11679
rect 20605 11639 20663 11645
rect 22005 11679 22063 11685
rect 22005 11645 22017 11679
rect 22051 11645 22063 11679
rect 22005 11639 22063 11645
rect 17828 11580 18092 11608
rect 17828 11568 17834 11580
rect 18506 11568 18512 11620
rect 18564 11608 18570 11620
rect 22020 11608 22048 11639
rect 18564 11580 22048 11608
rect 18564 11568 18570 11580
rect 16482 11540 16488 11552
rect 16408 11512 16488 11540
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 16574 11500 16580 11552
rect 16632 11500 16638 11552
rect 16942 11540 16948 11552
rect 16903 11512 16948 11540
rect 16942 11500 16948 11512
rect 17000 11500 17006 11552
rect 17310 11500 17316 11552
rect 17368 11500 17374 11552
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 17460 11512 17505 11540
rect 17460 11500 17466 11512
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 19429 11543 19487 11549
rect 19429 11540 19441 11543
rect 18104 11512 19441 11540
rect 18104 11500 18110 11512
rect 19429 11509 19441 11512
rect 19475 11509 19487 11543
rect 19429 11503 19487 11509
rect 1104 11450 22816 11472
rect 1104 11398 8246 11450
rect 8298 11398 8310 11450
rect 8362 11398 8374 11450
rect 8426 11398 8438 11450
rect 8490 11398 15510 11450
rect 15562 11398 15574 11450
rect 15626 11398 15638 11450
rect 15690 11398 15702 11450
rect 15754 11398 22816 11450
rect 1104 11376 22816 11398
rect 1397 11339 1455 11345
rect 1397 11305 1409 11339
rect 1443 11336 1455 11339
rect 1578 11336 1584 11348
rect 1443 11308 1584 11336
rect 1443 11305 1455 11308
rect 1397 11299 1455 11305
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 1854 11336 1860 11348
rect 1815 11308 1860 11336
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 2409 11339 2467 11345
rect 2409 11305 2421 11339
rect 2455 11336 2467 11339
rect 2682 11336 2688 11348
rect 2455 11308 2688 11336
rect 2455 11305 2467 11308
rect 2409 11299 2467 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 2866 11336 2872 11348
rect 2823 11308 2872 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 5166 11336 5172 11348
rect 3344 11308 5172 11336
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 3344 11268 3372 11308
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 5258 11296 5264 11348
rect 5316 11336 5322 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 5316 11308 6285 11336
rect 5316 11296 5322 11308
rect 6273 11305 6285 11308
rect 6319 11305 6331 11339
rect 6273 11299 6331 11305
rect 6549 11339 6607 11345
rect 6549 11305 6561 11339
rect 6595 11336 6607 11339
rect 6822 11336 6828 11348
rect 6595 11308 6828 11336
rect 6595 11305 6607 11308
rect 6549 11299 6607 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 8570 11336 8576 11348
rect 7300 11308 8576 11336
rect 7300 11268 7328 11308
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 11054 11336 11060 11348
rect 9364 11308 9987 11336
rect 11015 11308 11060 11336
rect 9364 11296 9370 11308
rect 1811 11240 3372 11268
rect 3436 11240 7328 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 2314 11160 2320 11212
rect 2372 11200 2378 11212
rect 3436 11209 3464 11240
rect 7374 11228 7380 11280
rect 7432 11268 7438 11280
rect 7990 11271 8048 11277
rect 7990 11268 8002 11271
rect 7432 11240 8002 11268
rect 7432 11228 7438 11240
rect 7990 11237 8002 11240
rect 8036 11268 8048 11271
rect 8202 11268 8208 11280
rect 8036 11240 8208 11268
rect 8036 11237 8048 11240
rect 7990 11231 8048 11237
rect 8202 11228 8208 11240
rect 8260 11228 8266 11280
rect 9959 11277 9987 11308
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 12713 11339 12771 11345
rect 12713 11336 12725 11339
rect 12360 11308 12725 11336
rect 9944 11271 10002 11277
rect 9600 11240 9904 11268
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2372 11172 2881 11200
rect 2372 11160 2378 11172
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 2869 11163 2927 11169
rect 3421 11203 3479 11209
rect 3421 11169 3433 11203
rect 3467 11169 3479 11203
rect 4338 11200 4344 11212
rect 4299 11172 4344 11200
rect 3421 11163 3479 11169
rect 4338 11160 4344 11172
rect 4396 11160 4402 11212
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 4893 11203 4951 11209
rect 4893 11200 4905 11203
rect 4764 11172 4905 11200
rect 4764 11160 4770 11172
rect 4893 11169 4905 11172
rect 4939 11169 4951 11203
rect 4893 11163 4951 11169
rect 5160 11203 5218 11209
rect 5160 11169 5172 11203
rect 5206 11200 5218 11203
rect 5902 11200 5908 11212
rect 5206 11172 5908 11200
rect 5206 11169 5218 11172
rect 5160 11163 5218 11169
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2682 11132 2688 11144
rect 2087 11104 2688 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11132 3111 11135
rect 4430 11132 4436 11144
rect 3099 11104 4436 11132
rect 3099 11101 3111 11104
rect 3053 11095 3111 11101
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3605 11067 3663 11073
rect 3605 11064 3617 11067
rect 3476 11036 3617 11064
rect 3476 11024 3482 11036
rect 3605 11033 3617 11036
rect 3651 11033 3663 11067
rect 3605 11027 3663 11033
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 4212 11036 4537 11064
rect 4212 11024 4218 11036
rect 4525 11033 4537 11036
rect 4571 11033 4583 11067
rect 4525 11027 4583 11033
rect 4908 10996 4936 11163
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6914 11200 6920 11212
rect 6875 11172 6920 11200
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7098 11200 7104 11212
rect 7055 11172 7104 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 7650 11160 7656 11212
rect 7708 11200 7714 11212
rect 7745 11203 7803 11209
rect 7745 11200 7757 11203
rect 7708 11172 7757 11200
rect 7708 11160 7714 11172
rect 7745 11169 7757 11172
rect 7791 11169 7803 11203
rect 9600 11200 9628 11240
rect 7745 11163 7803 11169
rect 7852 11172 9628 11200
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7852 11132 7880 11172
rect 9674 11160 9680 11212
rect 9732 11200 9738 11212
rect 9876 11200 9904 11240
rect 9944 11237 9956 11271
rect 9990 11268 10002 11271
rect 12360 11268 12388 11308
rect 12713 11305 12725 11308
rect 12759 11305 12771 11339
rect 13998 11336 14004 11348
rect 12713 11299 12771 11305
rect 13096 11308 14004 11336
rect 9990 11240 12388 11268
rect 9990 11237 10002 11240
rect 9944 11231 10002 11237
rect 12526 11228 12532 11280
rect 12584 11268 12590 11280
rect 13096 11268 13124 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14182 11296 14188 11348
rect 14240 11336 14246 11348
rect 15013 11339 15071 11345
rect 15013 11336 15025 11339
rect 14240 11308 15025 11336
rect 14240 11296 14246 11308
rect 15013 11305 15025 11308
rect 15059 11305 15071 11339
rect 15013 11299 15071 11305
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 16632 11308 16773 11336
rect 16632 11296 16638 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17681 11339 17739 11345
rect 17681 11336 17693 11339
rect 17000 11308 17693 11336
rect 17000 11296 17006 11308
rect 17681 11305 17693 11308
rect 17727 11305 17739 11339
rect 19886 11336 19892 11348
rect 17681 11299 17739 11305
rect 19260 11308 19892 11336
rect 18138 11268 18144 11280
rect 12584 11240 13124 11268
rect 13188 11240 14136 11268
rect 12584 11228 12590 11240
rect 10686 11200 10692 11212
rect 9732 11172 9777 11200
rect 9876 11172 10692 11200
rect 9732 11160 9738 11172
rect 10686 11160 10692 11172
rect 10744 11160 10750 11212
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11422 11200 11428 11212
rect 11379 11172 11428 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 11422 11160 11428 11172
rect 11480 11160 11486 11212
rect 11606 11209 11612 11212
rect 11600 11200 11612 11209
rect 11567 11172 11612 11200
rect 11600 11163 11612 11172
rect 11606 11160 11612 11163
rect 11664 11160 11670 11212
rect 12342 11160 12348 11212
rect 12400 11200 12406 11212
rect 13188 11200 13216 11240
rect 12400 11172 13216 11200
rect 13256 11203 13314 11209
rect 12400 11160 12406 11172
rect 13256 11169 13268 11203
rect 13302 11200 13314 11203
rect 13722 11200 13728 11212
rect 13302 11172 13728 11200
rect 13302 11169 13314 11172
rect 13256 11163 13314 11169
rect 13722 11160 13728 11172
rect 13780 11160 13786 11212
rect 13998 11160 14004 11212
rect 14056 11160 14062 11212
rect 12986 11132 12992 11144
rect 7760 11104 7880 11132
rect 12947 11104 12992 11132
rect 6178 11024 6184 11076
rect 6236 11064 6242 11076
rect 7760 11064 7788 11104
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 14016 11064 14044 11160
rect 14108 11132 14136 11240
rect 14476 11240 18144 11268
rect 14476 11209 14504 11240
rect 18138 11228 18144 11240
rect 18196 11228 18202 11280
rect 18690 11228 18696 11280
rect 18748 11268 18754 11280
rect 19260 11268 19288 11308
rect 19886 11296 19892 11308
rect 19944 11336 19950 11348
rect 19944 11308 20484 11336
rect 19944 11296 19950 11308
rect 18748 11240 19288 11268
rect 18748 11228 18754 11240
rect 19702 11228 19708 11280
rect 19760 11268 19766 11280
rect 19760 11240 20208 11268
rect 19760 11228 19766 11240
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11169 14519 11203
rect 14461 11163 14519 11169
rect 14829 11203 14887 11209
rect 14829 11169 14841 11203
rect 14875 11200 14887 11203
rect 15102 11200 15108 11212
rect 14875 11172 15108 11200
rect 14875 11169 14887 11172
rect 14829 11163 14887 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 15648 11203 15706 11209
rect 15648 11169 15660 11203
rect 15694 11200 15706 11203
rect 15694 11172 16436 11200
rect 15694 11169 15706 11172
rect 15648 11163 15706 11169
rect 14108 11104 14688 11132
rect 14660 11076 14688 11104
rect 15378 11092 15384 11144
rect 15436 11132 15442 11144
rect 15436 11104 15481 11132
rect 15436 11092 15442 11104
rect 14642 11064 14648 11076
rect 6236 11036 7788 11064
rect 9048 11036 9352 11064
rect 14016 11036 14504 11064
rect 14555 11036 14648 11064
rect 6236 11024 6242 11036
rect 5074 10996 5080 11008
rect 4908 10968 5080 10996
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 5166 10956 5172 11008
rect 5224 10996 5230 11008
rect 9048 10996 9076 11036
rect 5224 10968 9076 10996
rect 9125 10999 9183 11005
rect 5224 10956 5230 10968
rect 9125 10965 9137 10999
rect 9171 10996 9183 10999
rect 9214 10996 9220 11008
rect 9171 10968 9220 10996
rect 9171 10965 9183 10968
rect 9125 10959 9183 10965
rect 9214 10956 9220 10968
rect 9272 10956 9278 11008
rect 9324 10996 9352 11036
rect 11238 10996 11244 11008
rect 9324 10968 11244 10996
rect 11238 10956 11244 10968
rect 11296 10956 11302 11008
rect 11330 10956 11336 11008
rect 11388 10996 11394 11008
rect 13998 10996 14004 11008
rect 11388 10968 14004 10996
rect 11388 10956 11394 10968
rect 13998 10956 14004 10968
rect 14056 10956 14062 11008
rect 14090 10956 14096 11008
rect 14148 10996 14154 11008
rect 14369 10999 14427 11005
rect 14369 10996 14381 10999
rect 14148 10968 14381 10996
rect 14148 10956 14154 10968
rect 14369 10965 14381 10968
rect 14415 10965 14427 10999
rect 14476 10996 14504 11036
rect 14642 11024 14648 11036
rect 14700 11024 14706 11076
rect 14918 11024 14924 11076
rect 14976 11064 14982 11076
rect 16408 11064 16436 11172
rect 16666 11160 16672 11212
rect 16724 11200 16730 11212
rect 17589 11203 17647 11209
rect 17589 11200 17601 11203
rect 16724 11172 17601 11200
rect 16724 11160 16730 11172
rect 17589 11169 17601 11172
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 18500 11203 18558 11209
rect 17828 11172 18184 11200
rect 17828 11160 17834 11172
rect 17865 11135 17923 11141
rect 17865 11101 17877 11135
rect 17911 11132 17923 11135
rect 18046 11132 18052 11144
rect 17911 11104 18052 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 18046 11092 18052 11104
rect 18104 11092 18110 11144
rect 18156 11132 18184 11172
rect 18500 11169 18512 11203
rect 18546 11200 18558 11203
rect 18782 11200 18788 11212
rect 18546 11172 18788 11200
rect 18546 11169 18558 11172
rect 18500 11163 18558 11169
rect 18782 11160 18788 11172
rect 18840 11160 18846 11212
rect 19794 11160 19800 11212
rect 19852 11200 19858 11212
rect 20180 11209 20208 11240
rect 20073 11203 20131 11209
rect 20073 11200 20085 11203
rect 19852 11172 20085 11200
rect 19852 11160 19858 11172
rect 20073 11169 20085 11172
rect 20119 11169 20131 11203
rect 20073 11163 20131 11169
rect 20165 11203 20223 11209
rect 20165 11169 20177 11203
rect 20211 11169 20223 11203
rect 20456 11200 20484 11308
rect 20806 11296 20812 11348
rect 20864 11336 20870 11348
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 20864 11308 22293 11336
rect 20864 11296 20870 11308
rect 22281 11305 22293 11308
rect 22327 11305 22339 11339
rect 22281 11299 22339 11305
rect 20714 11228 20720 11280
rect 20772 11268 20778 11280
rect 21146 11271 21204 11277
rect 21146 11268 21158 11271
rect 20772 11240 21158 11268
rect 20772 11228 20778 11240
rect 21146 11237 21158 11240
rect 21192 11237 21204 11271
rect 21146 11231 21204 11237
rect 20898 11200 20904 11212
rect 20456 11172 20904 11200
rect 20165 11163 20223 11169
rect 20898 11160 20904 11172
rect 20956 11160 20962 11212
rect 18233 11135 18291 11141
rect 18233 11132 18245 11135
rect 18156 11104 18245 11132
rect 18233 11101 18245 11104
rect 18279 11101 18291 11135
rect 18233 11095 18291 11101
rect 16482 11064 16488 11076
rect 14976 11036 15424 11064
rect 16408 11036 16488 11064
rect 14976 11024 14982 11036
rect 14550 10996 14556 11008
rect 14463 10968 14556 10996
rect 14369 10959 14427 10965
rect 14550 10956 14556 10968
rect 14608 10996 14614 11008
rect 15102 10996 15108 11008
rect 14608 10968 15108 10996
rect 14608 10956 14614 10968
rect 15102 10956 15108 10968
rect 15160 10956 15166 11008
rect 15396 10996 15424 11036
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 16850 10996 16856 11008
rect 15396 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17221 10999 17279 11005
rect 17221 10965 17233 10999
rect 17267 10996 17279 10999
rect 17310 10996 17316 11008
rect 17267 10968 17316 10996
rect 17267 10965 17279 10968
rect 17221 10959 17279 10965
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 17770 10956 17776 11008
rect 17828 10996 17834 11008
rect 19426 10996 19432 11008
rect 17828 10968 19432 10996
rect 17828 10956 17834 10968
rect 19426 10956 19432 10968
rect 19484 10956 19490 11008
rect 19610 10996 19616 11008
rect 19571 10968 19616 10996
rect 19610 10956 19616 10968
rect 19668 10956 19674 11008
rect 19702 10956 19708 11008
rect 19760 10996 19766 11008
rect 20349 10999 20407 11005
rect 20349 10996 20361 10999
rect 19760 10968 20361 10996
rect 19760 10956 19766 10968
rect 20349 10965 20361 10968
rect 20395 10965 20407 10999
rect 20349 10959 20407 10965
rect 1104 10906 22816 10928
rect 1104 10854 4614 10906
rect 4666 10854 4678 10906
rect 4730 10854 4742 10906
rect 4794 10854 4806 10906
rect 4858 10854 11878 10906
rect 11930 10854 11942 10906
rect 11994 10854 12006 10906
rect 12058 10854 12070 10906
rect 12122 10854 19142 10906
rect 19194 10854 19206 10906
rect 19258 10854 19270 10906
rect 19322 10854 19334 10906
rect 19386 10854 22816 10906
rect 1104 10832 22816 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2593 10795 2651 10801
rect 2593 10792 2605 10795
rect 2464 10764 2605 10792
rect 2464 10752 2470 10764
rect 2593 10761 2605 10764
rect 2639 10761 2651 10795
rect 2593 10755 2651 10761
rect 3510 10752 3516 10804
rect 3568 10792 3574 10804
rect 3605 10795 3663 10801
rect 3605 10792 3617 10795
rect 3568 10764 3617 10792
rect 3568 10752 3574 10764
rect 3605 10761 3617 10764
rect 3651 10761 3663 10795
rect 3605 10755 3663 10761
rect 4433 10795 4491 10801
rect 4433 10761 4445 10795
rect 4479 10792 4491 10795
rect 7101 10795 7159 10801
rect 4479 10764 7052 10792
rect 4479 10761 4491 10764
rect 4433 10755 4491 10761
rect 7024 10724 7052 10764
rect 7101 10761 7113 10795
rect 7147 10792 7159 10795
rect 7190 10792 7196 10804
rect 7147 10764 7196 10792
rect 7147 10761 7159 10764
rect 7101 10755 7159 10761
rect 7190 10752 7196 10764
rect 7248 10752 7254 10804
rect 8110 10792 8116 10804
rect 7484 10764 8116 10792
rect 7484 10724 7512 10764
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 8260 10764 8861 10792
rect 8260 10752 8266 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9766 10752 9772 10804
rect 9824 10792 9830 10804
rect 10965 10795 11023 10801
rect 10965 10792 10977 10795
rect 9824 10764 10977 10792
rect 9824 10752 9830 10764
rect 10965 10761 10977 10764
rect 11011 10761 11023 10795
rect 10965 10755 11023 10761
rect 12434 10752 12440 10804
rect 12492 10792 12498 10804
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 12492 10764 14841 10792
rect 12492 10752 12498 10764
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 14829 10755 14887 10761
rect 14936 10764 20361 10792
rect 7024 10696 7512 10724
rect 10226 10684 10232 10736
rect 10284 10724 10290 10736
rect 10505 10727 10563 10733
rect 10505 10724 10517 10727
rect 10284 10696 10517 10724
rect 10284 10684 10290 10696
rect 10505 10693 10517 10696
rect 10551 10693 10563 10727
rect 11977 10727 12035 10733
rect 11977 10724 11989 10727
rect 10505 10687 10563 10693
rect 10796 10696 11989 10724
rect 10796 10668 10824 10696
rect 11977 10693 11989 10696
rect 12023 10693 12035 10727
rect 14936 10724 14964 10764
rect 20349 10761 20361 10764
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 11977 10687 12035 10693
rect 14016 10696 14964 10724
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2866 10656 2872 10668
rect 2271 10628 2872 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2866 10616 2872 10628
rect 2924 10616 2930 10668
rect 3142 10656 3148 10668
rect 3103 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10616 3206 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 4065 10659 4123 10665
rect 4065 10656 4077 10659
rect 3844 10628 4077 10656
rect 3844 10616 3850 10628
rect 4065 10625 4077 10628
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 4249 10659 4307 10665
rect 4249 10625 4261 10659
rect 4295 10656 4307 10659
rect 4430 10656 4436 10668
rect 4295 10628 4436 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4430 10616 4436 10628
rect 4488 10616 4494 10668
rect 4540 10628 5203 10656
rect 1762 10548 1768 10600
rect 1820 10588 1826 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1820 10560 1961 10588
rect 1820 10548 1826 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 2041 10591 2099 10597
rect 2041 10557 2053 10591
rect 2087 10588 2099 10591
rect 2958 10588 2964 10600
rect 2087 10560 2964 10588
rect 2087 10557 2099 10560
rect 2041 10551 2099 10557
rect 2958 10548 2964 10560
rect 3016 10548 3022 10600
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10588 3111 10591
rect 3694 10588 3700 10600
rect 3099 10560 3700 10588
rect 3099 10557 3111 10560
rect 3053 10551 3111 10557
rect 3694 10548 3700 10560
rect 3752 10548 3758 10600
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3936 10560 3985 10588
rect 3936 10548 3942 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 3973 10551 4031 10557
rect 2590 10480 2596 10532
rect 2648 10520 2654 10532
rect 4540 10520 4568 10628
rect 5074 10588 5080 10600
rect 5035 10560 5080 10588
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 5175 10588 5203 10628
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 10778 10656 10784 10668
rect 10376 10628 10784 10656
rect 10376 10616 10382 10628
rect 10778 10616 10784 10628
rect 10836 10616 10842 10668
rect 11609 10659 11667 10665
rect 11609 10625 11621 10659
rect 11655 10656 11667 10659
rect 12342 10656 12348 10668
rect 11655 10628 12348 10656
rect 11655 10625 11667 10628
rect 11609 10619 11667 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 5175 10560 5488 10588
rect 2648 10492 4568 10520
rect 4617 10523 4675 10529
rect 2648 10480 2654 10492
rect 4617 10489 4629 10523
rect 4663 10520 4675 10523
rect 5166 10520 5172 10532
rect 4663 10492 5172 10520
rect 4663 10489 4675 10492
rect 4617 10483 4675 10489
rect 5166 10480 5172 10492
rect 5224 10480 5230 10532
rect 5258 10480 5264 10532
rect 5316 10529 5322 10532
rect 5316 10523 5380 10529
rect 5316 10489 5334 10523
rect 5368 10489 5380 10523
rect 5460 10520 5488 10560
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6086 10588 6092 10600
rect 5868 10560 6092 10588
rect 5868 10548 5874 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7006 10588 7012 10600
rect 6963 10560 7012 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 7469 10591 7527 10597
rect 7469 10557 7481 10591
rect 7515 10588 7527 10591
rect 7558 10588 7564 10600
rect 7515 10560 7564 10588
rect 7515 10557 7527 10560
rect 7469 10551 7527 10557
rect 7558 10548 7564 10560
rect 7616 10548 7622 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 7668 10560 8953 10588
rect 7668 10520 7696 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9766 10588 9772 10600
rect 9171 10560 9772 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9766 10548 9772 10560
rect 9824 10548 9830 10600
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 11330 10588 11336 10600
rect 9916 10560 11336 10588
rect 9916 10548 9922 10560
rect 11330 10548 11336 10560
rect 11388 10548 11394 10600
rect 12158 10588 12164 10600
rect 12119 10560 12164 10588
rect 12158 10548 12164 10560
rect 12216 10548 12222 10600
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 12483 10560 12909 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 12986 10548 12992 10600
rect 13044 10588 13050 10600
rect 14016 10588 14044 10696
rect 15102 10684 15108 10736
rect 15160 10724 15166 10736
rect 17402 10724 17408 10736
rect 15160 10696 15608 10724
rect 17363 10696 17408 10724
rect 15160 10684 15166 10696
rect 14826 10616 14832 10668
rect 14884 10656 14890 10668
rect 15580 10665 15608 10696
rect 17402 10684 17408 10696
rect 17460 10684 17466 10736
rect 15565 10659 15623 10665
rect 14884 10628 15424 10656
rect 14884 10616 14890 10628
rect 13044 10560 13089 10588
rect 13188 10560 14044 10588
rect 14645 10591 14703 10597
rect 13044 10548 13050 10560
rect 5460 10492 7696 10520
rect 7736 10523 7794 10529
rect 5316 10483 5380 10489
rect 7736 10489 7748 10523
rect 7782 10489 7794 10523
rect 7736 10483 7794 10489
rect 5316 10480 5322 10483
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 2406 10452 2412 10464
rect 1627 10424 2412 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 2406 10412 2412 10424
rect 2464 10412 2470 10464
rect 2961 10455 3019 10461
rect 2961 10421 2973 10455
rect 3007 10452 3019 10455
rect 3970 10452 3976 10464
rect 3007 10424 3976 10452
rect 3007 10421 3019 10424
rect 2961 10415 3019 10421
rect 3970 10412 3976 10424
rect 4028 10412 4034 10464
rect 4430 10452 4436 10464
rect 4391 10424 4436 10452
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5442 10452 5448 10464
rect 5132 10424 5448 10452
rect 5132 10412 5138 10424
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5626 10412 5632 10464
rect 5684 10452 5690 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5684 10424 6469 10452
rect 5684 10412 5690 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6822 10412 6828 10464
rect 6880 10452 6886 10464
rect 7760 10452 7788 10483
rect 8018 10480 8024 10532
rect 8076 10520 8082 10532
rect 9214 10520 9220 10532
rect 8076 10492 9220 10520
rect 8076 10480 8082 10492
rect 9214 10480 9220 10492
rect 9272 10520 9278 10532
rect 9370 10523 9428 10529
rect 9370 10520 9382 10523
rect 9272 10492 9382 10520
rect 9272 10480 9278 10492
rect 9370 10489 9382 10492
rect 9416 10489 9428 10523
rect 13188 10520 13216 10560
rect 14645 10557 14657 10591
rect 14691 10588 14703 10591
rect 15286 10588 15292 10600
rect 14691 10560 15292 10588
rect 14691 10557 14703 10560
rect 14645 10551 14703 10557
rect 15286 10548 15292 10560
rect 15344 10548 15350 10600
rect 15396 10597 15424 10628
rect 15565 10625 15577 10659
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 15838 10616 15844 10668
rect 15896 10656 15902 10668
rect 16028 10659 16086 10665
rect 16028 10656 16040 10659
rect 15896 10628 16040 10656
rect 15896 10616 15902 10628
rect 16028 10625 16040 10628
rect 16074 10625 16086 10659
rect 17420 10656 17448 10684
rect 18555 10659 18613 10665
rect 16028 10619 16086 10625
rect 16224 10628 17364 10656
rect 17420 10628 18184 10656
rect 15381 10591 15439 10597
rect 15381 10557 15393 10591
rect 15427 10557 15439 10591
rect 16224 10588 16252 10628
rect 15381 10551 15439 10557
rect 15672 10560 16252 10588
rect 16301 10591 16359 10597
rect 9370 10483 9428 10489
rect 9508 10492 13216 10520
rect 13256 10523 13314 10529
rect 8754 10452 8760 10464
rect 6880 10424 8760 10452
rect 6880 10412 6886 10424
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8941 10455 8999 10461
rect 8941 10421 8953 10455
rect 8987 10452 8999 10455
rect 9508 10452 9536 10492
rect 13256 10489 13268 10523
rect 13302 10520 13314 10523
rect 14090 10520 14096 10532
rect 13302 10492 14096 10520
rect 13302 10489 13314 10492
rect 13256 10483 13314 10489
rect 14090 10480 14096 10492
rect 14148 10480 14154 10532
rect 15672 10520 15700 10560
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 16758 10588 16764 10600
rect 16347 10560 16764 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 16758 10548 16764 10560
rect 16816 10548 16822 10600
rect 14200 10492 15700 10520
rect 17336 10520 17364 10628
rect 17402 10548 17408 10600
rect 17460 10588 17466 10600
rect 17865 10591 17923 10597
rect 17865 10588 17877 10591
rect 17460 10560 17877 10588
rect 17460 10548 17466 10560
rect 17865 10557 17877 10560
rect 17911 10557 17923 10591
rect 18046 10588 18052 10600
rect 18007 10560 18052 10588
rect 17865 10551 17923 10557
rect 18046 10548 18052 10560
rect 18104 10548 18110 10600
rect 18156 10588 18184 10628
rect 18555 10625 18567 10659
rect 18601 10656 18613 10659
rect 18966 10656 18972 10668
rect 18601 10628 18972 10656
rect 18601 10625 18613 10628
rect 18555 10619 18613 10625
rect 18966 10616 18972 10628
rect 19024 10616 19030 10668
rect 20898 10656 20904 10668
rect 20859 10628 20904 10656
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 18785 10591 18843 10597
rect 18785 10588 18797 10591
rect 18156 10560 18797 10588
rect 18785 10557 18797 10560
rect 18831 10557 18843 10591
rect 20162 10588 20168 10600
rect 20123 10560 20168 10588
rect 18785 10551 18843 10557
rect 20162 10548 20168 10560
rect 20220 10548 20226 10600
rect 17336 10492 18184 10520
rect 8987 10424 9536 10452
rect 8987 10421 8999 10424
rect 8941 10415 8999 10421
rect 9582 10412 9588 10464
rect 9640 10452 9646 10464
rect 11333 10455 11391 10461
rect 11333 10452 11345 10455
rect 9640 10424 11345 10452
rect 9640 10412 9646 10424
rect 11333 10421 11345 10424
rect 11379 10421 11391 10455
rect 11333 10415 11391 10421
rect 11422 10412 11428 10464
rect 11480 10452 11486 10464
rect 11480 10424 11525 10452
rect 11480 10412 11486 10424
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 11756 10424 12633 10452
rect 11756 10412 11762 10424
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 12897 10455 12955 10461
rect 12897 10421 12909 10455
rect 12943 10452 12955 10455
rect 14200 10452 14228 10492
rect 14366 10452 14372 10464
rect 12943 10424 14228 10452
rect 14327 10424 14372 10452
rect 12943 10421 12955 10424
rect 12897 10415 12955 10421
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15194 10452 15200 10464
rect 15155 10424 15200 10452
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15930 10412 15936 10464
rect 15988 10452 15994 10464
rect 16031 10455 16089 10461
rect 16031 10452 16043 10455
rect 15988 10424 16043 10452
rect 15988 10412 15994 10424
rect 16031 10421 16043 10424
rect 16077 10421 16089 10455
rect 16031 10415 16089 10421
rect 16574 10412 16580 10464
rect 16632 10452 16638 10464
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 16632 10424 17693 10452
rect 16632 10412 16638 10424
rect 17681 10421 17693 10424
rect 17727 10421 17739 10455
rect 18156 10452 18184 10492
rect 20806 10480 20812 10532
rect 20864 10520 20870 10532
rect 21146 10523 21204 10529
rect 21146 10520 21158 10523
rect 20864 10492 21158 10520
rect 20864 10480 20870 10492
rect 21146 10489 21158 10492
rect 21192 10489 21204 10523
rect 21146 10483 21204 10489
rect 18414 10452 18420 10464
rect 18156 10424 18420 10452
rect 17681 10415 17739 10421
rect 18414 10412 18420 10424
rect 18472 10412 18478 10464
rect 18515 10455 18573 10461
rect 18515 10421 18527 10455
rect 18561 10452 18573 10455
rect 18690 10452 18696 10464
rect 18561 10424 18696 10452
rect 18561 10421 18573 10424
rect 18515 10415 18573 10421
rect 18690 10412 18696 10424
rect 18748 10412 18754 10464
rect 19058 10412 19064 10464
rect 19116 10452 19122 10464
rect 19889 10455 19947 10461
rect 19889 10452 19901 10455
rect 19116 10424 19901 10452
rect 19116 10412 19122 10424
rect 19889 10421 19901 10424
rect 19935 10452 19947 10455
rect 20530 10452 20536 10464
rect 19935 10424 20536 10452
rect 19935 10421 19947 10424
rect 19889 10415 19947 10421
rect 20530 10412 20536 10424
rect 20588 10412 20594 10464
rect 22278 10452 22284 10464
rect 22239 10424 22284 10452
rect 22278 10412 22284 10424
rect 22336 10412 22342 10464
rect 1104 10362 22816 10384
rect 1104 10310 8246 10362
rect 8298 10310 8310 10362
rect 8362 10310 8374 10362
rect 8426 10310 8438 10362
rect 8490 10310 15510 10362
rect 15562 10310 15574 10362
rect 15626 10310 15638 10362
rect 15690 10310 15702 10362
rect 15754 10310 22816 10362
rect 1104 10288 22816 10310
rect 1949 10251 2007 10257
rect 1949 10217 1961 10251
rect 1995 10248 2007 10251
rect 4246 10248 4252 10260
rect 1995 10220 4252 10248
rect 1995 10217 2007 10220
rect 1949 10211 2007 10217
rect 4246 10208 4252 10220
rect 4304 10208 4310 10260
rect 5350 10248 5356 10260
rect 5311 10220 5356 10248
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5442 10208 5448 10260
rect 5500 10248 5506 10260
rect 5721 10251 5779 10257
rect 5721 10248 5733 10251
rect 5500 10220 5733 10248
rect 5500 10208 5506 10220
rect 5721 10217 5733 10220
rect 5767 10217 5779 10251
rect 5721 10211 5779 10217
rect 5813 10251 5871 10257
rect 5813 10217 5825 10251
rect 5859 10248 5871 10251
rect 6546 10248 6552 10260
rect 5859 10220 6552 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7834 10208 7840 10260
rect 7892 10208 7898 10260
rect 8570 10208 8576 10260
rect 8628 10248 8634 10260
rect 10502 10248 10508 10260
rect 8628 10220 10508 10248
rect 8628 10208 8634 10220
rect 10502 10208 10508 10220
rect 10560 10248 10566 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 10560 10220 13369 10248
rect 10560 10208 10566 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 14090 10248 14096 10260
rect 14051 10220 14096 10248
rect 13357 10211 13415 10217
rect 14090 10208 14096 10220
rect 14148 10208 14154 10260
rect 16482 10208 16488 10260
rect 16540 10248 16546 10260
rect 16669 10251 16727 10257
rect 16669 10248 16681 10251
rect 16540 10220 16681 10248
rect 16540 10208 16546 10220
rect 16669 10217 16681 10220
rect 16715 10217 16727 10251
rect 16669 10211 16727 10217
rect 16850 10208 16856 10260
rect 16908 10248 16914 10260
rect 17129 10251 17187 10257
rect 17129 10248 17141 10251
rect 16908 10220 17141 10248
rect 16908 10208 16914 10220
rect 17129 10217 17141 10220
rect 17175 10217 17187 10251
rect 17129 10211 17187 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18049 10251 18107 10257
rect 18049 10248 18061 10251
rect 18012 10220 18061 10248
rect 18012 10208 18018 10220
rect 18049 10217 18061 10220
rect 18095 10217 18107 10251
rect 18049 10211 18107 10217
rect 18601 10251 18659 10257
rect 18601 10217 18613 10251
rect 18647 10248 18659 10251
rect 18874 10248 18880 10260
rect 18647 10220 18880 10248
rect 18647 10217 18659 10220
rect 18601 10211 18659 10217
rect 18874 10208 18880 10220
rect 18932 10208 18938 10260
rect 19058 10248 19064 10260
rect 19019 10220 19064 10248
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19150 10208 19156 10260
rect 19208 10248 19214 10260
rect 20073 10251 20131 10257
rect 20073 10248 20085 10251
rect 19208 10220 20085 10248
rect 19208 10208 19214 10220
rect 20073 10217 20085 10220
rect 20119 10217 20131 10251
rect 20073 10211 20131 10217
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10180 3479 10183
rect 4890 10180 4896 10192
rect 3467 10152 4896 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 4890 10140 4896 10152
rect 4948 10140 4954 10192
rect 4982 10140 4988 10192
rect 5040 10180 5046 10192
rect 5261 10183 5319 10189
rect 5261 10180 5273 10183
rect 5040 10152 5273 10180
rect 5040 10140 5046 10152
rect 5261 10149 5273 10152
rect 5307 10149 5319 10183
rect 7852 10180 7880 10208
rect 11422 10180 11428 10192
rect 5261 10143 5319 10149
rect 5368 10152 7880 10180
rect 8763 10152 11428 10180
rect 2317 10115 2375 10121
rect 2317 10081 2329 10115
rect 2363 10112 2375 10115
rect 3050 10112 3056 10124
rect 2363 10084 3056 10112
rect 2363 10081 2375 10084
rect 2317 10075 2375 10081
rect 3050 10072 3056 10084
rect 3108 10072 3114 10124
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 4341 10115 4399 10121
rect 3375 10084 4292 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10013 1547 10047
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 1489 10007 1547 10013
rect 1504 9976 1532 10007
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 2590 10044 2596 10056
rect 2551 10016 2596 10044
rect 2590 10004 2596 10016
rect 2648 10004 2654 10056
rect 2682 10004 2688 10056
rect 2740 10044 2746 10056
rect 3605 10047 3663 10053
rect 3605 10044 3617 10047
rect 2740 10016 3617 10044
rect 2740 10004 2746 10016
rect 3605 10013 3617 10016
rect 3651 10044 3663 10047
rect 3786 10044 3792 10056
rect 3651 10016 3792 10044
rect 3651 10013 3663 10016
rect 3605 10007 3663 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4264 10044 4292 10084
rect 4341 10081 4353 10115
rect 4387 10112 4399 10115
rect 4430 10112 4436 10124
rect 4387 10084 4436 10112
rect 4387 10081 4399 10084
rect 4341 10075 4399 10081
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 5368 10044 5396 10152
rect 6178 10121 6184 10124
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 5905 10115 5963 10121
rect 5905 10112 5917 10115
rect 5767 10084 5917 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 5905 10081 5917 10084
rect 5951 10081 5963 10115
rect 5905 10075 5963 10081
rect 6172 10075 6184 10121
rect 6236 10112 6242 10124
rect 7558 10112 7564 10124
rect 6236 10084 6272 10112
rect 7519 10084 7564 10112
rect 6178 10072 6184 10075
rect 6236 10072 6242 10084
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 7817 10115 7875 10121
rect 7817 10112 7829 10115
rect 7668 10084 7829 10112
rect 4264 10016 5396 10044
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 5537 10047 5595 10053
rect 5537 10044 5549 10047
rect 5500 10016 5549 10044
rect 5500 10004 5506 10016
rect 5537 10013 5549 10016
rect 5583 10044 5595 10047
rect 5813 10047 5871 10053
rect 5813 10044 5825 10047
rect 5583 10016 5825 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5813 10013 5825 10016
rect 5859 10013 5871 10047
rect 7668 10044 7696 10084
rect 7817 10081 7829 10084
rect 7863 10081 7875 10115
rect 7817 10075 7875 10081
rect 8386 10072 8392 10124
rect 8444 10112 8450 10124
rect 8763 10112 8791 10152
rect 11422 10140 11428 10152
rect 11480 10140 11486 10192
rect 14001 10183 14059 10189
rect 14001 10180 14013 10183
rect 11532 10152 14013 10180
rect 9398 10112 9404 10124
rect 8444 10084 8791 10112
rect 9359 10084 9404 10112
rect 8444 10072 8450 10084
rect 9398 10072 9404 10084
rect 9456 10072 9462 10124
rect 9766 10112 9772 10124
rect 9727 10084 9772 10112
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 10318 10112 10324 10124
rect 10279 10084 10324 10112
rect 10318 10072 10324 10084
rect 10376 10072 10382 10124
rect 10594 10121 10600 10124
rect 10588 10112 10600 10121
rect 10555 10084 10600 10112
rect 10588 10075 10600 10084
rect 10594 10072 10600 10075
rect 10652 10072 10658 10124
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 11532 10112 11560 10152
rect 14001 10149 14013 10152
rect 14047 10180 14059 10183
rect 14366 10180 14372 10192
rect 14047 10152 14372 10180
rect 14047 10149 14059 10152
rect 14001 10143 14059 10149
rect 14366 10140 14372 10152
rect 14424 10140 14430 10192
rect 19334 10180 19340 10192
rect 14660 10152 19340 10180
rect 14660 10121 14688 10152
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 21146 10183 21204 10189
rect 21146 10180 21158 10183
rect 19904 10152 21158 10180
rect 12233 10115 12291 10121
rect 12233 10112 12245 10115
rect 10928 10084 11560 10112
rect 11593 10084 12245 10112
rect 10928 10072 10934 10084
rect 5813 10007 5871 10013
rect 7576 10016 7696 10044
rect 1854 9976 1860 9988
rect 1504 9948 1860 9976
rect 1854 9936 1860 9948
rect 1912 9936 1918 9988
rect 2961 9979 3019 9985
rect 2961 9945 2973 9979
rect 3007 9976 3019 9979
rect 4062 9976 4068 9988
rect 3007 9948 4068 9976
rect 3007 9945 3019 9948
rect 2961 9939 3019 9945
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4893 9979 4951 9985
rect 4893 9945 4905 9979
rect 4939 9976 4951 9979
rect 5718 9976 5724 9988
rect 4939 9948 5724 9976
rect 4939 9945 4951 9948
rect 4893 9939 4951 9945
rect 5718 9936 5724 9948
rect 5776 9936 5782 9988
rect 7576 9976 7604 10016
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 10226 10044 10232 10056
rect 9272 10016 10232 10044
rect 9272 10004 9278 10016
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 11330 10004 11336 10056
rect 11388 10044 11394 10056
rect 11593 10044 11621 10084
rect 12233 10081 12245 10084
rect 12279 10081 12291 10115
rect 12233 10075 12291 10081
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10081 14703 10115
rect 15286 10112 15292 10124
rect 15247 10084 15292 10112
rect 14645 10075 14703 10081
rect 15286 10072 15292 10084
rect 15344 10072 15350 10124
rect 15378 10072 15384 10124
rect 15436 10072 15442 10124
rect 15556 10115 15614 10121
rect 15556 10081 15568 10115
rect 15602 10112 15614 10115
rect 16850 10112 16856 10124
rect 15602 10084 16856 10112
rect 15602 10081 15614 10084
rect 15556 10075 15614 10081
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 17957 10115 18015 10121
rect 17957 10081 17969 10115
rect 18003 10112 18015 10115
rect 18966 10112 18972 10124
rect 18003 10084 18184 10112
rect 18927 10084 18972 10112
rect 18003 10081 18015 10084
rect 17957 10075 18015 10081
rect 11388 10016 11621 10044
rect 11977 10047 12035 10053
rect 11388 10004 11394 10016
rect 11977 10013 11989 10047
rect 12023 10013 12035 10047
rect 14182 10044 14188 10056
rect 14143 10016 14188 10044
rect 11977 10007 12035 10013
rect 7300 9948 7604 9976
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3694 9908 3700 9920
rect 2924 9880 3700 9908
rect 2924 9868 2930 9880
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 4525 9911 4583 9917
rect 4525 9877 4537 9911
rect 4571 9908 4583 9911
rect 5350 9908 5356 9920
rect 4571 9880 5356 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 7300 9917 7328 9948
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8812 9948 8953 9976
rect 8812 9936 8818 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 9858 9976 9864 9988
rect 8941 9939 8999 9945
rect 9048 9948 9864 9976
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 6144 9880 7297 9908
rect 6144 9868 6150 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7466 9868 7472 9920
rect 7524 9908 7530 9920
rect 9048 9908 9076 9948
rect 9858 9936 9864 9948
rect 9916 9936 9922 9988
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10100 9948 10364 9976
rect 10100 9936 10106 9948
rect 7524 9880 9076 9908
rect 7524 9868 7530 9880
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 9180 9880 9229 9908
rect 9180 9868 9186 9880
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9217 9871 9275 9877
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10226 9908 10232 9920
rect 9999 9880 10232 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10226 9868 10232 9880
rect 10284 9868 10290 9920
rect 10336 9908 10364 9948
rect 11514 9936 11520 9988
rect 11572 9976 11578 9988
rect 11992 9976 12020 10007
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 15396 10044 15424 10072
rect 14292 10016 15424 10044
rect 14292 9976 14320 10016
rect 11572 9948 12020 9976
rect 11572 9936 11578 9948
rect 11606 9908 11612 9920
rect 10336 9880 11612 9908
rect 11606 9868 11612 9880
rect 11664 9908 11670 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 11664 9880 11713 9908
rect 11664 9868 11670 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11992 9908 12020 9948
rect 12912 9948 14320 9976
rect 14829 9979 14887 9985
rect 12912 9920 12940 9948
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 15102 9976 15108 9988
rect 14875 9948 15108 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 15102 9936 15108 9948
rect 15160 9936 15166 9988
rect 12250 9908 12256 9920
rect 11992 9880 12256 9908
rect 11701 9871 11759 9877
rect 12250 9868 12256 9880
rect 12308 9868 12314 9920
rect 12894 9868 12900 9920
rect 12952 9868 12958 9920
rect 13633 9911 13691 9917
rect 13633 9877 13645 9911
rect 13679 9908 13691 9911
rect 14734 9908 14740 9920
rect 13679 9880 14740 9908
rect 13679 9877 13691 9880
rect 13633 9871 13691 9877
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 16960 9908 16988 10075
rect 18156 9976 18184 10084
rect 18966 10072 18972 10084
rect 19024 10072 19030 10124
rect 19904 10112 19932 10152
rect 21146 10149 21158 10152
rect 21192 10180 21204 10183
rect 22278 10180 22284 10192
rect 21192 10152 22284 10180
rect 21192 10149 21204 10152
rect 21146 10143 21204 10149
rect 22278 10140 22284 10152
rect 22336 10140 22342 10192
rect 19076 10084 19932 10112
rect 18233 10047 18291 10053
rect 18233 10013 18245 10047
rect 18279 10044 18291 10047
rect 19076 10044 19104 10084
rect 19978 10072 19984 10124
rect 20036 10112 20042 10124
rect 20898 10112 20904 10124
rect 20036 10084 20081 10112
rect 20859 10084 20904 10112
rect 20036 10072 20042 10084
rect 20898 10072 20904 10084
rect 20956 10072 20962 10124
rect 18279 10016 19104 10044
rect 19153 10047 19211 10053
rect 18279 10013 18291 10016
rect 18233 10007 18291 10013
rect 19153 10013 19165 10047
rect 19199 10013 19211 10047
rect 20162 10044 20168 10056
rect 20123 10016 20168 10044
rect 19153 10007 19211 10013
rect 18156 9948 18276 9976
rect 14976 9880 16988 9908
rect 17589 9911 17647 9917
rect 14976 9868 14982 9880
rect 17589 9877 17601 9911
rect 17635 9908 17647 9911
rect 18138 9908 18144 9920
rect 17635 9880 18144 9908
rect 17635 9877 17647 9880
rect 17589 9871 17647 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 18248 9908 18276 9948
rect 18782 9936 18788 9988
rect 18840 9976 18846 9988
rect 19168 9976 19196 10007
rect 20162 10004 20168 10016
rect 20220 10004 20226 10056
rect 19702 9976 19708 9988
rect 18840 9948 19196 9976
rect 19260 9948 19708 9976
rect 18840 9936 18846 9948
rect 19260 9908 19288 9948
rect 19702 9936 19708 9948
rect 19760 9936 19766 9988
rect 18248 9880 19288 9908
rect 19518 9868 19524 9920
rect 19576 9908 19582 9920
rect 19613 9911 19671 9917
rect 19613 9908 19625 9911
rect 19576 9880 19625 9908
rect 19576 9868 19582 9880
rect 19613 9877 19625 9880
rect 19659 9908 19671 9911
rect 19886 9908 19892 9920
rect 19659 9880 19892 9908
rect 19659 9877 19671 9880
rect 19613 9871 19671 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 22278 9908 22284 9920
rect 22239 9880 22284 9908
rect 22278 9868 22284 9880
rect 22336 9868 22342 9920
rect 1104 9818 22816 9840
rect 1104 9766 4614 9818
rect 4666 9766 4678 9818
rect 4730 9766 4742 9818
rect 4794 9766 4806 9818
rect 4858 9766 11878 9818
rect 11930 9766 11942 9818
rect 11994 9766 12006 9818
rect 12058 9766 12070 9818
rect 12122 9766 19142 9818
rect 19194 9766 19206 9818
rect 19258 9766 19270 9818
rect 19322 9766 19334 9818
rect 19386 9766 22816 9818
rect 1104 9744 22816 9766
rect 2406 9664 2412 9716
rect 2464 9704 2470 9716
rect 9766 9704 9772 9716
rect 2464 9676 9772 9704
rect 2464 9664 2470 9676
rect 9766 9664 9772 9676
rect 9824 9664 9830 9716
rect 10244 9676 11192 9704
rect 2041 9639 2099 9645
rect 2041 9605 2053 9639
rect 2087 9636 2099 9639
rect 4338 9636 4344 9648
rect 2087 9608 4344 9636
rect 2087 9605 2099 9608
rect 2041 9599 2099 9605
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 7193 9639 7251 9645
rect 7193 9605 7205 9639
rect 7239 9636 7251 9639
rect 9217 9639 9275 9645
rect 7239 9608 9168 9636
rect 7239 9605 7251 9608
rect 7193 9599 7251 9605
rect 2498 9568 2504 9580
rect 2459 9540 2504 9568
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 2682 9568 2688 9580
rect 2643 9540 2688 9568
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 3694 9568 3700 9580
rect 3655 9540 3700 9568
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 4709 9571 4767 9577
rect 4709 9568 4721 9571
rect 3844 9540 4721 9568
rect 3844 9528 3850 9540
rect 4709 9537 4721 9540
rect 4755 9537 4767 9571
rect 5074 9568 5080 9580
rect 5035 9540 5080 9568
rect 4709 9531 4767 9537
rect 1578 9500 1584 9512
rect 1539 9472 1584 9500
rect 1578 9460 1584 9472
rect 1636 9460 1642 9512
rect 2038 9460 2044 9512
rect 2096 9500 2102 9512
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2096 9472 2421 9500
rect 2096 9460 2102 9472
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 3418 9500 3424 9512
rect 3379 9472 3424 9500
rect 2409 9463 2467 9469
rect 3418 9460 3424 9472
rect 3476 9460 3482 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9500 3571 9503
rect 4154 9500 4160 9512
rect 3559 9472 4160 9500
rect 3559 9469 3571 9472
rect 3513 9463 3571 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4724 9500 4752 9531
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8849 9571 8907 9577
rect 7883 9540 8708 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 4982 9500 4988 9512
rect 4724 9472 4988 9500
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 5344 9503 5402 9509
rect 5344 9469 5356 9503
rect 5390 9500 5402 9503
rect 5626 9500 5632 9512
rect 5390 9472 5632 9500
rect 5390 9469 5402 9472
rect 5344 9463 5402 9469
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 5359 9432 5387 9463
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 6270 9500 6276 9512
rect 5776 9472 6276 9500
rect 5776 9460 5782 9472
rect 6270 9460 6276 9472
rect 6328 9460 6334 9512
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9500 8171 9503
rect 8386 9500 8392 9512
rect 8159 9472 8392 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 8386 9460 8392 9472
rect 8444 9460 8450 9512
rect 8570 9500 8576 9512
rect 8531 9472 8576 9500
rect 8570 9460 8576 9472
rect 8628 9460 8634 9512
rect 8680 9500 8708 9540
rect 8849 9537 8861 9571
rect 8895 9537 8907 9571
rect 9140 9568 9168 9608
rect 9217 9605 9229 9639
rect 9263 9636 9275 9639
rect 9582 9636 9588 9648
rect 9263 9608 9588 9636
rect 9263 9605 9275 9608
rect 9217 9599 9275 9605
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10244 9636 10272 9676
rect 9784 9608 10272 9636
rect 11164 9636 11192 9676
rect 11238 9664 11244 9716
rect 11296 9704 11302 9716
rect 12894 9704 12900 9716
rect 11296 9676 12900 9704
rect 11296 9664 11302 9676
rect 12894 9664 12900 9676
rect 12952 9664 12958 9716
rect 13096 9676 14136 9704
rect 13096 9648 13124 9676
rect 11164 9608 13032 9636
rect 9784 9568 9812 9608
rect 9140 9540 9812 9568
rect 8849 9531 8907 9537
rect 8864 9500 8892 9531
rect 9858 9528 9864 9580
rect 9916 9568 9922 9580
rect 10134 9568 10140 9580
rect 9916 9540 10140 9568
rect 9916 9528 9922 9540
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 11480 9540 12817 9568
rect 11480 9528 11486 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 13004 9568 13032 9608
rect 13078 9596 13084 9648
rect 13136 9596 13142 9648
rect 14108 9636 14136 9676
rect 14752 9676 15056 9704
rect 14752 9636 14780 9676
rect 14108 9608 14780 9636
rect 14829 9639 14887 9645
rect 14829 9605 14841 9639
rect 14875 9636 14887 9639
rect 14918 9636 14924 9648
rect 14875 9608 14924 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 15028 9636 15056 9676
rect 15948 9676 16528 9704
rect 15948 9636 15976 9676
rect 15028 9608 15976 9636
rect 16025 9639 16083 9645
rect 16025 9605 16037 9639
rect 16071 9636 16083 9639
rect 16390 9636 16396 9648
rect 16071 9608 16396 9636
rect 16071 9605 16083 9608
rect 16025 9599 16083 9605
rect 16390 9596 16396 9608
rect 16448 9596 16454 9648
rect 16500 9636 16528 9676
rect 16850 9664 16856 9716
rect 16908 9704 16914 9716
rect 19610 9704 19616 9716
rect 16908 9676 19616 9704
rect 16908 9664 16914 9676
rect 19610 9664 19616 9676
rect 19668 9704 19674 9716
rect 20162 9704 20168 9716
rect 19668 9676 20168 9704
rect 19668 9664 19674 9676
rect 20162 9664 20168 9676
rect 20220 9664 20226 9716
rect 16666 9636 16672 9648
rect 16500 9608 16672 9636
rect 16666 9596 16672 9608
rect 16724 9596 16730 9648
rect 17221 9639 17279 9645
rect 17221 9605 17233 9639
rect 17267 9636 17279 9639
rect 18966 9636 18972 9648
rect 17267 9608 18972 9636
rect 17267 9605 17279 9608
rect 17221 9599 17279 9605
rect 18966 9596 18972 9608
rect 19024 9596 19030 9648
rect 13004 9540 13299 9568
rect 12805 9531 12863 9537
rect 9030 9500 9036 9512
rect 8680 9472 9036 9500
rect 9030 9460 9036 9472
rect 9088 9500 9094 9512
rect 9490 9500 9496 9512
rect 9088 9472 9496 9500
rect 9088 9460 9094 9472
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9500 9643 9503
rect 9766 9500 9772 9512
rect 9631 9472 9772 9500
rect 9631 9469 9643 9472
rect 9585 9463 9643 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10229 9503 10287 9509
rect 10229 9469 10241 9503
rect 10275 9500 10287 9503
rect 10318 9500 10324 9512
rect 10275 9472 10324 9500
rect 10275 9469 10287 9472
rect 10229 9463 10287 9469
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10502 9509 10508 9512
rect 10496 9500 10508 9509
rect 10463 9472 10508 9500
rect 10496 9463 10508 9472
rect 10502 9460 10508 9463
rect 10560 9460 10566 9512
rect 12434 9500 12440 9512
rect 12395 9472 12440 9500
rect 12434 9460 12440 9472
rect 12492 9460 12498 9512
rect 13173 9503 13231 9509
rect 13173 9469 13185 9503
rect 13219 9469 13231 9503
rect 13271 9500 13299 9540
rect 14642 9528 14648 9580
rect 14700 9568 14706 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 14700 9540 15393 9568
rect 14700 9528 14706 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 15381 9531 15439 9537
rect 16482 9528 16488 9580
rect 16540 9568 16546 9580
rect 16577 9571 16635 9577
rect 16577 9568 16589 9571
rect 16540 9540 16589 9568
rect 16540 9528 16546 9540
rect 16577 9537 16589 9540
rect 16623 9537 16635 9571
rect 16577 9531 16635 9537
rect 16868 9540 18000 9568
rect 13271 9472 13584 9500
rect 13173 9463 13231 9469
rect 7374 9432 7380 9444
rect 4479 9404 5387 9432
rect 6104 9404 7380 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 3050 9364 3056 9376
rect 3011 9336 3056 9364
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3510 9324 3516 9376
rect 3568 9364 3574 9376
rect 3694 9364 3700 9376
rect 3568 9336 3700 9364
rect 3568 9324 3574 9336
rect 3694 9324 3700 9336
rect 3752 9324 3758 9376
rect 4062 9364 4068 9376
rect 4023 9336 4068 9364
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 5258 9364 5264 9376
rect 4571 9336 5264 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5350 9324 5356 9376
rect 5408 9364 5414 9376
rect 6104 9364 6132 9404
rect 7374 9392 7380 9404
rect 7432 9392 7438 9444
rect 7650 9432 7656 9444
rect 7611 9404 7656 9432
rect 7650 9392 7656 9404
rect 7708 9392 7714 9444
rect 8665 9435 8723 9441
rect 8036 9404 8616 9432
rect 5408 9336 6132 9364
rect 5408 9324 5414 9336
rect 6178 9324 6184 9376
rect 6236 9364 6242 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 6236 9336 6469 9364
rect 6236 9324 6242 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8036 9364 8064 9404
rect 7607 9336 8064 9364
rect 8113 9367 8171 9373
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8113 9333 8125 9367
rect 8159 9364 8171 9367
rect 8205 9367 8263 9373
rect 8205 9364 8217 9367
rect 8159 9336 8217 9364
rect 8159 9333 8171 9336
rect 8113 9327 8171 9333
rect 8205 9333 8217 9336
rect 8251 9333 8263 9367
rect 8588 9364 8616 9404
rect 8665 9401 8677 9435
rect 8711 9432 8723 9435
rect 9122 9432 9128 9444
rect 8711 9404 9128 9432
rect 8711 9401 8723 9404
rect 8665 9395 8723 9401
rect 9122 9392 9128 9404
rect 9180 9392 9186 9444
rect 11238 9432 11244 9444
rect 9600 9404 11244 9432
rect 9600 9364 9628 9404
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 12621 9435 12679 9441
rect 12621 9432 12633 9435
rect 11848 9404 12633 9432
rect 11848 9392 11854 9404
rect 12621 9401 12633 9404
rect 12667 9401 12679 9435
rect 12621 9395 12679 9401
rect 12986 9392 12992 9444
rect 13044 9432 13050 9444
rect 13188 9432 13216 9463
rect 13044 9404 13216 9432
rect 13044 9392 13050 9404
rect 13354 9392 13360 9444
rect 13412 9441 13418 9444
rect 13412 9435 13476 9441
rect 13412 9401 13430 9435
rect 13464 9401 13476 9435
rect 13556 9432 13584 9472
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14550 9500 14556 9512
rect 14424 9472 14556 9500
rect 14424 9460 14430 9472
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 15197 9503 15255 9509
rect 15197 9500 15209 9503
rect 14792 9472 15209 9500
rect 14792 9460 14798 9472
rect 15197 9469 15209 9472
rect 15243 9469 15255 9503
rect 16868 9500 16896 9540
rect 15197 9463 15255 9469
rect 16132 9472 16896 9500
rect 15289 9435 15347 9441
rect 15289 9432 15301 9435
rect 13556 9404 15301 9432
rect 13412 9395 13476 9401
rect 15289 9401 15301 9404
rect 15335 9401 15347 9435
rect 15289 9395 15347 9401
rect 13412 9392 13418 9395
rect 8588 9336 9628 9364
rect 9677 9367 9735 9373
rect 8205 9327 8263 9333
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 10594 9364 10600 9376
rect 9723 9336 10600 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 10594 9324 10600 9336
rect 10652 9364 10658 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 10652 9336 11621 9364
rect 10652 9324 10658 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 11609 9327 11667 9333
rect 11885 9367 11943 9373
rect 11885 9333 11897 9367
rect 11931 9364 11943 9367
rect 13078 9364 13084 9376
rect 11931 9336 13084 9364
rect 11931 9333 11943 9336
rect 11885 9327 11943 9333
rect 13078 9324 13084 9336
rect 13136 9324 13142 9376
rect 14550 9364 14556 9376
rect 14511 9336 14556 9364
rect 14550 9324 14556 9336
rect 14608 9324 14614 9376
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 16132 9364 16160 9472
rect 16942 9460 16948 9512
rect 17000 9500 17006 9512
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 17000 9472 17049 9500
rect 17000 9460 17006 9472
rect 17037 9469 17049 9472
rect 17083 9469 17095 9503
rect 17773 9503 17831 9509
rect 17773 9500 17785 9503
rect 17037 9463 17095 9469
rect 17512 9472 17785 9500
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 16485 9435 16543 9441
rect 16485 9432 16497 9435
rect 16264 9404 16497 9432
rect 16264 9392 16270 9404
rect 16485 9401 16497 9404
rect 16531 9401 16543 9435
rect 17512 9432 17540 9472
rect 17773 9469 17785 9472
rect 17819 9469 17831 9503
rect 17972 9500 18000 9540
rect 18138 9528 18144 9580
rect 18196 9568 18202 9580
rect 18509 9571 18567 9577
rect 18509 9568 18521 9571
rect 18196 9540 18521 9568
rect 18196 9528 18202 9540
rect 18509 9537 18521 9540
rect 18555 9537 18567 9571
rect 18509 9531 18567 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9568 18751 9571
rect 19334 9568 19340 9580
rect 18739 9540 19340 9568
rect 18739 9537 18751 9540
rect 18693 9531 18751 9537
rect 19334 9528 19340 9540
rect 19392 9528 19398 9580
rect 19610 9577 19616 9580
rect 19567 9571 19616 9577
rect 19567 9537 19579 9571
rect 19613 9537 19616 9571
rect 19567 9531 19616 9537
rect 19610 9528 19616 9531
rect 19668 9528 19674 9580
rect 21634 9568 21640 9580
rect 21595 9540 21640 9568
rect 21634 9528 21640 9540
rect 21692 9528 21698 9580
rect 21821 9571 21879 9577
rect 21821 9537 21833 9571
rect 21867 9568 21879 9571
rect 22186 9568 22192 9580
rect 21867 9540 22192 9568
rect 21867 9537 21879 9540
rect 21821 9531 21879 9537
rect 22186 9528 22192 9540
rect 22244 9528 22250 9580
rect 18417 9503 18475 9509
rect 18417 9500 18429 9503
rect 17972 9472 18429 9500
rect 17773 9463 17831 9469
rect 18417 9469 18429 9472
rect 18463 9500 18475 9503
rect 18877 9503 18935 9509
rect 18877 9500 18889 9503
rect 18463 9472 18889 9500
rect 18463 9469 18475 9472
rect 18417 9463 18475 9469
rect 18877 9469 18889 9472
rect 18923 9469 18935 9503
rect 18877 9463 18935 9469
rect 18966 9460 18972 9512
rect 19024 9500 19030 9512
rect 19061 9503 19119 9509
rect 19061 9500 19073 9503
rect 19024 9472 19073 9500
rect 19024 9460 19030 9472
rect 19061 9469 19073 9472
rect 19107 9469 19119 9503
rect 19061 9463 19119 9469
rect 19150 9460 19156 9512
rect 19208 9500 19214 9512
rect 19426 9500 19432 9512
rect 19208 9472 19432 9500
rect 19208 9460 19214 9472
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19797 9503 19855 9509
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 20254 9500 20260 9512
rect 19843 9472 20260 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 20254 9460 20260 9472
rect 20312 9460 20318 9512
rect 16485 9395 16543 9401
rect 16592 9404 17540 9432
rect 17604 9404 19012 9432
rect 16592 9376 16620 9404
rect 16390 9364 16396 9376
rect 14792 9336 16160 9364
rect 16351 9336 16396 9364
rect 14792 9324 14798 9336
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16574 9324 16580 9376
rect 16632 9324 16638 9376
rect 17604 9373 17632 9404
rect 17589 9367 17647 9373
rect 17589 9333 17601 9367
rect 17635 9333 17647 9367
rect 17589 9327 17647 9333
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18598 9364 18604 9376
rect 18095 9336 18604 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18598 9324 18604 9336
rect 18656 9364 18662 9376
rect 18782 9364 18788 9376
rect 18656 9336 18788 9364
rect 18656 9324 18662 9336
rect 18782 9324 18788 9336
rect 18840 9324 18846 9376
rect 18984 9364 19012 9404
rect 20530 9392 20536 9444
rect 20588 9432 20594 9444
rect 21545 9435 21603 9441
rect 21545 9432 21557 9435
rect 20588 9404 21557 9432
rect 20588 9392 20594 9404
rect 21545 9401 21557 9404
rect 21591 9401 21603 9435
rect 21545 9395 21603 9401
rect 19426 9364 19432 9376
rect 18984 9336 19432 9364
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 19518 9324 19524 9376
rect 19576 9373 19582 9376
rect 19576 9364 19585 9373
rect 19576 9336 19621 9364
rect 19576 9327 19585 9336
rect 19576 9324 19582 9327
rect 20070 9324 20076 9376
rect 20128 9364 20134 9376
rect 20901 9367 20959 9373
rect 20901 9364 20913 9367
rect 20128 9336 20913 9364
rect 20128 9324 20134 9336
rect 20901 9333 20913 9336
rect 20947 9333 20959 9367
rect 21174 9364 21180 9376
rect 21135 9336 21180 9364
rect 20901 9327 20959 9333
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 1104 9274 22816 9296
rect 1104 9222 8246 9274
rect 8298 9222 8310 9274
rect 8362 9222 8374 9274
rect 8426 9222 8438 9274
rect 8490 9222 15510 9274
rect 15562 9222 15574 9274
rect 15626 9222 15638 9274
rect 15690 9222 15702 9274
rect 15754 9222 22816 9274
rect 1104 9200 22816 9222
rect 2498 9160 2504 9172
rect 2459 9132 2504 9160
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4488 9132 4537 9160
rect 4488 9120 4494 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 4525 9123 4583 9129
rect 4893 9163 4951 9169
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5350 9160 5356 9172
rect 4939 9132 5356 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5350 9120 5356 9132
rect 5408 9120 5414 9172
rect 5534 9160 5540 9172
rect 5495 9132 5540 9160
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 5902 9160 5908 9172
rect 5863 9132 5908 9160
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 5994 9120 6000 9172
rect 6052 9160 6058 9172
rect 6546 9160 6552 9172
rect 6052 9132 6097 9160
rect 6507 9132 6552 9160
rect 6052 9120 6058 9132
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 9401 9163 9459 9169
rect 7208 9132 9076 9160
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9092 3479 9095
rect 3878 9092 3884 9104
rect 3467 9064 3884 9092
rect 3467 9061 3479 9064
rect 3421 9055 3479 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 7098 9092 7104 9104
rect 4120 9064 7104 9092
rect 4120 9052 4126 9064
rect 7098 9052 7104 9064
rect 7156 9052 7162 9104
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3694 9024 3700 9036
rect 3375 8996 3700 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3694 8984 3700 8996
rect 3752 8984 3758 9036
rect 4985 9027 5043 9033
rect 3896 8996 4200 9024
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 3896 8956 3924 8996
rect 3651 8928 3924 8956
rect 4065 8959 4123 8965
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4172 8956 4200 8996
rect 4985 8993 4997 9027
rect 5031 9024 5043 9027
rect 6822 9024 6828 9036
rect 5031 8996 6828 9024
rect 5031 8993 5043 8996
rect 4985 8987 5043 8993
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 6963 8996 7144 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 5074 8956 5080 8968
rect 4172 8928 5080 8956
rect 4065 8919 4123 8925
rect 4080 8888 4108 8919
rect 5074 8916 5080 8928
rect 5132 8916 5138 8968
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8956 5322 8968
rect 5442 8956 5448 8968
rect 5316 8928 5448 8956
rect 5316 8916 5322 8928
rect 5442 8916 5448 8928
rect 5500 8956 5506 8968
rect 5994 8956 6000 8968
rect 5500 8928 6000 8956
rect 5500 8916 5506 8928
rect 5994 8916 6000 8928
rect 6052 8956 6058 8968
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 6052 8928 6101 8956
rect 6052 8916 6058 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 7006 8956 7012 8968
rect 6967 8928 7012 8956
rect 6089 8919 6147 8925
rect 7006 8916 7012 8928
rect 7064 8916 7070 8968
rect 4433 8891 4491 8897
rect 4433 8888 4445 8891
rect 4080 8860 4445 8888
rect 4433 8857 4445 8860
rect 4479 8888 4491 8891
rect 4479 8860 5120 8888
rect 4479 8857 4491 8860
rect 4433 8851 4491 8857
rect 5092 8832 5120 8860
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 5408 8860 6408 8888
rect 5408 8848 5414 8860
rect 2958 8820 2964 8832
rect 2919 8792 2964 8820
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 5074 8780 5080 8832
rect 5132 8780 5138 8832
rect 5442 8780 5448 8832
rect 5500 8820 5506 8832
rect 6270 8820 6276 8832
rect 5500 8792 6276 8820
rect 5500 8780 5506 8792
rect 6270 8780 6276 8792
rect 6328 8780 6334 8832
rect 6380 8820 6408 8860
rect 6822 8848 6828 8900
rect 6880 8888 6886 8900
rect 7116 8888 7144 8996
rect 7208 8965 7236 9132
rect 8021 9095 8079 9101
rect 8021 9092 8033 9095
rect 7852 9064 8033 9092
rect 7374 8984 7380 9036
rect 7432 9024 7438 9036
rect 7852 9024 7880 9064
rect 8021 9061 8033 9064
rect 8067 9061 8079 9095
rect 8021 9055 8079 9061
rect 8570 9052 8576 9104
rect 8628 9092 8634 9104
rect 8941 9095 8999 9101
rect 8941 9092 8953 9095
rect 8628 9064 8953 9092
rect 8628 9052 8634 9064
rect 8941 9061 8953 9064
rect 8987 9061 8999 9095
rect 9048 9092 9076 9132
rect 9401 9129 9413 9163
rect 9447 9160 9459 9163
rect 9766 9160 9772 9172
rect 9447 9132 9772 9160
rect 9447 9129 9459 9132
rect 9401 9123 9459 9129
rect 9766 9120 9772 9132
rect 9824 9120 9830 9172
rect 9876 9132 10180 9160
rect 9876 9092 9904 9132
rect 9048 9064 9904 9092
rect 9944 9095 10002 9101
rect 8941 9055 8999 9061
rect 9944 9061 9956 9095
rect 9990 9092 10002 9095
rect 10152 9092 10180 9132
rect 10778 9120 10784 9172
rect 10836 9160 10842 9172
rect 10836 9132 13369 9160
rect 10836 9120 10842 9132
rect 9990 9064 10088 9092
rect 10152 9064 12572 9092
rect 9990 9061 10002 9064
rect 9944 9055 10002 9061
rect 7432 8996 7880 9024
rect 7432 8984 7438 8996
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 7984 8996 8029 9024
rect 8128 8996 9413 9024
rect 7984 8984 7990 8996
rect 7193 8959 7251 8965
rect 7193 8925 7205 8959
rect 7239 8925 7251 8959
rect 7193 8919 7251 8925
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 8128 8956 8156 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9490 8984 9496 9036
rect 9548 8984 9554 9036
rect 9674 8984 9680 9036
rect 9732 9024 9738 9036
rect 10060 9024 10088 9064
rect 10870 9024 10876 9036
rect 9732 8996 9777 9024
rect 10060 8996 10876 9024
rect 9732 8984 9738 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 11425 9027 11483 9033
rect 11425 8993 11437 9027
rect 11471 9024 11483 9027
rect 11514 9024 11520 9036
rect 11471 8996 11520 9024
rect 11471 8993 11483 8996
rect 11425 8987 11483 8993
rect 11514 8984 11520 8996
rect 11572 8984 11578 9036
rect 11698 9033 11704 9036
rect 11692 9024 11704 9033
rect 11659 8996 11704 9024
rect 11692 8987 11704 8996
rect 11698 8984 11704 8987
rect 11756 8984 11762 9036
rect 12544 9024 12572 9064
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12894 9092 12900 9104
rect 12676 9064 12900 9092
rect 12676 9052 12682 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 13341 9101 13369 9132
rect 13446 9120 13452 9172
rect 13504 9160 13510 9172
rect 14642 9160 14648 9172
rect 13504 9132 14648 9160
rect 13504 9120 13510 9132
rect 14642 9120 14648 9132
rect 14700 9120 14706 9172
rect 14737 9163 14795 9169
rect 14737 9129 14749 9163
rect 14783 9160 14795 9163
rect 16298 9160 16304 9172
rect 14783 9132 16304 9160
rect 14783 9129 14795 9132
rect 14737 9123 14795 9129
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 16390 9120 16396 9172
rect 16448 9160 16454 9172
rect 16850 9160 16856 9172
rect 16448 9132 16856 9160
rect 16448 9120 16454 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 18230 9160 18236 9172
rect 18191 9132 18236 9160
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 18564 9132 20024 9160
rect 18564 9120 18570 9132
rect 13326 9095 13384 9101
rect 13326 9061 13338 9095
rect 13372 9092 13384 9095
rect 14550 9092 14556 9104
rect 13372 9064 14556 9092
rect 13372 9061 13384 9064
rect 13326 9055 13384 9061
rect 14550 9052 14556 9064
rect 14608 9052 14614 9104
rect 14918 9052 14924 9104
rect 14976 9092 14982 9104
rect 14976 9064 15424 9092
rect 14976 9052 14982 9064
rect 15286 9024 15292 9036
rect 12544 8996 15292 9024
rect 15286 8984 15292 8996
rect 15344 8984 15350 9036
rect 15396 9024 15424 9064
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 16638 9095 16696 9101
rect 16638 9092 16650 9095
rect 15528 9064 16650 9092
rect 15528 9052 15534 9064
rect 16638 9061 16650 9064
rect 16684 9092 16696 9095
rect 16758 9092 16764 9104
rect 16684 9064 16764 9092
rect 16684 9061 16696 9064
rect 16638 9055 16696 9061
rect 16758 9052 16764 9064
rect 16816 9052 16822 9104
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15396 8996 15669 9024
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 16393 9027 16451 9033
rect 16393 8993 16405 9027
rect 16439 9024 16451 9027
rect 16482 9024 16488 9036
rect 16439 8996 16488 9024
rect 16439 8993 16451 8996
rect 16393 8987 16451 8993
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 18049 9027 18107 9033
rect 18049 8993 18061 9027
rect 18095 9024 18107 9027
rect 18322 9024 18328 9036
rect 18095 8996 18328 9024
rect 18095 8993 18107 8996
rect 18049 8987 18107 8993
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 18924 9027 18982 9033
rect 18924 9024 18936 9027
rect 18748 8996 18936 9024
rect 18748 8984 18754 8996
rect 18924 8993 18936 8996
rect 18970 8993 18982 9027
rect 19702 9024 19708 9036
rect 18924 8987 18982 8993
rect 19260 8996 19708 9024
rect 7708 8928 8156 8956
rect 8205 8959 8263 8965
rect 7708 8916 7714 8928
rect 8205 8925 8217 8959
rect 8251 8956 8263 8959
rect 8846 8956 8852 8968
rect 8251 8928 8852 8956
rect 8251 8925 8263 8928
rect 8205 8919 8263 8925
rect 8846 8916 8852 8928
rect 8904 8916 8910 8968
rect 8938 8916 8944 8968
rect 8996 8956 9002 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8996 8928 9045 8956
rect 8996 8916 9002 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9508 8956 9536 8984
rect 9263 8928 9536 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 12434 8916 12440 8968
rect 12492 8956 12498 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12492 8928 13093 8956
rect 12492 8916 12498 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14550 8956 14556 8968
rect 14424 8928 14556 8956
rect 14424 8916 14430 8928
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14826 8916 14832 8968
rect 14884 8956 14890 8968
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 14884 8928 15761 8956
rect 14884 8916 14890 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 15838 8916 15844 8968
rect 15896 8956 15902 8968
rect 15896 8928 15941 8956
rect 15896 8916 15902 8928
rect 18138 8916 18144 8968
rect 18196 8956 18202 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18196 8928 18613 8956
rect 18196 8916 18202 8928
rect 18601 8925 18613 8928
rect 18647 8956 18659 8959
rect 18782 8956 18788 8968
rect 18647 8928 18788 8956
rect 18647 8925 18659 8928
rect 18601 8919 18659 8925
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 19107 8959 19165 8965
rect 19107 8925 19119 8959
rect 19153 8956 19165 8959
rect 19260 8956 19288 8996
rect 19702 8984 19708 8996
rect 19760 8984 19766 9036
rect 19996 9024 20024 9132
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20404 9132 20453 9160
rect 20404 9120 20410 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 20162 9052 20168 9104
rect 20220 9092 20226 9104
rect 21168 9095 21226 9101
rect 21168 9092 21180 9095
rect 20220 9064 21180 9092
rect 20220 9052 20226 9064
rect 21168 9061 21180 9064
rect 21214 9092 21226 9095
rect 22278 9092 22284 9104
rect 21214 9064 22284 9092
rect 21214 9061 21226 9064
rect 21168 9055 21226 9061
rect 22278 9052 22284 9064
rect 22336 9052 22342 9104
rect 20898 9024 20904 9036
rect 19996 8996 20904 9024
rect 20898 8984 20904 8996
rect 20956 8984 20962 9036
rect 19153 8928 19288 8956
rect 19337 8959 19395 8965
rect 19153 8925 19165 8928
rect 19107 8919 19165 8925
rect 19337 8925 19349 8959
rect 19383 8956 19395 8959
rect 20530 8956 20536 8968
rect 19383 8928 20536 8956
rect 19383 8925 19395 8928
rect 19337 8919 19395 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 7558 8888 7564 8900
rect 6880 8860 7144 8888
rect 7519 8860 7564 8888
rect 6880 8848 6886 8860
rect 7558 8848 7564 8860
rect 7616 8848 7622 8900
rect 9490 8888 9496 8900
rect 7668 8860 9496 8888
rect 7668 8820 7696 8860
rect 9490 8848 9496 8860
rect 9548 8848 9554 8900
rect 11330 8888 11336 8900
rect 11072 8860 11336 8888
rect 6380 8792 7696 8820
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9674 8820 9680 8832
rect 8619 8792 9680 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 10042 8780 10048 8832
rect 10100 8820 10106 8832
rect 11072 8829 11100 8860
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 14090 8848 14096 8900
rect 14148 8888 14154 8900
rect 14148 8860 15424 8888
rect 14148 8848 14154 8860
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10100 8792 11069 8820
rect 10100 8780 10106 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 12618 8820 12624 8832
rect 11296 8792 12624 8820
rect 11296 8780 11302 8792
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 12805 8823 12863 8829
rect 12805 8789 12817 8823
rect 12851 8820 12863 8823
rect 12986 8820 12992 8832
rect 12851 8792 12992 8820
rect 12851 8789 12863 8792
rect 12805 8783 12863 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 14182 8780 14188 8832
rect 14240 8820 14246 8832
rect 14461 8823 14519 8829
rect 14461 8820 14473 8823
rect 14240 8792 14473 8820
rect 14240 8780 14246 8792
rect 14461 8789 14473 8792
rect 14507 8789 14519 8823
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 14461 8783 14519 8789
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15396 8820 15424 8860
rect 15470 8848 15476 8900
rect 15528 8888 15534 8900
rect 16390 8888 16396 8900
rect 15528 8860 16396 8888
rect 15528 8848 15534 8860
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 17328 8860 17908 8888
rect 17328 8820 17356 8860
rect 17770 8820 17776 8832
rect 15396 8792 17356 8820
rect 17731 8792 17776 8820
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 17880 8820 17908 8860
rect 22186 8848 22192 8900
rect 22244 8888 22250 8900
rect 22281 8891 22339 8897
rect 22281 8888 22293 8891
rect 22244 8860 22293 8888
rect 22244 8848 22250 8860
rect 22281 8857 22293 8860
rect 22327 8857 22339 8891
rect 22281 8851 22339 8857
rect 19426 8820 19432 8832
rect 17880 8792 19432 8820
rect 19426 8780 19432 8792
rect 19484 8780 19490 8832
rect 1104 8730 22816 8752
rect 1104 8678 4614 8730
rect 4666 8678 4678 8730
rect 4730 8678 4742 8730
rect 4794 8678 4806 8730
rect 4858 8678 11878 8730
rect 11930 8678 11942 8730
rect 11994 8678 12006 8730
rect 12058 8678 12070 8730
rect 12122 8678 19142 8730
rect 19194 8678 19206 8730
rect 19258 8678 19270 8730
rect 19322 8678 19334 8730
rect 19386 8678 22816 8730
rect 1104 8656 22816 8678
rect 2685 8619 2743 8625
rect 2685 8585 2697 8619
rect 2731 8616 2743 8619
rect 4062 8616 4068 8628
rect 2731 8588 4068 8616
rect 2731 8585 2743 8588
rect 2685 8579 2743 8585
rect 2792 8489 2820 8588
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 6914 8616 6920 8628
rect 5767 8588 6920 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7285 8619 7343 8625
rect 7285 8585 7297 8619
rect 7331 8616 7343 8619
rect 11238 8616 11244 8628
rect 7331 8588 11244 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11698 8616 11704 8628
rect 11659 8588 11704 8616
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 15286 8616 15292 8628
rect 12299 8588 15292 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15930 8616 15936 8628
rect 15436 8588 15936 8616
rect 15436 8576 15442 8588
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16356 8588 17417 8616
rect 16356 8576 16362 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 17405 8579 17463 8585
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 21174 8616 21180 8628
rect 20272 8588 21180 8616
rect 4709 8551 4767 8557
rect 4709 8517 4721 8551
rect 4755 8548 4767 8551
rect 5442 8548 5448 8560
rect 4755 8520 5448 8548
rect 4755 8517 4767 8520
rect 4709 8511 4767 8517
rect 5442 8508 5448 8520
rect 5500 8508 5506 8560
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6052 8520 6408 8548
rect 6052 8508 6058 8520
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 2958 8440 2964 8492
rect 3016 8480 3022 8492
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3016 8452 3985 8480
rect 3016 8440 3022 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 3973 8443 4031 8449
rect 4080 8452 4169 8480
rect 4080 8424 4108 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 5350 8480 5356 8492
rect 5311 8452 5356 8480
rect 4157 8443 4215 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 6380 8489 6408 8520
rect 7466 8508 7472 8560
rect 7524 8548 7530 8560
rect 7653 8551 7711 8557
rect 7653 8548 7665 8551
rect 7524 8520 7665 8548
rect 7524 8508 7530 8520
rect 7653 8517 7665 8520
rect 7699 8517 7711 8551
rect 7653 8511 7711 8517
rect 8110 8508 8116 8560
rect 8168 8548 8174 8560
rect 8662 8548 8668 8560
rect 8168 8520 8668 8548
rect 8168 8508 8174 8520
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11480 8520 11989 8548
rect 11480 8508 11486 8520
rect 11977 8517 11989 8520
rect 12023 8548 12035 8551
rect 12158 8548 12164 8560
rect 12023 8520 12164 8548
rect 12023 8517 12035 8520
rect 11977 8511 12035 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 12268 8520 13124 8548
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 7926 8440 7932 8492
rect 7984 8480 7990 8492
rect 8202 8480 8208 8492
rect 7984 8452 8208 8480
rect 7984 8440 7990 8452
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8343 8452 8800 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 3881 8415 3939 8421
rect 3881 8412 3893 8415
rect 2096 8384 3893 8412
rect 2096 8372 2102 8384
rect 3881 8381 3893 8384
rect 3927 8381 3939 8415
rect 3881 8375 3939 8381
rect 4062 8372 4068 8424
rect 4120 8372 4126 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 5074 8412 5080 8424
rect 4663 8384 5080 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 5074 8372 5080 8384
rect 5132 8372 5138 8424
rect 6086 8412 6092 8424
rect 6047 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 8478 8412 8484 8424
rect 7147 8384 8484 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 8478 8372 8484 8384
rect 8536 8372 8542 8424
rect 8665 8415 8723 8421
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 8772 8412 8800 8452
rect 9950 8440 9956 8492
rect 10008 8480 10014 8492
rect 10318 8480 10324 8492
rect 10008 8452 10324 8480
rect 10008 8440 10014 8452
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 12268 8480 12296 8520
rect 12986 8480 12992 8492
rect 11348 8452 12296 8480
rect 12947 8452 12992 8480
rect 8772 8384 9076 8412
rect 8665 8375 8723 8381
rect 3237 8347 3295 8353
rect 3237 8313 3249 8347
rect 3283 8344 3295 8347
rect 4246 8344 4252 8356
rect 3283 8316 4252 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 5902 8344 5908 8356
rect 5215 8316 5908 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5902 8304 5908 8316
rect 5960 8304 5966 8356
rect 6178 8344 6184 8356
rect 6139 8316 6184 8344
rect 6178 8304 6184 8316
rect 6236 8304 6242 8356
rect 8018 8344 8024 8356
rect 7979 8316 8024 8344
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8680 8344 8708 8375
rect 8260 8316 8708 8344
rect 8260 8304 8266 8316
rect 8754 8304 8760 8356
rect 8812 8344 8818 8356
rect 8910 8347 8968 8353
rect 8910 8344 8922 8347
rect 8812 8316 8922 8344
rect 8812 8304 8818 8316
rect 8910 8313 8922 8316
rect 8956 8313 8968 8347
rect 9048 8344 9076 8384
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 10229 8415 10287 8421
rect 10229 8412 10241 8415
rect 9272 8384 10241 8412
rect 9272 8372 9278 8384
rect 10229 8381 10241 8384
rect 10275 8381 10287 8415
rect 11348 8412 11376 8452
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13096 8480 13124 8520
rect 14642 8508 14648 8560
rect 14700 8548 14706 8560
rect 14829 8551 14887 8557
rect 14829 8548 14841 8551
rect 14700 8520 14841 8548
rect 14700 8508 14706 8520
rect 14829 8517 14841 8520
rect 14875 8517 14887 8551
rect 14829 8511 14887 8517
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8517 17003 8551
rect 16945 8511 17003 8517
rect 13096 8452 13584 8480
rect 10229 8375 10287 8381
rect 10520 8384 11376 8412
rect 12161 8415 12219 8421
rect 10520 8344 10548 8384
rect 12161 8381 12173 8415
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8412 12863 8415
rect 13078 8412 13084 8424
rect 12851 8384 13084 8412
rect 12851 8381 12863 8384
rect 12805 8375 12863 8381
rect 9048 8316 10548 8344
rect 10588 8347 10646 8353
rect 8910 8307 8968 8313
rect 10588 8313 10600 8347
rect 10634 8344 10646 8347
rect 10870 8344 10876 8356
rect 10634 8316 10876 8344
rect 10634 8313 10646 8316
rect 10588 8307 10646 8313
rect 10870 8304 10876 8316
rect 10928 8304 10934 8356
rect 11054 8304 11060 8356
rect 11112 8344 11118 8356
rect 12176 8344 12204 8375
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13446 8412 13452 8424
rect 13407 8384 13452 8412
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 13556 8412 13584 8452
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 15105 8483 15163 8489
rect 15105 8480 15117 8483
rect 14608 8452 15117 8480
rect 14608 8440 14614 8452
rect 15105 8449 15117 8452
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15378 8440 15384 8492
rect 15436 8489 15442 8492
rect 15436 8483 15486 8489
rect 15436 8449 15440 8483
rect 15474 8449 15486 8483
rect 15436 8443 15486 8449
rect 15568 8483 15626 8489
rect 15568 8449 15580 8483
rect 15614 8480 15626 8483
rect 16298 8480 16304 8492
rect 15614 8452 16304 8480
rect 15614 8449 15626 8452
rect 15568 8443 15626 8449
rect 15436 8440 15442 8443
rect 13716 8415 13774 8421
rect 13716 8412 13728 8415
rect 13556 8384 13728 8412
rect 13716 8381 13728 8384
rect 13762 8412 13774 8415
rect 14090 8412 14096 8424
rect 13762 8384 14096 8412
rect 13762 8381 13774 8384
rect 13716 8375 13774 8381
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 15583 8412 15611 8443
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 16960 8480 16988 8511
rect 16408 8452 16988 8480
rect 14700 8384 15611 8412
rect 15841 8415 15899 8421
rect 14700 8372 14706 8384
rect 15841 8381 15853 8415
rect 15887 8412 15899 8415
rect 15930 8412 15936 8424
rect 15887 8384 15936 8412
rect 15887 8381 15899 8384
rect 15841 8375 15899 8381
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 16206 8372 16212 8424
rect 16264 8412 16270 8424
rect 16408 8412 16436 8452
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 20070 8480 20076 8492
rect 18012 8452 20076 8480
rect 18012 8440 18018 8452
rect 20070 8440 20076 8452
rect 20128 8440 20134 8492
rect 20165 8483 20223 8489
rect 20165 8449 20177 8483
rect 20211 8480 20223 8483
rect 20272 8480 20300 8588
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8548 20775 8551
rect 20806 8548 20812 8560
rect 20763 8520 20812 8548
rect 20763 8517 20775 8520
rect 20717 8511 20775 8517
rect 20806 8508 20812 8520
rect 20864 8508 20870 8560
rect 22278 8548 22284 8560
rect 22239 8520 22284 8548
rect 22278 8508 22284 8520
rect 22336 8508 22342 8560
rect 20211 8452 20300 8480
rect 20349 8483 20407 8489
rect 20211 8449 20223 8452
rect 20165 8443 20223 8449
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20898 8480 20904 8492
rect 20859 8452 20904 8480
rect 20349 8443 20407 8449
rect 16264 8384 16436 8412
rect 16264 8372 16270 8384
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17221 8415 17279 8421
rect 17221 8412 17233 8415
rect 16632 8384 17233 8412
rect 16632 8372 16638 8384
rect 17221 8381 17233 8384
rect 17267 8381 17279 8415
rect 17221 8375 17279 8381
rect 18877 8415 18935 8421
rect 18877 8381 18889 8415
rect 18923 8412 18935 8415
rect 19610 8412 19616 8424
rect 18923 8384 19616 8412
rect 18923 8381 18935 8384
rect 18877 8375 18935 8381
rect 19610 8372 19616 8384
rect 19668 8372 19674 8424
rect 14826 8344 14832 8356
rect 11112 8316 12204 8344
rect 12452 8316 14832 8344
rect 11112 8304 11118 8316
rect 3513 8279 3571 8285
rect 3513 8245 3525 8279
rect 3559 8276 3571 8279
rect 5718 8276 5724 8288
rect 3559 8248 5724 8276
rect 3559 8245 3571 8248
rect 3513 8239 3571 8245
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 7742 8236 7748 8288
rect 7800 8276 7806 8288
rect 8113 8279 8171 8285
rect 8113 8276 8125 8279
rect 7800 8248 8125 8276
rect 7800 8236 7806 8248
rect 8113 8245 8125 8248
rect 8159 8276 8171 8279
rect 9214 8276 9220 8288
rect 8159 8248 9220 8276
rect 8159 8245 8171 8248
rect 8113 8239 8171 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 12452 8285 12480 8316
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 17954 8344 17960 8356
rect 17184 8316 17960 8344
rect 17184 8304 17190 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 19518 8344 19524 8356
rect 19479 8316 19524 8344
rect 19518 8304 19524 8316
rect 19576 8344 19582 8356
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 19576 8316 20085 8344
rect 19576 8304 19582 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20364 8344 20392 8443
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 20533 8415 20591 8421
rect 20533 8381 20545 8415
rect 20579 8412 20591 8415
rect 20622 8412 20628 8424
rect 20579 8384 20628 8412
rect 20579 8381 20591 8384
rect 20533 8375 20591 8381
rect 20622 8372 20628 8384
rect 20680 8372 20686 8424
rect 21168 8415 21226 8421
rect 21168 8381 21180 8415
rect 21214 8412 21226 8415
rect 22186 8412 22192 8424
rect 21214 8384 22192 8412
rect 21214 8381 21226 8384
rect 21168 8375 21226 8381
rect 22186 8372 22192 8384
rect 22244 8372 22250 8424
rect 22278 8344 22284 8356
rect 20364 8316 22284 8344
rect 20073 8307 20131 8313
rect 22278 8304 22284 8316
rect 22336 8304 22342 8356
rect 10229 8279 10287 8285
rect 10229 8245 10241 8279
rect 10275 8276 10287 8279
rect 12253 8279 12311 8285
rect 12253 8276 12265 8279
rect 10275 8248 12265 8276
rect 10275 8245 10287 8248
rect 10229 8239 10287 8245
rect 12253 8245 12265 8248
rect 12299 8245 12311 8279
rect 12253 8239 12311 8245
rect 12437 8279 12495 8285
rect 12437 8245 12449 8279
rect 12483 8245 12495 8279
rect 12437 8239 12495 8245
rect 12897 8279 12955 8285
rect 12897 8245 12909 8279
rect 12943 8276 12955 8279
rect 13722 8276 13728 8288
rect 12943 8248 13728 8276
rect 12943 8245 12955 8248
rect 12897 8239 12955 8245
rect 13722 8236 13728 8248
rect 13780 8236 13786 8288
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 15194 8276 15200 8288
rect 14608 8248 15200 8276
rect 14608 8236 14614 8248
rect 15194 8236 15200 8248
rect 15252 8236 15258 8288
rect 18690 8276 18696 8288
rect 18651 8248 18696 8276
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 1104 8186 22816 8208
rect 1104 8134 8246 8186
rect 8298 8134 8310 8186
rect 8362 8134 8374 8186
rect 8426 8134 8438 8186
rect 8490 8134 15510 8186
rect 15562 8134 15574 8186
rect 15626 8134 15638 8186
rect 15690 8134 15702 8186
rect 15754 8134 22816 8186
rect 1104 8112 22816 8134
rect 5258 8072 5264 8084
rect 5219 8044 5264 8072
rect 5258 8032 5264 8044
rect 5316 8032 5322 8084
rect 5902 8072 5908 8084
rect 5863 8044 5908 8072
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6638 8072 6644 8084
rect 6411 8044 6644 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6638 8032 6644 8044
rect 6696 8032 6702 8084
rect 6917 8075 6975 8081
rect 6917 8041 6929 8075
rect 6963 8072 6975 8075
rect 7374 8072 7380 8084
rect 6963 8044 7380 8072
rect 6963 8041 6975 8044
rect 6917 8035 6975 8041
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8812 8044 9321 8072
rect 8812 8032 8818 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 11701 8075 11759 8081
rect 9309 8035 9367 8041
rect 9876 8044 11652 8072
rect 3513 8007 3571 8013
rect 3513 7973 3525 8007
rect 3559 8004 3571 8007
rect 7190 8004 7196 8016
rect 3559 7976 7196 8004
rect 3559 7973 3571 7976
rect 3513 7967 3571 7973
rect 7190 7964 7196 7976
rect 7248 7964 7254 8016
rect 7285 8007 7343 8013
rect 7285 7973 7297 8007
rect 7331 8004 7343 8007
rect 9876 8004 9904 8044
rect 7331 7976 9904 8004
rect 9944 8007 10002 8013
rect 7331 7973 7343 7976
rect 7285 7967 7343 7973
rect 9944 7973 9956 8007
rect 9990 8004 10002 8007
rect 10042 8004 10048 8016
rect 9990 7976 10048 8004
rect 9990 7973 10002 7976
rect 9944 7967 10002 7973
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 5353 7939 5411 7945
rect 5353 7905 5365 7939
rect 5399 7936 5411 7939
rect 6270 7936 6276 7948
rect 5399 7908 6276 7936
rect 5399 7905 5411 7908
rect 5353 7899 5411 7905
rect 6270 7896 6276 7908
rect 6328 7896 6334 7948
rect 8196 7939 8254 7945
rect 8196 7905 8208 7939
rect 8242 7936 8254 7939
rect 9030 7936 9036 7948
rect 8242 7908 9036 7936
rect 8242 7905 8254 7908
rect 8196 7899 8254 7905
rect 9030 7896 9036 7908
rect 9088 7936 9094 7948
rect 9582 7936 9588 7948
rect 9088 7908 9588 7936
rect 9088 7896 9094 7908
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 9677 7939 9735 7945
rect 9677 7905 9689 7939
rect 9723 7936 9735 7939
rect 10502 7936 10508 7948
rect 9723 7908 10508 7936
rect 9723 7905 9735 7908
rect 9677 7899 9735 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 11330 7936 11336 7948
rect 11291 7908 11336 7936
rect 11330 7896 11336 7908
rect 11388 7896 11394 7948
rect 11624 7936 11652 8044
rect 11701 8041 11713 8075
rect 11747 8072 11759 8075
rect 14734 8072 14740 8084
rect 11747 8044 14740 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 14734 8032 14740 8044
rect 14792 8032 14798 8084
rect 16758 8072 16764 8084
rect 16719 8044 16764 8072
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 18414 8072 18420 8084
rect 18375 8044 18420 8072
rect 18414 8032 18420 8044
rect 18472 8032 18478 8084
rect 19426 8032 19432 8084
rect 19484 8072 19490 8084
rect 19889 8075 19947 8081
rect 19889 8072 19901 8075
rect 19484 8044 19901 8072
rect 19484 8032 19490 8044
rect 19889 8041 19901 8044
rect 19935 8041 19947 8075
rect 19889 8035 19947 8041
rect 19978 8032 19984 8084
rect 20036 8072 20042 8084
rect 20162 8072 20168 8084
rect 20036 8044 20168 8072
rect 20036 8032 20042 8044
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 12152 8007 12210 8013
rect 12152 7973 12164 8007
rect 12198 8004 12210 8007
rect 12986 8004 12992 8016
rect 12198 7976 12992 8004
rect 12198 7973 12210 7976
rect 12152 7967 12210 7973
rect 12986 7964 12992 7976
rect 13044 7964 13050 8016
rect 13357 8007 13415 8013
rect 13357 7973 13369 8007
rect 13403 8004 13415 8007
rect 13808 8007 13866 8013
rect 13808 8004 13820 8007
rect 13403 7976 13820 8004
rect 13403 7973 13415 7976
rect 13357 7967 13415 7973
rect 13808 7973 13820 7976
rect 13854 8004 13866 8007
rect 15838 8004 15844 8016
rect 13854 7976 15844 8004
rect 13854 7973 13866 7976
rect 13808 7967 13866 7973
rect 15838 7964 15844 7976
rect 15896 7964 15902 8016
rect 16298 7964 16304 8016
rect 16356 8004 16362 8016
rect 18432 8004 18460 8032
rect 18754 8007 18812 8013
rect 18754 8004 18766 8007
rect 16356 7976 17908 8004
rect 18432 7976 18766 8004
rect 16356 7964 16362 7976
rect 14642 7936 14648 7948
rect 11624 7908 14648 7936
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 15289 7939 15347 7945
rect 15289 7905 15301 7939
rect 15335 7936 15347 7939
rect 15637 7939 15695 7945
rect 15637 7936 15649 7939
rect 15335 7908 15649 7936
rect 15335 7905 15347 7908
rect 15289 7899 15347 7905
rect 15637 7905 15649 7908
rect 15683 7905 15695 7939
rect 17293 7939 17351 7945
rect 17293 7936 17305 7939
rect 15637 7899 15695 7905
rect 16408 7908 17305 7936
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4430 7868 4436 7880
rect 4387 7840 4436 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 5442 7828 5448 7880
rect 5500 7868 5506 7880
rect 6454 7868 6460 7880
rect 5500 7840 5545 7868
rect 6415 7840 6460 7868
rect 5500 7828 5506 7840
rect 6454 7828 6460 7840
rect 6512 7828 6518 7880
rect 7374 7868 7380 7880
rect 7335 7840 7380 7868
rect 7374 7828 7380 7840
rect 7432 7828 7438 7880
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 7607 7840 7880 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7732 4951 7735
rect 6178 7732 6184 7744
rect 4939 7704 6184 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 7852 7732 7880 7840
rect 7926 7828 7932 7880
rect 7984 7868 7990 7880
rect 7984 7840 8029 7868
rect 7984 7828 7990 7840
rect 9122 7828 9128 7880
rect 9180 7868 9186 7880
rect 9490 7868 9496 7880
rect 9180 7840 9496 7868
rect 9180 7828 9186 7840
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 11514 7828 11520 7880
rect 11572 7868 11578 7880
rect 11885 7871 11943 7877
rect 11885 7868 11897 7871
rect 11572 7840 11897 7868
rect 11572 7828 11578 7840
rect 11885 7837 11897 7840
rect 11931 7837 11943 7871
rect 13538 7868 13544 7880
rect 13499 7840 13544 7868
rect 11885 7831 11943 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15381 7871 15439 7877
rect 15381 7868 15393 7871
rect 15252 7840 15393 7868
rect 15252 7828 15258 7840
rect 15381 7837 15393 7840
rect 15427 7837 15439 7871
rect 15381 7831 15439 7837
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9306 7800 9312 7812
rect 8996 7772 9312 7800
rect 8996 7760 9002 7772
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 11701 7803 11759 7809
rect 11701 7800 11713 7803
rect 10612 7772 11713 7800
rect 10612 7732 10640 7772
rect 11701 7769 11713 7772
rect 11747 7769 11759 7803
rect 11701 7763 11759 7769
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 13357 7803 13415 7809
rect 13357 7800 13369 7803
rect 13311 7772 13369 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 13357 7769 13369 7772
rect 13403 7769 13415 7803
rect 13357 7763 13415 7769
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 14792 7772 15424 7800
rect 14792 7760 14798 7772
rect 7852 7704 10640 7732
rect 10870 7692 10876 7744
rect 10928 7732 10934 7744
rect 11057 7735 11115 7741
rect 11057 7732 11069 7735
rect 10928 7704 11069 7732
rect 10928 7692 10934 7704
rect 11057 7701 11069 7704
rect 11103 7701 11115 7735
rect 11057 7695 11115 7701
rect 11517 7735 11575 7741
rect 11517 7701 11529 7735
rect 11563 7732 11575 7735
rect 12986 7732 12992 7744
rect 11563 7704 12992 7732
rect 11563 7701 11575 7704
rect 11517 7695 11575 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 13814 7732 13820 7744
rect 13136 7704 13820 7732
rect 13136 7692 13142 7704
rect 13814 7692 13820 7704
rect 13872 7692 13878 7744
rect 13906 7692 13912 7744
rect 13964 7732 13970 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 13964 7704 14933 7732
rect 13964 7692 13970 7704
rect 14921 7701 14933 7704
rect 14967 7732 14979 7735
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 14967 7704 15301 7732
rect 14967 7701 14979 7704
rect 14921 7695 14979 7701
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15396 7732 15424 7772
rect 16408 7732 16436 7908
rect 17293 7905 17305 7908
rect 17339 7936 17351 7939
rect 17770 7936 17776 7948
rect 17339 7908 17776 7936
rect 17339 7905 17351 7908
rect 17293 7899 17351 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 17880 7936 17908 7976
rect 18754 7973 18766 7976
rect 18800 7973 18812 8007
rect 18754 7967 18812 7973
rect 20254 7964 20260 8016
rect 20312 8004 20318 8016
rect 21269 8007 21327 8013
rect 21269 8004 21281 8007
rect 20312 7976 21281 8004
rect 20312 7964 20318 7976
rect 21269 7973 21281 7976
rect 21315 7973 21327 8007
rect 21269 7967 21327 7973
rect 17880 7908 19564 7936
rect 17037 7871 17095 7877
rect 17037 7837 17049 7871
rect 17083 7837 17095 7871
rect 18506 7868 18512 7880
rect 18467 7840 18512 7868
rect 17037 7831 17095 7837
rect 15396 7704 16436 7732
rect 17052 7732 17080 7831
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 19536 7868 19564 7908
rect 19610 7896 19616 7948
rect 19668 7936 19674 7948
rect 20349 7939 20407 7945
rect 20349 7936 20361 7939
rect 19668 7908 20361 7936
rect 19668 7896 19674 7908
rect 20349 7905 20361 7908
rect 20395 7905 20407 7939
rect 21910 7936 21916 7948
rect 21871 7908 21916 7936
rect 20349 7899 20407 7905
rect 21910 7896 21916 7908
rect 21968 7896 21974 7948
rect 20070 7868 20076 7880
rect 19536 7840 20076 7868
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20438 7868 20444 7880
rect 20399 7840 20444 7868
rect 20438 7828 20444 7840
rect 20496 7828 20502 7880
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 21361 7871 21419 7877
rect 20588 7840 20633 7868
rect 20588 7828 20594 7840
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21542 7868 21548 7880
rect 21503 7840 21548 7868
rect 21361 7831 21419 7837
rect 18414 7732 18420 7744
rect 17052 7704 18420 7732
rect 15289 7695 15347 7701
rect 18414 7692 18420 7704
rect 18472 7732 18478 7744
rect 18524 7732 18552 7828
rect 20088 7800 20116 7828
rect 21376 7800 21404 7831
rect 21542 7828 21548 7840
rect 21600 7828 21606 7880
rect 20088 7772 21404 7800
rect 18472 7704 18552 7732
rect 18472 7692 18478 7704
rect 19978 7692 19984 7744
rect 20036 7732 20042 7744
rect 20901 7735 20959 7741
rect 20036 7704 20081 7732
rect 20036 7692 20042 7704
rect 20901 7701 20913 7735
rect 20947 7732 20959 7735
rect 21634 7732 21640 7744
rect 20947 7704 21640 7732
rect 20947 7701 20959 7704
rect 20901 7695 20959 7701
rect 21634 7692 21640 7704
rect 21692 7692 21698 7744
rect 22097 7735 22155 7741
rect 22097 7701 22109 7735
rect 22143 7732 22155 7735
rect 22370 7732 22376 7744
rect 22143 7704 22376 7732
rect 22143 7701 22155 7704
rect 22097 7695 22155 7701
rect 22370 7692 22376 7704
rect 22428 7692 22434 7744
rect 1104 7642 22816 7664
rect 1104 7590 4614 7642
rect 4666 7590 4678 7642
rect 4730 7590 4742 7642
rect 4794 7590 4806 7642
rect 4858 7590 11878 7642
rect 11930 7590 11942 7642
rect 11994 7590 12006 7642
rect 12058 7590 12070 7642
rect 12122 7590 19142 7642
rect 19194 7590 19206 7642
rect 19258 7590 19270 7642
rect 19322 7590 19334 7642
rect 19386 7590 22816 7642
rect 1104 7568 22816 7590
rect 5721 7531 5779 7537
rect 5721 7497 5733 7531
rect 5767 7528 5779 7531
rect 6730 7528 6736 7540
rect 5767 7500 6736 7528
rect 5767 7497 5779 7500
rect 5721 7491 5779 7497
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7193 7531 7251 7537
rect 7193 7528 7205 7531
rect 7064 7500 7205 7528
rect 7064 7488 7070 7500
rect 7193 7497 7205 7500
rect 7239 7497 7251 7531
rect 9582 7528 9588 7540
rect 7193 7491 7251 7497
rect 7668 7500 9444 7528
rect 9543 7500 9588 7528
rect 7558 7460 7564 7472
rect 5276 7432 7564 7460
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7324 5135 7327
rect 5276 7324 5304 7432
rect 7558 7420 7564 7432
rect 7616 7420 7622 7472
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7392 5411 7395
rect 6178 7392 6184 7404
rect 5399 7364 6040 7392
rect 6139 7364 6184 7392
rect 5399 7361 5411 7364
rect 5353 7355 5411 7361
rect 5123 7296 5304 7324
rect 5123 7293 5135 7296
rect 5077 7287 5135 7293
rect 4246 7256 4252 7268
rect 4207 7228 4252 7256
rect 4246 7216 4252 7228
rect 4304 7216 4310 7268
rect 5169 7259 5227 7265
rect 5169 7225 5181 7259
rect 5215 7256 5227 7259
rect 5258 7256 5264 7268
rect 5215 7228 5264 7256
rect 5215 7225 5227 7228
rect 5169 7219 5227 7225
rect 5258 7216 5264 7228
rect 5316 7216 5322 7268
rect 4706 7188 4712 7200
rect 4667 7160 4712 7188
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 6012 7188 6040 7364
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6362 7392 6368 7404
rect 6323 7364 6368 7392
rect 6362 7352 6368 7364
rect 6420 7352 6426 7404
rect 7668 7401 7696 7500
rect 9416 7460 9444 7500
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 9674 7488 9680 7540
rect 9732 7528 9738 7540
rect 10410 7528 10416 7540
rect 9732 7500 10416 7528
rect 9732 7488 9738 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 12250 7528 12256 7540
rect 10888 7500 12256 7528
rect 10888 7460 10916 7500
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 12483 7500 16129 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 16117 7497 16129 7500
rect 16163 7497 16175 7531
rect 16390 7528 16396 7540
rect 16351 7500 16396 7528
rect 16117 7491 16175 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 19610 7528 19616 7540
rect 18156 7500 19616 7528
rect 9416 7432 10916 7460
rect 10965 7463 11023 7469
rect 10965 7429 10977 7463
rect 11011 7460 11023 7463
rect 12710 7460 12716 7472
rect 11011 7432 12716 7460
rect 11011 7429 11023 7432
rect 10965 7423 11023 7429
rect 12710 7420 12716 7432
rect 12768 7420 12774 7472
rect 13906 7460 13912 7472
rect 12820 7432 13912 7460
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 7883 7364 8340 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 7561 7327 7619 7333
rect 7561 7293 7573 7327
rect 7607 7324 7619 7327
rect 7742 7324 7748 7336
rect 7607 7296 7748 7324
rect 7607 7293 7619 7296
rect 7561 7287 7619 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 7984 7296 8217 7324
rect 7984 7284 7990 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8312 7324 8340 7364
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 10100 7364 10333 7392
rect 10100 7352 10106 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10410 7352 10416 7404
rect 10468 7392 10474 7404
rect 11514 7392 11520 7404
rect 10468 7364 10513 7392
rect 11475 7364 11520 7392
rect 10468 7352 10474 7364
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 12820 7392 12848 7432
rect 13906 7420 13912 7432
rect 13964 7420 13970 7472
rect 15470 7420 15476 7472
rect 15528 7460 15534 7472
rect 15930 7460 15936 7472
rect 15528 7432 15936 7460
rect 15528 7420 15534 7432
rect 15930 7420 15936 7432
rect 15988 7420 15994 7472
rect 16025 7463 16083 7469
rect 16025 7429 16037 7463
rect 16071 7460 16083 7463
rect 16298 7460 16304 7472
rect 16071 7432 16304 7460
rect 16071 7429 16083 7432
rect 16025 7423 16083 7429
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 12986 7392 12992 7404
rect 11624 7364 12848 7392
rect 12947 7364 12992 7392
rect 11624 7324 11652 7364
rect 12986 7352 12992 7364
rect 13044 7352 13050 7404
rect 13262 7352 13268 7404
rect 13320 7392 13326 7404
rect 14556 7395 14614 7401
rect 14556 7392 14568 7395
rect 13320 7364 14568 7392
rect 13320 7352 13326 7364
rect 14556 7361 14568 7364
rect 14602 7361 14614 7395
rect 14556 7355 14614 7361
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 14792 7364 16335 7392
rect 14792 7352 14798 7364
rect 8312 7296 11652 7324
rect 8205 7287 8263 7293
rect 11698 7284 11704 7336
rect 11756 7324 11762 7336
rect 12158 7324 12164 7336
rect 11756 7296 12164 7324
rect 11756 7284 11762 7296
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12342 7324 12348 7336
rect 12299 7296 12348 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 13449 7327 13507 7333
rect 13449 7324 13461 7327
rect 12860 7296 13461 7324
rect 12860 7284 12866 7296
rect 13449 7293 13461 7296
rect 13495 7293 13507 7327
rect 13449 7287 13507 7293
rect 13630 7284 13636 7336
rect 13688 7324 13694 7336
rect 13688 7296 13952 7324
rect 13688 7284 13694 7296
rect 6089 7259 6147 7265
rect 6089 7225 6101 7259
rect 6135 7256 6147 7259
rect 8110 7256 8116 7268
rect 6135 7228 8116 7256
rect 6135 7225 6147 7228
rect 6089 7219 6147 7225
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 8472 7259 8530 7265
rect 8472 7225 8484 7259
rect 8518 7256 8530 7259
rect 8570 7256 8576 7268
rect 8518 7228 8576 7256
rect 8518 7225 8530 7228
rect 8472 7219 8530 7225
rect 8570 7216 8576 7228
rect 8628 7216 8634 7268
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 10229 7259 10287 7265
rect 9548 7228 10180 7256
rect 9548 7216 9554 7228
rect 7558 7188 7564 7200
rect 6012 7160 7564 7188
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 9861 7191 9919 7197
rect 9861 7157 9873 7191
rect 9907 7188 9919 7191
rect 10042 7188 10048 7200
rect 9907 7160 10048 7188
rect 9907 7157 9919 7160
rect 9861 7151 9919 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 10152 7188 10180 7228
rect 10229 7225 10241 7259
rect 10275 7256 10287 7259
rect 10870 7256 10876 7268
rect 10275 7228 10876 7256
rect 10275 7225 10287 7228
rect 10229 7219 10287 7225
rect 10870 7216 10876 7228
rect 10928 7216 10934 7268
rect 11425 7259 11483 7265
rect 11425 7225 11437 7259
rect 11471 7256 11483 7259
rect 13924 7256 13952 7296
rect 13998 7284 14004 7336
rect 14056 7324 14062 7336
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 14056 7296 14105 7324
rect 14056 7284 14062 7296
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14829 7327 14887 7333
rect 14829 7324 14841 7327
rect 14093 7287 14151 7293
rect 14200 7296 14841 7324
rect 14200 7256 14228 7296
rect 14829 7293 14841 7296
rect 14875 7324 14887 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 14875 7296 16037 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16025 7287 16083 7293
rect 16117 7327 16175 7333
rect 16117 7293 16129 7327
rect 16163 7324 16175 7327
rect 16209 7327 16267 7333
rect 16209 7324 16221 7327
rect 16163 7296 16221 7324
rect 16163 7293 16175 7296
rect 16117 7287 16175 7293
rect 16209 7293 16221 7296
rect 16255 7293 16267 7327
rect 16307 7324 16335 7364
rect 16850 7352 16856 7404
rect 16908 7392 16914 7404
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 16908 7364 17509 7392
rect 16908 7352 16914 7364
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 18156 7333 18184 7500
rect 19610 7488 19616 7500
rect 19668 7488 19674 7540
rect 20346 7488 20352 7540
rect 20404 7528 20410 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 20404 7500 21189 7528
rect 20404 7488 20410 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 20070 7420 20076 7472
rect 20128 7460 20134 7472
rect 20533 7463 20591 7469
rect 20533 7460 20545 7463
rect 20128 7432 20545 7460
rect 20128 7420 20134 7432
rect 20533 7429 20545 7432
rect 20579 7429 20591 7463
rect 20533 7423 20591 7429
rect 19199 7395 19257 7401
rect 19199 7361 19211 7395
rect 19245 7361 19257 7395
rect 19426 7392 19432 7404
rect 19339 7364 19432 7392
rect 19199 7355 19257 7361
rect 17313 7327 17371 7333
rect 17313 7324 17325 7327
rect 16307 7296 17325 7324
rect 16209 7287 16267 7293
rect 17313 7293 17325 7296
rect 17359 7293 17371 7327
rect 17313 7287 17371 7293
rect 18141 7327 18199 7333
rect 18141 7293 18153 7327
rect 18187 7293 18199 7327
rect 18141 7287 18199 7293
rect 18693 7327 18751 7333
rect 18693 7293 18705 7327
rect 18739 7293 18751 7327
rect 18693 7287 18751 7293
rect 17405 7259 17463 7265
rect 17405 7256 17417 7259
rect 11471 7228 13676 7256
rect 13924 7228 14228 7256
rect 15488 7228 17417 7256
rect 11471 7225 11483 7228
rect 11425 7219 11483 7225
rect 10410 7188 10416 7200
rect 10152 7160 10416 7188
rect 10410 7148 10416 7160
rect 10468 7148 10474 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11112 7160 11345 7188
rect 11112 7148 11118 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 12069 7191 12127 7197
rect 12069 7157 12081 7191
rect 12115 7188 12127 7191
rect 12618 7188 12624 7200
rect 12115 7160 12624 7188
rect 12115 7157 12127 7160
rect 12069 7151 12127 7157
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 12805 7191 12863 7197
rect 12805 7188 12817 7191
rect 12768 7160 12817 7188
rect 12768 7148 12774 7160
rect 12805 7157 12817 7160
rect 12851 7157 12863 7191
rect 12805 7151 12863 7157
rect 12897 7191 12955 7197
rect 12897 7157 12909 7191
rect 12943 7188 12955 7191
rect 13170 7188 13176 7200
rect 12943 7160 13176 7188
rect 12943 7157 12955 7160
rect 12897 7151 12955 7157
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13648 7197 13676 7228
rect 13633 7191 13691 7197
rect 13633 7157 13645 7191
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 14550 7148 14556 7200
rect 14608 7197 14614 7200
rect 14608 7188 14617 7197
rect 14608 7160 14653 7188
rect 14608 7151 14617 7160
rect 14608 7148 14614 7151
rect 14826 7148 14832 7200
rect 14884 7188 14890 7200
rect 15488 7188 15516 7228
rect 17405 7225 17417 7228
rect 17451 7225 17463 7259
rect 17405 7219 17463 7225
rect 18046 7216 18052 7268
rect 18104 7256 18110 7268
rect 18708 7256 18736 7287
rect 18782 7284 18788 7336
rect 18840 7324 18846 7336
rect 19016 7327 19074 7333
rect 19016 7324 19028 7327
rect 18840 7296 19028 7324
rect 18840 7284 18846 7296
rect 19016 7293 19028 7296
rect 19062 7293 19074 7327
rect 19214 7324 19242 7355
rect 19426 7352 19432 7364
rect 19484 7392 19490 7404
rect 20438 7392 20444 7404
rect 19484 7364 20444 7392
rect 19484 7352 19490 7364
rect 20438 7352 20444 7364
rect 20496 7352 20502 7404
rect 21726 7392 21732 7404
rect 21687 7364 21732 7392
rect 21726 7352 21732 7364
rect 21784 7352 21790 7404
rect 20254 7324 20260 7336
rect 19214 7296 20260 7324
rect 19016 7287 19074 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 21634 7324 21640 7336
rect 21595 7296 21640 7324
rect 21634 7284 21640 7296
rect 21692 7284 21698 7336
rect 18104 7228 18736 7256
rect 18104 7216 18110 7228
rect 16942 7188 16948 7200
rect 14884 7160 15516 7188
rect 16903 7160 16948 7188
rect 14884 7148 14890 7160
rect 16942 7148 16948 7160
rect 17000 7148 17006 7200
rect 18325 7191 18383 7197
rect 18325 7157 18337 7191
rect 18371 7188 18383 7191
rect 18966 7188 18972 7200
rect 18371 7160 18972 7188
rect 18371 7157 18383 7160
rect 18325 7151 18383 7157
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 19794 7148 19800 7200
rect 19852 7188 19858 7200
rect 20070 7188 20076 7200
rect 19852 7160 20076 7188
rect 19852 7148 19858 7160
rect 20070 7148 20076 7160
rect 20128 7148 20134 7200
rect 20898 7148 20904 7200
rect 20956 7188 20962 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 20956 7160 21557 7188
rect 20956 7148 20962 7160
rect 21545 7157 21557 7160
rect 21591 7157 21603 7191
rect 21545 7151 21603 7157
rect 1104 7098 22816 7120
rect 1104 7046 8246 7098
rect 8298 7046 8310 7098
rect 8362 7046 8374 7098
rect 8426 7046 8438 7098
rect 8490 7046 15510 7098
rect 15562 7046 15574 7098
rect 15626 7046 15638 7098
rect 15690 7046 15702 7098
rect 15754 7046 22816 7098
rect 1104 7024 22816 7046
rect 6825 6987 6883 6993
rect 6825 6953 6837 6987
rect 6871 6984 6883 6987
rect 7282 6984 7288 6996
rect 6871 6956 7288 6984
rect 6871 6953 6883 6956
rect 6825 6947 6883 6953
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 9674 6984 9680 6996
rect 7616 6956 9680 6984
rect 7616 6944 7622 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 10042 6984 10048 6996
rect 10003 6956 10048 6984
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 12250 6984 12256 6996
rect 11164 6956 12256 6984
rect 7374 6876 7380 6928
rect 7432 6916 7438 6928
rect 11164 6916 11192 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12345 6987 12403 6993
rect 12345 6953 12357 6987
rect 12391 6984 12403 6987
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12391 6956 13093 6984
rect 12391 6953 12403 6956
rect 12345 6947 12403 6953
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 16574 6984 16580 6996
rect 13081 6947 13139 6953
rect 13188 6956 16580 6984
rect 7432 6888 11192 6916
rect 11241 6919 11299 6925
rect 7432 6876 7438 6888
rect 11241 6885 11253 6919
rect 11287 6916 11299 6919
rect 12158 6916 12164 6928
rect 11287 6888 12164 6916
rect 11287 6885 11299 6888
rect 11241 6879 11299 6885
rect 12158 6876 12164 6888
rect 12216 6876 12222 6928
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 13188 6916 13216 6956
rect 16574 6944 16580 6956
rect 16632 6944 16638 6996
rect 17402 6984 17408 6996
rect 17144 6956 17408 6984
rect 15534 6919 15592 6925
rect 15534 6916 15546 6919
rect 12768 6888 13216 6916
rect 13464 6888 15546 6916
rect 12768 6876 12774 6888
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 6089 6851 6147 6857
rect 6089 6848 6101 6851
rect 5491 6820 6101 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 6089 6817 6101 6820
rect 6135 6817 6147 6851
rect 7650 6848 7656 6860
rect 6089 6811 6147 6817
rect 6380 6820 7656 6848
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 6380 6789 6408 6820
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8196 6851 8254 6857
rect 8196 6817 8208 6851
rect 8242 6848 8254 6851
rect 9214 6848 9220 6860
rect 8242 6820 9220 6848
rect 8242 6817 8254 6820
rect 8196 6811 8254 6817
rect 9214 6808 9220 6820
rect 9272 6808 9278 6860
rect 9766 6808 9772 6860
rect 9824 6848 9830 6860
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 9824 6820 10149 6848
rect 9824 6808 9830 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10137 6811 10195 6817
rect 10336 6820 11560 6848
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 4396 6752 6193 6780
rect 4396 6740 4402 6752
rect 6181 6749 6193 6752
rect 6227 6749 6239 6783
rect 6181 6743 6239 6749
rect 6365 6783 6423 6789
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 7377 6743 7435 6749
rect 5721 6715 5779 6721
rect 5721 6681 5733 6715
rect 5767 6712 5779 6715
rect 6546 6712 6552 6724
rect 5767 6684 6552 6712
rect 5767 6681 5779 6684
rect 5721 6675 5779 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 7392 6712 7420 6743
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7926 6780 7932 6792
rect 7887 6752 7932 6780
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 9858 6740 9864 6792
rect 9916 6780 9922 6792
rect 10336 6789 10364 6820
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 9916 6752 10333 6780
rect 9916 6740 9922 6752
rect 10321 6749 10333 6752
rect 10367 6749 10379 6783
rect 11330 6780 11336 6792
rect 11291 6752 11336 6780
rect 10321 6743 10379 6749
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11532 6789 11560 6820
rect 11606 6808 11612 6860
rect 11664 6848 11670 6860
rect 11664 6820 12204 6848
rect 11664 6808 11670 6820
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 12066 6780 12072 6792
rect 11563 6752 12072 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 12066 6740 12072 6752
rect 12124 6740 12130 6792
rect 12176 6780 12204 6820
rect 12250 6808 12256 6860
rect 12308 6848 12314 6860
rect 12894 6848 12900 6860
rect 12308 6820 12353 6848
rect 12855 6820 12900 6848
rect 12308 6808 12314 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 12437 6783 12495 6789
rect 12437 6780 12449 6783
rect 12176 6752 12449 6780
rect 12437 6749 12449 6752
rect 12483 6749 12495 6783
rect 12437 6743 12495 6749
rect 12526 6740 12532 6792
rect 12584 6780 12590 6792
rect 13464 6780 13492 6888
rect 15534 6885 15546 6888
rect 15580 6916 15592 6919
rect 17144 6916 17172 6956
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 17503 6987 17561 6993
rect 17503 6953 17515 6987
rect 17549 6984 17561 6987
rect 18782 6984 18788 6996
rect 17549 6956 18788 6984
rect 17549 6953 17561 6956
rect 17503 6947 17561 6953
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 15580 6888 17172 6916
rect 19420 6919 19478 6925
rect 15580 6885 15592 6888
rect 15534 6879 15592 6885
rect 19420 6885 19432 6919
rect 19466 6916 19478 6919
rect 19794 6916 19800 6928
rect 19466 6888 19800 6916
rect 19466 6885 19478 6888
rect 19420 6879 19478 6885
rect 19794 6876 19800 6888
rect 19852 6916 19858 6928
rect 20530 6916 20536 6928
rect 19852 6888 20536 6916
rect 19852 6876 19858 6888
rect 20530 6876 20536 6888
rect 20588 6876 20594 6928
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13630 6848 13636 6860
rect 13587 6820 13636 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 13808 6851 13866 6857
rect 13808 6817 13820 6851
rect 13854 6848 13866 6851
rect 13854 6820 15148 6848
rect 13854 6817 13866 6820
rect 13808 6811 13866 6817
rect 12584 6752 13492 6780
rect 12584 6740 12590 6752
rect 7742 6712 7748 6724
rect 7392 6684 7748 6712
rect 7742 6672 7748 6684
rect 7800 6672 7806 6724
rect 11885 6715 11943 6721
rect 9140 6684 11468 6712
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 9140 6644 9168 6684
rect 9306 6644 9312 6656
rect 6963 6616 9168 6644
rect 9267 6616 9312 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 10042 6644 10048 6656
rect 9723 6616 10048 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 10870 6644 10876 6656
rect 10831 6616 10876 6644
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 11440 6644 11468 6684
rect 11885 6681 11897 6715
rect 11931 6712 11943 6715
rect 13170 6712 13176 6724
rect 11931 6684 13176 6712
rect 11931 6681 11943 6684
rect 11885 6675 11943 6681
rect 13170 6672 13176 6684
rect 13228 6672 13234 6724
rect 13078 6644 13084 6656
rect 11440 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14642 6644 14648 6656
rect 13872 6616 14648 6644
rect 13872 6604 13878 6616
rect 14642 6604 14648 6616
rect 14700 6644 14706 6656
rect 14921 6647 14979 6653
rect 14921 6644 14933 6647
rect 14700 6616 14933 6644
rect 14700 6604 14706 6616
rect 14921 6613 14933 6616
rect 14967 6613 14979 6647
rect 15120 6644 15148 6820
rect 16942 6808 16948 6860
rect 17000 6848 17006 6860
rect 17000 6820 17540 6848
rect 17000 6808 17006 6820
rect 15194 6740 15200 6792
rect 15252 6780 15258 6792
rect 15289 6783 15347 6789
rect 15289 6780 15301 6783
rect 15252 6752 15301 6780
rect 15252 6740 15258 6752
rect 15289 6749 15301 6752
rect 15335 6749 15347 6783
rect 15289 6743 15347 6749
rect 16666 6740 16672 6792
rect 16724 6780 16730 6792
rect 17512 6789 17540 6820
rect 17678 6808 17684 6860
rect 17736 6848 17742 6860
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 17736 6820 17785 6848
rect 17736 6808 17742 6820
rect 17773 6817 17785 6820
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 18690 6808 18696 6860
rect 18748 6848 18754 6860
rect 19153 6851 19211 6857
rect 19153 6848 19165 6851
rect 18748 6820 19165 6848
rect 18748 6808 18754 6820
rect 19153 6817 19165 6820
rect 19199 6848 19211 6851
rect 20625 6851 20683 6857
rect 19199 6820 20300 6848
rect 19199 6817 19211 6820
rect 19153 6811 19211 6817
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16724 6752 17049 6780
rect 16724 6740 16730 6752
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 17500 6783 17558 6789
rect 17500 6749 17512 6783
rect 17546 6749 17558 6783
rect 20272 6780 20300 6820
rect 20625 6817 20637 6851
rect 20671 6848 20683 6851
rect 21157 6851 21215 6857
rect 21157 6848 21169 6851
rect 20671 6820 21169 6848
rect 20671 6817 20683 6820
rect 20625 6811 20683 6817
rect 21157 6817 21169 6820
rect 21203 6817 21215 6851
rect 21157 6811 21215 6817
rect 20714 6780 20720 6792
rect 20272 6752 20720 6780
rect 17500 6743 17558 6749
rect 20714 6740 20720 6752
rect 20772 6780 20778 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20772 6752 20913 6780
rect 20772 6740 20778 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 16850 6712 16856 6724
rect 16316 6684 16856 6712
rect 16316 6644 16344 6684
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 15120 6616 16344 6644
rect 14921 6607 14979 6613
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 16669 6647 16727 6653
rect 16669 6644 16681 6647
rect 16448 6616 16681 6644
rect 16448 6604 16454 6616
rect 16669 6613 16681 6616
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 18877 6647 18935 6653
rect 18877 6613 18889 6647
rect 18923 6644 18935 6647
rect 19426 6644 19432 6656
rect 18923 6616 19432 6644
rect 18923 6613 18935 6616
rect 18877 6607 18935 6613
rect 19426 6604 19432 6616
rect 19484 6604 19490 6656
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 20346 6644 20352 6656
rect 20128 6616 20352 6644
rect 20128 6604 20134 6616
rect 20346 6604 20352 6616
rect 20404 6604 20410 6656
rect 20530 6644 20536 6656
rect 20491 6616 20536 6644
rect 20530 6604 20536 6616
rect 20588 6644 20594 6656
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20588 6616 20637 6644
rect 20588 6604 20594 6616
rect 20625 6613 20637 6616
rect 20671 6613 20683 6647
rect 20625 6607 20683 6613
rect 21634 6604 21640 6656
rect 21692 6644 21698 6656
rect 22281 6647 22339 6653
rect 22281 6644 22293 6647
rect 21692 6616 22293 6644
rect 21692 6604 21698 6616
rect 22281 6613 22293 6616
rect 22327 6613 22339 6647
rect 22281 6607 22339 6613
rect 1104 6554 22816 6576
rect 1104 6502 4614 6554
rect 4666 6502 4678 6554
rect 4730 6502 4742 6554
rect 4794 6502 4806 6554
rect 4858 6502 11878 6554
rect 11930 6502 11942 6554
rect 11994 6502 12006 6554
rect 12058 6502 12070 6554
rect 12122 6502 19142 6554
rect 19194 6502 19206 6554
rect 19258 6502 19270 6554
rect 19322 6502 19334 6554
rect 19386 6502 22816 6554
rect 1104 6480 22816 6502
rect 8570 6440 8576 6452
rect 8220 6412 8576 6440
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 8018 6372 8024 6384
rect 3108 6344 8024 6372
rect 3108 6332 3114 6344
rect 8018 6332 8024 6344
rect 8076 6332 8082 6384
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6304 6331 6307
rect 7098 6304 7104 6316
rect 6319 6276 7104 6304
rect 6319 6273 6331 6276
rect 6273 6267 6331 6273
rect 7098 6264 7104 6276
rect 7156 6264 7162 6316
rect 7929 6307 7987 6313
rect 7929 6273 7941 6307
rect 7975 6304 7987 6307
rect 8110 6304 8116 6316
rect 7975 6276 8116 6304
rect 7975 6273 7987 6276
rect 7929 6267 7987 6273
rect 8110 6264 8116 6276
rect 8168 6264 8174 6316
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 8220 6236 8248 6412
rect 8570 6400 8576 6412
rect 8628 6440 8634 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 8628 6412 9689 6440
rect 8628 6400 8634 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 10870 6400 10876 6452
rect 10928 6440 10934 6452
rect 11698 6440 11704 6452
rect 10928 6412 11704 6440
rect 10928 6400 10934 6412
rect 11698 6400 11704 6412
rect 11756 6400 11762 6452
rect 12250 6400 12256 6452
rect 12308 6440 12314 6452
rect 12621 6443 12679 6449
rect 12621 6440 12633 6443
rect 12308 6412 12633 6440
rect 12308 6400 12314 6412
rect 12621 6409 12633 6412
rect 12667 6409 12679 6443
rect 12621 6403 12679 6409
rect 12894 6400 12900 6452
rect 12952 6440 12958 6452
rect 14737 6443 14795 6449
rect 14737 6440 14749 6443
rect 12952 6412 14749 6440
rect 12952 6400 12958 6412
rect 14737 6409 14749 6412
rect 14783 6409 14795 6443
rect 14737 6403 14795 6409
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 15933 6443 15991 6449
rect 15933 6440 15945 6443
rect 15344 6412 15945 6440
rect 15344 6400 15350 6412
rect 15933 6409 15945 6412
rect 15979 6440 15991 6443
rect 16114 6440 16120 6452
rect 15979 6412 16120 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16114 6400 16120 6412
rect 16172 6400 16178 6452
rect 19794 6440 19800 6452
rect 16224 6412 19380 6440
rect 19755 6412 19800 6440
rect 13078 6372 13084 6384
rect 11716 6344 13084 6372
rect 11716 6304 11744 6344
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 14090 6332 14096 6384
rect 14148 6372 14154 6384
rect 16224 6372 16252 6412
rect 14148 6344 16252 6372
rect 19352 6372 19380 6412
rect 19794 6400 19800 6412
rect 19852 6400 19858 6452
rect 20254 6440 20260 6452
rect 20215 6412 20260 6440
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 20898 6440 20904 6452
rect 20364 6412 20904 6440
rect 20364 6372 20392 6412
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 19352 6344 20392 6372
rect 14148 6332 14154 6344
rect 11624 6276 11744 6304
rect 7699 6208 8248 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 8564 6239 8622 6245
rect 8564 6236 8576 6239
rect 8352 6208 8397 6236
rect 8496 6208 8576 6236
rect 8352 6196 8358 6208
rect 7745 6171 7803 6177
rect 7745 6137 7757 6171
rect 7791 6168 7803 6171
rect 8496 6168 8524 6208
rect 8564 6205 8576 6208
rect 8610 6236 8622 6239
rect 9306 6236 9312 6248
rect 8610 6208 9312 6236
rect 8610 6205 8622 6208
rect 8564 6199 8622 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 10042 6236 10048 6248
rect 10003 6208 10048 6236
rect 10042 6196 10048 6208
rect 10100 6196 10106 6248
rect 10502 6196 10508 6248
rect 10560 6236 10566 6248
rect 10597 6239 10655 6245
rect 10597 6236 10609 6239
rect 10560 6208 10609 6236
rect 10560 6196 10566 6208
rect 10597 6205 10609 6208
rect 10643 6205 10655 6239
rect 11624 6236 11652 6276
rect 11790 6264 11796 6316
rect 11848 6304 11854 6316
rect 11848 6276 13216 6304
rect 11848 6264 11854 6276
rect 10597 6199 10655 6205
rect 10704 6208 11652 6236
rect 10704 6168 10732 6208
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 12437 6239 12495 6245
rect 12437 6236 12449 6239
rect 11756 6208 12449 6236
rect 11756 6196 11762 6208
rect 12437 6205 12449 6208
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13188 6236 13216 6276
rect 14274 6264 14280 6316
rect 14332 6304 14338 6316
rect 14826 6304 14832 6316
rect 14332 6276 14832 6304
rect 14332 6264 14338 6276
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 15102 6264 15108 6316
rect 15160 6304 15166 6316
rect 15289 6307 15347 6313
rect 15289 6304 15301 6307
rect 15160 6276 15301 6304
rect 15160 6264 15166 6276
rect 15289 6273 15301 6276
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 18309 6276 18552 6304
rect 15749 6239 15807 6245
rect 15749 6236 15761 6239
rect 13188 6208 15761 6236
rect 13081 6199 13139 6205
rect 15749 6205 15761 6208
rect 15795 6205 15807 6239
rect 16298 6236 16304 6248
rect 16259 6208 16304 6236
rect 15749 6199 15807 6205
rect 7791 6140 8524 6168
rect 8588 6140 10732 6168
rect 10864 6171 10922 6177
rect 7791 6137 7803 6140
rect 7745 6131 7803 6137
rect 6822 6100 6828 6112
rect 6783 6072 6828 6100
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 7282 6100 7288 6112
rect 7243 6072 7288 6100
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 8588 6100 8616 6140
rect 10864 6137 10876 6171
rect 10910 6168 10922 6171
rect 11514 6168 11520 6180
rect 10910 6140 11520 6168
rect 10910 6137 10922 6140
rect 10864 6131 10922 6137
rect 11514 6128 11520 6140
rect 11572 6128 11578 6180
rect 7616 6072 8616 6100
rect 10229 6103 10287 6109
rect 7616 6060 7622 6072
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 11054 6100 11060 6112
rect 10275 6072 11060 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11977 6103 12035 6109
rect 11977 6100 11989 6103
rect 11296 6072 11989 6100
rect 11296 6060 11302 6072
rect 11977 6069 11989 6072
rect 12023 6069 12035 6103
rect 11977 6063 12035 6069
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13096 6100 13124 6199
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 18309 6236 18337 6276
rect 18414 6236 18420 6248
rect 16500 6208 18337 6236
rect 18375 6208 18420 6236
rect 13348 6171 13406 6177
rect 13348 6137 13360 6171
rect 13394 6168 13406 6171
rect 13814 6168 13820 6180
rect 13394 6140 13820 6168
rect 13394 6137 13406 6140
rect 13348 6131 13406 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 15197 6171 15255 6177
rect 15197 6168 15209 6171
rect 14240 6140 15209 6168
rect 14240 6128 14246 6140
rect 15197 6137 15209 6140
rect 15243 6137 15255 6171
rect 15197 6131 15255 6137
rect 15930 6128 15936 6180
rect 15988 6168 15994 6180
rect 16500 6168 16528 6208
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18524 6236 18552 6276
rect 19702 6236 19708 6248
rect 18524 6208 19708 6236
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 20070 6236 20076 6248
rect 20031 6208 20076 6236
rect 20070 6196 20076 6208
rect 20128 6196 20134 6248
rect 20625 6239 20683 6245
rect 20625 6205 20637 6239
rect 20671 6236 20683 6239
rect 20714 6236 20720 6248
rect 20671 6208 20720 6236
rect 20671 6205 20683 6208
rect 20625 6199 20683 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 20892 6239 20950 6245
rect 20892 6205 20904 6239
rect 20938 6236 20950 6239
rect 21634 6236 21640 6248
rect 20938 6208 21640 6236
rect 20938 6205 20950 6208
rect 20892 6199 20950 6205
rect 21634 6196 21640 6208
rect 21692 6196 21698 6248
rect 15988 6140 16528 6168
rect 16568 6171 16626 6177
rect 15988 6128 15994 6140
rect 16568 6137 16580 6171
rect 16614 6168 16626 6171
rect 18684 6171 18742 6177
rect 16614 6140 18644 6168
rect 16614 6137 16626 6140
rect 16568 6131 16626 6137
rect 13722 6100 13728 6112
rect 13044 6072 13728 6100
rect 13044 6060 13050 6072
rect 13722 6060 13728 6072
rect 13780 6060 13786 6112
rect 14458 6100 14464 6112
rect 14419 6072 14464 6100
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15102 6100 15108 6112
rect 15063 6072 15108 6100
rect 15102 6060 15108 6072
rect 15160 6060 15166 6112
rect 17678 6100 17684 6112
rect 17639 6072 17684 6100
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 18616 6100 18644 6140
rect 18684 6137 18696 6171
rect 18730 6168 18742 6171
rect 19426 6168 19432 6180
rect 18730 6140 19432 6168
rect 18730 6137 18742 6140
rect 18684 6131 18742 6137
rect 19426 6128 19432 6140
rect 19484 6128 19490 6180
rect 21726 6100 21732 6112
rect 18616 6072 21732 6100
rect 21726 6060 21732 6072
rect 21784 6100 21790 6112
rect 22005 6103 22063 6109
rect 22005 6100 22017 6103
rect 21784 6072 22017 6100
rect 21784 6060 21790 6072
rect 22005 6069 22017 6072
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 1104 6010 22816 6032
rect 1104 5958 8246 6010
rect 8298 5958 8310 6010
rect 8362 5958 8374 6010
rect 8426 5958 8438 6010
rect 8490 5958 15510 6010
rect 15562 5958 15574 6010
rect 15626 5958 15638 6010
rect 15690 5958 15702 6010
rect 15754 5958 22816 6010
rect 1104 5936 22816 5958
rect 6270 5856 6276 5908
rect 6328 5896 6334 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 6328 5868 6929 5896
rect 6328 5856 6334 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 10045 5899 10103 5905
rect 10045 5896 10057 5899
rect 7340 5868 10057 5896
rect 7340 5856 7346 5868
rect 10045 5865 10057 5868
rect 10091 5865 10103 5899
rect 13814 5896 13820 5908
rect 10045 5859 10103 5865
rect 10152 5868 13820 5896
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 10152 5828 10180 5868
rect 13814 5856 13820 5868
rect 13872 5856 13878 5908
rect 13906 5856 13912 5908
rect 13964 5896 13970 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 13964 5868 14841 5896
rect 13964 5856 13970 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 16850 5856 16856 5908
rect 16908 5896 16914 5908
rect 17497 5899 17555 5905
rect 17497 5896 17509 5899
rect 16908 5868 17509 5896
rect 16908 5856 16914 5868
rect 17497 5865 17509 5868
rect 17543 5865 17555 5899
rect 17497 5859 17555 5865
rect 19978 5856 19984 5908
rect 20036 5896 20042 5908
rect 20257 5899 20315 5905
rect 20257 5896 20269 5899
rect 20036 5868 20269 5896
rect 20036 5856 20042 5868
rect 20257 5865 20269 5868
rect 20303 5865 20315 5899
rect 20257 5859 20315 5865
rect 12250 5828 12256 5840
rect 6880 5800 10180 5828
rect 10327 5800 12256 5828
rect 6880 5788 6886 5800
rect 7190 5720 7196 5772
rect 7248 5760 7254 5772
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 7248 5732 7297 5760
rect 7248 5720 7254 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7377 5763 7435 5769
rect 7377 5729 7389 5763
rect 7423 5760 7435 5763
rect 8018 5760 8024 5772
rect 7423 5732 8024 5760
rect 7423 5729 7435 5732
rect 7377 5723 7435 5729
rect 8018 5720 8024 5732
rect 8076 5720 8082 5772
rect 8196 5763 8254 5769
rect 8196 5729 8208 5763
rect 8242 5760 8254 5763
rect 9582 5760 9588 5772
rect 8242 5732 9588 5760
rect 8242 5729 8254 5732
rect 8196 5723 8254 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 9916 5732 10272 5760
rect 9916 5720 9922 5732
rect 7561 5695 7619 5701
rect 7561 5661 7573 5695
rect 7607 5692 7619 5695
rect 7607 5664 7880 5692
rect 7607 5661 7619 5664
rect 7561 5655 7619 5661
rect 7852 5556 7880 5664
rect 7926 5652 7932 5704
rect 7984 5692 7990 5704
rect 7984 5664 8029 5692
rect 7984 5652 7990 5664
rect 9122 5652 9128 5704
rect 9180 5692 9186 5704
rect 10244 5701 10272 5732
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9180 5664 10149 5692
rect 9180 5652 9186 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10229 5695 10287 5701
rect 10229 5661 10241 5695
rect 10275 5661 10287 5695
rect 10229 5655 10287 5661
rect 10327 5624 10355 5800
rect 12250 5788 12256 5800
rect 12308 5788 12314 5840
rect 12434 5788 12440 5840
rect 12492 5828 12498 5840
rect 18785 5831 18843 5837
rect 18785 5828 18797 5831
rect 12492 5800 18797 5828
rect 12492 5788 12498 5800
rect 18785 5797 18797 5800
rect 18831 5797 18843 5831
rect 18785 5791 18843 5797
rect 11232 5763 11290 5769
rect 11232 5729 11244 5763
rect 11278 5760 11290 5763
rect 11698 5760 11704 5772
rect 11278 5732 11704 5760
rect 11278 5729 11290 5732
rect 11232 5723 11290 5729
rect 11698 5720 11704 5732
rect 11756 5720 11762 5772
rect 12618 5720 12624 5772
rect 12676 5760 12682 5772
rect 12897 5763 12955 5769
rect 12897 5760 12909 5763
rect 12676 5732 12909 5760
rect 12676 5720 12682 5732
rect 12897 5729 12909 5732
rect 12943 5729 12955 5763
rect 12897 5723 12955 5729
rect 12986 5720 12992 5772
rect 13044 5760 13050 5772
rect 13256 5763 13314 5769
rect 13044 5732 13089 5760
rect 13044 5720 13050 5732
rect 13256 5729 13268 5763
rect 13302 5760 13314 5763
rect 14458 5760 14464 5772
rect 13302 5732 14464 5760
rect 13302 5729 13314 5732
rect 13256 5723 13314 5729
rect 14458 5720 14464 5732
rect 14516 5720 14522 5772
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15565 5763 15623 5769
rect 15565 5729 15577 5763
rect 15611 5760 15623 5763
rect 15930 5760 15936 5772
rect 15611 5732 15936 5760
rect 15611 5729 15623 5732
rect 15565 5723 15623 5729
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 10560 5664 10977 5692
rect 10560 5652 10566 5664
rect 10965 5661 10977 5664
rect 11011 5661 11023 5695
rect 10965 5655 11023 5661
rect 12802 5624 12808 5636
rect 8864 5596 10355 5624
rect 11900 5596 12808 5624
rect 8864 5556 8892 5596
rect 7852 5528 8892 5556
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 9309 5559 9367 5565
rect 9309 5556 9321 5559
rect 9272 5528 9321 5556
rect 9272 5516 9278 5528
rect 9309 5525 9321 5528
rect 9355 5525 9367 5559
rect 9309 5519 9367 5525
rect 9677 5559 9735 5565
rect 9677 5525 9689 5559
rect 9723 5556 9735 5559
rect 11900 5556 11928 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 14660 5624 14688 5723
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16373 5763 16431 5769
rect 16373 5760 16385 5763
rect 16040 5732 16385 5760
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 16040 5692 16068 5732
rect 16373 5729 16385 5732
rect 16419 5760 16431 5763
rect 17678 5760 17684 5772
rect 16419 5732 17684 5760
rect 16419 5729 16431 5732
rect 16373 5723 16431 5729
rect 17678 5720 17684 5732
rect 17736 5720 17742 5772
rect 17862 5760 17868 5772
rect 17823 5732 17868 5760
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 20165 5763 20223 5769
rect 20165 5760 20177 5763
rect 19576 5732 20177 5760
rect 19576 5720 19582 5732
rect 20165 5729 20177 5732
rect 20211 5729 20223 5763
rect 20165 5723 20223 5729
rect 21168 5763 21226 5769
rect 21168 5729 21180 5763
rect 21214 5760 21226 5763
rect 22094 5760 22100 5772
rect 21214 5732 22100 5760
rect 21214 5729 21226 5732
rect 21168 5723 21226 5729
rect 22094 5720 22100 5732
rect 22152 5720 22158 5772
rect 14884 5664 16068 5692
rect 14884 5652 14890 5664
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 18874 5692 18880 5704
rect 16172 5664 16217 5692
rect 18835 5664 18880 5692
rect 16172 5652 16178 5664
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5692 19119 5695
rect 19426 5692 19432 5704
rect 19107 5664 19432 5692
rect 19107 5661 19119 5664
rect 19061 5655 19119 5661
rect 19426 5652 19432 5664
rect 19484 5652 19490 5704
rect 20441 5695 20499 5701
rect 20441 5661 20453 5695
rect 20487 5692 20499 5695
rect 20530 5692 20536 5704
rect 20487 5664 20536 5692
rect 20487 5661 20499 5664
rect 20441 5655 20499 5661
rect 20530 5652 20536 5664
rect 20588 5652 20594 5704
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 19334 5624 19340 5636
rect 13924 5596 14688 5624
rect 18432 5596 19340 5624
rect 12342 5556 12348 5568
rect 9723 5528 11928 5556
rect 12303 5528 12348 5556
rect 9723 5525 9735 5528
rect 9677 5519 9735 5525
rect 12342 5516 12348 5528
rect 12400 5516 12406 5568
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 12894 5556 12900 5568
rect 12759 5528 12900 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13170 5516 13176 5568
rect 13228 5556 13234 5568
rect 13924 5556 13952 5596
rect 18432 5568 18460 5596
rect 19334 5584 19340 5596
rect 19392 5584 19398 5636
rect 19797 5627 19855 5633
rect 19797 5593 19809 5627
rect 19843 5624 19855 5627
rect 20162 5624 20168 5636
rect 19843 5596 20168 5624
rect 19843 5593 19855 5596
rect 19797 5587 19855 5593
rect 20162 5584 20168 5596
rect 20220 5624 20226 5636
rect 20220 5596 20576 5624
rect 20220 5584 20226 5596
rect 20548 5568 20576 5596
rect 14366 5556 14372 5568
rect 13228 5528 13952 5556
rect 14327 5528 14372 5556
rect 13228 5516 13234 5528
rect 14366 5516 14372 5528
rect 14424 5516 14430 5568
rect 15749 5559 15807 5565
rect 15749 5525 15761 5559
rect 15795 5556 15807 5559
rect 17402 5556 17408 5568
rect 15795 5528 17408 5556
rect 15795 5525 15807 5528
rect 15749 5519 15807 5525
rect 17402 5516 17408 5528
rect 17460 5516 17466 5568
rect 18046 5556 18052 5568
rect 18007 5528 18052 5556
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 20530 5516 20536 5568
rect 20588 5516 20594 5568
rect 22278 5556 22284 5568
rect 22239 5528 22284 5556
rect 22278 5516 22284 5528
rect 22336 5516 22342 5568
rect 1104 5466 22816 5488
rect 1104 5414 4614 5466
rect 4666 5414 4678 5466
rect 4730 5414 4742 5466
rect 4794 5414 4806 5466
rect 4858 5414 11878 5466
rect 11930 5414 11942 5466
rect 11994 5414 12006 5466
rect 12058 5414 12070 5466
rect 12122 5414 19142 5466
rect 19194 5414 19206 5466
rect 19258 5414 19270 5466
rect 19322 5414 19334 5466
rect 19386 5414 22816 5466
rect 1104 5392 22816 5414
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 9582 5352 9588 5364
rect 7892 5324 9260 5352
rect 9543 5324 9588 5352
rect 7892 5312 7898 5324
rect 9232 5216 9260 5324
rect 9582 5312 9588 5324
rect 9640 5312 9646 5364
rect 11422 5352 11428 5364
rect 10428 5324 11428 5352
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 9232 5188 10241 5216
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8205 5151 8263 5157
rect 8205 5148 8217 5151
rect 7984 5120 8217 5148
rect 7984 5108 7990 5120
rect 8205 5117 8217 5120
rect 8251 5117 8263 5151
rect 8205 5111 8263 5117
rect 10045 5151 10103 5157
rect 10045 5117 10057 5151
rect 10091 5148 10103 5151
rect 10428 5148 10456 5324
rect 11422 5312 11428 5324
rect 11480 5312 11486 5364
rect 11698 5312 11704 5364
rect 11756 5352 11762 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 11756 5324 12081 5352
rect 11756 5312 11762 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12618 5312 12624 5364
rect 12676 5352 12682 5364
rect 12676 5324 16252 5352
rect 12676 5312 12682 5324
rect 13906 5244 13912 5296
rect 13964 5284 13970 5296
rect 15010 5284 15016 5296
rect 13964 5256 15016 5284
rect 13964 5244 13970 5256
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 16224 5284 16252 5324
rect 17402 5312 17408 5364
rect 17460 5352 17466 5364
rect 19426 5352 19432 5364
rect 17460 5324 19104 5352
rect 19387 5324 19432 5352
rect 17460 5312 17466 5324
rect 16224 5256 17724 5284
rect 12894 5216 12900 5228
rect 12855 5188 12900 5216
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 17586 5216 17592 5228
rect 14292 5188 15424 5216
rect 17547 5188 17592 5216
rect 10091 5120 10456 5148
rect 10091 5117 10103 5120
rect 10045 5111 10103 5117
rect 8220 5012 8248 5111
rect 10502 5108 10508 5160
rect 10560 5148 10566 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10560 5120 10701 5148
rect 10560 5108 10566 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 10956 5151 11014 5157
rect 10956 5117 10968 5151
rect 11002 5148 11014 5151
rect 11238 5148 11244 5160
rect 11002 5120 11244 5148
rect 11002 5117 11014 5120
rect 10956 5111 11014 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 12986 5108 12992 5160
rect 13044 5148 13050 5160
rect 14292 5148 14320 5188
rect 13044 5120 14320 5148
rect 14737 5151 14795 5157
rect 13044 5108 13050 5120
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 8472 5083 8530 5089
rect 8472 5049 8484 5083
rect 8518 5080 8530 5083
rect 12342 5080 12348 5092
rect 8518 5052 12348 5080
rect 8518 5049 8530 5052
rect 8472 5043 8530 5049
rect 12342 5040 12348 5052
rect 12400 5040 12406 5092
rect 13164 5083 13222 5089
rect 13164 5049 13176 5083
rect 13210 5080 13222 5083
rect 14366 5080 14372 5092
rect 13210 5052 14372 5080
rect 13210 5049 13222 5052
rect 13164 5043 13222 5049
rect 14366 5040 14372 5052
rect 14424 5040 14430 5092
rect 14752 5080 14780 5111
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 15252 5120 15301 5148
rect 15252 5108 15258 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15396 5148 15424 5188
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17696 5216 17724 5256
rect 19076 5216 19104 5324
rect 19426 5312 19432 5324
rect 19484 5312 19490 5364
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 20070 5352 20076 5364
rect 19751 5324 20076 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20257 5219 20315 5225
rect 20257 5216 20269 5219
rect 17696 5188 18184 5216
rect 19076 5188 20269 5216
rect 17405 5151 17463 5157
rect 17405 5148 17417 5151
rect 15396 5120 17417 5148
rect 15289 5111 15347 5117
rect 17405 5117 17417 5120
rect 17451 5117 17463 5151
rect 17405 5111 17463 5117
rect 18049 5151 18107 5157
rect 18049 5117 18061 5151
rect 18095 5117 18107 5151
rect 18156 5148 18184 5188
rect 20257 5185 20269 5188
rect 20303 5185 20315 5219
rect 20257 5179 20315 5185
rect 19518 5148 19524 5160
rect 18156 5120 19524 5148
rect 18049 5111 18107 5117
rect 15562 5089 15568 5092
rect 14752 5052 15516 5080
rect 9861 5015 9919 5021
rect 9861 5012 9873 5015
rect 8220 4984 9873 5012
rect 9861 4981 9873 4984
rect 9907 5012 9919 5015
rect 10502 5012 10508 5024
rect 9907 4984 10508 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 12437 5015 12495 5021
rect 12437 4981 12449 5015
rect 12483 5012 12495 5015
rect 13446 5012 13452 5024
rect 12483 4984 13452 5012
rect 12483 4981 12495 4984
rect 12437 4975 12495 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 14277 5015 14335 5021
rect 14277 5012 14289 5015
rect 13596 4984 14289 5012
rect 13596 4972 13602 4984
rect 14277 4981 14289 4984
rect 14323 4981 14335 5015
rect 14277 4975 14335 4981
rect 14921 5015 14979 5021
rect 14921 4981 14933 5015
rect 14967 5012 14979 5015
rect 15010 5012 15016 5024
rect 14967 4984 15016 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15010 4972 15016 4984
rect 15068 4972 15074 5024
rect 15488 5012 15516 5052
rect 15556 5043 15568 5089
rect 15620 5080 15626 5092
rect 16390 5080 16396 5092
rect 15620 5052 16396 5080
rect 15562 5040 15568 5043
rect 15620 5040 15626 5052
rect 16390 5040 16396 5052
rect 16448 5040 16454 5092
rect 18064 5080 18092 5111
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 20898 5148 20904 5160
rect 20859 5120 20904 5148
rect 20898 5108 20904 5120
rect 20956 5108 20962 5160
rect 18316 5083 18374 5089
rect 18064 5052 18184 5080
rect 16482 5012 16488 5024
rect 15488 4984 16488 5012
rect 16482 4972 16488 4984
rect 16540 4972 16546 5024
rect 16666 5012 16672 5024
rect 16627 4984 16672 5012
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17034 4972 17040 5024
rect 17092 5012 17098 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 17092 4984 17325 5012
rect 17092 4972 17098 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 18156 5012 18184 5052
rect 18316 5049 18328 5083
rect 18362 5080 18374 5083
rect 19242 5080 19248 5092
rect 18362 5052 19248 5080
rect 18362 5049 18374 5052
rect 18316 5043 18374 5049
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 20073 5083 20131 5089
rect 20073 5049 20085 5083
rect 20119 5080 20131 5083
rect 20254 5080 20260 5092
rect 20119 5052 20260 5080
rect 20119 5049 20131 5052
rect 20073 5043 20131 5049
rect 20254 5040 20260 5052
rect 20312 5040 20318 5092
rect 20714 5040 20720 5092
rect 20772 5080 20778 5092
rect 21146 5083 21204 5089
rect 21146 5080 21158 5083
rect 20772 5052 21158 5080
rect 20772 5040 20778 5052
rect 21146 5049 21158 5052
rect 21192 5049 21204 5083
rect 21146 5043 21204 5049
rect 18690 5012 18696 5024
rect 18156 4984 18696 5012
rect 17313 4975 17371 4981
rect 18690 4972 18696 4984
rect 18748 4972 18754 5024
rect 20162 4972 20168 5024
rect 20220 5012 20226 5024
rect 20220 4984 20265 5012
rect 20220 4972 20226 4984
rect 22094 4972 22100 5024
rect 22152 5012 22158 5024
rect 22281 5015 22339 5021
rect 22281 5012 22293 5015
rect 22152 4984 22293 5012
rect 22152 4972 22158 4984
rect 22281 4981 22293 4984
rect 22327 4981 22339 5015
rect 22281 4975 22339 4981
rect 1104 4922 22816 4944
rect 1104 4870 8246 4922
rect 8298 4870 8310 4922
rect 8362 4870 8374 4922
rect 8426 4870 8438 4922
rect 8490 4870 15510 4922
rect 15562 4870 15574 4922
rect 15626 4870 15638 4922
rect 15690 4870 15702 4922
rect 15754 4870 22816 4922
rect 1104 4848 22816 4870
rect 10042 4808 10048 4820
rect 10003 4780 10048 4808
rect 10042 4768 10048 4780
rect 10100 4768 10106 4820
rect 11698 4768 11704 4820
rect 11756 4808 11762 4820
rect 12621 4811 12679 4817
rect 12621 4808 12633 4811
rect 11756 4780 12633 4808
rect 11756 4768 11762 4780
rect 12621 4777 12633 4780
rect 12667 4777 12679 4811
rect 12621 4771 12679 4777
rect 13081 4811 13139 4817
rect 13081 4777 13093 4811
rect 13127 4808 13139 4811
rect 13173 4811 13231 4817
rect 13173 4808 13185 4811
rect 13127 4780 13185 4808
rect 13127 4777 13139 4780
rect 13081 4771 13139 4777
rect 13173 4777 13185 4780
rect 13219 4777 13231 4811
rect 13538 4808 13544 4820
rect 13499 4780 13544 4808
rect 13173 4771 13231 4777
rect 13538 4768 13544 4780
rect 13596 4768 13602 4820
rect 13633 4811 13691 4817
rect 13633 4777 13645 4811
rect 13679 4808 13691 4811
rect 14366 4808 14372 4820
rect 13679 4780 14372 4808
rect 13679 4777 13691 4780
rect 13633 4771 13691 4777
rect 14366 4768 14372 4780
rect 14424 4768 14430 4820
rect 14458 4768 14464 4820
rect 14516 4808 14522 4820
rect 14553 4811 14611 4817
rect 14553 4808 14565 4811
rect 14516 4780 14565 4808
rect 14516 4768 14522 4780
rect 14553 4777 14565 4780
rect 14599 4777 14611 4811
rect 14553 4771 14611 4777
rect 14642 4768 14648 4820
rect 14700 4808 14706 4820
rect 15841 4811 15899 4817
rect 14700 4780 14745 4808
rect 14700 4768 14706 4780
rect 15841 4777 15853 4811
rect 15887 4808 15899 4811
rect 17865 4811 17923 4817
rect 17865 4808 17877 4811
rect 15887 4780 17877 4808
rect 15887 4777 15899 4780
rect 15841 4771 15899 4777
rect 17865 4777 17877 4780
rect 17911 4777 17923 4811
rect 17865 4771 17923 4777
rect 18693 4811 18751 4817
rect 18693 4777 18705 4811
rect 18739 4808 18751 4811
rect 18874 4808 18880 4820
rect 18739 4780 18880 4808
rect 18739 4777 18751 4780
rect 18693 4771 18751 4777
rect 18874 4768 18880 4780
rect 18932 4768 18938 4820
rect 18966 4768 18972 4820
rect 19024 4808 19030 4820
rect 19153 4811 19211 4817
rect 19153 4808 19165 4811
rect 19024 4780 19165 4808
rect 19024 4768 19030 4780
rect 19153 4777 19165 4780
rect 19199 4777 19211 4811
rect 19153 4771 19211 4777
rect 19610 4768 19616 4820
rect 19668 4808 19674 4820
rect 19705 4811 19763 4817
rect 19705 4808 19717 4811
rect 19668 4780 19717 4808
rect 19668 4768 19674 4780
rect 19705 4777 19717 4780
rect 19751 4777 19763 4811
rect 20070 4808 20076 4820
rect 20031 4780 20076 4808
rect 19705 4771 19763 4777
rect 20070 4768 20076 4780
rect 20128 4768 20134 4820
rect 22278 4808 22284 4820
rect 20180 4780 22284 4808
rect 10772 4743 10830 4749
rect 10772 4709 10784 4743
rect 10818 4740 10830 4743
rect 13556 4740 13584 4768
rect 10818 4712 13584 4740
rect 10818 4709 10830 4712
rect 10772 4703 10830 4709
rect 13722 4700 13728 4752
rect 13780 4740 13786 4752
rect 14918 4740 14924 4752
rect 13780 4712 14924 4740
rect 13780 4700 13786 4712
rect 14918 4700 14924 4712
rect 14976 4740 14982 4752
rect 15194 4740 15200 4752
rect 14976 4712 15200 4740
rect 14976 4700 14982 4712
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 16942 4740 16948 4752
rect 15672 4712 16948 4740
rect 9125 4675 9183 4681
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9171 4644 11560 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 10502 4604 10508 4616
rect 10463 4576 10508 4604
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 11532 4604 11560 4644
rect 11606 4632 11612 4684
rect 11664 4672 11670 4684
rect 11977 4675 12035 4681
rect 11977 4672 11989 4675
rect 11664 4644 11989 4672
rect 11664 4632 11670 4644
rect 11977 4641 11989 4644
rect 12023 4641 12035 4675
rect 11977 4635 12035 4641
rect 12342 4632 12348 4684
rect 12400 4672 12406 4684
rect 12529 4675 12587 4681
rect 12529 4672 12541 4675
rect 12400 4644 12541 4672
rect 12400 4632 12406 4644
rect 12529 4641 12541 4644
rect 12575 4641 12587 4675
rect 12529 4635 12587 4641
rect 13081 4675 13139 4681
rect 13081 4641 13093 4675
rect 13127 4672 13139 4675
rect 15102 4672 15108 4684
rect 13127 4644 15108 4672
rect 13127 4641 13139 4644
rect 13081 4635 13139 4641
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 15672 4681 15700 4712
rect 16942 4700 16948 4712
rect 17000 4700 17006 4752
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 19061 4743 19119 4749
rect 19061 4740 19073 4743
rect 18104 4712 19073 4740
rect 18104 4700 18110 4712
rect 19061 4709 19073 4712
rect 19107 4709 19119 4743
rect 19242 4740 19248 4752
rect 19155 4712 19248 4740
rect 19061 4703 19119 4709
rect 19242 4700 19248 4712
rect 19300 4740 19306 4752
rect 20180 4740 20208 4780
rect 22278 4768 22284 4780
rect 22336 4768 22342 4820
rect 19300 4712 20208 4740
rect 21168 4743 21226 4749
rect 19300 4700 19306 4712
rect 21168 4709 21180 4743
rect 21214 4740 21226 4743
rect 21266 4740 21272 4752
rect 21214 4712 21272 4740
rect 21214 4709 21226 4712
rect 21168 4703 21226 4709
rect 21266 4700 21272 4712
rect 21324 4700 21330 4752
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4641 15715 4675
rect 16574 4672 16580 4684
rect 16535 4644 16580 4672
rect 15657 4635 15715 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 17586 4672 17592 4684
rect 16868 4644 17592 4672
rect 12618 4604 12624 4616
rect 11532 4576 12624 4604
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 12802 4604 12808 4616
rect 12715 4576 12808 4604
rect 12802 4564 12808 4576
rect 12860 4604 12866 4616
rect 13817 4607 13875 4613
rect 13817 4604 13829 4607
rect 12860 4576 13829 4604
rect 12860 4564 12866 4576
rect 13817 4573 13829 4576
rect 13863 4573 13875 4607
rect 13817 4567 13875 4573
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 13078 4496 13084 4548
rect 13136 4536 13142 4548
rect 13722 4536 13728 4548
rect 13136 4508 13728 4536
rect 13136 4496 13142 4508
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 13832 4536 13860 4567
rect 14752 4536 14780 4567
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 16868 4613 16896 4644
rect 17586 4632 17592 4644
rect 17644 4632 17650 4684
rect 17773 4675 17831 4681
rect 17773 4641 17785 4675
rect 17819 4672 17831 4675
rect 18230 4672 18236 4684
rect 17819 4644 18236 4672
rect 17819 4641 17831 4644
rect 17773 4635 17831 4641
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 16669 4607 16727 4613
rect 16669 4604 16681 4607
rect 15252 4576 16681 4604
rect 15252 4564 15258 4576
rect 16669 4573 16681 4576
rect 16715 4573 16727 4607
rect 16669 4567 16727 4573
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 17402 4564 17408 4616
rect 17460 4604 17466 4616
rect 19260 4613 19288 4700
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17460 4576 17969 4604
rect 17460 4564 17466 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 19521 4607 19579 4613
rect 19521 4573 19533 4607
rect 19567 4604 19579 4607
rect 20165 4607 20223 4613
rect 20165 4604 20177 4607
rect 19567 4576 20177 4604
rect 19567 4573 19579 4576
rect 19521 4567 19579 4573
rect 20165 4573 20177 4576
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 20257 4607 20315 4613
rect 20257 4573 20269 4607
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 13832 4508 14780 4536
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 20272 4536 20300 4567
rect 20438 4564 20444 4616
rect 20496 4604 20502 4616
rect 20898 4604 20904 4616
rect 20496 4576 20904 4604
rect 20496 4564 20502 4576
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 20806 4536 20812 4548
rect 15068 4508 20300 4536
rect 20364 4508 20812 4536
rect 15068 4496 15074 4508
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11931 4440 11989 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 11977 4431 12035 4437
rect 12161 4471 12219 4477
rect 12161 4437 12173 4471
rect 12207 4468 12219 4471
rect 12250 4468 12256 4480
rect 12207 4440 12256 4468
rect 12207 4437 12219 4440
rect 12161 4431 12219 4437
rect 12250 4428 12256 4440
rect 12308 4428 12314 4480
rect 14182 4468 14188 4480
rect 14143 4440 14188 4468
rect 14182 4428 14188 4440
rect 14240 4428 14246 4480
rect 14366 4428 14372 4480
rect 14424 4468 14430 4480
rect 14918 4468 14924 4480
rect 14424 4440 14924 4468
rect 14424 4428 14430 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 16209 4471 16267 4477
rect 16209 4437 16221 4471
rect 16255 4468 16267 4471
rect 17310 4468 17316 4480
rect 16255 4440 17316 4468
rect 16255 4437 16267 4440
rect 16209 4431 16267 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 17405 4471 17463 4477
rect 17405 4437 17417 4471
rect 17451 4468 17463 4471
rect 17862 4468 17868 4480
rect 17451 4440 17868 4468
rect 17451 4437 17463 4440
rect 17405 4431 17463 4437
rect 17862 4428 17868 4440
rect 17920 4468 17926 4480
rect 19521 4471 19579 4477
rect 19521 4468 19533 4471
rect 17920 4440 19533 4468
rect 17920 4428 17926 4440
rect 19521 4437 19533 4440
rect 19567 4437 19579 4471
rect 19521 4431 19579 4437
rect 19702 4428 19708 4480
rect 19760 4468 19766 4480
rect 20364 4468 20392 4508
rect 20806 4496 20812 4508
rect 20864 4496 20870 4548
rect 19760 4440 20392 4468
rect 19760 4428 19766 4440
rect 20714 4428 20720 4480
rect 20772 4468 20778 4480
rect 22281 4471 22339 4477
rect 22281 4468 22293 4471
rect 20772 4440 22293 4468
rect 20772 4428 20778 4440
rect 22281 4437 22293 4440
rect 22327 4437 22339 4471
rect 22281 4431 22339 4437
rect 1104 4378 22816 4400
rect 1104 4326 4614 4378
rect 4666 4326 4678 4378
rect 4730 4326 4742 4378
rect 4794 4326 4806 4378
rect 4858 4326 11878 4378
rect 11930 4326 11942 4378
rect 11994 4326 12006 4378
rect 12058 4326 12070 4378
rect 12122 4326 19142 4378
rect 19194 4326 19206 4378
rect 19258 4326 19270 4378
rect 19322 4326 19334 4378
rect 19386 4326 22816 4378
rect 1104 4304 22816 4326
rect 13078 4264 13084 4276
rect 10980 4236 13084 4264
rect 9490 4156 9496 4208
rect 9548 4196 9554 4208
rect 10980 4196 11008 4236
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 13262 4264 13268 4276
rect 13223 4236 13268 4264
rect 13262 4224 13268 4236
rect 13320 4224 13326 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 14550 4264 14556 4276
rect 13596 4236 14556 4264
rect 13596 4224 13602 4236
rect 14550 4224 14556 4236
rect 14608 4264 14614 4276
rect 16666 4264 16672 4276
rect 14608 4236 16672 4264
rect 14608 4224 14614 4236
rect 16666 4224 16672 4236
rect 16724 4224 16730 4276
rect 20254 4264 20260 4276
rect 20215 4236 20260 4264
rect 20254 4224 20260 4236
rect 20312 4224 20318 4276
rect 22370 4264 22376 4276
rect 20364 4236 22376 4264
rect 12802 4196 12808 4208
rect 9548 4168 10824 4196
rect 9548 4156 9554 4168
rect 9582 4128 9588 4140
rect 9543 4100 9588 4128
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 9784 4137 9812 4168
rect 9769 4131 9827 4137
rect 9769 4097 9781 4131
rect 9815 4097 9827 4131
rect 10686 4128 10692 4140
rect 10647 4100 10692 4128
rect 9769 4091 9827 4097
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 9214 4020 9220 4072
rect 9272 4060 9278 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9272 4032 9505 4060
rect 9272 4020 9278 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 10226 4020 10232 4072
rect 10284 4060 10290 4072
rect 10597 4063 10655 4069
rect 10597 4060 10609 4063
rect 10284 4032 10609 4060
rect 10284 4020 10290 4032
rect 10597 4029 10609 4032
rect 10643 4029 10655 4063
rect 10796 4060 10824 4168
rect 10888 4168 11008 4196
rect 11072 4168 12808 4196
rect 10888 4137 10916 4168
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 11072 4128 11100 4168
rect 10873 4091 10931 4097
rect 10980 4100 11100 4128
rect 10980 4060 11008 4100
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 11808 4137 11836 4168
rect 12802 4156 12808 4168
rect 12860 4156 12866 4208
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 13412 4168 13768 4196
rect 13412 4156 13418 4168
rect 11701 4131 11759 4137
rect 11701 4128 11713 4131
rect 11572 4100 11713 4128
rect 11572 4088 11578 4100
rect 11701 4097 11713 4100
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 11882 4088 11888 4140
rect 11940 4128 11946 4140
rect 13538 4128 13544 4140
rect 11940 4100 13544 4128
rect 11940 4088 11946 4100
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 13740 4128 13768 4168
rect 17586 4156 17592 4208
rect 17644 4196 17650 4208
rect 20364 4196 20392 4236
rect 22370 4224 22376 4236
rect 22428 4224 22434 4276
rect 17644 4168 20392 4196
rect 17644 4156 17650 4168
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13740 4100 13829 4128
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 13817 4091 13875 4097
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 18138 4088 18144 4140
rect 18196 4128 18202 4140
rect 18708 4137 18736 4168
rect 18693 4131 18751 4137
rect 18196 4100 18644 4128
rect 18196 4088 18202 4100
rect 10796 4032 11008 4060
rect 10597 4023 10655 4029
rect 11238 4020 11244 4072
rect 11296 4060 11302 4072
rect 11609 4063 11667 4069
rect 11609 4060 11621 4063
rect 11296 4032 11621 4060
rect 11296 4020 11302 4032
rect 11609 4029 11621 4032
rect 11655 4029 11667 4063
rect 12710 4060 12716 4072
rect 12671 4032 12716 4060
rect 11609 4023 11667 4029
rect 12710 4020 12716 4032
rect 12768 4020 12774 4072
rect 13446 4020 13452 4072
rect 13504 4060 13510 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13504 4032 13645 4060
rect 13504 4020 13510 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 14277 4063 14335 4069
rect 14277 4029 14289 4063
rect 14323 4060 14335 4063
rect 14366 4060 14372 4072
rect 14323 4032 14372 4060
rect 14323 4029 14335 4032
rect 14277 4023 14335 4029
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 16574 4060 16580 4072
rect 15948 4032 16580 4060
rect 8570 3952 8576 4004
rect 8628 3992 8634 4004
rect 8628 3964 10272 3992
rect 8628 3952 8634 3964
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 10244 3933 10272 3964
rect 13170 3952 13176 4004
rect 13228 3992 13234 4004
rect 14550 4001 14556 4004
rect 14544 3992 14556 4001
rect 13228 3964 13860 3992
rect 14511 3964 14556 3992
rect 13228 3952 13234 3964
rect 10229 3927 10287 3933
rect 10229 3893 10241 3927
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 11241 3927 11299 3933
rect 11241 3893 11253 3927
rect 11287 3924 11299 3927
rect 11330 3924 11336 3936
rect 11287 3896 11336 3924
rect 11287 3893 11299 3896
rect 11241 3887 11299 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11422 3884 11428 3936
rect 11480 3924 11486 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 11480 3896 12909 3924
rect 11480 3884 11486 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 13722 3924 13728 3936
rect 13683 3896 13728 3924
rect 12897 3887 12955 3893
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 13832 3924 13860 3964
rect 14544 3955 14556 3964
rect 14550 3952 14556 3955
rect 14608 3952 14614 4004
rect 15948 3992 15976 4032
rect 16574 4020 16580 4032
rect 16632 4020 16638 4072
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 18509 4063 18567 4069
rect 18509 4060 18521 4063
rect 16724 4032 18521 4060
rect 16724 4020 16730 4032
rect 18509 4029 18521 4032
rect 18555 4029 18567 4063
rect 18616 4060 18644 4100
rect 18693 4097 18705 4131
rect 18739 4097 18751 4131
rect 19702 4128 19708 4140
rect 19663 4100 19708 4128
rect 18693 4091 18751 4097
rect 19702 4088 19708 4100
rect 19760 4088 19766 4140
rect 20070 4060 20076 4072
rect 18616 4032 19932 4060
rect 20031 4032 20076 4060
rect 18509 4023 18567 4029
rect 14752 3964 15976 3992
rect 14752 3924 14780 3964
rect 16114 3952 16120 4004
rect 16172 4001 16178 4004
rect 16172 3995 16236 4001
rect 16172 3961 16190 3995
rect 16224 3992 16236 3995
rect 16850 3992 16856 4004
rect 16224 3964 16856 3992
rect 16224 3961 16236 3964
rect 16172 3955 16236 3961
rect 16172 3952 16178 3955
rect 16850 3952 16856 3964
rect 16908 3952 16914 4004
rect 18417 3995 18475 4001
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 19429 3995 19487 4001
rect 18463 3964 19104 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 13832 3896 14780 3924
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15160 3896 15669 3924
rect 15160 3884 15166 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 16356 3896 17325 3924
rect 16356 3884 16362 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 18046 3924 18052 3936
rect 18007 3896 18052 3924
rect 17313 3887 17371 3893
rect 18046 3884 18052 3896
rect 18104 3884 18110 3936
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 18874 3924 18880 3936
rect 18380 3896 18880 3924
rect 18380 3884 18386 3896
rect 18874 3884 18880 3896
rect 18932 3884 18938 3936
rect 19076 3933 19104 3964
rect 19429 3961 19441 3995
rect 19475 3992 19487 3995
rect 19794 3992 19800 4004
rect 19475 3964 19800 3992
rect 19475 3961 19487 3964
rect 19429 3955 19487 3961
rect 19794 3952 19800 3964
rect 19852 3952 19858 4004
rect 19904 3992 19932 4032
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20438 4020 20444 4072
rect 20496 4060 20502 4072
rect 20717 4063 20775 4069
rect 20717 4060 20729 4063
rect 20496 4032 20729 4060
rect 20496 4020 20502 4032
rect 20717 4029 20729 4032
rect 20763 4029 20775 4063
rect 20717 4023 20775 4029
rect 20962 3995 21020 4001
rect 20962 3992 20974 3995
rect 19904 3964 20974 3992
rect 20962 3961 20974 3964
rect 21008 3992 21020 3995
rect 22278 3992 22284 4004
rect 21008 3964 22284 3992
rect 21008 3961 21020 3964
rect 20962 3955 21020 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 19521 3927 19579 3933
rect 19521 3893 19533 3927
rect 19567 3924 19579 3927
rect 19978 3924 19984 3936
rect 19567 3896 19984 3924
rect 19567 3893 19579 3896
rect 19521 3887 19579 3893
rect 19978 3884 19984 3896
rect 20036 3884 20042 3936
rect 21266 3884 21272 3936
rect 21324 3924 21330 3936
rect 22097 3927 22155 3933
rect 22097 3924 22109 3927
rect 21324 3896 22109 3924
rect 21324 3884 21330 3896
rect 22097 3893 22109 3896
rect 22143 3893 22155 3927
rect 22097 3887 22155 3893
rect 1104 3834 22816 3856
rect 1104 3782 8246 3834
rect 8298 3782 8310 3834
rect 8362 3782 8374 3834
rect 8426 3782 8438 3834
rect 8490 3782 15510 3834
rect 15562 3782 15574 3834
rect 15626 3782 15638 3834
rect 15690 3782 15702 3834
rect 15754 3782 22816 3834
rect 1104 3760 22816 3782
rect 11149 3723 11207 3729
rect 11149 3689 11161 3723
rect 11195 3720 11207 3723
rect 12986 3720 12992 3732
rect 11195 3692 12992 3720
rect 11195 3689 11207 3692
rect 11149 3683 11207 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13170 3720 13176 3732
rect 13131 3692 13176 3720
rect 13170 3680 13176 3692
rect 13228 3680 13234 3732
rect 13541 3723 13599 3729
rect 13541 3689 13553 3723
rect 13587 3720 13599 3723
rect 13587 3692 16436 3720
rect 13587 3689 13599 3692
rect 13541 3683 13599 3689
rect 3510 3612 3516 3664
rect 3568 3652 3574 3664
rect 11422 3652 11428 3664
rect 3568 3624 11428 3652
rect 3568 3612 3574 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 11517 3655 11575 3661
rect 11517 3621 11529 3655
rect 11563 3652 11575 3655
rect 11882 3652 11888 3664
rect 11563 3624 11888 3652
rect 11563 3621 11575 3624
rect 11517 3615 11575 3621
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 12526 3652 12532 3664
rect 12487 3624 12532 3652
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13633 3655 13691 3661
rect 13633 3621 13645 3655
rect 13679 3652 13691 3655
rect 13906 3652 13912 3664
rect 13679 3624 13912 3652
rect 13679 3621 13691 3624
rect 13633 3615 13691 3621
rect 13906 3612 13912 3624
rect 13964 3612 13970 3664
rect 14550 3652 14556 3664
rect 14463 3624 14556 3652
rect 14550 3612 14556 3624
rect 14608 3652 14614 3664
rect 16206 3652 16212 3664
rect 14608 3624 16212 3652
rect 14608 3612 14614 3624
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 16408 3652 16436 3692
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 19886 3720 19892 3732
rect 18840 3692 19892 3720
rect 18840 3680 18846 3692
rect 19886 3680 19892 3692
rect 19944 3680 19950 3732
rect 20162 3680 20168 3732
rect 20220 3720 20226 3732
rect 20441 3723 20499 3729
rect 20441 3720 20453 3723
rect 20220 3692 20453 3720
rect 20220 3680 20226 3692
rect 20441 3689 20453 3692
rect 20487 3689 20499 3723
rect 22278 3720 22284 3732
rect 22239 3692 22284 3720
rect 20441 3683 20499 3689
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 17190 3655 17248 3661
rect 17190 3652 17202 3655
rect 16408 3624 17202 3652
rect 17190 3621 17202 3624
rect 17236 3652 17248 3655
rect 17402 3652 17408 3664
rect 17236 3624 17408 3652
rect 17236 3621 17248 3624
rect 17190 3615 17248 3621
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 18046 3612 18052 3664
rect 18104 3652 18110 3664
rect 18104 3624 20300 3652
rect 18104 3612 18110 3624
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 12434 3584 12440 3596
rect 10735 3556 12440 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 12621 3587 12679 3593
rect 12621 3553 12633 3587
rect 12667 3584 12679 3587
rect 12667 3556 14412 3584
rect 12667 3553 12679 3556
rect 12621 3547 12679 3553
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3516 11851 3519
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 11839 3488 12817 3516
rect 11839 3485 11851 3488
rect 11793 3479 11851 3485
rect 12805 3485 12817 3488
rect 12851 3516 12863 3519
rect 13630 3516 13636 3528
rect 12851 3488 13636 3516
rect 12851 3485 12863 3488
rect 12805 3479 12863 3485
rect 11624 3448 11652 3479
rect 13630 3476 13636 3488
rect 13688 3516 13694 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 12434 3448 12440 3460
rect 11624 3420 12440 3448
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 14185 3451 14243 3457
rect 14185 3417 14197 3451
rect 14231 3448 14243 3451
rect 14274 3448 14280 3460
rect 14231 3420 14280 3448
rect 14231 3417 14243 3420
rect 14185 3411 14243 3417
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 12161 3383 12219 3389
rect 12161 3349 12173 3383
rect 12207 3380 12219 3383
rect 12250 3380 12256 3392
rect 12207 3352 12256 3380
rect 12207 3349 12219 3352
rect 12161 3343 12219 3349
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 14384 3380 14412 3556
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 14700 3556 14745 3584
rect 14700 3544 14706 3556
rect 15010 3544 15016 3596
rect 15068 3584 15074 3596
rect 15562 3593 15568 3596
rect 15545 3587 15568 3593
rect 15545 3584 15557 3587
rect 15068 3556 15557 3584
rect 15068 3544 15074 3556
rect 15545 3553 15557 3556
rect 15620 3584 15626 3596
rect 15620 3556 15693 3584
rect 15545 3547 15568 3553
rect 15562 3544 15568 3547
rect 15620 3544 15626 3556
rect 15838 3544 15844 3596
rect 15896 3584 15902 3596
rect 18414 3584 18420 3596
rect 15896 3556 18420 3584
rect 15896 3544 15902 3556
rect 18414 3544 18420 3556
rect 18472 3544 18478 3596
rect 18598 3584 18604 3596
rect 18559 3556 18604 3584
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 20272 3593 20300 3624
rect 21174 3593 21180 3596
rect 18857 3587 18915 3593
rect 18857 3584 18869 3587
rect 18748 3556 18869 3584
rect 18748 3544 18754 3556
rect 18857 3553 18869 3556
rect 18903 3553 18915 3587
rect 18857 3547 18915 3553
rect 20257 3587 20315 3593
rect 20257 3553 20269 3587
rect 20303 3553 20315 3587
rect 21168 3584 21180 3593
rect 21135 3556 21180 3584
rect 20257 3547 20315 3553
rect 21168 3547 21180 3556
rect 21174 3544 21180 3547
rect 21232 3544 21238 3596
rect 14826 3516 14832 3528
rect 14787 3488 14832 3516
rect 14826 3476 14832 3488
rect 14884 3476 14890 3528
rect 14918 3476 14924 3528
rect 14976 3516 14982 3528
rect 15289 3519 15347 3525
rect 15289 3516 15301 3519
rect 14976 3488 15301 3516
rect 14976 3476 14982 3488
rect 15289 3485 15301 3488
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 16390 3408 16396 3460
rect 16448 3448 16454 3460
rect 16960 3448 16988 3479
rect 20162 3476 20168 3528
rect 20220 3516 20226 3528
rect 20438 3516 20444 3528
rect 20220 3488 20444 3516
rect 20220 3476 20226 3488
rect 20438 3476 20444 3488
rect 20496 3516 20502 3528
rect 20901 3519 20959 3525
rect 20901 3516 20913 3519
rect 20496 3488 20913 3516
rect 20496 3476 20502 3488
rect 20901 3485 20913 3488
rect 20947 3485 20959 3519
rect 20901 3479 20959 3485
rect 18598 3448 18604 3460
rect 16448 3420 16988 3448
rect 16448 3408 16454 3420
rect 15930 3380 15936 3392
rect 14384 3352 15936 3380
rect 15930 3340 15936 3352
rect 15988 3380 15994 3392
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 15988 3352 16681 3380
rect 15988 3340 15994 3352
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16960 3380 16988 3420
rect 17880 3420 18604 3448
rect 17880 3380 17908 3420
rect 18598 3408 18604 3420
rect 18656 3408 18662 3460
rect 18322 3380 18328 3392
rect 16960 3352 17908 3380
rect 18283 3352 18328 3380
rect 16669 3343 16727 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 1104 3290 22816 3312
rect 1104 3238 4614 3290
rect 4666 3238 4678 3290
rect 4730 3238 4742 3290
rect 4794 3238 4806 3290
rect 4858 3238 11878 3290
rect 11930 3238 11942 3290
rect 11994 3238 12006 3290
rect 12058 3238 12070 3290
rect 12122 3238 19142 3290
rect 19194 3238 19206 3290
rect 19258 3238 19270 3290
rect 19322 3238 19334 3290
rect 19386 3238 22816 3290
rect 1104 3216 22816 3238
rect 7466 3136 7472 3188
rect 7524 3176 7530 3188
rect 13722 3176 13728 3188
rect 7524 3148 13728 3176
rect 7524 3136 7530 3148
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 16666 3176 16672 3188
rect 14200 3148 16672 3176
rect 13173 3111 13231 3117
rect 13173 3077 13185 3111
rect 13219 3108 13231 3111
rect 14200 3108 14228 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 17402 3176 17408 3188
rect 17363 3148 17408 3176
rect 17402 3136 17408 3148
rect 17460 3136 17466 3188
rect 18230 3176 18236 3188
rect 18191 3148 18236 3176
rect 18230 3136 18236 3148
rect 18288 3136 18294 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18656 3148 19748 3176
rect 18656 3136 18662 3148
rect 15562 3108 15568 3120
rect 13219 3080 14228 3108
rect 15523 3080 15568 3108
rect 13219 3077 13231 3080
rect 13173 3071 13231 3077
rect 15562 3068 15568 3080
rect 15620 3068 15626 3120
rect 19720 3108 19748 3148
rect 19794 3136 19800 3188
rect 19852 3176 19858 3188
rect 19981 3179 20039 3185
rect 19981 3176 19993 3179
rect 19852 3148 19993 3176
rect 19852 3136 19858 3148
rect 19981 3145 19993 3148
rect 20027 3176 20039 3179
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 20027 3148 20085 3176
rect 20027 3145 20039 3148
rect 19981 3139 20039 3145
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 20162 3108 20168 3120
rect 19720 3080 20168 3108
rect 20162 3068 20168 3080
rect 20220 3068 20226 3120
rect 6914 3000 6920 3052
rect 6972 3040 6978 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 6972 3012 12725 3040
rect 6972 3000 6978 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 13722 3040 13728 3052
rect 13683 3012 13728 3040
rect 12713 3003 12771 3009
rect 13722 3000 13728 3012
rect 13780 3000 13786 3052
rect 20073 3043 20131 3049
rect 17236 3012 18736 3040
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 4028 2944 11713 2972
rect 4028 2932 4034 2944
rect 11701 2941 11713 2944
rect 11747 2972 11759 2975
rect 14090 2972 14096 2984
rect 11747 2944 14096 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 14090 2932 14096 2944
rect 14148 2932 14154 2984
rect 14185 2975 14243 2981
rect 14185 2941 14197 2975
rect 14231 2972 14243 2975
rect 14274 2972 14280 2984
rect 14231 2944 14280 2972
rect 14231 2941 14243 2944
rect 14185 2935 14243 2941
rect 14274 2932 14280 2944
rect 14332 2932 14338 2984
rect 16025 2975 16083 2981
rect 14384 2944 15976 2972
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 14384 2904 14412 2944
rect 13679 2876 14412 2904
rect 14452 2907 14510 2913
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 14452 2873 14464 2907
rect 14498 2904 14510 2907
rect 15102 2904 15108 2916
rect 14498 2876 15108 2904
rect 14498 2873 14510 2876
rect 14452 2867 14510 2873
rect 15102 2864 15108 2876
rect 15160 2864 15166 2916
rect 15948 2904 15976 2944
rect 16025 2941 16037 2975
rect 16071 2972 16083 2975
rect 16114 2972 16120 2984
rect 16071 2944 16120 2972
rect 16071 2941 16083 2944
rect 16025 2935 16083 2941
rect 16114 2932 16120 2944
rect 16172 2932 16178 2984
rect 16298 2981 16304 2984
rect 16292 2972 16304 2981
rect 16259 2944 16304 2972
rect 16292 2935 16304 2944
rect 16298 2932 16304 2935
rect 16356 2932 16362 2984
rect 16574 2932 16580 2984
rect 16632 2972 16638 2984
rect 17236 2972 17264 3012
rect 16632 2944 17264 2972
rect 16632 2932 16638 2944
rect 17310 2932 17316 2984
rect 17368 2972 17374 2984
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 17368 2944 18061 2972
rect 17368 2932 17374 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18598 2972 18604 2984
rect 18559 2944 18604 2972
rect 18049 2935 18107 2941
rect 18598 2932 18604 2944
rect 18656 2932 18662 2984
rect 18322 2904 18328 2916
rect 15212 2876 15884 2904
rect 15948 2876 18328 2904
rect 11885 2839 11943 2845
rect 11885 2805 11897 2839
rect 11931 2836 11943 2839
rect 12158 2836 12164 2848
rect 11931 2808 12164 2836
rect 11931 2805 11943 2808
rect 11885 2799 11943 2805
rect 12158 2796 12164 2808
rect 12216 2796 12222 2848
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 15212 2836 15240 2876
rect 13587 2808 15240 2836
rect 15856 2836 15884 2876
rect 18322 2864 18328 2876
rect 18380 2864 18386 2916
rect 18708 2904 18736 3012
rect 20073 3009 20085 3043
rect 20119 3040 20131 3043
rect 20119 3012 20392 3040
rect 20119 3009 20131 3012
rect 20073 3003 20131 3009
rect 18868 2975 18926 2981
rect 18868 2941 18880 2975
rect 18914 2972 18926 2975
rect 19978 2972 19984 2984
rect 18914 2944 19984 2972
rect 18914 2941 18926 2944
rect 18868 2935 18926 2941
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20165 2975 20223 2981
rect 20165 2941 20177 2975
rect 20211 2972 20223 2975
rect 20257 2975 20315 2981
rect 20257 2972 20269 2975
rect 20211 2944 20269 2972
rect 20211 2941 20223 2944
rect 20165 2935 20223 2941
rect 20257 2941 20269 2944
rect 20303 2941 20315 2975
rect 20364 2972 20392 3012
rect 20513 2975 20571 2981
rect 20513 2972 20525 2975
rect 20364 2944 20525 2972
rect 20257 2935 20315 2941
rect 20513 2941 20525 2944
rect 20559 2941 20571 2975
rect 20513 2935 20571 2941
rect 21913 2975 21971 2981
rect 21913 2941 21925 2975
rect 21959 2972 21971 2975
rect 22002 2972 22008 2984
rect 21959 2944 22008 2972
rect 21959 2941 21971 2944
rect 21913 2935 21971 2941
rect 22002 2932 22008 2944
rect 22060 2932 22066 2984
rect 22094 2932 22100 2984
rect 22152 2972 22158 2984
rect 22152 2944 22197 2972
rect 22152 2932 22158 2944
rect 22281 2907 22339 2913
rect 22281 2904 22293 2907
rect 18708 2876 22293 2904
rect 22281 2873 22293 2876
rect 22327 2873 22339 2907
rect 22281 2867 22339 2873
rect 18690 2836 18696 2848
rect 15856 2808 18696 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 21174 2836 21180 2848
rect 19300 2808 21180 2836
rect 19300 2796 19306 2808
rect 21174 2796 21180 2808
rect 21232 2836 21238 2848
rect 21637 2839 21695 2845
rect 21637 2836 21649 2839
rect 21232 2808 21649 2836
rect 21232 2796 21238 2808
rect 21637 2805 21649 2808
rect 21683 2805 21695 2839
rect 21637 2799 21695 2805
rect 1104 2746 22816 2768
rect 1104 2694 8246 2746
rect 8298 2694 8310 2746
rect 8362 2694 8374 2746
rect 8426 2694 8438 2746
rect 8490 2694 15510 2746
rect 15562 2694 15574 2746
rect 15626 2694 15638 2746
rect 15690 2694 15702 2746
rect 15754 2694 22816 2746
rect 1104 2672 22816 2694
rect 13814 2592 13820 2644
rect 13872 2632 13878 2644
rect 14369 2635 14427 2641
rect 14369 2632 14381 2635
rect 13872 2604 14381 2632
rect 13872 2592 13878 2604
rect 14369 2601 14381 2604
rect 14415 2601 14427 2635
rect 14369 2595 14427 2601
rect 14550 2592 14556 2644
rect 14608 2632 14614 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 14608 2604 14841 2632
rect 14608 2592 14614 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 15197 2635 15255 2641
rect 15197 2601 15209 2635
rect 15243 2632 15255 2635
rect 16850 2632 16856 2644
rect 15243 2604 16068 2632
rect 16811 2604 16856 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2564 12955 2567
rect 14642 2564 14648 2576
rect 12943 2536 14648 2564
rect 12943 2533 12955 2536
rect 12897 2527 12955 2533
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 14737 2567 14795 2573
rect 14737 2533 14749 2567
rect 14783 2564 14795 2567
rect 15286 2564 15292 2576
rect 14783 2536 15292 2564
rect 14783 2533 14795 2536
rect 14737 2527 14795 2533
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 15740 2567 15798 2573
rect 15740 2533 15752 2567
rect 15786 2564 15798 2567
rect 15930 2564 15936 2576
rect 15786 2536 15936 2564
rect 15786 2533 15798 2536
rect 15740 2527 15798 2533
rect 15930 2524 15936 2536
rect 15988 2524 15994 2576
rect 16040 2564 16068 2604
rect 16850 2592 16856 2604
rect 16908 2592 16914 2644
rect 17589 2635 17647 2641
rect 17589 2601 17601 2635
rect 17635 2632 17647 2635
rect 18138 2632 18144 2644
rect 17635 2604 18144 2632
rect 17635 2601 17647 2604
rect 17589 2595 17647 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18690 2592 18696 2644
rect 18748 2632 18754 2644
rect 19705 2635 19763 2641
rect 19705 2632 19717 2635
rect 18748 2604 19717 2632
rect 18748 2592 18754 2604
rect 19705 2601 19717 2604
rect 19751 2601 19763 2635
rect 19705 2595 19763 2601
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2632 20499 2635
rect 20714 2632 20720 2644
rect 20487 2604 20720 2632
rect 20487 2601 20499 2604
rect 20441 2595 20499 2601
rect 17034 2564 17040 2576
rect 16040 2536 17040 2564
rect 17034 2524 17040 2536
rect 17092 2524 17098 2576
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 18570 2567 18628 2573
rect 18570 2564 18582 2567
rect 18380 2536 18582 2564
rect 18380 2524 18386 2536
rect 18570 2533 18582 2536
rect 18616 2533 18628 2567
rect 18570 2527 18628 2533
rect 19242 2524 19248 2576
rect 19300 2524 19306 2576
rect 20088 2564 20116 2595
rect 20714 2592 20720 2604
rect 20772 2592 20778 2644
rect 21545 2567 21603 2573
rect 21545 2564 21557 2567
rect 20088 2536 21557 2564
rect 21545 2533 21557 2536
rect 21591 2533 21603 2567
rect 21545 2527 21603 2533
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 15010 2496 15016 2508
rect 13771 2468 15016 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 15473 2499 15531 2505
rect 15473 2465 15485 2499
rect 15519 2496 15531 2499
rect 16114 2496 16120 2508
rect 15519 2468 16120 2496
rect 15519 2465 15531 2468
rect 15473 2459 15531 2465
rect 16114 2456 16120 2468
rect 16172 2456 16178 2508
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 19260 2496 19288 2524
rect 17727 2468 19288 2496
rect 20533 2499 20591 2505
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 20533 2465 20545 2499
rect 20579 2496 20591 2499
rect 21266 2496 21272 2508
rect 20579 2468 21272 2496
rect 20579 2465 20591 2468
rect 20533 2459 20591 2465
rect 21266 2456 21272 2468
rect 21324 2456 21330 2508
rect 13817 2431 13875 2437
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 13832 2360 13860 2391
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14921 2431 14979 2437
rect 13964 2400 14009 2428
rect 13964 2388 13970 2400
rect 14921 2397 14933 2431
rect 14967 2428 14979 2431
rect 17770 2428 17776 2440
rect 14967 2400 15516 2428
rect 17731 2400 17776 2428
rect 14967 2397 14979 2400
rect 14921 2391 14979 2397
rect 15102 2360 15108 2372
rect 13832 2332 15108 2360
rect 15102 2320 15108 2332
rect 15160 2320 15166 2372
rect 13357 2295 13415 2301
rect 13357 2261 13369 2295
rect 13403 2292 13415 2295
rect 15197 2295 15255 2301
rect 15197 2292 15209 2295
rect 13403 2264 15209 2292
rect 13403 2261 13415 2264
rect 13357 2255 13415 2261
rect 15197 2261 15209 2264
rect 15243 2261 15255 2295
rect 15488 2292 15516 2400
rect 17770 2388 17776 2400
rect 17828 2388 17834 2440
rect 18322 2428 18328 2440
rect 18283 2400 18328 2428
rect 18322 2388 18328 2400
rect 18380 2388 18386 2440
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2428 20683 2431
rect 20714 2428 20720 2440
rect 20671 2400 20720 2428
rect 20671 2397 20683 2400
rect 20625 2391 20683 2397
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 21637 2431 21695 2437
rect 21637 2397 21649 2431
rect 21683 2397 21695 2431
rect 21637 2391 21695 2397
rect 21821 2431 21879 2437
rect 21821 2397 21833 2431
rect 21867 2428 21879 2431
rect 22094 2428 22100 2440
rect 21867 2400 22100 2428
rect 21867 2397 21879 2400
rect 21821 2391 21879 2397
rect 20070 2320 20076 2372
rect 20128 2360 20134 2372
rect 21177 2363 21235 2369
rect 21177 2360 21189 2363
rect 20128 2332 21189 2360
rect 20128 2320 20134 2332
rect 21177 2329 21189 2332
rect 21223 2329 21235 2363
rect 21177 2323 21235 2329
rect 16942 2292 16948 2304
rect 15488 2264 16948 2292
rect 15197 2255 15255 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2292 17279 2295
rect 21652 2292 21680 2391
rect 22094 2388 22100 2400
rect 22152 2388 22158 2440
rect 17267 2264 21680 2292
rect 17267 2261 17279 2264
rect 17221 2255 17279 2261
rect 1104 2202 22816 2224
rect 1104 2150 4614 2202
rect 4666 2150 4678 2202
rect 4730 2150 4742 2202
rect 4794 2150 4806 2202
rect 4858 2150 11878 2202
rect 11930 2150 11942 2202
rect 11994 2150 12006 2202
rect 12058 2150 12070 2202
rect 12122 2150 19142 2202
rect 19194 2150 19206 2202
rect 19258 2150 19270 2202
rect 19322 2150 19334 2202
rect 19386 2150 22816 2202
rect 1104 2128 22816 2150
rect 13722 2048 13728 2100
rect 13780 2088 13786 2100
rect 17770 2088 17776 2100
rect 13780 2060 17776 2088
rect 13780 2048 13786 2060
rect 17770 2048 17776 2060
rect 17828 2088 17834 2100
rect 20714 2088 20720 2100
rect 17828 2060 20720 2088
rect 17828 2048 17834 2060
rect 20714 2048 20720 2060
rect 20772 2048 20778 2100
<< via1 >>
rect 14280 22788 14332 22840
rect 19432 22788 19484 22840
rect 10508 22312 10560 22364
rect 17868 22312 17920 22364
rect 12164 22244 12216 22296
rect 17224 22244 17276 22296
rect 16580 22176 16632 22228
rect 19340 22176 19392 22228
rect 19616 22040 19668 22092
rect 14924 21972 14976 22024
rect 8668 21904 8720 21956
rect 18604 21904 18656 21956
rect 12716 21836 12768 21888
rect 21732 21836 21784 21888
rect 4614 21734 4666 21786
rect 4678 21734 4730 21786
rect 4742 21734 4794 21786
rect 4806 21734 4858 21786
rect 11878 21734 11930 21786
rect 11942 21734 11994 21786
rect 12006 21734 12058 21786
rect 12070 21734 12122 21786
rect 19142 21734 19194 21786
rect 19206 21734 19258 21786
rect 19270 21734 19322 21786
rect 19334 21734 19386 21786
rect 296 21632 348 21684
rect 3240 21496 3292 21548
rect 4344 21632 4396 21684
rect 3608 21564 3660 21616
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 3700 21496 3752 21548
rect 4988 21564 5040 21616
rect 8116 21632 8168 21684
rect 9680 21564 9732 21616
rect 14832 21607 14884 21616
rect 3884 21428 3936 21480
rect 4160 21428 4212 21480
rect 4896 21428 4948 21480
rect 6828 21496 6880 21548
rect 7932 21496 7984 21548
rect 14832 21573 14841 21607
rect 14841 21573 14875 21607
rect 14875 21573 14884 21607
rect 14832 21564 14884 21573
rect 6644 21428 6696 21480
rect 1400 21292 1452 21344
rect 2596 21292 2648 21344
rect 2964 21335 3016 21344
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 3332 21335 3384 21344
rect 3332 21301 3341 21335
rect 3341 21301 3375 21335
rect 3375 21301 3384 21335
rect 3332 21292 3384 21301
rect 8576 21428 8628 21480
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9588 21428 9640 21480
rect 12532 21496 12584 21548
rect 14464 21496 14516 21548
rect 17316 21632 17368 21684
rect 12624 21471 12676 21480
rect 12624 21437 12633 21471
rect 12633 21437 12667 21471
rect 12667 21437 12676 21471
rect 12624 21428 12676 21437
rect 16212 21428 16264 21480
rect 16396 21428 16448 21480
rect 17684 21471 17736 21480
rect 17684 21437 17693 21471
rect 17693 21437 17727 21471
rect 17727 21437 17736 21471
rect 17684 21428 17736 21437
rect 5080 21335 5132 21344
rect 5080 21301 5089 21335
rect 5089 21301 5123 21335
rect 5123 21301 5132 21335
rect 5080 21292 5132 21301
rect 5264 21292 5316 21344
rect 9956 21360 10008 21412
rect 8116 21292 8168 21344
rect 8668 21292 8720 21344
rect 9036 21335 9088 21344
rect 9036 21301 9045 21335
rect 9045 21301 9079 21335
rect 9079 21301 9088 21335
rect 9036 21292 9088 21301
rect 11060 21292 11112 21344
rect 12164 21292 12216 21344
rect 12808 21335 12860 21344
rect 12808 21301 12817 21335
rect 12817 21301 12851 21335
rect 12851 21301 12860 21335
rect 12808 21292 12860 21301
rect 13912 21360 13964 21412
rect 14648 21360 14700 21412
rect 15384 21292 15436 21344
rect 17224 21360 17276 21412
rect 20536 21496 20588 21548
rect 21732 21539 21784 21548
rect 21732 21505 21741 21539
rect 21741 21505 21775 21539
rect 21775 21505 21784 21539
rect 21732 21496 21784 21505
rect 19064 21428 19116 21480
rect 19984 21360 20036 21412
rect 20720 21360 20772 21412
rect 21732 21360 21784 21412
rect 15936 21335 15988 21344
rect 15936 21301 15945 21335
rect 15945 21301 15979 21335
rect 15979 21301 15988 21335
rect 15936 21292 15988 21301
rect 16028 21292 16080 21344
rect 16856 21335 16908 21344
rect 16856 21301 16865 21335
rect 16865 21301 16899 21335
rect 16899 21301 16908 21335
rect 16856 21292 16908 21301
rect 17132 21292 17184 21344
rect 19432 21292 19484 21344
rect 20812 21292 20864 21344
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 8246 21190 8298 21242
rect 8310 21190 8362 21242
rect 8374 21190 8426 21242
rect 8438 21190 8490 21242
rect 15510 21190 15562 21242
rect 15574 21190 15626 21242
rect 15638 21190 15690 21242
rect 15702 21190 15754 21242
rect 3608 21088 3660 21140
rect 5080 21088 5132 21140
rect 8576 21088 8628 21140
rect 9312 21088 9364 21140
rect 12256 21088 12308 21140
rect 14464 21088 14516 21140
rect 14924 21088 14976 21140
rect 16580 21088 16632 21140
rect 17224 21131 17276 21140
rect 17224 21097 17233 21131
rect 17233 21097 17267 21131
rect 17267 21097 17276 21131
rect 17224 21088 17276 21097
rect 17684 21088 17736 21140
rect 19708 21088 19760 21140
rect 2780 21020 2832 21072
rect 3700 21020 3752 21072
rect 2136 20927 2188 20936
rect 2136 20893 2145 20927
rect 2145 20893 2179 20927
rect 2179 20893 2188 20927
rect 2136 20884 2188 20893
rect 6184 20952 6236 21004
rect 7932 21020 7984 21072
rect 13820 21020 13872 21072
rect 6920 20952 6972 21004
rect 4252 20884 4304 20936
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 6276 20884 6328 20936
rect 7104 20952 7156 21004
rect 7748 20952 7800 21004
rect 10416 20995 10468 21004
rect 10416 20961 10425 20995
rect 10425 20961 10459 20995
rect 10459 20961 10468 20995
rect 10416 20952 10468 20961
rect 12256 20952 12308 21004
rect 14556 20952 14608 21004
rect 16764 21020 16816 21072
rect 17868 21020 17920 21072
rect 19064 21020 19116 21072
rect 16120 20995 16172 21004
rect 16120 20961 16154 20995
rect 16154 20961 16172 20995
rect 16120 20952 16172 20961
rect 18328 20952 18380 21004
rect 20812 20952 20864 21004
rect 20904 20952 20956 21004
rect 1952 20748 2004 20800
rect 3884 20748 3936 20800
rect 5356 20748 5408 20800
rect 6644 20791 6696 20800
rect 6644 20757 6653 20791
rect 6653 20757 6687 20791
rect 6687 20757 6696 20791
rect 6644 20748 6696 20757
rect 9772 20884 9824 20936
rect 10968 20884 11020 20936
rect 10600 20816 10652 20868
rect 12532 20884 12584 20936
rect 8576 20748 8628 20800
rect 9496 20748 9548 20800
rect 10784 20748 10836 20800
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 13912 20748 13964 20800
rect 15476 20748 15528 20800
rect 16948 20748 17000 20800
rect 18972 20884 19024 20936
rect 18696 20816 18748 20868
rect 18420 20748 18472 20800
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 21272 20816 21324 20868
rect 20720 20748 20772 20800
rect 20996 20748 21048 20800
rect 22100 20791 22152 20800
rect 22100 20757 22109 20791
rect 22109 20757 22143 20791
rect 22143 20757 22152 20791
rect 22100 20748 22152 20757
rect 4614 20646 4666 20698
rect 4678 20646 4730 20698
rect 4742 20646 4794 20698
rect 4806 20646 4858 20698
rect 11878 20646 11930 20698
rect 11942 20646 11994 20698
rect 12006 20646 12058 20698
rect 12070 20646 12122 20698
rect 19142 20646 19194 20698
rect 19206 20646 19258 20698
rect 19270 20646 19322 20698
rect 19334 20646 19386 20698
rect 2780 20587 2832 20596
rect 2780 20553 2789 20587
rect 2789 20553 2823 20587
rect 2823 20553 2832 20587
rect 2780 20544 2832 20553
rect 2964 20544 3016 20596
rect 3792 20544 3844 20596
rect 4068 20544 4120 20596
rect 4252 20544 4304 20596
rect 5908 20544 5960 20596
rect 4804 20476 4856 20528
rect 1492 20340 1544 20392
rect 2136 20340 2188 20392
rect 4896 20340 4948 20392
rect 5356 20340 5408 20392
rect 5448 20340 5500 20392
rect 8024 20544 8076 20596
rect 8116 20544 8168 20596
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 7104 20383 7156 20392
rect 7104 20349 7138 20383
rect 7138 20349 7156 20383
rect 7104 20340 7156 20349
rect 2964 20272 3016 20324
rect 3608 20272 3660 20324
rect 4436 20272 4488 20324
rect 11336 20544 11388 20596
rect 11612 20544 11664 20596
rect 12256 20544 12308 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 14740 20476 14792 20528
rect 16120 20476 16172 20528
rect 16396 20476 16448 20528
rect 9680 20408 9732 20460
rect 20812 20544 20864 20596
rect 18972 20476 19024 20528
rect 8576 20383 8628 20392
rect 8576 20349 8585 20383
rect 8585 20349 8619 20383
rect 8619 20349 8628 20383
rect 8576 20340 8628 20349
rect 9128 20340 9180 20392
rect 9588 20340 9640 20392
rect 10600 20340 10652 20392
rect 9496 20272 9548 20324
rect 12164 20340 12216 20392
rect 12532 20340 12584 20392
rect 17316 20408 17368 20460
rect 17500 20408 17552 20460
rect 18696 20408 18748 20460
rect 19340 20408 19392 20460
rect 20536 20408 20588 20460
rect 21456 20408 21508 20460
rect 14924 20383 14976 20392
rect 14924 20349 14933 20383
rect 14933 20349 14967 20383
rect 14967 20349 14976 20383
rect 14924 20340 14976 20349
rect 15016 20340 15068 20392
rect 15200 20383 15252 20392
rect 15200 20349 15234 20383
rect 15234 20349 15252 20383
rect 15200 20340 15252 20349
rect 15476 20340 15528 20392
rect 18512 20340 18564 20392
rect 19432 20340 19484 20392
rect 10968 20315 11020 20324
rect 2412 20204 2464 20256
rect 4160 20204 4212 20256
rect 5356 20204 5408 20256
rect 6184 20247 6236 20256
rect 6184 20213 6193 20247
rect 6193 20213 6227 20247
rect 6227 20213 6236 20247
rect 6184 20204 6236 20213
rect 8668 20204 8720 20256
rect 10968 20281 11002 20315
rect 11002 20281 11020 20315
rect 10968 20272 11020 20281
rect 12716 20315 12768 20324
rect 12716 20281 12750 20315
rect 12750 20281 12768 20315
rect 12716 20272 12768 20281
rect 16856 20272 16908 20324
rect 19984 20272 20036 20324
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 11336 20204 11388 20256
rect 12808 20204 12860 20256
rect 14280 20204 14332 20256
rect 16396 20204 16448 20256
rect 18788 20204 18840 20256
rect 21548 20247 21600 20256
rect 21548 20213 21557 20247
rect 21557 20213 21591 20247
rect 21591 20213 21600 20247
rect 21548 20204 21600 20213
rect 21640 20247 21692 20256
rect 21640 20213 21649 20247
rect 21649 20213 21683 20247
rect 21683 20213 21692 20247
rect 21640 20204 21692 20213
rect 8246 20102 8298 20154
rect 8310 20102 8362 20154
rect 8374 20102 8426 20154
rect 8438 20102 8490 20154
rect 15510 20102 15562 20154
rect 15574 20102 15626 20154
rect 15638 20102 15690 20154
rect 15702 20102 15754 20154
rect 2412 20043 2464 20052
rect 2412 20009 2421 20043
rect 2421 20009 2455 20043
rect 2455 20009 2464 20043
rect 2412 20000 2464 20009
rect 3240 20000 3292 20052
rect 6184 20000 6236 20052
rect 4252 19932 4304 19984
rect 4804 19932 4856 19984
rect 6092 19932 6144 19984
rect 9036 20000 9088 20052
rect 15200 20000 15252 20052
rect 1768 19907 1820 19916
rect 1768 19873 1777 19907
rect 1777 19873 1811 19907
rect 1811 19873 1820 19907
rect 1768 19864 1820 19873
rect 2872 19907 2924 19916
rect 2872 19873 2881 19907
rect 2881 19873 2915 19907
rect 2915 19873 2924 19907
rect 2872 19864 2924 19873
rect 3424 19907 3476 19916
rect 3424 19873 3433 19907
rect 3433 19873 3467 19907
rect 3467 19873 3476 19907
rect 3424 19864 3476 19873
rect 3608 19864 3660 19916
rect 1860 19839 1912 19848
rect 1860 19805 1869 19839
rect 1869 19805 1903 19839
rect 1903 19805 1912 19839
rect 1860 19796 1912 19805
rect 1952 19839 2004 19848
rect 1952 19805 1961 19839
rect 1961 19805 1995 19839
rect 1995 19805 2004 19839
rect 1952 19796 2004 19805
rect 2412 19796 2464 19848
rect 2964 19839 3016 19848
rect 2964 19805 2973 19839
rect 2973 19805 3007 19839
rect 3007 19805 3016 19839
rect 2964 19796 3016 19805
rect 3700 19796 3752 19848
rect 4620 19839 4672 19848
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 5080 19796 5132 19848
rect 5356 19796 5408 19848
rect 6552 19796 6604 19848
rect 6736 19796 6788 19848
rect 8668 19864 8720 19916
rect 8852 19907 8904 19916
rect 8852 19873 8861 19907
rect 8861 19873 8895 19907
rect 8895 19873 8904 19907
rect 8852 19864 8904 19873
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 12164 19932 12216 19984
rect 15384 20000 15436 20052
rect 15936 20000 15988 20052
rect 15844 19932 15896 19984
rect 12072 19864 12124 19916
rect 7104 19796 7156 19805
rect 3516 19660 3568 19712
rect 5264 19660 5316 19712
rect 8668 19660 8720 19712
rect 10324 19839 10376 19848
rect 10324 19805 10333 19839
rect 10333 19805 10367 19839
rect 10367 19805 10376 19839
rect 10324 19796 10376 19805
rect 10600 19796 10652 19848
rect 11060 19796 11112 19848
rect 11244 19796 11296 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 11612 19796 11664 19848
rect 12900 19864 12952 19916
rect 14832 19864 14884 19916
rect 16488 20000 16540 20052
rect 18328 20043 18380 20052
rect 17224 19975 17276 19984
rect 17224 19941 17258 19975
rect 17258 19941 17276 19975
rect 17224 19932 17276 19941
rect 18328 20009 18337 20043
rect 18337 20009 18371 20043
rect 18371 20009 18380 20043
rect 18328 20000 18380 20009
rect 19524 20000 19576 20052
rect 21548 20000 21600 20052
rect 20260 19932 20312 19984
rect 20720 19932 20772 19984
rect 18604 19907 18656 19916
rect 12532 19796 12584 19848
rect 13452 19796 13504 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14648 19796 14700 19848
rect 15568 19796 15620 19848
rect 16948 19839 17000 19848
rect 9220 19728 9272 19780
rect 10508 19728 10560 19780
rect 16948 19805 16957 19839
rect 16957 19805 16991 19839
rect 16991 19805 17000 19839
rect 16948 19796 17000 19805
rect 9772 19660 9824 19712
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 12624 19660 12676 19712
rect 14740 19660 14792 19712
rect 16580 19660 16632 19712
rect 18604 19873 18613 19907
rect 18613 19873 18647 19907
rect 18647 19873 18656 19907
rect 18604 19864 18656 19873
rect 19248 19864 19300 19916
rect 20812 19864 20864 19916
rect 20352 19796 20404 19848
rect 4614 19558 4666 19610
rect 4678 19558 4730 19610
rect 4742 19558 4794 19610
rect 4806 19558 4858 19610
rect 11878 19558 11930 19610
rect 11942 19558 11994 19610
rect 12006 19558 12058 19610
rect 12070 19558 12122 19610
rect 19142 19558 19194 19610
rect 19206 19558 19258 19610
rect 19270 19558 19322 19610
rect 19334 19558 19386 19610
rect 2320 19456 2372 19508
rect 2964 19456 3016 19508
rect 3056 19456 3108 19508
rect 4160 19456 4212 19508
rect 4436 19456 4488 19508
rect 4988 19456 5040 19508
rect 5172 19456 5224 19508
rect 6184 19456 6236 19508
rect 6368 19456 6420 19508
rect 8668 19456 8720 19508
rect 8852 19456 8904 19508
rect 10140 19456 10192 19508
rect 2412 19320 2464 19372
rect 4068 19320 4120 19372
rect 1492 19252 1544 19304
rect 3056 19252 3108 19304
rect 4528 19252 4580 19304
rect 4988 19320 5040 19372
rect 6092 19320 6144 19372
rect 6920 19320 6972 19372
rect 7564 19320 7616 19372
rect 8576 19320 8628 19372
rect 13176 19456 13228 19508
rect 12348 19388 12400 19440
rect 13268 19388 13320 19440
rect 12808 19320 12860 19372
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 5264 19252 5316 19304
rect 3240 19184 3292 19236
rect 2964 19116 3016 19168
rect 3148 19116 3200 19168
rect 6828 19252 6880 19304
rect 8208 19295 8260 19304
rect 7380 19184 7432 19236
rect 6644 19116 6696 19168
rect 7840 19116 7892 19168
rect 8208 19261 8217 19295
rect 8217 19261 8251 19295
rect 8251 19261 8260 19295
rect 8208 19252 8260 19261
rect 8116 19184 8168 19236
rect 9680 19252 9732 19304
rect 10600 19252 10652 19304
rect 12440 19252 12492 19304
rect 20812 19499 20864 19508
rect 13544 19388 13596 19440
rect 13636 19320 13688 19372
rect 15200 19388 15252 19440
rect 14188 19295 14240 19304
rect 14188 19261 14197 19295
rect 14197 19261 14231 19295
rect 14231 19261 14240 19295
rect 14188 19252 14240 19261
rect 12256 19184 12308 19236
rect 12532 19184 12584 19236
rect 13636 19227 13688 19236
rect 9588 19116 9640 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 10324 19159 10376 19168
rect 10324 19125 10333 19159
rect 10333 19125 10367 19159
rect 10367 19125 10376 19159
rect 10324 19116 10376 19125
rect 10416 19116 10468 19168
rect 10968 19116 11020 19168
rect 12808 19159 12860 19168
rect 12808 19125 12817 19159
rect 12817 19125 12851 19159
rect 12851 19125 12860 19159
rect 12808 19116 12860 19125
rect 12900 19159 12952 19168
rect 12900 19125 12909 19159
rect 12909 19125 12943 19159
rect 12943 19125 12952 19159
rect 13636 19193 13645 19227
rect 13645 19193 13679 19227
rect 13679 19193 13688 19227
rect 13636 19184 13688 19193
rect 14648 19184 14700 19236
rect 17868 19388 17920 19440
rect 18052 19431 18104 19440
rect 18052 19397 18061 19431
rect 18061 19397 18095 19431
rect 18095 19397 18104 19431
rect 18052 19388 18104 19397
rect 20812 19465 20821 19499
rect 20821 19465 20855 19499
rect 20855 19465 20864 19499
rect 20812 19456 20864 19465
rect 21640 19456 21692 19508
rect 17500 19320 17552 19372
rect 17592 19363 17644 19372
rect 17592 19329 17601 19363
rect 17601 19329 17635 19363
rect 17635 19329 17644 19363
rect 17592 19320 17644 19329
rect 18328 19320 18380 19372
rect 21180 19388 21232 19440
rect 21456 19363 21508 19372
rect 21456 19329 21465 19363
rect 21465 19329 21499 19363
rect 21499 19329 21508 19363
rect 21456 19320 21508 19329
rect 18236 19252 18288 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 19340 19252 19392 19304
rect 12900 19116 12952 19125
rect 14280 19116 14332 19168
rect 15384 19116 15436 19168
rect 18880 19184 18932 19236
rect 16120 19116 16172 19168
rect 21364 19252 21416 19304
rect 20536 19184 20588 19236
rect 20904 19159 20956 19168
rect 20904 19125 20913 19159
rect 20913 19125 20947 19159
rect 20947 19125 20956 19159
rect 21364 19159 21416 19168
rect 20904 19116 20956 19125
rect 21364 19125 21373 19159
rect 21373 19125 21407 19159
rect 21407 19125 21416 19159
rect 21364 19116 21416 19125
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 21916 19116 21968 19125
rect 8246 19014 8298 19066
rect 8310 19014 8362 19066
rect 8374 19014 8426 19066
rect 8438 19014 8490 19066
rect 15510 19014 15562 19066
rect 15574 19014 15626 19066
rect 15638 19014 15690 19066
rect 15702 19014 15754 19066
rect 2872 18912 2924 18964
rect 3240 18912 3292 18964
rect 4252 18955 4304 18964
rect 4252 18921 4261 18955
rect 4261 18921 4295 18955
rect 4295 18921 4304 18955
rect 4252 18912 4304 18921
rect 5172 18912 5224 18964
rect 1768 18844 1820 18896
rect 2228 18887 2280 18896
rect 2228 18853 2240 18887
rect 2240 18853 2280 18887
rect 2228 18844 2280 18853
rect 5448 18844 5500 18896
rect 6552 18912 6604 18964
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 8116 18912 8168 18964
rect 6460 18887 6512 18896
rect 1400 18819 1452 18828
rect 1400 18785 1409 18819
rect 1409 18785 1443 18819
rect 1443 18785 1452 18819
rect 1400 18776 1452 18785
rect 2504 18776 2556 18828
rect 6092 18819 6144 18828
rect 6092 18785 6101 18819
rect 6101 18785 6135 18819
rect 6135 18785 6144 18819
rect 6092 18776 6144 18785
rect 6460 18853 6494 18887
rect 6494 18853 6512 18887
rect 6460 18844 6512 18853
rect 6736 18776 6788 18828
rect 7012 18776 7064 18828
rect 7196 18776 7248 18828
rect 1492 18708 1544 18760
rect 4988 18708 5040 18760
rect 5724 18708 5776 18760
rect 8576 18912 8628 18964
rect 8576 18776 8628 18828
rect 12164 18844 12216 18896
rect 12808 18912 12860 18964
rect 16488 18912 16540 18964
rect 18880 18955 18932 18964
rect 10416 18819 10468 18828
rect 10416 18785 10425 18819
rect 10425 18785 10459 18819
rect 10459 18785 10468 18819
rect 10416 18776 10468 18785
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 11520 18776 11572 18828
rect 12440 18776 12492 18828
rect 12716 18776 12768 18828
rect 13636 18776 13688 18828
rect 4344 18572 4396 18624
rect 5356 18572 5408 18624
rect 10600 18751 10652 18760
rect 10600 18717 10609 18751
rect 10609 18717 10643 18751
rect 10643 18717 10652 18751
rect 12164 18751 12216 18760
rect 10600 18708 10652 18717
rect 12164 18717 12173 18751
rect 12173 18717 12207 18751
rect 12207 18717 12216 18751
rect 12164 18708 12216 18717
rect 11060 18640 11112 18692
rect 7564 18615 7616 18624
rect 7564 18581 7573 18615
rect 7573 18581 7607 18615
rect 7607 18581 7616 18615
rect 7564 18572 7616 18581
rect 8944 18572 8996 18624
rect 11244 18615 11296 18624
rect 11244 18581 11253 18615
rect 11253 18581 11287 18615
rect 11287 18581 11296 18615
rect 12624 18640 12676 18692
rect 11244 18572 11296 18581
rect 12348 18572 12400 18624
rect 12532 18572 12584 18624
rect 15936 18844 15988 18896
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 19156 18912 19208 18964
rect 19340 18912 19392 18964
rect 20352 18912 20404 18964
rect 20536 18955 20588 18964
rect 20536 18921 20545 18955
rect 20545 18921 20579 18955
rect 20579 18921 20588 18955
rect 20536 18912 20588 18921
rect 14280 18819 14332 18828
rect 14280 18785 14289 18819
rect 14289 18785 14323 18819
rect 14323 18785 14332 18819
rect 14280 18776 14332 18785
rect 14740 18776 14792 18828
rect 18420 18844 18472 18896
rect 21364 18844 21416 18896
rect 16580 18776 16632 18828
rect 21088 18776 21140 18828
rect 14188 18708 14240 18760
rect 14924 18708 14976 18760
rect 19156 18751 19208 18760
rect 14464 18683 14516 18692
rect 14464 18649 14473 18683
rect 14473 18649 14507 18683
rect 14507 18649 14516 18683
rect 14464 18640 14516 18649
rect 16948 18640 17000 18692
rect 19156 18717 19165 18751
rect 19165 18717 19199 18751
rect 19199 18717 19208 18751
rect 19156 18708 19208 18717
rect 21824 18708 21876 18760
rect 21548 18640 21600 18692
rect 15936 18572 15988 18624
rect 16672 18615 16724 18624
rect 16672 18581 16681 18615
rect 16681 18581 16715 18615
rect 16715 18581 16724 18615
rect 16672 18572 16724 18581
rect 16856 18572 16908 18624
rect 20628 18572 20680 18624
rect 20904 18615 20956 18624
rect 20904 18581 20913 18615
rect 20913 18581 20947 18615
rect 20947 18581 20956 18615
rect 20904 18572 20956 18581
rect 20996 18572 21048 18624
rect 4614 18470 4666 18522
rect 4678 18470 4730 18522
rect 4742 18470 4794 18522
rect 4806 18470 4858 18522
rect 11878 18470 11930 18522
rect 11942 18470 11994 18522
rect 12006 18470 12058 18522
rect 12070 18470 12122 18522
rect 19142 18470 19194 18522
rect 19206 18470 19258 18522
rect 19270 18470 19322 18522
rect 19334 18470 19386 18522
rect 2228 18368 2280 18420
rect 3424 18368 3476 18420
rect 6460 18411 6512 18420
rect 3240 18232 3292 18284
rect 6460 18377 6469 18411
rect 6469 18377 6503 18411
rect 6503 18377 6512 18411
rect 6460 18368 6512 18377
rect 6736 18368 6788 18420
rect 9864 18368 9916 18420
rect 11612 18368 11664 18420
rect 6644 18300 6696 18352
rect 10048 18300 10100 18352
rect 11428 18300 11480 18352
rect 11520 18300 11572 18352
rect 11796 18300 11848 18352
rect 1492 18164 1544 18216
rect 1860 18207 1912 18216
rect 1860 18173 1894 18207
rect 1894 18173 1912 18207
rect 1860 18164 1912 18173
rect 4344 18164 4396 18216
rect 6552 18232 6604 18284
rect 10600 18232 10652 18284
rect 12164 18232 12216 18284
rect 12256 18232 12308 18284
rect 12716 18368 12768 18420
rect 13636 18368 13688 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 14464 18368 14516 18420
rect 14648 18368 14700 18420
rect 16672 18368 16724 18420
rect 19616 18368 19668 18420
rect 21364 18368 21416 18420
rect 18696 18300 18748 18352
rect 17132 18275 17184 18284
rect 17132 18241 17141 18275
rect 17141 18241 17175 18275
rect 17175 18241 17184 18275
rect 17132 18232 17184 18241
rect 17224 18275 17276 18284
rect 17224 18241 17233 18275
rect 17233 18241 17267 18275
rect 17267 18241 17276 18275
rect 17224 18232 17276 18241
rect 6736 18164 6788 18216
rect 7564 18164 7616 18216
rect 9128 18164 9180 18216
rect 10324 18164 10376 18216
rect 13176 18164 13228 18216
rect 13268 18164 13320 18216
rect 14188 18164 14240 18216
rect 5172 18096 5224 18148
rect 5724 18096 5776 18148
rect 7748 18096 7800 18148
rect 4344 18028 4396 18080
rect 5080 18028 5132 18080
rect 8116 18028 8168 18080
rect 8944 18096 8996 18148
rect 11152 18096 11204 18148
rect 12348 18096 12400 18148
rect 12532 18096 12584 18148
rect 12716 18139 12768 18148
rect 12716 18105 12750 18139
rect 12750 18105 12768 18139
rect 12716 18096 12768 18105
rect 18052 18164 18104 18216
rect 18420 18164 18472 18216
rect 21180 18232 21232 18284
rect 21824 18232 21876 18284
rect 20628 18164 20680 18216
rect 15200 18139 15252 18148
rect 15200 18105 15234 18139
rect 15234 18105 15252 18139
rect 15200 18096 15252 18105
rect 10600 18071 10652 18080
rect 10600 18037 10609 18071
rect 10609 18037 10643 18071
rect 10643 18037 10652 18071
rect 11336 18071 11388 18080
rect 10600 18028 10652 18037
rect 11336 18037 11345 18071
rect 11345 18037 11379 18071
rect 11379 18037 11388 18071
rect 11336 18028 11388 18037
rect 11428 18028 11480 18080
rect 13268 18028 13320 18080
rect 13728 18028 13780 18080
rect 14924 18028 14976 18080
rect 15016 18028 15068 18080
rect 16120 18028 16172 18080
rect 16672 18071 16724 18080
rect 16672 18037 16681 18071
rect 16681 18037 16715 18071
rect 16715 18037 16724 18071
rect 16672 18028 16724 18037
rect 18236 18096 18288 18148
rect 19248 18096 19300 18148
rect 21456 18096 21508 18148
rect 19892 18028 19944 18080
rect 20168 18028 20220 18080
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 20812 18071 20864 18080
rect 20812 18037 20821 18071
rect 20821 18037 20855 18071
rect 20855 18037 20864 18071
rect 21364 18071 21416 18080
rect 20812 18028 20864 18037
rect 21364 18037 21373 18071
rect 21373 18037 21407 18071
rect 21407 18037 21416 18071
rect 21364 18028 21416 18037
rect 21732 18071 21784 18080
rect 21732 18037 21741 18071
rect 21741 18037 21775 18071
rect 21775 18037 21784 18071
rect 21732 18028 21784 18037
rect 8246 17926 8298 17978
rect 8310 17926 8362 17978
rect 8374 17926 8426 17978
rect 8438 17926 8490 17978
rect 15510 17926 15562 17978
rect 15574 17926 15626 17978
rect 15638 17926 15690 17978
rect 15702 17926 15754 17978
rect 1860 17824 1912 17876
rect 3332 17824 3384 17876
rect 5172 17824 5224 17876
rect 5724 17867 5776 17876
rect 5724 17833 5733 17867
rect 5733 17833 5767 17867
rect 5767 17833 5776 17867
rect 5724 17824 5776 17833
rect 6184 17867 6236 17876
rect 6184 17833 6193 17867
rect 6193 17833 6227 17867
rect 6227 17833 6236 17867
rect 6184 17824 6236 17833
rect 2136 17756 2188 17808
rect 3976 17756 4028 17808
rect 2228 17688 2280 17740
rect 3516 17688 3568 17740
rect 5356 17756 5408 17808
rect 5172 17688 5224 17740
rect 5908 17688 5960 17740
rect 6460 17688 6512 17740
rect 6552 17688 6604 17740
rect 7012 17824 7064 17876
rect 7288 17824 7340 17876
rect 10600 17824 10652 17876
rect 12716 17824 12768 17876
rect 9772 17756 9824 17808
rect 6828 17688 6880 17740
rect 8852 17731 8904 17740
rect 8852 17697 8861 17731
rect 8861 17697 8895 17731
rect 8895 17697 8904 17731
rect 8852 17688 8904 17697
rect 10508 17688 10560 17740
rect 11704 17756 11756 17808
rect 12256 17756 12308 17808
rect 12440 17756 12492 17808
rect 16396 17824 16448 17876
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 16028 17756 16080 17808
rect 17224 17824 17276 17876
rect 19248 17824 19300 17876
rect 21364 17824 21416 17876
rect 22100 17867 22152 17876
rect 22100 17833 22109 17867
rect 22109 17833 22143 17867
rect 22143 17833 22152 17867
rect 22100 17824 22152 17833
rect 13820 17688 13872 17740
rect 14004 17688 14056 17740
rect 1492 17620 1544 17672
rect 7196 17663 7248 17672
rect 7196 17629 7208 17663
rect 7208 17629 7242 17663
rect 7242 17629 7248 17663
rect 7472 17663 7524 17672
rect 7196 17620 7248 17629
rect 7472 17629 7481 17663
rect 7481 17629 7515 17663
rect 7515 17629 7524 17663
rect 7472 17620 7524 17629
rect 7840 17620 7892 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10183 17663
rect 10183 17629 10192 17663
rect 10140 17620 10192 17629
rect 11704 17620 11756 17672
rect 12164 17620 12216 17672
rect 14096 17620 14148 17672
rect 14740 17663 14792 17672
rect 14740 17629 14749 17663
rect 14749 17629 14783 17663
rect 14783 17629 14792 17663
rect 14740 17620 14792 17629
rect 15016 17620 15068 17672
rect 17040 17756 17092 17808
rect 18880 17756 18932 17808
rect 18972 17756 19024 17808
rect 23572 17756 23624 17808
rect 20168 17731 20220 17740
rect 2320 17484 2372 17536
rect 4068 17484 4120 17536
rect 11796 17552 11848 17604
rect 20168 17697 20177 17731
rect 20177 17697 20211 17731
rect 20211 17697 20220 17731
rect 20168 17688 20220 17697
rect 20904 17688 20956 17740
rect 16856 17663 16908 17672
rect 16856 17629 16865 17663
rect 16865 17629 16899 17663
rect 16899 17629 16908 17663
rect 16856 17620 16908 17629
rect 18144 17620 18196 17672
rect 18420 17620 18472 17672
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 12348 17484 12400 17536
rect 12624 17484 12676 17536
rect 14648 17484 14700 17536
rect 17132 17484 17184 17536
rect 18696 17484 18748 17536
rect 21180 17552 21232 17604
rect 21364 17552 21416 17604
rect 20352 17527 20404 17536
rect 20352 17493 20361 17527
rect 20361 17493 20395 17527
rect 20395 17493 20404 17527
rect 20352 17484 20404 17493
rect 20536 17484 20588 17536
rect 4614 17382 4666 17434
rect 4678 17382 4730 17434
rect 4742 17382 4794 17434
rect 4806 17382 4858 17434
rect 11878 17382 11930 17434
rect 11942 17382 11994 17434
rect 12006 17382 12058 17434
rect 12070 17382 12122 17434
rect 19142 17382 19194 17434
rect 19206 17382 19258 17434
rect 19270 17382 19322 17434
rect 19334 17382 19386 17434
rect 940 17280 992 17332
rect 2228 17280 2280 17332
rect 3608 17323 3660 17332
rect 3608 17289 3617 17323
rect 3617 17289 3651 17323
rect 3651 17289 3660 17323
rect 3608 17280 3660 17289
rect 10508 17323 10560 17332
rect 2136 17076 2188 17128
rect 2228 17119 2280 17128
rect 2228 17085 2237 17119
rect 2237 17085 2271 17119
rect 2271 17085 2280 17119
rect 2228 17076 2280 17085
rect 3700 17076 3752 17128
rect 3792 17076 3844 17128
rect 4344 17144 4396 17196
rect 5264 17144 5316 17196
rect 7472 17212 7524 17264
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 11428 17280 11480 17332
rect 12440 17280 12492 17332
rect 13820 17323 13872 17332
rect 13820 17289 13829 17323
rect 13829 17289 13863 17323
rect 13863 17289 13872 17323
rect 13820 17280 13872 17289
rect 20812 17280 20864 17332
rect 12164 17212 12216 17264
rect 14188 17212 14240 17264
rect 14280 17212 14332 17264
rect 17960 17212 18012 17264
rect 6644 17144 6696 17196
rect 4620 17119 4672 17128
rect 4620 17085 4629 17119
rect 4629 17085 4663 17119
rect 4663 17085 4672 17119
rect 4620 17076 4672 17085
rect 6368 17076 6420 17128
rect 6552 17076 6604 17128
rect 7012 17076 7064 17128
rect 6736 17008 6788 17060
rect 8024 17076 8076 17128
rect 2504 16940 2556 16992
rect 4436 16940 4488 16992
rect 6828 16940 6880 16992
rect 6920 16940 6972 16992
rect 9128 17008 9180 17060
rect 11704 17144 11756 17196
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 8576 16940 8628 16992
rect 10140 17076 10192 17128
rect 10784 17119 10836 17128
rect 10784 17085 10793 17119
rect 10793 17085 10827 17119
rect 10827 17085 10836 17119
rect 10784 17076 10836 17085
rect 9588 17008 9640 17060
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 12532 17008 12584 17060
rect 12808 17008 12860 17060
rect 12624 16940 12676 16992
rect 13176 17076 13228 17128
rect 17500 17144 17552 17196
rect 19708 17144 19760 17196
rect 20812 17144 20864 17196
rect 21824 17144 21876 17196
rect 13544 17076 13596 17128
rect 14188 17076 14240 17128
rect 14924 17076 14976 17128
rect 16856 17076 16908 17128
rect 17868 17119 17920 17128
rect 14740 17008 14792 17060
rect 15384 17008 15436 17060
rect 16120 17008 16172 17060
rect 16488 17008 16540 17060
rect 15200 16940 15252 16992
rect 17040 16940 17092 16992
rect 17868 17085 17877 17119
rect 17877 17085 17911 17119
rect 17911 17085 17920 17119
rect 17868 17076 17920 17085
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 19064 17076 19116 17128
rect 18144 16940 18196 16992
rect 20444 17076 20496 17128
rect 20996 16940 21048 16992
rect 21180 16983 21232 16992
rect 21180 16949 21189 16983
rect 21189 16949 21223 16983
rect 21223 16949 21232 16983
rect 21180 16940 21232 16949
rect 21824 16983 21876 16992
rect 21824 16949 21833 16983
rect 21833 16949 21867 16983
rect 21867 16949 21876 16983
rect 21824 16940 21876 16949
rect 8246 16838 8298 16890
rect 8310 16838 8362 16890
rect 8374 16838 8426 16890
rect 8438 16838 8490 16890
rect 15510 16838 15562 16890
rect 15574 16838 15626 16890
rect 15638 16838 15690 16890
rect 15702 16838 15754 16890
rect 1676 16736 1728 16788
rect 2136 16736 2188 16788
rect 4068 16736 4120 16788
rect 4252 16779 4304 16788
rect 4252 16745 4261 16779
rect 4261 16745 4295 16779
rect 4295 16745 4304 16779
rect 4252 16736 4304 16745
rect 4896 16736 4948 16788
rect 9680 16736 9732 16788
rect 10784 16736 10836 16788
rect 1860 16668 1912 16720
rect 1584 16643 1636 16652
rect 1584 16609 1593 16643
rect 1593 16609 1627 16643
rect 1627 16609 1636 16643
rect 1584 16600 1636 16609
rect 2228 16600 2280 16652
rect 3148 16668 3200 16720
rect 5264 16668 5316 16720
rect 7840 16668 7892 16720
rect 8668 16711 8720 16720
rect 8668 16677 8677 16711
rect 8677 16677 8711 16711
rect 8711 16677 8720 16711
rect 8668 16668 8720 16677
rect 9128 16668 9180 16720
rect 6000 16643 6052 16652
rect 6000 16609 6009 16643
rect 6009 16609 6043 16643
rect 6043 16609 6052 16643
rect 6000 16600 6052 16609
rect 6368 16600 6420 16652
rect 6552 16600 6604 16652
rect 6736 16600 6788 16652
rect 5172 16575 5224 16584
rect 5172 16541 5181 16575
rect 5181 16541 5215 16575
rect 5215 16541 5224 16575
rect 6184 16575 6236 16584
rect 5172 16532 5224 16541
rect 6184 16541 6193 16575
rect 6193 16541 6227 16575
rect 6227 16541 6236 16575
rect 6184 16532 6236 16541
rect 9220 16600 9272 16652
rect 10508 16668 10560 16720
rect 12808 16668 12860 16720
rect 8116 16532 8168 16584
rect 9588 16532 9640 16584
rect 11152 16600 11204 16652
rect 11704 16643 11756 16652
rect 3700 16464 3752 16516
rect 8024 16507 8076 16516
rect 8024 16473 8033 16507
rect 8033 16473 8067 16507
rect 8067 16473 8076 16507
rect 8024 16464 8076 16473
rect 8576 16464 8628 16516
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 12440 16643 12492 16652
rect 12440 16609 12449 16643
rect 12449 16609 12483 16643
rect 12483 16609 12492 16643
rect 12440 16600 12492 16609
rect 13728 16600 13780 16652
rect 11612 16532 11664 16584
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 11888 16532 11940 16541
rect 14004 16668 14056 16720
rect 14188 16668 14240 16720
rect 18880 16736 18932 16788
rect 21824 16736 21876 16788
rect 13912 16600 13964 16652
rect 15936 16600 15988 16652
rect 22284 16668 22336 16720
rect 16212 16600 16264 16652
rect 16856 16643 16908 16652
rect 14004 16532 14056 16584
rect 14832 16532 14884 16584
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 16396 16532 16448 16584
rect 16856 16609 16865 16643
rect 16865 16609 16899 16643
rect 16899 16609 16908 16643
rect 16856 16600 16908 16609
rect 18696 16600 18748 16652
rect 20444 16600 20496 16652
rect 20996 16600 21048 16652
rect 21180 16643 21232 16652
rect 21180 16609 21214 16643
rect 21214 16609 21232 16643
rect 21180 16600 21232 16609
rect 18144 16532 18196 16584
rect 19064 16532 19116 16584
rect 1400 16396 1452 16448
rect 6552 16396 6604 16448
rect 6644 16396 6696 16448
rect 7932 16396 7984 16448
rect 11520 16396 11572 16448
rect 12348 16396 12400 16448
rect 17776 16464 17828 16516
rect 14280 16396 14332 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 17868 16396 17920 16448
rect 22284 16439 22336 16448
rect 22284 16405 22293 16439
rect 22293 16405 22327 16439
rect 22327 16405 22336 16439
rect 22284 16396 22336 16405
rect 4614 16294 4666 16346
rect 4678 16294 4730 16346
rect 4742 16294 4794 16346
rect 4806 16294 4858 16346
rect 11878 16294 11930 16346
rect 11942 16294 11994 16346
rect 12006 16294 12058 16346
rect 12070 16294 12122 16346
rect 19142 16294 19194 16346
rect 19206 16294 19258 16346
rect 19270 16294 19322 16346
rect 19334 16294 19386 16346
rect 3148 16192 3200 16244
rect 5264 16192 5316 16244
rect 6736 16192 6788 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 7932 16192 7984 16244
rect 5724 16124 5776 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 3976 16056 4028 16108
rect 6276 16099 6328 16108
rect 6276 16065 6285 16099
rect 6285 16065 6319 16099
rect 6319 16065 6328 16099
rect 6276 16056 6328 16065
rect 6828 16056 6880 16108
rect 1676 15988 1728 16040
rect 3608 15988 3660 16040
rect 4436 15988 4488 16040
rect 5356 15988 5408 16040
rect 8668 16056 8720 16108
rect 11060 16192 11112 16244
rect 11704 16192 11756 16244
rect 12440 16192 12492 16244
rect 10416 16124 10468 16176
rect 13820 16192 13872 16244
rect 14096 16192 14148 16244
rect 16856 16192 16908 16244
rect 18236 16192 18288 16244
rect 20444 16192 20496 16244
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 3056 15920 3108 15972
rect 3700 15920 3752 15972
rect 6184 15920 6236 15972
rect 6920 15920 6972 15972
rect 10784 15988 10836 16040
rect 3884 15852 3936 15904
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 4804 15852 4856 15904
rect 5264 15852 5316 15904
rect 6368 15852 6420 15904
rect 7196 15895 7248 15904
rect 7196 15861 7205 15895
rect 7205 15861 7239 15895
rect 7239 15861 7248 15895
rect 7196 15852 7248 15861
rect 8852 15895 8904 15904
rect 8852 15861 8861 15895
rect 8861 15861 8895 15895
rect 8895 15861 8904 15895
rect 8852 15852 8904 15861
rect 9772 15920 9824 15972
rect 12440 15988 12492 16040
rect 13912 15988 13964 16040
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 11520 15852 11572 15904
rect 13544 15920 13596 15972
rect 16120 16056 16172 16108
rect 20996 16192 21048 16244
rect 15016 16031 15068 16040
rect 15016 15997 15025 16031
rect 15025 15997 15059 16031
rect 15059 15997 15068 16031
rect 15016 15988 15068 15997
rect 14280 15852 14332 15904
rect 15016 15852 15068 15904
rect 16304 15988 16356 16040
rect 16120 15920 16172 15972
rect 16488 15920 16540 15972
rect 18236 15988 18288 16040
rect 20260 16031 20312 16040
rect 16580 15895 16632 15904
rect 16580 15861 16589 15895
rect 16589 15861 16623 15895
rect 16623 15861 16632 15895
rect 16580 15852 16632 15861
rect 17316 15895 17368 15904
rect 17316 15861 17325 15895
rect 17325 15861 17359 15895
rect 17359 15861 17368 15895
rect 17316 15852 17368 15861
rect 18052 15852 18104 15904
rect 18512 15852 18564 15904
rect 19432 15920 19484 15972
rect 20260 15997 20269 16031
rect 20269 15997 20303 16031
rect 20303 15997 20312 16031
rect 20260 15988 20312 15997
rect 22284 15988 22336 16040
rect 19892 15852 19944 15904
rect 19984 15852 20036 15904
rect 20260 15852 20312 15904
rect 21364 15920 21416 15972
rect 21548 15852 21600 15904
rect 8246 15750 8298 15802
rect 8310 15750 8362 15802
rect 8374 15750 8426 15802
rect 8438 15750 8490 15802
rect 15510 15750 15562 15802
rect 15574 15750 15626 15802
rect 15638 15750 15690 15802
rect 15702 15750 15754 15802
rect 3056 15691 3108 15700
rect 3056 15657 3065 15691
rect 3065 15657 3099 15691
rect 3099 15657 3108 15691
rect 3056 15648 3108 15657
rect 4160 15648 4212 15700
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 6828 15691 6880 15700
rect 6828 15657 6837 15691
rect 6837 15657 6871 15691
rect 6871 15657 6880 15691
rect 6828 15648 6880 15657
rect 1676 15555 1728 15564
rect 1676 15521 1685 15555
rect 1685 15521 1719 15555
rect 1719 15521 1728 15555
rect 1676 15512 1728 15521
rect 1952 15555 2004 15564
rect 1952 15521 1986 15555
rect 1986 15521 2004 15555
rect 1952 15512 2004 15521
rect 3516 15512 3568 15564
rect 4804 15555 4856 15564
rect 4804 15521 4813 15555
rect 4813 15521 4847 15555
rect 4847 15521 4856 15555
rect 4804 15512 4856 15521
rect 3976 15308 4028 15360
rect 8300 15512 8352 15564
rect 7104 15444 7156 15496
rect 8484 15580 8536 15632
rect 10416 15648 10468 15700
rect 11152 15648 11204 15700
rect 13912 15691 13964 15700
rect 13912 15657 13921 15691
rect 13921 15657 13955 15691
rect 13955 15657 13964 15691
rect 13912 15648 13964 15657
rect 18328 15648 18380 15700
rect 20720 15648 20772 15700
rect 21180 15648 21232 15700
rect 11060 15580 11112 15632
rect 14004 15580 14056 15632
rect 16488 15580 16540 15632
rect 22284 15580 22336 15632
rect 10232 15512 10284 15564
rect 11704 15555 11756 15564
rect 11704 15521 11713 15555
rect 11713 15521 11747 15555
rect 11747 15521 11756 15555
rect 11704 15512 11756 15521
rect 13912 15512 13964 15564
rect 14372 15512 14424 15564
rect 15200 15512 15252 15564
rect 15568 15555 15620 15564
rect 15568 15521 15602 15555
rect 15602 15521 15620 15555
rect 15568 15512 15620 15521
rect 17224 15512 17276 15564
rect 17684 15512 17736 15564
rect 19432 15512 19484 15564
rect 21364 15512 21416 15564
rect 21916 15555 21968 15564
rect 21916 15521 21925 15555
rect 21925 15521 21959 15555
rect 21959 15521 21968 15555
rect 21916 15512 21968 15521
rect 8668 15308 8720 15360
rect 9864 15308 9916 15360
rect 10784 15308 10836 15360
rect 11612 15376 11664 15428
rect 12440 15444 12492 15496
rect 14924 15444 14976 15496
rect 18512 15444 18564 15496
rect 18972 15444 19024 15496
rect 15016 15376 15068 15428
rect 16948 15376 17000 15428
rect 19984 15444 20036 15496
rect 20996 15444 21048 15496
rect 21180 15444 21232 15496
rect 16856 15308 16908 15360
rect 17316 15308 17368 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 20720 15376 20772 15428
rect 20812 15308 20864 15360
rect 21180 15308 21232 15360
rect 4614 15206 4666 15258
rect 4678 15206 4730 15258
rect 4742 15206 4794 15258
rect 4806 15206 4858 15258
rect 11878 15206 11930 15258
rect 11942 15206 11994 15258
rect 12006 15206 12058 15258
rect 12070 15206 12122 15258
rect 19142 15206 19194 15258
rect 19206 15206 19258 15258
rect 19270 15206 19322 15258
rect 19334 15206 19386 15258
rect 3700 15104 3752 15156
rect 4988 15104 5040 15156
rect 6920 15104 6972 15156
rect 8300 15104 8352 15156
rect 11060 15104 11112 15156
rect 11704 15104 11756 15156
rect 12348 15104 12400 15156
rect 14004 15104 14056 15156
rect 14188 15147 14240 15156
rect 14188 15113 14197 15147
rect 14197 15113 14231 15147
rect 14231 15113 14240 15147
rect 14188 15104 14240 15113
rect 15384 15104 15436 15156
rect 15568 15104 15620 15156
rect 15936 15104 15988 15156
rect 17684 15147 17736 15156
rect 3792 15036 3844 15088
rect 17684 15113 17693 15147
rect 17693 15113 17727 15147
rect 17727 15113 17736 15147
rect 17684 15104 17736 15113
rect 17960 15036 18012 15088
rect 3608 14968 3660 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 1584 14900 1636 14952
rect 4160 14900 4212 14952
rect 4436 14900 4488 14952
rect 6368 14900 6420 14952
rect 10324 14968 10376 15020
rect 2044 14832 2096 14884
rect 4068 14832 4120 14884
rect 6828 14832 6880 14884
rect 9404 14832 9456 14884
rect 10784 14900 10836 14952
rect 11704 14900 11756 14952
rect 12440 14943 12492 14952
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12716 14943 12768 14952
rect 12440 14900 12492 14909
rect 12716 14909 12750 14943
rect 12750 14909 12768 14943
rect 12716 14900 12768 14909
rect 9772 14832 9824 14884
rect 15752 14968 15804 15020
rect 17316 14968 17368 15020
rect 18236 15104 18288 15156
rect 19432 15147 19484 15156
rect 19432 15113 19441 15147
rect 19441 15113 19475 15147
rect 19475 15113 19484 15147
rect 19432 15104 19484 15113
rect 19708 15104 19760 15156
rect 20352 15011 20404 15020
rect 20352 14977 20361 15011
rect 20361 14977 20395 15011
rect 20395 14977 20404 15011
rect 20352 14968 20404 14977
rect 20720 15104 20772 15156
rect 21088 15104 21140 15156
rect 15016 14900 15068 14952
rect 14188 14832 14240 14884
rect 17132 14900 17184 14952
rect 17408 14900 17460 14952
rect 18328 14943 18380 14952
rect 17316 14832 17368 14884
rect 18328 14909 18362 14943
rect 18362 14909 18380 14943
rect 18328 14900 18380 14909
rect 18880 14900 18932 14952
rect 20720 14900 20772 14952
rect 21548 14900 21600 14952
rect 1952 14764 2004 14816
rect 3700 14807 3752 14816
rect 3700 14773 3709 14807
rect 3709 14773 3743 14807
rect 3743 14773 3752 14807
rect 3700 14764 3752 14773
rect 4252 14764 4304 14816
rect 4344 14764 4396 14816
rect 7472 14764 7524 14816
rect 8116 14764 8168 14816
rect 11152 14764 11204 14816
rect 11612 14764 11664 14816
rect 12164 14764 12216 14816
rect 15384 14764 15436 14816
rect 16488 14764 16540 14816
rect 19064 14764 19116 14816
rect 19892 14807 19944 14816
rect 19892 14773 19901 14807
rect 19901 14773 19935 14807
rect 19935 14773 19944 14807
rect 19892 14764 19944 14773
rect 8246 14662 8298 14714
rect 8310 14662 8362 14714
rect 8374 14662 8426 14714
rect 8438 14662 8490 14714
rect 15510 14662 15562 14714
rect 15574 14662 15626 14714
rect 15638 14662 15690 14714
rect 15702 14662 15754 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2688 14560 2740 14612
rect 3240 14560 3292 14612
rect 3608 14560 3660 14612
rect 4068 14560 4120 14612
rect 3700 14492 3752 14544
rect 4436 14492 4488 14544
rect 2964 14467 3016 14476
rect 2964 14433 2973 14467
rect 2973 14433 3007 14467
rect 3007 14433 3016 14467
rect 2964 14424 3016 14433
rect 6092 14560 6144 14612
rect 7196 14560 7248 14612
rect 7472 14560 7524 14612
rect 12624 14560 12676 14612
rect 11060 14492 11112 14544
rect 11336 14492 11388 14544
rect 12808 14560 12860 14612
rect 17408 14560 17460 14612
rect 14004 14492 14056 14544
rect 15108 14492 15160 14544
rect 17316 14492 17368 14544
rect 18052 14603 18104 14612
rect 18052 14569 18061 14603
rect 18061 14569 18095 14603
rect 18095 14569 18104 14603
rect 18052 14560 18104 14569
rect 18144 14560 18196 14612
rect 18512 14560 18564 14612
rect 19064 14603 19116 14612
rect 19064 14569 19073 14603
rect 19073 14569 19107 14603
rect 19107 14569 19116 14603
rect 19064 14560 19116 14569
rect 20812 14560 20864 14612
rect 21456 14560 21508 14612
rect 17684 14492 17736 14544
rect 18972 14492 19024 14544
rect 2044 14399 2096 14408
rect 2044 14365 2053 14399
rect 2053 14365 2087 14399
rect 2087 14365 2096 14399
rect 2044 14356 2096 14365
rect 2688 14356 2740 14408
rect 3056 14399 3108 14408
rect 3056 14365 3065 14399
rect 3065 14365 3099 14399
rect 3099 14365 3108 14399
rect 3056 14356 3108 14365
rect 3240 14399 3292 14408
rect 3240 14365 3249 14399
rect 3249 14365 3283 14399
rect 3283 14365 3292 14399
rect 3240 14356 3292 14365
rect 3700 14356 3752 14408
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 7472 14424 7524 14476
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 8760 14424 8812 14476
rect 9404 14467 9456 14476
rect 9404 14433 9413 14467
rect 9413 14433 9447 14467
rect 9447 14433 9456 14467
rect 9404 14424 9456 14433
rect 9772 14424 9824 14476
rect 14648 14467 14700 14476
rect 7104 14399 7156 14408
rect 7104 14365 7113 14399
rect 7113 14365 7147 14399
rect 7147 14365 7156 14399
rect 7104 14356 7156 14365
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 7564 14356 7616 14408
rect 8208 14399 8260 14408
rect 8208 14365 8217 14399
rect 8217 14365 8251 14399
rect 8251 14365 8260 14399
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 15936 14424 15988 14476
rect 16488 14424 16540 14476
rect 8208 14356 8260 14365
rect 12440 14356 12492 14408
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 9220 14331 9272 14340
rect 2320 14220 2372 14272
rect 3424 14220 3476 14272
rect 3700 14263 3752 14272
rect 3700 14229 3709 14263
rect 3709 14229 3743 14263
rect 3743 14229 3752 14263
rect 3700 14220 3752 14229
rect 9220 14297 9229 14331
rect 9229 14297 9263 14331
rect 9263 14297 9272 14331
rect 9220 14288 9272 14297
rect 5080 14220 5132 14272
rect 6276 14263 6328 14272
rect 6276 14229 6285 14263
rect 6285 14229 6319 14263
rect 6319 14229 6328 14263
rect 6276 14220 6328 14229
rect 7288 14220 7340 14272
rect 7748 14220 7800 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 11520 14220 11572 14272
rect 15936 14288 15988 14340
rect 13176 14220 13228 14272
rect 16120 14220 16172 14272
rect 18972 14356 19024 14408
rect 19524 14399 19576 14408
rect 19524 14365 19533 14399
rect 19533 14365 19567 14399
rect 19567 14365 19576 14399
rect 19524 14356 19576 14365
rect 20352 14492 20404 14544
rect 20536 14492 20588 14544
rect 21088 14492 21140 14544
rect 20260 14467 20312 14476
rect 20260 14433 20269 14467
rect 20269 14433 20303 14467
rect 20303 14433 20312 14467
rect 20260 14424 20312 14433
rect 20720 14424 20772 14476
rect 17960 14220 18012 14272
rect 19708 14220 19760 14272
rect 4614 14118 4666 14170
rect 4678 14118 4730 14170
rect 4742 14118 4794 14170
rect 4806 14118 4858 14170
rect 11878 14118 11930 14170
rect 11942 14118 11994 14170
rect 12006 14118 12058 14170
rect 12070 14118 12122 14170
rect 19142 14118 19194 14170
rect 19206 14118 19258 14170
rect 19270 14118 19322 14170
rect 19334 14118 19386 14170
rect 3608 14016 3660 14068
rect 4160 14016 4212 14068
rect 4436 14016 4488 14068
rect 5080 14016 5132 14068
rect 6828 14016 6880 14068
rect 9772 14016 9824 14068
rect 11336 14016 11388 14068
rect 13084 14016 13136 14068
rect 13176 14016 13228 14068
rect 3240 13948 3292 14000
rect 2688 13880 2740 13932
rect 5908 13948 5960 14000
rect 6368 13948 6420 14000
rect 7012 13948 7064 14000
rect 6276 13880 6328 13932
rect 7564 13880 7616 13932
rect 12900 13948 12952 14000
rect 10968 13880 11020 13932
rect 2136 13744 2188 13796
rect 2780 13676 2832 13728
rect 3240 13855 3292 13864
rect 3240 13821 3249 13855
rect 3249 13821 3283 13855
rect 3283 13821 3292 13855
rect 3240 13812 3292 13821
rect 4252 13812 4304 13864
rect 4988 13812 5040 13864
rect 4896 13744 4948 13796
rect 6552 13812 6604 13864
rect 7748 13812 7800 13864
rect 9680 13855 9732 13864
rect 9680 13821 9689 13855
rect 9689 13821 9723 13855
rect 9723 13821 9732 13855
rect 9680 13812 9732 13821
rect 11060 13812 11112 13864
rect 11428 13812 11480 13864
rect 12992 13812 13044 13864
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 13728 13812 13780 13864
rect 15200 14016 15252 14068
rect 18972 14016 19024 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 20720 14016 20772 14068
rect 21732 14016 21784 14068
rect 15108 13855 15160 13864
rect 15108 13821 15142 13855
rect 15142 13821 15160 13855
rect 15108 13812 15160 13821
rect 16488 13812 16540 13864
rect 17224 13812 17276 13864
rect 17960 13812 18012 13864
rect 19524 13812 19576 13864
rect 20076 13948 20128 14000
rect 21180 13812 21232 13864
rect 6920 13744 6972 13796
rect 7932 13744 7984 13796
rect 8852 13744 8904 13796
rect 12532 13744 12584 13796
rect 18236 13744 18288 13796
rect 20812 13787 20864 13796
rect 20812 13753 20846 13787
rect 20846 13753 20864 13787
rect 20812 13744 20864 13753
rect 3240 13676 3292 13728
rect 4436 13676 4488 13728
rect 5356 13676 5408 13728
rect 7012 13676 7064 13728
rect 8760 13676 8812 13728
rect 11796 13676 11848 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16488 13719 16540 13728
rect 16488 13685 16497 13719
rect 16497 13685 16531 13719
rect 16531 13685 16540 13719
rect 16488 13676 16540 13685
rect 17684 13676 17736 13728
rect 8246 13574 8298 13626
rect 8310 13574 8362 13626
rect 8374 13574 8426 13626
rect 8438 13574 8490 13626
rect 15510 13574 15562 13626
rect 15574 13574 15626 13626
rect 15638 13574 15690 13626
rect 15702 13574 15754 13626
rect 1860 13472 1912 13524
rect 2688 13472 2740 13524
rect 2964 13472 3016 13524
rect 3608 13472 3660 13524
rect 4252 13472 4304 13524
rect 4528 13472 4580 13524
rect 6920 13472 6972 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 7932 13472 7984 13524
rect 10968 13472 11020 13524
rect 11152 13515 11204 13524
rect 11152 13481 11161 13515
rect 11161 13481 11195 13515
rect 11195 13481 11204 13515
rect 11152 13472 11204 13481
rect 3056 13404 3108 13456
rect 1768 13336 1820 13388
rect 9312 13404 9364 13456
rect 13728 13472 13780 13524
rect 16580 13472 16632 13524
rect 16948 13472 17000 13524
rect 17408 13472 17460 13524
rect 17684 13515 17736 13524
rect 17684 13481 17693 13515
rect 17693 13481 17727 13515
rect 17727 13481 17736 13515
rect 17684 13472 17736 13481
rect 18052 13472 18104 13524
rect 19248 13472 19300 13524
rect 19524 13472 19576 13524
rect 19800 13472 19852 13524
rect 14372 13404 14424 13456
rect 16488 13404 16540 13456
rect 21732 13404 21784 13456
rect 6828 13336 6880 13388
rect 7288 13379 7340 13388
rect 7288 13345 7297 13379
rect 7297 13345 7331 13379
rect 7331 13345 7340 13379
rect 7288 13336 7340 13345
rect 7932 13336 7984 13388
rect 11796 13379 11848 13388
rect 11796 13345 11805 13379
rect 11805 13345 11839 13379
rect 11839 13345 11848 13379
rect 11796 13336 11848 13345
rect 1676 13268 1728 13320
rect 4252 13268 4304 13320
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5172 13268 5224 13320
rect 7748 13268 7800 13320
rect 9772 13268 9824 13320
rect 10324 13311 10376 13320
rect 10324 13277 10333 13311
rect 10333 13277 10367 13311
rect 10367 13277 10376 13311
rect 10324 13268 10376 13277
rect 10416 13268 10468 13320
rect 12348 13268 12400 13320
rect 12624 13268 12676 13320
rect 13176 13268 13228 13320
rect 7104 13200 7156 13252
rect 7288 13200 7340 13252
rect 9680 13200 9732 13252
rect 12716 13200 12768 13252
rect 1768 13175 1820 13184
rect 1768 13141 1777 13175
rect 1777 13141 1811 13175
rect 1811 13141 1820 13175
rect 1768 13132 1820 13141
rect 5356 13132 5408 13184
rect 10692 13132 10744 13184
rect 11428 13132 11480 13184
rect 11704 13132 11756 13184
rect 15292 13175 15344 13184
rect 15292 13141 15301 13175
rect 15301 13141 15335 13175
rect 15335 13141 15344 13175
rect 15292 13132 15344 13141
rect 15752 13336 15804 13388
rect 17316 13336 17368 13388
rect 18236 13379 18288 13388
rect 18236 13345 18270 13379
rect 18270 13345 18288 13379
rect 18236 13336 18288 13345
rect 19432 13336 19484 13388
rect 20720 13336 20772 13388
rect 20904 13379 20956 13388
rect 20904 13345 20913 13379
rect 20913 13345 20947 13379
rect 20947 13345 20956 13379
rect 20904 13336 20956 13345
rect 16212 13268 16264 13320
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 18236 13132 18288 13184
rect 20812 13132 20864 13184
rect 21180 13132 21232 13184
rect 4614 13030 4666 13082
rect 4678 13030 4730 13082
rect 4742 13030 4794 13082
rect 4806 13030 4858 13082
rect 11878 13030 11930 13082
rect 11942 13030 11994 13082
rect 12006 13030 12058 13082
rect 12070 13030 12122 13082
rect 19142 13030 19194 13082
rect 19206 13030 19258 13082
rect 19270 13030 19322 13082
rect 19334 13030 19386 13082
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 4252 12928 4304 12980
rect 5264 12928 5316 12980
rect 5724 12928 5776 12980
rect 7012 12971 7064 12980
rect 7012 12937 7021 12971
rect 7021 12937 7055 12971
rect 7055 12937 7064 12971
rect 7012 12928 7064 12937
rect 7932 12928 7984 12980
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 11888 12860 11940 12912
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 9680 12835 9732 12844
rect 9680 12801 9689 12835
rect 9689 12801 9723 12835
rect 9723 12801 9732 12835
rect 9680 12792 9732 12801
rect 9772 12835 9824 12844
rect 9772 12801 9781 12835
rect 9781 12801 9815 12835
rect 9815 12801 9824 12835
rect 9772 12792 9824 12801
rect 11060 12792 11112 12844
rect 12716 12928 12768 12980
rect 3608 12767 3660 12776
rect 3608 12733 3642 12767
rect 3642 12733 3660 12767
rect 2780 12656 2832 12708
rect 3608 12724 3660 12733
rect 5172 12724 5224 12776
rect 5356 12767 5408 12776
rect 5356 12733 5390 12767
rect 5390 12733 5408 12767
rect 5356 12724 5408 12733
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7564 12724 7616 12776
rect 4068 12656 4120 12708
rect 8760 12724 8812 12776
rect 9128 12724 9180 12776
rect 9864 12724 9916 12776
rect 10600 12724 10652 12776
rect 10692 12724 10744 12776
rect 12348 12792 12400 12844
rect 14924 12792 14976 12844
rect 8024 12699 8076 12708
rect 8024 12665 8058 12699
rect 8058 12665 8076 12699
rect 8024 12656 8076 12665
rect 4988 12588 5040 12640
rect 11336 12656 11388 12708
rect 12532 12724 12584 12776
rect 16764 12903 16816 12912
rect 16764 12869 16773 12903
rect 16773 12869 16807 12903
rect 16807 12869 16816 12903
rect 16764 12860 16816 12869
rect 16580 12792 16632 12844
rect 17316 12860 17368 12912
rect 17500 12928 17552 12980
rect 19432 12971 19484 12980
rect 19432 12937 19441 12971
rect 19441 12937 19475 12971
rect 19475 12937 19484 12971
rect 19432 12928 19484 12937
rect 19708 12928 19760 12980
rect 19892 12928 19944 12980
rect 21088 12928 21140 12980
rect 18052 12860 18104 12912
rect 15476 12724 15528 12776
rect 16212 12724 16264 12776
rect 17868 12792 17920 12844
rect 20720 12792 20772 12844
rect 20904 12835 20956 12844
rect 20904 12801 20913 12835
rect 20913 12801 20947 12835
rect 20947 12801 20956 12835
rect 20904 12792 20956 12801
rect 17408 12767 17460 12776
rect 17408 12733 17417 12767
rect 17417 12733 17451 12767
rect 17451 12733 17460 12767
rect 17408 12724 17460 12733
rect 17960 12724 18012 12776
rect 21180 12767 21232 12776
rect 21180 12733 21214 12767
rect 21214 12733 21232 12767
rect 21180 12724 21232 12733
rect 12164 12656 12216 12708
rect 11060 12588 11112 12640
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 15016 12656 15068 12708
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 14280 12588 14332 12597
rect 14924 12631 14976 12640
rect 14924 12597 14933 12631
rect 14933 12597 14967 12631
rect 14967 12597 14976 12631
rect 14924 12588 14976 12597
rect 15844 12588 15896 12640
rect 16212 12588 16264 12640
rect 17316 12588 17368 12640
rect 17684 12656 17736 12708
rect 20812 12656 20864 12708
rect 21640 12656 21692 12708
rect 19340 12588 19392 12640
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 20352 12631 20404 12640
rect 20352 12597 20361 12631
rect 20361 12597 20395 12631
rect 20395 12597 20404 12631
rect 20352 12588 20404 12597
rect 8246 12486 8298 12538
rect 8310 12486 8362 12538
rect 8374 12486 8426 12538
rect 8438 12486 8490 12538
rect 15510 12486 15562 12538
rect 15574 12486 15626 12538
rect 15638 12486 15690 12538
rect 15702 12486 15754 12538
rect 1584 12384 1636 12436
rect 2136 12384 2188 12436
rect 2964 12384 3016 12436
rect 4160 12384 4212 12436
rect 5264 12384 5316 12436
rect 6092 12384 6144 12436
rect 10416 12384 10468 12436
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 1492 12248 1544 12300
rect 3056 12248 3108 12300
rect 1400 12223 1452 12232
rect 1400 12189 1409 12223
rect 1409 12189 1443 12223
rect 1443 12189 1452 12223
rect 1400 12180 1452 12189
rect 4344 12248 4396 12300
rect 8852 12316 8904 12368
rect 4988 12291 5040 12300
rect 4988 12257 5022 12291
rect 5022 12257 5040 12291
rect 4988 12248 5040 12257
rect 5540 12248 5592 12300
rect 14372 12427 14424 12436
rect 14372 12393 14381 12427
rect 14381 12393 14415 12427
rect 14415 12393 14424 12427
rect 14372 12384 14424 12393
rect 16304 12384 16356 12436
rect 16396 12384 16448 12436
rect 18788 12384 18840 12436
rect 19340 12384 19392 12436
rect 11060 12316 11112 12368
rect 13820 12316 13872 12368
rect 15108 12316 15160 12368
rect 1400 12044 1452 12096
rect 4344 12112 4396 12164
rect 5724 12180 5776 12232
rect 5816 12112 5868 12164
rect 7196 12180 7248 12232
rect 7472 12180 7524 12232
rect 8116 12223 8168 12232
rect 8116 12189 8125 12223
rect 8125 12189 8159 12223
rect 8159 12189 8168 12223
rect 8116 12180 8168 12189
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9404 12180 9456 12232
rect 17132 12316 17184 12368
rect 17224 12316 17276 12368
rect 19616 12316 19668 12368
rect 19892 12384 19944 12436
rect 20444 12384 20496 12436
rect 21088 12316 21140 12368
rect 15660 12291 15712 12300
rect 10140 12180 10192 12232
rect 10232 12180 10284 12232
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 16212 12291 16264 12300
rect 16212 12257 16221 12291
rect 16221 12257 16255 12291
rect 16255 12257 16264 12291
rect 16212 12248 16264 12257
rect 16304 12248 16356 12300
rect 16764 12248 16816 12300
rect 17316 12248 17368 12300
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 18052 12248 18104 12300
rect 18788 12248 18840 12300
rect 12532 12180 12584 12232
rect 14648 12180 14700 12232
rect 15200 12180 15252 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15936 12223 15988 12232
rect 15752 12180 15804 12189
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 9312 12112 9364 12164
rect 19892 12248 19944 12300
rect 20076 12248 20128 12300
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 20812 12180 20864 12232
rect 6000 12044 6052 12096
rect 7104 12044 7156 12096
rect 8576 12044 8628 12096
rect 15660 12044 15712 12096
rect 16856 12044 16908 12096
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 17592 12044 17644 12053
rect 20536 12044 20588 12096
rect 4614 11942 4666 11994
rect 4678 11942 4730 11994
rect 4742 11942 4794 11994
rect 4806 11942 4858 11994
rect 11878 11942 11930 11994
rect 11942 11942 11994 11994
rect 12006 11942 12058 11994
rect 12070 11942 12122 11994
rect 19142 11942 19194 11994
rect 19206 11942 19258 11994
rect 19270 11942 19322 11994
rect 19334 11942 19386 11994
rect 2780 11883 2832 11892
rect 2780 11849 2789 11883
rect 2789 11849 2823 11883
rect 2823 11849 2832 11883
rect 2780 11840 2832 11849
rect 3240 11840 3292 11892
rect 4160 11840 4212 11892
rect 5816 11840 5868 11892
rect 6184 11840 6236 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 4344 11772 4396 11824
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 3332 11704 3384 11756
rect 4068 11704 4120 11756
rect 4436 11704 4488 11756
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 5816 11704 5868 11756
rect 8024 11840 8076 11892
rect 11336 11840 11388 11892
rect 13820 11883 13872 11892
rect 12440 11772 12492 11824
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 9680 11704 9732 11756
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 11428 11704 11480 11756
rect 2136 11636 2188 11688
rect 3424 11679 3476 11688
rect 3424 11645 3433 11679
rect 3433 11645 3467 11679
rect 3467 11645 3476 11679
rect 3424 11636 3476 11645
rect 4252 11636 4304 11688
rect 7104 11679 7156 11688
rect 1860 11568 1912 11620
rect 4804 11568 4856 11620
rect 5632 11568 5684 11620
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 9128 11636 9180 11688
rect 9772 11636 9824 11688
rect 11704 11679 11756 11688
rect 11704 11645 11713 11679
rect 11713 11645 11747 11679
rect 11747 11645 11756 11679
rect 11704 11636 11756 11645
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12440 11636 12492 11645
rect 12716 11679 12768 11688
rect 12716 11645 12750 11679
rect 12750 11645 12768 11679
rect 12716 11636 12768 11645
rect 4896 11500 4948 11552
rect 5172 11500 5224 11552
rect 5908 11500 5960 11552
rect 7840 11568 7892 11620
rect 10140 11611 10192 11620
rect 10140 11577 10174 11611
rect 10174 11577 10192 11611
rect 10140 11568 10192 11577
rect 11060 11568 11112 11620
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14280 11840 14332 11892
rect 15384 11840 15436 11892
rect 18420 11840 18472 11892
rect 19984 11883 20036 11892
rect 19984 11849 19993 11883
rect 19993 11849 20027 11883
rect 20027 11849 20036 11883
rect 19984 11840 20036 11849
rect 20720 11840 20772 11892
rect 15016 11772 15068 11824
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 15476 11704 15528 11756
rect 16764 11772 16816 11824
rect 21364 11772 21416 11824
rect 17592 11747 17644 11756
rect 13728 11636 13780 11688
rect 14464 11636 14516 11688
rect 15016 11636 15068 11688
rect 8024 11500 8076 11552
rect 14924 11568 14976 11620
rect 12440 11500 12492 11552
rect 15752 11568 15804 11620
rect 15384 11500 15436 11552
rect 15844 11500 15896 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 17592 11713 17601 11747
rect 17601 11713 17635 11747
rect 17635 11713 17644 11747
rect 17592 11704 17644 11713
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 19800 11679 19852 11688
rect 17776 11568 17828 11620
rect 19800 11645 19809 11679
rect 19809 11645 19843 11679
rect 19843 11645 19852 11679
rect 19800 11636 19852 11645
rect 19892 11636 19944 11688
rect 20444 11636 20496 11688
rect 18512 11568 18564 11620
rect 16488 11500 16540 11552
rect 16580 11500 16632 11552
rect 16948 11543 17000 11552
rect 16948 11509 16957 11543
rect 16957 11509 16991 11543
rect 16991 11509 17000 11543
rect 16948 11500 17000 11509
rect 17316 11500 17368 11552
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 18052 11500 18104 11552
rect 8246 11398 8298 11450
rect 8310 11398 8362 11450
rect 8374 11398 8426 11450
rect 8438 11398 8490 11450
rect 15510 11398 15562 11450
rect 15574 11398 15626 11450
rect 15638 11398 15690 11450
rect 15702 11398 15754 11450
rect 1584 11296 1636 11348
rect 1860 11339 1912 11348
rect 1860 11305 1869 11339
rect 1869 11305 1903 11339
rect 1903 11305 1912 11339
rect 1860 11296 1912 11305
rect 2688 11296 2740 11348
rect 2872 11296 2924 11348
rect 5172 11296 5224 11348
rect 5264 11296 5316 11348
rect 6828 11296 6880 11348
rect 8576 11296 8628 11348
rect 9312 11296 9364 11348
rect 11060 11339 11112 11348
rect 2320 11160 2372 11212
rect 7380 11228 7432 11280
rect 8208 11228 8260 11280
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 4344 11203 4396 11212
rect 4344 11169 4353 11203
rect 4353 11169 4387 11203
rect 4387 11169 4396 11203
rect 4344 11160 4396 11169
rect 4712 11160 4764 11212
rect 2688 11092 2740 11144
rect 4436 11092 4488 11144
rect 3424 11024 3476 11076
rect 4160 11024 4212 11076
rect 5908 11160 5960 11212
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 7104 11160 7156 11212
rect 7656 11160 7708 11212
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 9680 11203 9732 11212
rect 9680 11169 9689 11203
rect 9689 11169 9723 11203
rect 9723 11169 9732 11203
rect 12532 11228 12584 11280
rect 14004 11296 14056 11348
rect 14188 11296 14240 11348
rect 16580 11296 16632 11348
rect 16948 11296 17000 11348
rect 19892 11339 19944 11348
rect 9680 11160 9732 11169
rect 10692 11160 10744 11212
rect 11428 11160 11480 11212
rect 11612 11203 11664 11212
rect 11612 11169 11646 11203
rect 11646 11169 11664 11203
rect 11612 11160 11664 11169
rect 12348 11160 12400 11212
rect 13728 11160 13780 11212
rect 14004 11160 14056 11212
rect 12992 11135 13044 11144
rect 6184 11024 6236 11076
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 18144 11228 18196 11280
rect 18696 11228 18748 11280
rect 19892 11305 19901 11339
rect 19901 11305 19935 11339
rect 19935 11305 19944 11339
rect 19892 11296 19944 11305
rect 19708 11228 19760 11280
rect 15108 11160 15160 11212
rect 15384 11135 15436 11144
rect 15384 11101 15393 11135
rect 15393 11101 15427 11135
rect 15427 11101 15436 11135
rect 15384 11092 15436 11101
rect 14648 11067 14700 11076
rect 5080 10956 5132 11008
rect 5172 10956 5224 11008
rect 9220 10956 9272 11008
rect 11244 10956 11296 11008
rect 11336 10956 11388 11008
rect 14004 10956 14056 11008
rect 14096 10956 14148 11008
rect 14648 11033 14657 11067
rect 14657 11033 14691 11067
rect 14691 11033 14700 11067
rect 14648 11024 14700 11033
rect 14924 11024 14976 11076
rect 16672 11160 16724 11212
rect 17776 11160 17828 11212
rect 18052 11092 18104 11144
rect 18788 11160 18840 11212
rect 19800 11160 19852 11212
rect 20812 11296 20864 11348
rect 20720 11228 20772 11280
rect 20904 11203 20956 11212
rect 20904 11169 20913 11203
rect 20913 11169 20947 11203
rect 20947 11169 20956 11203
rect 20904 11160 20956 11169
rect 14556 10956 14608 11008
rect 15108 10956 15160 11008
rect 16488 11024 16540 11076
rect 16856 10956 16908 11008
rect 17316 10956 17368 11008
rect 17776 10956 17828 11008
rect 19432 10956 19484 11008
rect 19616 10999 19668 11008
rect 19616 10965 19625 10999
rect 19625 10965 19659 10999
rect 19659 10965 19668 10999
rect 19616 10956 19668 10965
rect 19708 10956 19760 11008
rect 4614 10854 4666 10906
rect 4678 10854 4730 10906
rect 4742 10854 4794 10906
rect 4806 10854 4858 10906
rect 11878 10854 11930 10906
rect 11942 10854 11994 10906
rect 12006 10854 12058 10906
rect 12070 10854 12122 10906
rect 19142 10854 19194 10906
rect 19206 10854 19258 10906
rect 19270 10854 19322 10906
rect 19334 10854 19386 10906
rect 2412 10752 2464 10804
rect 3516 10752 3568 10804
rect 7196 10752 7248 10804
rect 8116 10752 8168 10804
rect 8208 10752 8260 10804
rect 9772 10752 9824 10804
rect 12440 10752 12492 10804
rect 10232 10684 10284 10736
rect 2872 10616 2924 10668
rect 3148 10659 3200 10668
rect 3148 10625 3157 10659
rect 3157 10625 3191 10659
rect 3191 10625 3200 10659
rect 3148 10616 3200 10625
rect 3792 10616 3844 10668
rect 4436 10616 4488 10668
rect 1768 10548 1820 10600
rect 2964 10548 3016 10600
rect 3700 10548 3752 10600
rect 3884 10548 3936 10600
rect 2596 10480 2648 10532
rect 5080 10591 5132 10600
rect 5080 10557 5089 10591
rect 5089 10557 5123 10591
rect 5123 10557 5132 10591
rect 5080 10548 5132 10557
rect 10324 10616 10376 10668
rect 10784 10616 10836 10668
rect 12348 10616 12400 10668
rect 5172 10480 5224 10532
rect 5264 10480 5316 10532
rect 5816 10548 5868 10600
rect 6092 10548 6144 10600
rect 7012 10548 7064 10600
rect 7564 10548 7616 10600
rect 9772 10548 9824 10600
rect 9864 10548 9916 10600
rect 11336 10548 11388 10600
rect 12164 10591 12216 10600
rect 12164 10557 12173 10591
rect 12173 10557 12207 10591
rect 12207 10557 12216 10591
rect 12164 10548 12216 10557
rect 12992 10591 13044 10600
rect 12992 10557 13001 10591
rect 13001 10557 13035 10591
rect 13035 10557 13044 10591
rect 15108 10684 15160 10736
rect 17408 10727 17460 10736
rect 14832 10616 14884 10668
rect 17408 10693 17417 10727
rect 17417 10693 17451 10727
rect 17451 10693 17460 10727
rect 17408 10684 17460 10693
rect 12992 10548 13044 10557
rect 2412 10412 2464 10464
rect 3976 10412 4028 10464
rect 4436 10455 4488 10464
rect 4436 10421 4445 10455
rect 4445 10421 4479 10455
rect 4479 10421 4488 10455
rect 4436 10412 4488 10421
rect 5080 10412 5132 10464
rect 5448 10412 5500 10464
rect 5632 10412 5684 10464
rect 6828 10412 6880 10464
rect 8024 10480 8076 10532
rect 9220 10480 9272 10532
rect 15292 10548 15344 10600
rect 15844 10616 15896 10668
rect 8760 10412 8812 10464
rect 14096 10480 14148 10532
rect 16764 10548 16816 10600
rect 17408 10548 17460 10600
rect 18052 10591 18104 10600
rect 18052 10557 18061 10591
rect 18061 10557 18095 10591
rect 18095 10557 18104 10591
rect 18052 10548 18104 10557
rect 18972 10616 19024 10668
rect 20904 10659 20956 10668
rect 20904 10625 20913 10659
rect 20913 10625 20947 10659
rect 20947 10625 20956 10659
rect 20904 10616 20956 10625
rect 20168 10591 20220 10600
rect 20168 10557 20177 10591
rect 20177 10557 20211 10591
rect 20211 10557 20220 10591
rect 20168 10548 20220 10557
rect 9588 10412 9640 10464
rect 11428 10455 11480 10464
rect 11428 10421 11437 10455
rect 11437 10421 11471 10455
rect 11471 10421 11480 10455
rect 11428 10412 11480 10421
rect 11704 10412 11756 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 15936 10412 15988 10464
rect 16580 10412 16632 10464
rect 20812 10480 20864 10532
rect 18420 10412 18472 10464
rect 18696 10412 18748 10464
rect 19064 10412 19116 10464
rect 20536 10412 20588 10464
rect 22284 10455 22336 10464
rect 22284 10421 22293 10455
rect 22293 10421 22327 10455
rect 22327 10421 22336 10455
rect 22284 10412 22336 10421
rect 8246 10310 8298 10362
rect 8310 10310 8362 10362
rect 8374 10310 8426 10362
rect 8438 10310 8490 10362
rect 15510 10310 15562 10362
rect 15574 10310 15626 10362
rect 15638 10310 15690 10362
rect 15702 10310 15754 10362
rect 4252 10208 4304 10260
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 5448 10208 5500 10260
rect 6552 10208 6604 10260
rect 7840 10208 7892 10260
rect 8576 10208 8628 10260
rect 10508 10208 10560 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 16488 10208 16540 10260
rect 16856 10208 16908 10260
rect 17960 10208 18012 10260
rect 18880 10208 18932 10260
rect 19064 10251 19116 10260
rect 19064 10217 19073 10251
rect 19073 10217 19107 10251
rect 19107 10217 19116 10251
rect 19064 10208 19116 10217
rect 19156 10208 19208 10260
rect 4896 10140 4948 10192
rect 4988 10140 5040 10192
rect 3056 10072 3108 10124
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 2596 10047 2648 10056
rect 2596 10013 2605 10047
rect 2605 10013 2639 10047
rect 2639 10013 2648 10047
rect 2596 10004 2648 10013
rect 2688 10004 2740 10056
rect 3792 10004 3844 10056
rect 4436 10072 4488 10124
rect 6184 10115 6236 10124
rect 6184 10081 6218 10115
rect 6218 10081 6236 10115
rect 7564 10115 7616 10124
rect 6184 10072 6236 10081
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 5448 10004 5500 10056
rect 8392 10072 8444 10124
rect 11428 10140 11480 10192
rect 9404 10115 9456 10124
rect 9404 10081 9413 10115
rect 9413 10081 9447 10115
rect 9447 10081 9456 10115
rect 9404 10072 9456 10081
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 10600 10115 10652 10124
rect 10600 10081 10634 10115
rect 10634 10081 10652 10115
rect 10600 10072 10652 10081
rect 10876 10072 10928 10124
rect 14372 10140 14424 10192
rect 19340 10140 19392 10192
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 4068 9936 4120 9988
rect 5724 9936 5776 9988
rect 9220 10004 9272 10056
rect 10232 10004 10284 10056
rect 11336 10004 11388 10056
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 15384 10072 15436 10124
rect 16856 10072 16908 10124
rect 18972 10115 19024 10124
rect 14188 10047 14240 10056
rect 2872 9868 2924 9920
rect 3700 9868 3752 9920
rect 5356 9868 5408 9920
rect 6092 9868 6144 9920
rect 8760 9936 8812 9988
rect 7472 9868 7524 9920
rect 9864 9936 9916 9988
rect 10048 9936 10100 9988
rect 9128 9868 9180 9920
rect 10232 9868 10284 9920
rect 11520 9936 11572 9988
rect 14188 10013 14197 10047
rect 14197 10013 14231 10047
rect 14231 10013 14240 10047
rect 14188 10004 14240 10013
rect 11612 9868 11664 9920
rect 15108 9936 15160 9988
rect 12256 9868 12308 9920
rect 12900 9868 12952 9920
rect 14740 9868 14792 9920
rect 14924 9868 14976 9920
rect 18972 10081 18981 10115
rect 18981 10081 19015 10115
rect 19015 10081 19024 10115
rect 18972 10072 19024 10081
rect 22284 10140 22336 10192
rect 19984 10115 20036 10124
rect 19984 10081 19993 10115
rect 19993 10081 20027 10115
rect 20027 10081 20036 10115
rect 20904 10115 20956 10124
rect 19984 10072 20036 10081
rect 20904 10081 20913 10115
rect 20913 10081 20947 10115
rect 20947 10081 20956 10115
rect 20904 10072 20956 10081
rect 20168 10047 20220 10056
rect 18144 9868 18196 9920
rect 18788 9936 18840 9988
rect 20168 10013 20177 10047
rect 20177 10013 20211 10047
rect 20211 10013 20220 10047
rect 20168 10004 20220 10013
rect 19708 9936 19760 9988
rect 19524 9868 19576 9920
rect 19892 9868 19944 9920
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 4614 9766 4666 9818
rect 4678 9766 4730 9818
rect 4742 9766 4794 9818
rect 4806 9766 4858 9818
rect 11878 9766 11930 9818
rect 11942 9766 11994 9818
rect 12006 9766 12058 9818
rect 12070 9766 12122 9818
rect 19142 9766 19194 9818
rect 19206 9766 19258 9818
rect 19270 9766 19322 9818
rect 19334 9766 19386 9818
rect 2412 9664 2464 9716
rect 9772 9664 9824 9716
rect 4344 9596 4396 9648
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 3700 9571 3752 9580
rect 3700 9537 3709 9571
rect 3709 9537 3743 9571
rect 3743 9537 3752 9571
rect 3700 9528 3752 9537
rect 3792 9528 3844 9580
rect 5080 9571 5132 9580
rect 1584 9503 1636 9512
rect 1584 9469 1593 9503
rect 1593 9469 1627 9503
rect 1627 9469 1636 9503
rect 1584 9460 1636 9469
rect 2044 9460 2096 9512
rect 3424 9503 3476 9512
rect 3424 9469 3433 9503
rect 3433 9469 3467 9503
rect 3467 9469 3476 9503
rect 3424 9460 3476 9469
rect 4160 9460 4212 9512
rect 5080 9537 5089 9571
rect 5089 9537 5123 9571
rect 5123 9537 5132 9571
rect 5080 9528 5132 9537
rect 4988 9460 5040 9512
rect 5632 9460 5684 9512
rect 5724 9460 5776 9512
rect 6276 9460 6328 9512
rect 8392 9460 8444 9512
rect 8576 9503 8628 9512
rect 8576 9469 8585 9503
rect 8585 9469 8619 9503
rect 8619 9469 8628 9503
rect 8576 9460 8628 9469
rect 9588 9596 9640 9648
rect 11244 9664 11296 9716
rect 12900 9664 12952 9716
rect 9864 9571 9916 9580
rect 9864 9537 9873 9571
rect 9873 9537 9907 9571
rect 9907 9537 9916 9571
rect 9864 9528 9916 9537
rect 10140 9528 10192 9580
rect 11428 9528 11480 9580
rect 13084 9596 13136 9648
rect 14924 9596 14976 9648
rect 16396 9596 16448 9648
rect 16856 9664 16908 9716
rect 19616 9664 19668 9716
rect 20168 9664 20220 9716
rect 16672 9596 16724 9648
rect 18972 9596 19024 9648
rect 9036 9460 9088 9512
rect 9496 9460 9548 9512
rect 9772 9460 9824 9512
rect 10324 9460 10376 9512
rect 10508 9503 10560 9512
rect 10508 9469 10542 9503
rect 10542 9469 10560 9503
rect 10508 9460 10560 9469
rect 12440 9503 12492 9512
rect 12440 9469 12449 9503
rect 12449 9469 12483 9503
rect 12483 9469 12492 9503
rect 12440 9460 12492 9469
rect 14648 9528 14700 9580
rect 16488 9528 16540 9580
rect 3056 9367 3108 9376
rect 3056 9333 3065 9367
rect 3065 9333 3099 9367
rect 3099 9333 3108 9367
rect 3056 9324 3108 9333
rect 3516 9324 3568 9376
rect 3700 9324 3752 9376
rect 4068 9367 4120 9376
rect 4068 9333 4077 9367
rect 4077 9333 4111 9367
rect 4111 9333 4120 9367
rect 4068 9324 4120 9333
rect 5264 9324 5316 9376
rect 5356 9324 5408 9376
rect 7380 9392 7432 9444
rect 7656 9435 7708 9444
rect 7656 9401 7665 9435
rect 7665 9401 7699 9435
rect 7699 9401 7708 9435
rect 7656 9392 7708 9401
rect 6184 9324 6236 9376
rect 9128 9392 9180 9444
rect 11244 9392 11296 9444
rect 11796 9392 11848 9444
rect 12992 9392 13044 9444
rect 13360 9392 13412 9444
rect 14372 9460 14424 9512
rect 14556 9460 14608 9512
rect 14740 9460 14792 9512
rect 10600 9324 10652 9376
rect 13084 9324 13136 9376
rect 14556 9367 14608 9376
rect 14556 9333 14565 9367
rect 14565 9333 14599 9367
rect 14599 9333 14608 9367
rect 14556 9324 14608 9333
rect 14740 9324 14792 9376
rect 16948 9460 17000 9512
rect 16212 9392 16264 9444
rect 18144 9528 18196 9580
rect 19340 9528 19392 9580
rect 19616 9528 19668 9580
rect 21640 9571 21692 9580
rect 21640 9537 21649 9571
rect 21649 9537 21683 9571
rect 21683 9537 21692 9571
rect 21640 9528 21692 9537
rect 22192 9528 22244 9580
rect 18972 9460 19024 9512
rect 19156 9460 19208 9512
rect 19432 9460 19484 9512
rect 20260 9460 20312 9512
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 16580 9324 16632 9376
rect 18604 9324 18656 9376
rect 18788 9324 18840 9376
rect 20536 9392 20588 9444
rect 19432 9324 19484 9376
rect 19524 9367 19576 9376
rect 19524 9333 19539 9367
rect 19539 9333 19573 9367
rect 19573 9333 19576 9367
rect 19524 9324 19576 9333
rect 20076 9324 20128 9376
rect 21180 9367 21232 9376
rect 21180 9333 21189 9367
rect 21189 9333 21223 9367
rect 21223 9333 21232 9367
rect 21180 9324 21232 9333
rect 8246 9222 8298 9274
rect 8310 9222 8362 9274
rect 8374 9222 8426 9274
rect 8438 9222 8490 9274
rect 15510 9222 15562 9274
rect 15574 9222 15626 9274
rect 15638 9222 15690 9274
rect 15702 9222 15754 9274
rect 2504 9163 2556 9172
rect 2504 9129 2513 9163
rect 2513 9129 2547 9163
rect 2547 9129 2556 9163
rect 2504 9120 2556 9129
rect 4436 9120 4488 9172
rect 5356 9120 5408 9172
rect 5540 9163 5592 9172
rect 5540 9129 5549 9163
rect 5549 9129 5583 9163
rect 5583 9129 5592 9163
rect 5540 9120 5592 9129
rect 5908 9163 5960 9172
rect 5908 9129 5917 9163
rect 5917 9129 5951 9163
rect 5951 9129 5960 9163
rect 5908 9120 5960 9129
rect 6000 9163 6052 9172
rect 6000 9129 6009 9163
rect 6009 9129 6043 9163
rect 6043 9129 6052 9163
rect 6552 9163 6604 9172
rect 6000 9120 6052 9129
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 3884 9052 3936 9104
rect 4068 9052 4120 9104
rect 7104 9052 7156 9104
rect 3700 8984 3752 9036
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 6828 8984 6880 9036
rect 5080 8916 5132 8968
rect 5264 8916 5316 8968
rect 5448 8916 5500 8968
rect 6000 8916 6052 8968
rect 7012 8959 7064 8968
rect 7012 8925 7021 8959
rect 7021 8925 7055 8959
rect 7055 8925 7064 8959
rect 7012 8916 7064 8925
rect 5356 8848 5408 8900
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 5080 8780 5132 8832
rect 5448 8780 5500 8832
rect 6276 8780 6328 8832
rect 6828 8848 6880 8900
rect 7380 8984 7432 9036
rect 8576 9052 8628 9104
rect 9772 9120 9824 9172
rect 10784 9120 10836 9172
rect 7932 9027 7984 9036
rect 7932 8993 7941 9027
rect 7941 8993 7975 9027
rect 7975 8993 7984 9027
rect 7932 8984 7984 8993
rect 7656 8916 7708 8968
rect 9496 8984 9548 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10876 8984 10928 9036
rect 11520 8984 11572 9036
rect 11704 9027 11756 9036
rect 11704 8993 11738 9027
rect 11738 8993 11756 9027
rect 11704 8984 11756 8993
rect 12624 9052 12676 9104
rect 12900 9052 12952 9104
rect 13452 9120 13504 9172
rect 14648 9120 14700 9172
rect 16304 9120 16356 9172
rect 16396 9120 16448 9172
rect 16856 9120 16908 9172
rect 18236 9163 18288 9172
rect 18236 9129 18245 9163
rect 18245 9129 18279 9163
rect 18279 9129 18288 9163
rect 18236 9120 18288 9129
rect 18512 9120 18564 9172
rect 14556 9052 14608 9104
rect 14924 9052 14976 9104
rect 15292 8984 15344 9036
rect 15476 9052 15528 9104
rect 16764 9052 16816 9104
rect 16488 8984 16540 9036
rect 18328 8984 18380 9036
rect 18696 8984 18748 9036
rect 8852 8916 8904 8968
rect 8944 8916 8996 8968
rect 12440 8916 12492 8968
rect 14372 8916 14424 8968
rect 14556 8916 14608 8968
rect 14832 8916 14884 8968
rect 15844 8959 15896 8968
rect 15844 8925 15853 8959
rect 15853 8925 15887 8959
rect 15887 8925 15896 8959
rect 15844 8916 15896 8925
rect 18144 8916 18196 8968
rect 18788 8916 18840 8968
rect 19708 8984 19760 9036
rect 20352 9120 20404 9172
rect 20168 9052 20220 9104
rect 22284 9052 22336 9104
rect 20904 9027 20956 9036
rect 20904 8993 20913 9027
rect 20913 8993 20947 9027
rect 20947 8993 20956 9027
rect 20904 8984 20956 8993
rect 20536 8916 20588 8968
rect 7564 8891 7616 8900
rect 7564 8857 7573 8891
rect 7573 8857 7607 8891
rect 7607 8857 7616 8891
rect 7564 8848 7616 8857
rect 9496 8848 9548 8900
rect 9680 8780 9732 8832
rect 10048 8780 10100 8832
rect 11336 8848 11388 8900
rect 14096 8848 14148 8900
rect 11244 8780 11296 8832
rect 12624 8780 12676 8832
rect 12992 8780 13044 8832
rect 14188 8780 14240 8832
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 15476 8848 15528 8900
rect 16396 8848 16448 8900
rect 17776 8823 17828 8832
rect 17776 8789 17785 8823
rect 17785 8789 17819 8823
rect 17819 8789 17828 8823
rect 17776 8780 17828 8789
rect 22192 8848 22244 8900
rect 19432 8780 19484 8832
rect 4614 8678 4666 8730
rect 4678 8678 4730 8730
rect 4742 8678 4794 8730
rect 4806 8678 4858 8730
rect 11878 8678 11930 8730
rect 11942 8678 11994 8730
rect 12006 8678 12058 8730
rect 12070 8678 12122 8730
rect 19142 8678 19194 8730
rect 19206 8678 19258 8730
rect 19270 8678 19322 8730
rect 19334 8678 19386 8730
rect 4068 8576 4120 8628
rect 6920 8576 6972 8628
rect 11244 8576 11296 8628
rect 11704 8619 11756 8628
rect 11704 8585 11713 8619
rect 11713 8585 11747 8619
rect 11747 8585 11756 8619
rect 11704 8576 11756 8585
rect 15292 8576 15344 8628
rect 15384 8576 15436 8628
rect 15936 8576 15988 8628
rect 16304 8576 16356 8628
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 5448 8508 5500 8560
rect 6000 8508 6052 8560
rect 2964 8440 3016 8492
rect 5356 8483 5408 8492
rect 5356 8449 5365 8483
rect 5365 8449 5399 8483
rect 5399 8449 5408 8483
rect 5356 8440 5408 8449
rect 7472 8508 7524 8560
rect 8116 8508 8168 8560
rect 8668 8508 8720 8560
rect 11428 8508 11480 8560
rect 12164 8508 12216 8560
rect 7932 8440 7984 8492
rect 8208 8440 8260 8492
rect 2044 8372 2096 8424
rect 4068 8372 4120 8424
rect 5080 8415 5132 8424
rect 5080 8381 5089 8415
rect 5089 8381 5123 8415
rect 5123 8381 5132 8415
rect 5080 8372 5132 8381
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 8484 8372 8536 8424
rect 9956 8440 10008 8492
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 12992 8483 13044 8492
rect 4252 8304 4304 8356
rect 5908 8304 5960 8356
rect 6184 8347 6236 8356
rect 6184 8313 6193 8347
rect 6193 8313 6227 8347
rect 6227 8313 6236 8347
rect 6184 8304 6236 8313
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 8208 8304 8260 8356
rect 8760 8304 8812 8356
rect 9220 8372 9272 8424
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 14648 8508 14700 8560
rect 10876 8304 10928 8356
rect 11060 8304 11112 8356
rect 13084 8372 13136 8424
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 14556 8440 14608 8492
rect 15384 8440 15436 8492
rect 14096 8372 14148 8424
rect 14648 8372 14700 8424
rect 16304 8440 16356 8492
rect 15936 8372 15988 8424
rect 16212 8372 16264 8424
rect 17960 8440 18012 8492
rect 20076 8440 20128 8492
rect 21180 8576 21232 8628
rect 20812 8508 20864 8560
rect 22284 8551 22336 8560
rect 22284 8517 22293 8551
rect 22293 8517 22327 8551
rect 22327 8517 22336 8551
rect 22284 8508 22336 8517
rect 20904 8483 20956 8492
rect 16580 8372 16632 8424
rect 19616 8372 19668 8424
rect 5724 8236 5776 8288
rect 7748 8236 7800 8288
rect 9220 8236 9272 8288
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 14832 8304 14884 8356
rect 17132 8304 17184 8356
rect 17960 8304 18012 8356
rect 19524 8347 19576 8356
rect 19524 8313 19533 8347
rect 19533 8313 19567 8347
rect 19567 8313 19576 8347
rect 19524 8304 19576 8313
rect 20904 8449 20913 8483
rect 20913 8449 20947 8483
rect 20947 8449 20956 8483
rect 20904 8440 20956 8449
rect 20628 8372 20680 8424
rect 22192 8372 22244 8424
rect 22284 8304 22336 8356
rect 13728 8236 13780 8288
rect 14556 8236 14608 8288
rect 15200 8236 15252 8288
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 8246 8134 8298 8186
rect 8310 8134 8362 8186
rect 8374 8134 8426 8186
rect 8438 8134 8490 8186
rect 15510 8134 15562 8186
rect 15574 8134 15626 8186
rect 15638 8134 15690 8186
rect 15702 8134 15754 8186
rect 5264 8075 5316 8084
rect 5264 8041 5273 8075
rect 5273 8041 5307 8075
rect 5307 8041 5316 8075
rect 5264 8032 5316 8041
rect 5908 8075 5960 8084
rect 5908 8041 5917 8075
rect 5917 8041 5951 8075
rect 5951 8041 5960 8075
rect 5908 8032 5960 8041
rect 6644 8032 6696 8084
rect 7380 8032 7432 8084
rect 8760 8032 8812 8084
rect 7196 7964 7248 8016
rect 10048 7964 10100 8016
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 9036 7896 9088 7948
rect 9588 7896 9640 7948
rect 10508 7896 10560 7948
rect 11336 7939 11388 7948
rect 11336 7905 11345 7939
rect 11345 7905 11379 7939
rect 11379 7905 11388 7939
rect 11336 7896 11388 7905
rect 14740 8032 14792 8084
rect 16764 8075 16816 8084
rect 16764 8041 16773 8075
rect 16773 8041 16807 8075
rect 16807 8041 16816 8075
rect 16764 8032 16816 8041
rect 18420 8075 18472 8084
rect 18420 8041 18429 8075
rect 18429 8041 18463 8075
rect 18463 8041 18472 8075
rect 18420 8032 18472 8041
rect 19432 8032 19484 8084
rect 19984 8032 20036 8084
rect 20168 8032 20220 8084
rect 12992 7964 13044 8016
rect 15844 7964 15896 8016
rect 16304 7964 16356 8016
rect 14648 7896 14700 7948
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 6460 7871 6512 7880
rect 5448 7828 5500 7837
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 6184 7692 6236 7744
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 9128 7828 9180 7880
rect 9496 7828 9548 7880
rect 11520 7828 11572 7880
rect 13544 7871 13596 7880
rect 13544 7837 13553 7871
rect 13553 7837 13587 7871
rect 13587 7837 13596 7871
rect 13544 7828 13596 7837
rect 15200 7828 15252 7880
rect 8944 7760 8996 7812
rect 9312 7760 9364 7812
rect 14740 7760 14792 7812
rect 10876 7692 10928 7744
rect 12992 7692 13044 7744
rect 13084 7692 13136 7744
rect 13820 7692 13872 7744
rect 13912 7692 13964 7744
rect 17776 7896 17828 7948
rect 20260 7964 20312 8016
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 19616 7896 19668 7948
rect 21916 7939 21968 7948
rect 21916 7905 21925 7939
rect 21925 7905 21959 7939
rect 21959 7905 21968 7939
rect 21916 7896 21968 7905
rect 20076 7828 20128 7880
rect 20444 7871 20496 7880
rect 20444 7837 20453 7871
rect 20453 7837 20487 7871
rect 20487 7837 20496 7871
rect 20444 7828 20496 7837
rect 20536 7871 20588 7880
rect 20536 7837 20545 7871
rect 20545 7837 20579 7871
rect 20579 7837 20588 7871
rect 20536 7828 20588 7837
rect 21548 7871 21600 7880
rect 18420 7692 18472 7744
rect 21548 7837 21557 7871
rect 21557 7837 21591 7871
rect 21591 7837 21600 7871
rect 21548 7828 21600 7837
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 21640 7692 21692 7744
rect 22376 7692 22428 7744
rect 4614 7590 4666 7642
rect 4678 7590 4730 7642
rect 4742 7590 4794 7642
rect 4806 7590 4858 7642
rect 11878 7590 11930 7642
rect 11942 7590 11994 7642
rect 12006 7590 12058 7642
rect 12070 7590 12122 7642
rect 19142 7590 19194 7642
rect 19206 7590 19258 7642
rect 19270 7590 19322 7642
rect 19334 7590 19386 7642
rect 6736 7488 6788 7540
rect 7012 7488 7064 7540
rect 9588 7531 9640 7540
rect 7564 7420 7616 7472
rect 6184 7395 6236 7404
rect 4252 7259 4304 7268
rect 4252 7225 4261 7259
rect 4261 7225 4295 7259
rect 4295 7225 4304 7259
rect 4252 7216 4304 7225
rect 5264 7216 5316 7268
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 9680 7488 9732 7540
rect 10416 7488 10468 7540
rect 12256 7488 12308 7540
rect 16396 7531 16448 7540
rect 16396 7497 16405 7531
rect 16405 7497 16439 7531
rect 16439 7497 16448 7531
rect 16396 7488 16448 7497
rect 12716 7420 12768 7472
rect 7748 7284 7800 7336
rect 7932 7284 7984 7336
rect 10048 7352 10100 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 11520 7395 11572 7404
rect 10416 7352 10468 7361
rect 11520 7361 11529 7395
rect 11529 7361 11563 7395
rect 11563 7361 11572 7395
rect 11520 7352 11572 7361
rect 13912 7420 13964 7472
rect 15476 7420 15528 7472
rect 15936 7463 15988 7472
rect 15936 7429 15945 7463
rect 15945 7429 15979 7463
rect 15979 7429 15988 7463
rect 15936 7420 15988 7429
rect 16304 7420 16356 7472
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 13268 7352 13320 7404
rect 14740 7352 14792 7404
rect 11704 7284 11756 7336
rect 12164 7284 12216 7336
rect 12348 7284 12400 7336
rect 12808 7284 12860 7336
rect 13636 7284 13688 7336
rect 8116 7216 8168 7268
rect 8576 7216 8628 7268
rect 9496 7216 9548 7268
rect 7564 7148 7616 7200
rect 10048 7148 10100 7200
rect 10876 7216 10928 7268
rect 14004 7284 14056 7336
rect 16856 7352 16908 7404
rect 19616 7488 19668 7540
rect 20352 7488 20404 7540
rect 20076 7420 20128 7472
rect 19432 7395 19484 7404
rect 10416 7148 10468 7200
rect 11060 7148 11112 7200
rect 12624 7148 12676 7200
rect 12716 7148 12768 7200
rect 13176 7148 13228 7200
rect 14556 7191 14608 7200
rect 14556 7157 14571 7191
rect 14571 7157 14605 7191
rect 14605 7157 14608 7191
rect 14556 7148 14608 7157
rect 14832 7148 14884 7200
rect 18052 7216 18104 7268
rect 18788 7284 18840 7336
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 20444 7352 20496 7404
rect 21732 7395 21784 7404
rect 21732 7361 21741 7395
rect 21741 7361 21775 7395
rect 21775 7361 21784 7395
rect 21732 7352 21784 7361
rect 20260 7284 20312 7336
rect 21640 7327 21692 7336
rect 21640 7293 21649 7327
rect 21649 7293 21683 7327
rect 21683 7293 21692 7327
rect 21640 7284 21692 7293
rect 16948 7191 17000 7200
rect 16948 7157 16957 7191
rect 16957 7157 16991 7191
rect 16991 7157 17000 7191
rect 16948 7148 17000 7157
rect 18972 7148 19024 7200
rect 19800 7148 19852 7200
rect 20076 7148 20128 7200
rect 20904 7148 20956 7200
rect 8246 7046 8298 7098
rect 8310 7046 8362 7098
rect 8374 7046 8426 7098
rect 8438 7046 8490 7098
rect 15510 7046 15562 7098
rect 15574 7046 15626 7098
rect 15638 7046 15690 7098
rect 15702 7046 15754 7098
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 7564 6944 7616 6996
rect 9680 6944 9732 6996
rect 10048 6987 10100 6996
rect 10048 6953 10057 6987
rect 10057 6953 10091 6987
rect 10091 6953 10100 6987
rect 10048 6944 10100 6953
rect 7380 6876 7432 6928
rect 12256 6944 12308 6996
rect 12164 6876 12216 6928
rect 12716 6876 12768 6928
rect 16580 6944 16632 6996
rect 4344 6740 4396 6792
rect 7656 6808 7708 6860
rect 9220 6808 9272 6860
rect 9772 6808 9824 6860
rect 7564 6783 7616 6792
rect 6552 6672 6604 6724
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 9864 6740 9916 6792
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11612 6808 11664 6860
rect 12072 6740 12124 6792
rect 12256 6851 12308 6860
rect 12256 6817 12265 6851
rect 12265 6817 12299 6851
rect 12299 6817 12308 6851
rect 12900 6851 12952 6860
rect 12256 6808 12308 6817
rect 12900 6817 12909 6851
rect 12909 6817 12943 6851
rect 12943 6817 12952 6851
rect 12900 6808 12952 6817
rect 12532 6740 12584 6792
rect 17408 6944 17460 6996
rect 18788 6944 18840 6996
rect 19800 6876 19852 6928
rect 20536 6876 20588 6928
rect 13636 6808 13688 6860
rect 7748 6672 7800 6724
rect 9312 6647 9364 6656
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 10048 6604 10100 6656
rect 10876 6647 10928 6656
rect 10876 6613 10885 6647
rect 10885 6613 10919 6647
rect 10919 6613 10928 6647
rect 10876 6604 10928 6613
rect 13176 6672 13228 6724
rect 13084 6604 13136 6656
rect 13820 6604 13872 6656
rect 14648 6604 14700 6656
rect 16948 6808 17000 6860
rect 15200 6740 15252 6792
rect 16672 6740 16724 6792
rect 17684 6808 17736 6860
rect 18696 6808 18748 6860
rect 20720 6740 20772 6792
rect 16856 6672 16908 6724
rect 16396 6604 16448 6656
rect 19432 6604 19484 6656
rect 20076 6604 20128 6656
rect 20352 6604 20404 6656
rect 20536 6647 20588 6656
rect 20536 6613 20545 6647
rect 20545 6613 20579 6647
rect 20579 6613 20588 6647
rect 20536 6604 20588 6613
rect 21640 6604 21692 6656
rect 4614 6502 4666 6554
rect 4678 6502 4730 6554
rect 4742 6502 4794 6554
rect 4806 6502 4858 6554
rect 11878 6502 11930 6554
rect 11942 6502 11994 6554
rect 12006 6502 12058 6554
rect 12070 6502 12122 6554
rect 19142 6502 19194 6554
rect 19206 6502 19258 6554
rect 19270 6502 19322 6554
rect 19334 6502 19386 6554
rect 3056 6332 3108 6384
rect 8024 6332 8076 6384
rect 7104 6264 7156 6316
rect 8116 6264 8168 6316
rect 8576 6400 8628 6452
rect 10876 6400 10928 6452
rect 11704 6400 11756 6452
rect 12256 6400 12308 6452
rect 12900 6400 12952 6452
rect 15292 6400 15344 6452
rect 16120 6400 16172 6452
rect 19800 6443 19852 6452
rect 13084 6332 13136 6384
rect 14096 6332 14148 6384
rect 19800 6409 19809 6443
rect 19809 6409 19843 6443
rect 19843 6409 19852 6443
rect 19800 6400 19852 6409
rect 20260 6443 20312 6452
rect 20260 6409 20269 6443
rect 20269 6409 20303 6443
rect 20303 6409 20312 6443
rect 20260 6400 20312 6409
rect 20904 6400 20956 6452
rect 8300 6239 8352 6248
rect 8300 6205 8309 6239
rect 8309 6205 8343 6239
rect 8343 6205 8352 6239
rect 8300 6196 8352 6205
rect 9312 6196 9364 6248
rect 10048 6239 10100 6248
rect 10048 6205 10057 6239
rect 10057 6205 10091 6239
rect 10091 6205 10100 6239
rect 10048 6196 10100 6205
rect 10508 6196 10560 6248
rect 11796 6264 11848 6316
rect 11704 6196 11756 6248
rect 14280 6264 14332 6316
rect 14832 6264 14884 6316
rect 15108 6264 15160 6316
rect 16304 6239 16356 6248
rect 6828 6103 6880 6112
rect 6828 6069 6837 6103
rect 6837 6069 6871 6103
rect 6871 6069 6880 6103
rect 6828 6060 6880 6069
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 7564 6060 7616 6112
rect 11520 6128 11572 6180
rect 11060 6060 11112 6112
rect 11244 6060 11296 6112
rect 12992 6060 13044 6112
rect 16304 6205 16313 6239
rect 16313 6205 16347 6239
rect 16347 6205 16356 6239
rect 16304 6196 16356 6205
rect 18420 6239 18472 6248
rect 13820 6128 13872 6180
rect 14188 6128 14240 6180
rect 15936 6128 15988 6180
rect 18420 6205 18429 6239
rect 18429 6205 18463 6239
rect 18463 6205 18472 6239
rect 18420 6196 18472 6205
rect 19708 6196 19760 6248
rect 20076 6239 20128 6248
rect 20076 6205 20085 6239
rect 20085 6205 20119 6239
rect 20119 6205 20128 6239
rect 20076 6196 20128 6205
rect 20720 6196 20772 6248
rect 21640 6196 21692 6248
rect 13728 6060 13780 6112
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 15108 6103 15160 6112
rect 15108 6069 15117 6103
rect 15117 6069 15151 6103
rect 15151 6069 15160 6103
rect 15108 6060 15160 6069
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 19432 6128 19484 6180
rect 21732 6060 21784 6112
rect 8246 5958 8298 6010
rect 8310 5958 8362 6010
rect 8374 5958 8426 6010
rect 8438 5958 8490 6010
rect 15510 5958 15562 6010
rect 15574 5958 15626 6010
rect 15638 5958 15690 6010
rect 15702 5958 15754 6010
rect 6276 5856 6328 5908
rect 7288 5856 7340 5908
rect 6828 5788 6880 5840
rect 13820 5856 13872 5908
rect 13912 5856 13964 5908
rect 16856 5856 16908 5908
rect 19984 5856 20036 5908
rect 7196 5720 7248 5772
rect 8024 5720 8076 5772
rect 9588 5720 9640 5772
rect 9864 5720 9916 5772
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 9128 5652 9180 5704
rect 12256 5788 12308 5840
rect 12440 5788 12492 5840
rect 11704 5720 11756 5772
rect 12624 5720 12676 5772
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 14464 5720 14516 5772
rect 10508 5652 10560 5704
rect 9220 5516 9272 5568
rect 12808 5584 12860 5636
rect 15936 5720 15988 5772
rect 14832 5652 14884 5704
rect 17684 5720 17736 5772
rect 17868 5763 17920 5772
rect 17868 5729 17877 5763
rect 17877 5729 17911 5763
rect 17911 5729 17920 5763
rect 17868 5720 17920 5729
rect 19524 5720 19576 5772
rect 22100 5720 22152 5772
rect 16120 5695 16172 5704
rect 16120 5661 16129 5695
rect 16129 5661 16163 5695
rect 16163 5661 16172 5695
rect 18880 5695 18932 5704
rect 16120 5652 16172 5661
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 19432 5652 19484 5704
rect 20536 5652 20588 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 12348 5559 12400 5568
rect 12348 5525 12357 5559
rect 12357 5525 12391 5559
rect 12391 5525 12400 5559
rect 12348 5516 12400 5525
rect 12900 5516 12952 5568
rect 13176 5516 13228 5568
rect 19340 5584 19392 5636
rect 20168 5584 20220 5636
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 17408 5516 17460 5568
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 20536 5516 20588 5568
rect 22284 5559 22336 5568
rect 22284 5525 22293 5559
rect 22293 5525 22327 5559
rect 22327 5525 22336 5559
rect 22284 5516 22336 5525
rect 4614 5414 4666 5466
rect 4678 5414 4730 5466
rect 4742 5414 4794 5466
rect 4806 5414 4858 5466
rect 11878 5414 11930 5466
rect 11942 5414 11994 5466
rect 12006 5414 12058 5466
rect 12070 5414 12122 5466
rect 19142 5414 19194 5466
rect 19206 5414 19258 5466
rect 19270 5414 19322 5466
rect 19334 5414 19386 5466
rect 7840 5312 7892 5364
rect 9588 5355 9640 5364
rect 9588 5321 9597 5355
rect 9597 5321 9631 5355
rect 9631 5321 9640 5355
rect 9588 5312 9640 5321
rect 7932 5108 7984 5160
rect 11428 5312 11480 5364
rect 11704 5312 11756 5364
rect 12624 5312 12676 5364
rect 13912 5244 13964 5296
rect 15016 5244 15068 5296
rect 17408 5312 17460 5364
rect 19432 5355 19484 5364
rect 12900 5219 12952 5228
rect 12900 5185 12909 5219
rect 12909 5185 12943 5219
rect 12943 5185 12952 5219
rect 12900 5176 12952 5185
rect 17592 5219 17644 5228
rect 10508 5108 10560 5160
rect 11244 5108 11296 5160
rect 12992 5108 13044 5160
rect 12348 5040 12400 5092
rect 14372 5040 14424 5092
rect 15200 5108 15252 5160
rect 17592 5185 17601 5219
rect 17601 5185 17635 5219
rect 17635 5185 17644 5219
rect 17592 5176 17644 5185
rect 19432 5321 19441 5355
rect 19441 5321 19475 5355
rect 19475 5321 19484 5355
rect 19432 5312 19484 5321
rect 20076 5312 20128 5364
rect 10508 4972 10560 5024
rect 13452 4972 13504 5024
rect 13544 4972 13596 5024
rect 15016 4972 15068 5024
rect 15568 5083 15620 5092
rect 15568 5049 15602 5083
rect 15602 5049 15620 5083
rect 15568 5040 15620 5049
rect 16396 5040 16448 5092
rect 19524 5108 19576 5160
rect 20904 5151 20956 5160
rect 20904 5117 20913 5151
rect 20913 5117 20947 5151
rect 20947 5117 20956 5151
rect 20904 5108 20956 5117
rect 16488 4972 16540 5024
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17040 4972 17092 5024
rect 19248 5040 19300 5092
rect 20260 5040 20312 5092
rect 20720 5040 20772 5092
rect 18696 4972 18748 5024
rect 20168 5015 20220 5024
rect 20168 4981 20177 5015
rect 20177 4981 20211 5015
rect 20211 4981 20220 5015
rect 20168 4972 20220 4981
rect 22100 4972 22152 5024
rect 8246 4870 8298 4922
rect 8310 4870 8362 4922
rect 8374 4870 8426 4922
rect 8438 4870 8490 4922
rect 15510 4870 15562 4922
rect 15574 4870 15626 4922
rect 15638 4870 15690 4922
rect 15702 4870 15754 4922
rect 10048 4811 10100 4820
rect 10048 4777 10057 4811
rect 10057 4777 10091 4811
rect 10091 4777 10100 4811
rect 10048 4768 10100 4777
rect 11704 4768 11756 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14372 4768 14424 4820
rect 14464 4768 14516 4820
rect 14648 4811 14700 4820
rect 14648 4777 14657 4811
rect 14657 4777 14691 4811
rect 14691 4777 14700 4811
rect 14648 4768 14700 4777
rect 18880 4768 18932 4820
rect 18972 4768 19024 4820
rect 19616 4768 19668 4820
rect 20076 4811 20128 4820
rect 20076 4777 20085 4811
rect 20085 4777 20119 4811
rect 20119 4777 20128 4811
rect 20076 4768 20128 4777
rect 13728 4700 13780 4752
rect 14924 4700 14976 4752
rect 15200 4700 15252 4752
rect 10508 4607 10560 4616
rect 10508 4573 10517 4607
rect 10517 4573 10551 4607
rect 10551 4573 10560 4607
rect 10508 4564 10560 4573
rect 11612 4632 11664 4684
rect 12348 4632 12400 4684
rect 15108 4632 15160 4684
rect 16948 4700 17000 4752
rect 18052 4700 18104 4752
rect 19248 4700 19300 4752
rect 22284 4768 22336 4820
rect 21272 4700 21324 4752
rect 16580 4675 16632 4684
rect 16580 4641 16589 4675
rect 16589 4641 16623 4675
rect 16623 4641 16632 4675
rect 16580 4632 16632 4641
rect 12624 4564 12676 4616
rect 12808 4607 12860 4616
rect 12808 4573 12817 4607
rect 12817 4573 12851 4607
rect 12851 4573 12860 4607
rect 12808 4564 12860 4573
rect 13084 4496 13136 4548
rect 13728 4496 13780 4548
rect 15200 4564 15252 4616
rect 17592 4632 17644 4684
rect 18236 4632 18288 4684
rect 17408 4564 17460 4616
rect 15016 4496 15068 4548
rect 20444 4564 20496 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 12256 4428 12308 4480
rect 14188 4471 14240 4480
rect 14188 4437 14197 4471
rect 14197 4437 14231 4471
rect 14231 4437 14240 4471
rect 14188 4428 14240 4437
rect 14372 4428 14424 4480
rect 14924 4428 14976 4480
rect 17316 4428 17368 4480
rect 17868 4428 17920 4480
rect 19708 4428 19760 4480
rect 20812 4496 20864 4548
rect 20720 4428 20772 4480
rect 4614 4326 4666 4378
rect 4678 4326 4730 4378
rect 4742 4326 4794 4378
rect 4806 4326 4858 4378
rect 11878 4326 11930 4378
rect 11942 4326 11994 4378
rect 12006 4326 12058 4378
rect 12070 4326 12122 4378
rect 19142 4326 19194 4378
rect 19206 4326 19258 4378
rect 19270 4326 19322 4378
rect 19334 4326 19386 4378
rect 9496 4156 9548 4208
rect 13084 4224 13136 4276
rect 13268 4267 13320 4276
rect 13268 4233 13277 4267
rect 13277 4233 13311 4267
rect 13311 4233 13320 4267
rect 13268 4224 13320 4233
rect 13544 4224 13596 4276
rect 14556 4224 14608 4276
rect 16672 4224 16724 4276
rect 20260 4267 20312 4276
rect 20260 4233 20269 4267
rect 20269 4233 20303 4267
rect 20303 4233 20312 4267
rect 20260 4224 20312 4233
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 9220 4020 9272 4072
rect 10232 4020 10284 4072
rect 11520 4088 11572 4140
rect 12808 4156 12860 4208
rect 13360 4156 13412 4208
rect 11888 4088 11940 4140
rect 13544 4088 13596 4140
rect 17592 4156 17644 4208
rect 22376 4224 22428 4276
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 18144 4088 18196 4140
rect 11244 4020 11296 4072
rect 12716 4063 12768 4072
rect 12716 4029 12725 4063
rect 12725 4029 12759 4063
rect 12759 4029 12768 4063
rect 12716 4020 12768 4029
rect 13452 4020 13504 4072
rect 14372 4020 14424 4072
rect 8576 3952 8628 4004
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 13176 3952 13228 4004
rect 14556 3995 14608 4004
rect 11336 3884 11388 3936
rect 11428 3884 11480 3936
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14556 3961 14590 3995
rect 14590 3961 14608 3995
rect 14556 3952 14608 3961
rect 16580 4020 16632 4072
rect 16672 4020 16724 4072
rect 19708 4131 19760 4140
rect 19708 4097 19717 4131
rect 19717 4097 19751 4131
rect 19751 4097 19760 4131
rect 19708 4088 19760 4097
rect 20076 4063 20128 4072
rect 16120 3952 16172 4004
rect 16856 3952 16908 4004
rect 15108 3884 15160 3936
rect 16304 3884 16356 3936
rect 18052 3927 18104 3936
rect 18052 3893 18061 3927
rect 18061 3893 18095 3927
rect 18095 3893 18104 3927
rect 18052 3884 18104 3893
rect 18328 3884 18380 3936
rect 18880 3884 18932 3936
rect 19800 3952 19852 4004
rect 20076 4029 20085 4063
rect 20085 4029 20119 4063
rect 20119 4029 20128 4063
rect 20076 4020 20128 4029
rect 20444 4020 20496 4072
rect 22284 3952 22336 4004
rect 19984 3884 20036 3936
rect 21272 3884 21324 3936
rect 8246 3782 8298 3834
rect 8310 3782 8362 3834
rect 8374 3782 8426 3834
rect 8438 3782 8490 3834
rect 15510 3782 15562 3834
rect 15574 3782 15626 3834
rect 15638 3782 15690 3834
rect 15702 3782 15754 3834
rect 12992 3680 13044 3732
rect 13176 3723 13228 3732
rect 13176 3689 13185 3723
rect 13185 3689 13219 3723
rect 13219 3689 13228 3723
rect 13176 3680 13228 3689
rect 3516 3612 3568 3664
rect 11428 3612 11480 3664
rect 11888 3612 11940 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 13912 3612 13964 3664
rect 14556 3655 14608 3664
rect 14556 3621 14565 3655
rect 14565 3621 14599 3655
rect 14599 3621 14608 3655
rect 14556 3612 14608 3621
rect 16212 3612 16264 3664
rect 18788 3680 18840 3732
rect 19892 3680 19944 3732
rect 20168 3680 20220 3732
rect 22284 3723 22336 3732
rect 22284 3689 22293 3723
rect 22293 3689 22327 3723
rect 22327 3689 22336 3723
rect 22284 3680 22336 3689
rect 17408 3612 17460 3664
rect 18052 3612 18104 3664
rect 12440 3544 12492 3596
rect 13636 3476 13688 3528
rect 12440 3408 12492 3460
rect 14280 3408 14332 3460
rect 12256 3340 12308 3392
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15016 3544 15068 3596
rect 15568 3587 15620 3596
rect 15568 3553 15591 3587
rect 15591 3553 15620 3587
rect 15568 3544 15620 3553
rect 15844 3544 15896 3596
rect 18420 3544 18472 3596
rect 18604 3587 18656 3596
rect 18604 3553 18613 3587
rect 18613 3553 18647 3587
rect 18647 3553 18656 3587
rect 18604 3544 18656 3553
rect 18696 3544 18748 3596
rect 21180 3587 21232 3596
rect 21180 3553 21214 3587
rect 21214 3553 21232 3587
rect 21180 3544 21232 3553
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 14924 3476 14976 3528
rect 16396 3408 16448 3460
rect 20168 3476 20220 3528
rect 20444 3476 20496 3528
rect 15936 3340 15988 3392
rect 18604 3408 18656 3460
rect 18328 3383 18380 3392
rect 18328 3349 18337 3383
rect 18337 3349 18371 3383
rect 18371 3349 18380 3383
rect 18328 3340 18380 3349
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 4614 3238 4666 3290
rect 4678 3238 4730 3290
rect 4742 3238 4794 3290
rect 4806 3238 4858 3290
rect 11878 3238 11930 3290
rect 11942 3238 11994 3290
rect 12006 3238 12058 3290
rect 12070 3238 12122 3290
rect 19142 3238 19194 3290
rect 19206 3238 19258 3290
rect 19270 3238 19322 3290
rect 19334 3238 19386 3290
rect 7472 3136 7524 3188
rect 13728 3136 13780 3188
rect 16672 3136 16724 3188
rect 17408 3179 17460 3188
rect 17408 3145 17417 3179
rect 17417 3145 17451 3179
rect 17451 3145 17460 3179
rect 17408 3136 17460 3145
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 18604 3136 18656 3188
rect 15568 3111 15620 3120
rect 15568 3077 15577 3111
rect 15577 3077 15611 3111
rect 15611 3077 15620 3111
rect 15568 3068 15620 3077
rect 19800 3136 19852 3188
rect 20168 3111 20220 3120
rect 20168 3077 20177 3111
rect 20177 3077 20211 3111
rect 20211 3077 20220 3111
rect 20168 3068 20220 3077
rect 6920 3000 6972 3052
rect 13728 3043 13780 3052
rect 13728 3009 13737 3043
rect 13737 3009 13771 3043
rect 13771 3009 13780 3043
rect 13728 3000 13780 3009
rect 3976 2932 4028 2984
rect 14096 2932 14148 2984
rect 14280 2932 14332 2984
rect 15108 2864 15160 2916
rect 16120 2932 16172 2984
rect 16304 2975 16356 2984
rect 16304 2941 16338 2975
rect 16338 2941 16356 2975
rect 16304 2932 16356 2941
rect 16580 2932 16632 2984
rect 17316 2932 17368 2984
rect 18604 2975 18656 2984
rect 18604 2941 18613 2975
rect 18613 2941 18647 2975
rect 18647 2941 18656 2975
rect 18604 2932 18656 2941
rect 12164 2796 12216 2848
rect 18328 2864 18380 2916
rect 19984 2932 20036 2984
rect 22008 2932 22060 2984
rect 22100 2975 22152 2984
rect 22100 2941 22109 2975
rect 22109 2941 22143 2975
rect 22143 2941 22152 2975
rect 22100 2932 22152 2941
rect 18696 2796 18748 2848
rect 19248 2796 19300 2848
rect 21180 2796 21232 2848
rect 8246 2694 8298 2746
rect 8310 2694 8362 2746
rect 8374 2694 8426 2746
rect 8438 2694 8490 2746
rect 15510 2694 15562 2746
rect 15574 2694 15626 2746
rect 15638 2694 15690 2746
rect 15702 2694 15754 2746
rect 13820 2592 13872 2644
rect 14556 2592 14608 2644
rect 16856 2635 16908 2644
rect 14648 2524 14700 2576
rect 15292 2524 15344 2576
rect 15936 2524 15988 2576
rect 16856 2601 16865 2635
rect 16865 2601 16899 2635
rect 16899 2601 16908 2635
rect 16856 2592 16908 2601
rect 18144 2592 18196 2644
rect 18696 2592 18748 2644
rect 17040 2524 17092 2576
rect 18328 2524 18380 2576
rect 19248 2524 19300 2576
rect 20720 2592 20772 2644
rect 15016 2456 15068 2508
rect 16120 2456 16172 2508
rect 21272 2456 21324 2508
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 17776 2431 17828 2440
rect 15108 2320 15160 2372
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 18328 2431 18380 2440
rect 18328 2397 18337 2431
rect 18337 2397 18371 2431
rect 18371 2397 18380 2431
rect 18328 2388 18380 2397
rect 20720 2388 20772 2440
rect 20076 2320 20128 2372
rect 16948 2252 17000 2304
rect 22100 2388 22152 2440
rect 4614 2150 4666 2202
rect 4678 2150 4730 2202
rect 4742 2150 4794 2202
rect 4806 2150 4858 2202
rect 11878 2150 11930 2202
rect 11942 2150 11994 2202
rect 12006 2150 12058 2202
rect 12070 2150 12122 2202
rect 19142 2150 19194 2202
rect 19206 2150 19258 2202
rect 19270 2150 19322 2202
rect 19334 2150 19386 2202
rect 13728 2048 13780 2100
rect 17776 2048 17828 2100
rect 20720 2048 20772 2100
<< metal2 >>
rect 294 23520 350 24000
rect 938 23520 994 24000
rect 1674 23520 1730 24000
rect 2410 23520 2466 24000
rect 3054 23520 3110 24000
rect 3790 23520 3846 24000
rect 4526 23520 4582 24000
rect 5170 23520 5226 24000
rect 5906 23520 5962 24000
rect 6642 23520 6698 24000
rect 7286 23520 7342 24000
rect 8022 23520 8078 24000
rect 8758 23520 8814 24000
rect 9402 23520 9458 24000
rect 10138 23520 10194 24000
rect 10874 23520 10930 24000
rect 11518 23520 11574 24000
rect 12254 23520 12310 24000
rect 12990 23520 13046 24000
rect 13634 23520 13690 24000
rect 14370 23520 14426 24000
rect 15106 23520 15162 24000
rect 15750 23520 15806 24000
rect 16486 23520 16542 24000
rect 17222 23520 17278 24000
rect 17866 23520 17922 24000
rect 18602 23520 18658 24000
rect 19338 23520 19394 24000
rect 19982 23520 20038 24000
rect 20718 23520 20774 24000
rect 21454 23520 21510 24000
rect 22098 23520 22154 24000
rect 22834 23520 22890 24000
rect 23570 23520 23626 24000
rect 308 21690 336 23520
rect 296 21684 348 21690
rect 296 21626 348 21632
rect 952 17338 980 23520
rect 1400 21480 1452 21486
rect 1398 21448 1400 21457
rect 1452 21448 1454 21457
rect 1398 21383 1454 21392
rect 1400 21344 1452 21350
rect 1400 21286 1452 21292
rect 1412 18834 1440 21286
rect 1492 20392 1544 20398
rect 1492 20334 1544 20340
rect 1504 19310 1532 20334
rect 1492 19304 1544 19310
rect 1492 19246 1544 19252
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1504 18766 1532 19246
rect 1492 18760 1544 18766
rect 1492 18702 1544 18708
rect 1582 18728 1638 18737
rect 1504 18222 1532 18702
rect 1582 18663 1638 18672
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1504 17678 1532 18158
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 940 17332 992 17338
rect 940 17274 992 17280
rect 1596 16658 1624 18663
rect 1688 16794 1716 23520
rect 2424 23474 2452 23520
rect 2332 23446 2452 23474
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 1952 20800 2004 20806
rect 1952 20742 2004 20748
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1780 18902 1808 19858
rect 1964 19854 1992 20742
rect 2148 20398 2176 20878
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1872 18222 1900 19790
rect 2332 19514 2360 23446
rect 2596 21344 2648 21350
rect 2596 21286 2648 21292
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 20058 2452 20198
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2412 19848 2464 19854
rect 2412 19790 2464 19796
rect 2320 19508 2372 19514
rect 2320 19450 2372 19456
rect 2424 19378 2452 19790
rect 2412 19372 2464 19378
rect 2412 19314 2464 19320
rect 2608 19292 2636 21286
rect 2780 21072 2832 21078
rect 2780 21014 2832 21020
rect 2792 20602 2820 21014
rect 2976 20602 3004 21286
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2964 20324 3016 20330
rect 2964 20266 3016 20272
rect 2778 19952 2834 19961
rect 2778 19887 2834 19896
rect 2872 19916 2924 19922
rect 2516 19264 2636 19292
rect 2228 18896 2280 18902
rect 2228 18838 2280 18844
rect 2240 18426 2268 18838
rect 2516 18834 2544 19264
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2516 18714 2544 18770
rect 2424 18686 2544 18714
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 1860 18216 1912 18222
rect 1766 18184 1822 18193
rect 1860 18158 1912 18164
rect 1766 18119 1822 18128
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 1400 16448 1452 16454
rect 1400 16390 1452 16396
rect 1412 16114 1440 16390
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15570 1716 15982
rect 1676 15564 1728 15570
rect 1676 15506 1728 15512
rect 1584 14952 1636 14958
rect 1688 14940 1716 15506
rect 1636 14912 1716 14940
rect 1584 14894 1636 14900
rect 1688 13841 1716 14912
rect 1674 13832 1730 13841
rect 1674 13767 1730 13776
rect 1688 13326 1716 13767
rect 1780 13394 1808 18119
rect 1872 17882 1900 18158
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 2136 17808 2188 17814
rect 2136 17750 2188 17756
rect 2148 17134 2176 17750
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2240 17338 2268 17682
rect 2320 17536 2372 17542
rect 2320 17478 2372 17484
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2228 17128 2280 17134
rect 2332 17116 2360 17478
rect 2280 17088 2360 17116
rect 2228 17070 2280 17076
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 1872 13530 1900 16662
rect 1952 15564 2004 15570
rect 1952 15506 2004 15512
rect 1964 14822 1992 15506
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14618 1992 14758
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2056 14414 2084 14826
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2148 14226 2176 16730
rect 2240 16658 2268 17070
rect 2228 16652 2280 16658
rect 2228 16594 2280 16600
rect 2056 14198 2176 14226
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1768 13388 1820 13394
rect 1768 13330 1820 13336
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12850 1716 13262
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1492 12300 1544 12306
rect 1492 12242 1544 12248
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 12102 1440 12174
rect 1400 12096 1452 12102
rect 1400 12038 1452 12044
rect 1412 11762 1440 12038
rect 1504 11937 1532 12242
rect 1490 11928 1546 11937
rect 1490 11863 1546 11872
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1596 11354 1624 12378
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1780 10606 1808 13126
rect 1860 11620 1912 11626
rect 1860 11562 1912 11568
rect 1872 11354 1900 11562
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1858 10024 1914 10033
rect 1858 9959 1860 9968
rect 1912 9959 1914 9968
rect 1860 9930 1912 9936
rect 2056 9518 2084 14198
rect 2136 13796 2188 13802
rect 2136 13738 2188 13744
rect 2148 12442 2176 13738
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 2148 11694 2176 12378
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2332 11218 2360 14214
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2424 10810 2452 18686
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2424 10062 2452 10406
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2424 9722 2452 9998
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9586 2544 16934
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2700 14414 2728 14554
rect 2792 14521 2820 19887
rect 2872 19858 2924 19864
rect 2884 18970 2912 19858
rect 2976 19854 3004 20266
rect 2964 19848 3016 19854
rect 2964 19790 3016 19796
rect 2976 19514 3004 19790
rect 3068 19514 3096 23520
rect 3804 22794 3832 23520
rect 4540 22794 4568 23520
rect 3804 22766 4108 22794
rect 3608 21616 3660 21622
rect 3608 21558 3660 21564
rect 3240 21548 3292 21554
rect 3240 21490 3292 21496
rect 3252 20058 3280 21490
rect 3332 21344 3384 21350
rect 3332 21286 3384 21292
rect 3240 20052 3292 20058
rect 3240 19994 3292 20000
rect 2964 19508 3016 19514
rect 2964 19450 3016 19456
rect 3056 19508 3108 19514
rect 3056 19450 3108 19456
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2976 15858 3004 19110
rect 3068 15978 3096 19246
rect 3240 19236 3292 19242
rect 3240 19178 3292 19184
rect 3148 19168 3200 19174
rect 3148 19110 3200 19116
rect 3160 16726 3188 19110
rect 3252 18970 3280 19178
rect 3240 18964 3292 18970
rect 3240 18906 3292 18912
rect 3252 18290 3280 18906
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3344 17882 3372 21286
rect 3620 21146 3648 21558
rect 3700 21548 3752 21554
rect 3700 21490 3752 21496
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3620 20330 3648 21082
rect 3712 21078 3740 21490
rect 3884 21480 3936 21486
rect 3884 21422 3936 21428
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3896 20806 3924 21422
rect 3884 20800 3936 20806
rect 3884 20742 3936 20748
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3608 20324 3660 20330
rect 3608 20266 3660 20272
rect 3424 19916 3476 19922
rect 3424 19858 3476 19864
rect 3608 19916 3660 19922
rect 3608 19858 3660 19864
rect 3436 18426 3464 19858
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3528 17746 3556 19654
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3620 17338 3648 19858
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3712 17134 3740 19790
rect 3804 17134 3832 20538
rect 3700 17128 3752 17134
rect 3700 17070 3752 17076
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3160 16250 3188 16662
rect 3712 16522 3740 17070
rect 3700 16516 3752 16522
rect 3700 16458 3752 16464
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3896 16130 3924 20742
rect 4080 20602 4108 22766
rect 4448 22766 4568 22794
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 4172 20262 4200 21422
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4264 20602 4292 20878
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4252 19984 4304 19990
rect 4252 19926 4304 19932
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4080 19378 4108 19751
rect 4160 19508 4212 19514
rect 4160 19450 4212 19456
rect 4068 19372 4120 19378
rect 4068 19314 4120 19320
rect 3974 17912 4030 17921
rect 3974 17847 4030 17856
rect 3988 17814 4016 17847
rect 3976 17808 4028 17814
rect 3976 17750 4028 17756
rect 4080 17626 4108 19314
rect 3160 16102 3924 16130
rect 3988 17598 4108 17626
rect 3988 16114 4016 17598
rect 4068 17536 4120 17542
rect 4068 17478 4120 17484
rect 4080 16794 4108 17478
rect 4068 16788 4120 16794
rect 4068 16730 4120 16736
rect 3976 16108 4028 16114
rect 3056 15972 3108 15978
rect 3056 15914 3108 15920
rect 2884 15830 3004 15858
rect 2778 14512 2834 14521
rect 2778 14447 2834 14456
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2700 13938 2728 14350
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2780 13728 2832 13734
rect 2780 13670 2832 13676
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2700 11354 2728 13466
rect 2792 12714 2820 13670
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 11898 2820 12650
rect 2780 11892 2832 11898
rect 2780 11834 2832 11840
rect 2884 11354 2912 15830
rect 3068 15706 3096 15914
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2976 13530 3004 14418
rect 3056 14408 3108 14414
rect 3056 14350 3108 14356
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 3068 13462 3096 14350
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3068 12986 3096 13398
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2688 11144 2740 11150
rect 2688 11086 2740 11092
rect 2596 10532 2648 10538
rect 2596 10474 2648 10480
rect 2608 10062 2636 10474
rect 2700 10062 2728 11086
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 2596 10056 2648 10062
rect 2596 9998 2648 10004
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2884 9926 2912 10610
rect 2976 10606 3004 12378
rect 3054 12336 3110 12345
rect 3054 12271 3056 12280
rect 3108 12271 3110 12280
rect 3056 12242 3108 12248
rect 3160 10674 3188 16102
rect 3976 16050 4028 16056
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3516 15564 3568 15570
rect 3516 15506 3568 15512
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3252 14414 3280 14554
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3240 14000 3292 14006
rect 3292 13948 3372 13954
rect 3240 13942 3372 13948
rect 3252 13926 3372 13942
rect 3240 13864 3292 13870
rect 3238 13832 3240 13841
rect 3292 13832 3294 13841
rect 3238 13767 3294 13776
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3252 11898 3280 13670
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3344 11762 3372 13926
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3436 11694 3464 14214
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 2964 10600 3016 10606
rect 2964 10542 3016 10548
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2686 9616 2742 9625
rect 2504 9580 2556 9586
rect 2686 9551 2688 9560
rect 2504 9522 2556 9528
rect 2740 9551 2742 9560
rect 2688 9522 2740 9528
rect 1584 9512 1636 9518
rect 1582 9480 1584 9489
rect 2044 9512 2096 9518
rect 1636 9480 1638 9489
rect 2044 9454 2096 9460
rect 1582 9415 1638 9424
rect 3068 9382 3096 10066
rect 3436 9518 3464 11018
rect 3528 10810 3556 15506
rect 3620 15026 3648 15982
rect 3700 15972 3752 15978
rect 3700 15914 3752 15920
rect 3712 15162 3740 15914
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3620 14618 3648 14962
rect 3700 14816 3752 14822
rect 3700 14758 3752 14764
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3712 14550 3740 14758
rect 3700 14544 3752 14550
rect 3700 14486 3752 14492
rect 3700 14408 3752 14414
rect 3700 14350 3752 14356
rect 3712 14278 3740 14350
rect 3700 14272 3752 14278
rect 3700 14214 3752 14220
rect 3712 14113 3740 14214
rect 3698 14104 3754 14113
rect 3608 14068 3660 14074
rect 3698 14039 3754 14048
rect 3608 14010 3660 14016
rect 3620 13954 3648 14010
rect 3620 13926 3740 13954
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3620 12782 3648 13466
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 3606 12200 3662 12209
rect 3606 12135 3662 12144
rect 3516 10804 3568 10810
rect 3516 10746 3568 10752
rect 3424 9512 3476 9518
rect 3424 9454 3476 9460
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2502 9208 2558 9217
rect 2502 9143 2504 9152
rect 2556 9143 2558 9152
rect 2504 9114 2556 9120
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2056 8430 2084 8910
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8498 3004 8774
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 3068 6390 3096 9318
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 3528 3670 3556 9318
rect 3620 4049 3648 12135
rect 3712 10606 3740 13926
rect 3804 10674 3832 15030
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 3896 10606 3924 15846
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3700 10600 3752 10606
rect 3700 10542 3752 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3988 10470 4016 15302
rect 4080 14890 4108 15846
rect 4172 15706 4200 19450
rect 4264 18970 4292 19926
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4356 18850 4384 21626
rect 4448 20330 4476 22766
rect 4588 21788 4884 21808
rect 4644 21786 4668 21788
rect 4724 21786 4748 21788
rect 4804 21786 4828 21788
rect 4666 21734 4668 21786
rect 4730 21734 4742 21786
rect 4804 21734 4806 21786
rect 4644 21732 4668 21734
rect 4724 21732 4748 21734
rect 4804 21732 4828 21734
rect 4588 21712 4884 21732
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 4896 21480 4948 21486
rect 4896 21422 4948 21428
rect 4908 20924 4936 21422
rect 5000 21026 5028 21558
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 5092 21146 5120 21286
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5000 20998 5120 21026
rect 4988 20936 5040 20942
rect 4908 20896 4988 20924
rect 4988 20878 5040 20884
rect 4588 20700 4884 20720
rect 4644 20698 4668 20700
rect 4724 20698 4748 20700
rect 4804 20698 4828 20700
rect 4666 20646 4668 20698
rect 4730 20646 4742 20698
rect 4804 20646 4806 20698
rect 4644 20644 4668 20646
rect 4724 20644 4748 20646
rect 4804 20644 4828 20646
rect 4588 20624 4884 20644
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4436 20324 4488 20330
rect 4436 20266 4488 20272
rect 4816 19990 4844 20470
rect 4896 20392 4948 20398
rect 5000 20380 5028 20878
rect 4948 20352 5028 20380
rect 4896 20334 4948 20340
rect 4804 19984 4856 19990
rect 4804 19926 4856 19932
rect 4620 19848 4672 19854
rect 4618 19816 4620 19825
rect 4672 19816 4674 19825
rect 4618 19751 4674 19760
rect 5000 19700 5028 20352
rect 5092 19854 5120 20998
rect 5080 19848 5132 19854
rect 5080 19790 5132 19796
rect 5000 19672 5120 19700
rect 4588 19612 4884 19632
rect 4644 19610 4668 19612
rect 4724 19610 4748 19612
rect 4804 19610 4828 19612
rect 4666 19558 4668 19610
rect 4730 19558 4742 19610
rect 4804 19558 4806 19610
rect 4644 19556 4668 19558
rect 4724 19556 4748 19558
rect 4804 19556 4828 19558
rect 4588 19536 4884 19556
rect 4986 19544 5042 19553
rect 4436 19508 4488 19514
rect 4986 19479 4988 19488
rect 4436 19450 4488 19456
rect 5040 19479 5042 19488
rect 4988 19450 5040 19456
rect 4264 18822 4384 18850
rect 4264 16794 4292 18822
rect 4344 18624 4396 18630
rect 4344 18566 4396 18572
rect 4356 18222 4384 18566
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4344 18080 4396 18086
rect 4344 18022 4396 18028
rect 4356 17202 4384 18022
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4448 16998 4476 19450
rect 5000 19378 5028 19450
rect 5092 19394 5120 19672
rect 5184 19514 5212 23520
rect 5264 21344 5316 21350
rect 5264 21286 5316 21292
rect 5276 19718 5304 21286
rect 5356 20800 5408 20806
rect 5356 20742 5408 20748
rect 5368 20398 5396 20742
rect 5538 20632 5594 20641
rect 5920 20602 5948 23520
rect 6656 21486 6684 23520
rect 7300 22794 7328 23520
rect 6932 22766 7328 22794
rect 6828 21548 6880 21554
rect 6828 21490 6880 21496
rect 6644 21480 6696 21486
rect 6644 21422 6696 21428
rect 6184 21004 6236 21010
rect 6184 20946 6236 20952
rect 5538 20567 5594 20576
rect 5908 20596 5960 20602
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 5448 20392 5500 20398
rect 5448 20334 5500 20340
rect 5368 20262 5396 20334
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 4988 19372 5040 19378
rect 5092 19366 5212 19394
rect 4988 19314 5040 19320
rect 4528 19304 4580 19310
rect 4526 19272 4528 19281
rect 4580 19272 4582 19281
rect 4526 19207 4582 19216
rect 5184 18970 5212 19366
rect 5276 19310 5304 19654
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5368 19145 5396 19790
rect 5354 19136 5410 19145
rect 5354 19071 5410 19080
rect 5460 18986 5488 20334
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5368 18958 5488 18986
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 4588 18524 4884 18544
rect 4644 18522 4668 18524
rect 4724 18522 4748 18524
rect 4804 18522 4828 18524
rect 4666 18470 4668 18522
rect 4730 18470 4742 18522
rect 4804 18470 4806 18522
rect 4644 18468 4668 18470
rect 4724 18468 4748 18470
rect 4804 18468 4828 18470
rect 4588 18448 4884 18468
rect 4588 17436 4884 17456
rect 4644 17434 4668 17436
rect 4724 17434 4748 17436
rect 4804 17434 4828 17436
rect 4666 17382 4668 17434
rect 4730 17382 4742 17434
rect 4804 17382 4806 17434
rect 4644 17380 4668 17382
rect 4724 17380 4748 17382
rect 4804 17380 4828 17382
rect 4588 17360 4884 17380
rect 4618 17232 4674 17241
rect 4618 17167 4674 17176
rect 4632 17134 4660 17167
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 5000 16810 5028 18702
rect 5184 18154 5212 18906
rect 5368 18630 5396 18958
rect 5448 18896 5500 18902
rect 5448 18838 5500 18844
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4908 16794 5028 16810
rect 4252 16788 4304 16794
rect 4252 16730 4304 16736
rect 4896 16788 5028 16794
rect 4948 16782 5028 16788
rect 4896 16730 4948 16736
rect 4588 16348 4884 16368
rect 4644 16346 4668 16348
rect 4724 16346 4748 16348
rect 4804 16346 4828 16348
rect 4666 16294 4668 16346
rect 4730 16294 4742 16346
rect 4804 16294 4806 16346
rect 4644 16292 4668 16294
rect 4724 16292 4748 16294
rect 4804 16292 4828 16294
rect 4588 16272 4884 16292
rect 4436 16040 4488 16046
rect 4436 15982 4488 15988
rect 4160 15700 4212 15706
rect 4160 15642 4212 15648
rect 4448 14958 4476 15982
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15570 4844 15846
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4588 15260 4884 15280
rect 4644 15258 4668 15260
rect 4724 15258 4748 15260
rect 4804 15258 4828 15260
rect 4666 15206 4668 15258
rect 4730 15206 4742 15258
rect 4804 15206 4806 15258
rect 4644 15204 4668 15206
rect 4724 15204 4748 15206
rect 4804 15204 4828 15206
rect 4588 15184 4884 15204
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4160 14952 4212 14958
rect 4160 14894 4212 14900
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 4080 14618 4108 14826
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4066 14512 4122 14521
rect 4066 14447 4122 14456
rect 4080 12714 4108 14447
rect 4172 14113 4200 14894
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4158 14104 4214 14113
rect 4158 14039 4160 14048
rect 4212 14039 4214 14048
rect 4160 14010 4212 14016
rect 4172 13979 4200 14010
rect 4264 13870 4292 14758
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4264 13530 4292 13806
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4356 13410 4384 14758
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4448 14074 4476 14486
rect 4588 14172 4884 14192
rect 4644 14170 4668 14172
rect 4724 14170 4748 14172
rect 4804 14170 4828 14172
rect 4666 14118 4668 14170
rect 4730 14118 4742 14170
rect 4804 14118 4806 14170
rect 4644 14116 4668 14118
rect 4724 14116 4748 14118
rect 4804 14116 4828 14118
rect 4588 14096 4884 14116
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 5000 13870 5028 15098
rect 5092 14362 5120 18022
rect 5184 17882 5212 18090
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5356 17808 5408 17814
rect 5356 17750 5408 17756
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 16590 5212 17682
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 5276 16726 5304 17138
rect 5264 16720 5316 16726
rect 5264 16662 5316 16668
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5184 16232 5212 16526
rect 5264 16244 5316 16250
rect 5184 16204 5264 16232
rect 5264 16186 5316 16192
rect 5368 16130 5396 17750
rect 5276 16102 5396 16130
rect 5276 15910 5304 16102
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5264 15904 5316 15910
rect 5264 15846 5316 15852
rect 5092 14334 5212 14362
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5092 14074 5120 14214
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5184 13954 5212 14334
rect 5092 13926 5212 13954
rect 4988 13864 5040 13870
rect 4988 13806 5040 13812
rect 4896 13796 4948 13802
rect 4896 13738 4948 13744
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4172 13382 4384 13410
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4172 12442 4200 13382
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12986 4292 13262
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4448 12764 4476 13670
rect 4526 13560 4582 13569
rect 4526 13495 4528 13504
rect 4580 13495 4582 13504
rect 4528 13466 4580 13472
rect 4908 13326 4936 13738
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4588 13084 4884 13104
rect 4644 13082 4668 13084
rect 4724 13082 4748 13084
rect 4804 13082 4828 13084
rect 4666 13030 4668 13082
rect 4730 13030 4742 13082
rect 4804 13030 4806 13082
rect 4644 13028 4668 13030
rect 4724 13028 4748 13030
rect 4804 13028 4828 13030
rect 4588 13008 4884 13028
rect 4356 12736 4476 12764
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4356 12306 4384 12736
rect 4988 12640 5040 12646
rect 4988 12582 5040 12588
rect 5000 12306 5028 12582
rect 4344 12300 4396 12306
rect 4344 12242 4396 12248
rect 4988 12300 5040 12306
rect 4988 12242 5040 12248
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 4066 11792 4122 11801
rect 4066 11727 4068 11736
rect 4120 11727 4122 11736
rect 4068 11698 4120 11704
rect 4172 11200 4200 11834
rect 4356 11830 4384 12106
rect 4588 11996 4884 12016
rect 4644 11994 4668 11996
rect 4724 11994 4748 11996
rect 4804 11994 4828 11996
rect 4666 11942 4668 11994
rect 4730 11942 4742 11994
rect 4804 11942 4806 11994
rect 4644 11940 4668 11942
rect 4724 11940 4748 11942
rect 4804 11940 4828 11942
rect 4588 11920 4884 11940
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4436 11756 4488 11762
rect 4436 11698 4488 11704
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4252 11688 4304 11694
rect 4252 11630 4304 11636
rect 4080 11172 4200 11200
rect 3976 10464 4028 10470
rect 3976 10406 4028 10412
rect 3882 10160 3938 10169
rect 3882 10095 3938 10104
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 9586 3740 9862
rect 3804 9586 3832 9998
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3712 9382 3740 9522
rect 3700 9376 3752 9382
rect 3700 9318 3752 9324
rect 3896 9110 3924 10095
rect 4080 9994 4108 11172
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4172 9518 4200 11018
rect 4264 10266 4292 11630
rect 4342 11248 4398 11257
rect 4342 11183 4344 11192
rect 4396 11183 4398 11192
rect 4344 11154 4396 11160
rect 4448 11150 4476 11698
rect 4724 11218 4752 11698
rect 4802 11656 4858 11665
rect 4802 11591 4804 11600
rect 4856 11591 4858 11600
rect 4804 11562 4856 11568
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 11393 4936 11494
rect 4894 11384 4950 11393
rect 4894 11319 4950 11328
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4436 11144 4488 11150
rect 4342 11112 4398 11121
rect 4436 11086 4488 11092
rect 4342 11047 4398 11056
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4356 9738 4384 11047
rect 4448 10674 4476 11086
rect 4588 10908 4884 10928
rect 4644 10906 4668 10908
rect 4724 10906 4748 10908
rect 4804 10906 4828 10908
rect 4666 10854 4668 10906
rect 4730 10854 4742 10906
rect 4804 10854 4806 10906
rect 4644 10852 4668 10854
rect 4724 10852 4748 10854
rect 4804 10852 4828 10854
rect 4588 10832 4884 10852
rect 4526 10704 4582 10713
rect 4436 10668 4488 10674
rect 4526 10639 4582 10648
rect 4436 10610 4488 10616
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4448 10130 4476 10406
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4540 10010 4568 10639
rect 4894 10296 4950 10305
rect 4894 10231 4950 10240
rect 4908 10198 4936 10231
rect 5000 10198 5028 12242
rect 5092 11121 5120 13926
rect 5368 13734 5396 15982
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5184 12782 5212 13262
rect 5356 13184 5408 13190
rect 5356 13126 5408 13132
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5172 12776 5224 12782
rect 5172 12718 5224 12724
rect 5276 12442 5304 12922
rect 5368 12782 5396 13126
rect 5356 12776 5408 12782
rect 5356 12718 5408 12724
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11354 5212 11494
rect 5172 11348 5224 11354
rect 5172 11290 5224 11296
rect 5264 11348 5316 11354
rect 5264 11290 5316 11296
rect 5078 11112 5134 11121
rect 5078 11047 5134 11056
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5092 10606 5120 10950
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10470 5120 10542
rect 5184 10538 5212 10950
rect 5276 10538 5304 11290
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5264 10532 5316 10538
rect 5264 10474 5316 10480
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 5170 10432 5226 10441
rect 4896 10192 4948 10198
rect 4896 10134 4948 10140
rect 4988 10192 5040 10198
rect 4988 10134 5040 10140
rect 4264 9710 4384 9738
rect 4448 9982 4568 10010
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4068 9376 4120 9382
rect 3974 9344 4030 9353
rect 4068 9318 4120 9324
rect 3974 9279 4030 9288
rect 3884 9104 3936 9110
rect 3698 9072 3754 9081
rect 3884 9046 3936 9052
rect 3698 9007 3700 9016
rect 3752 9007 3754 9016
rect 3700 8978 3752 8984
rect 3988 8514 4016 9279
rect 4080 9110 4108 9318
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 4066 8936 4122 8945
rect 4066 8871 4122 8880
rect 4080 8634 4108 8871
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3988 8486 4108 8514
rect 4080 8430 4108 8486
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4264 8362 4292 9710
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4250 7304 4306 7313
rect 4250 7239 4252 7248
rect 4304 7239 4306 7248
rect 4252 7210 4304 7216
rect 4356 6798 4384 9590
rect 4448 9178 4476 9982
rect 4588 9820 4884 9840
rect 4644 9818 4668 9820
rect 4724 9818 4748 9820
rect 4804 9818 4828 9820
rect 4666 9766 4668 9818
rect 4730 9766 4742 9818
rect 4804 9766 4806 9818
rect 4644 9764 4668 9766
rect 4724 9764 4748 9766
rect 4804 9764 4828 9766
rect 4588 9744 4884 9764
rect 5092 9586 5120 10406
rect 5170 10367 5226 10376
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9512 5040 9518
rect 5184 9489 5212 10367
rect 4988 9454 5040 9460
rect 5170 9480 5226 9489
rect 5000 9194 5028 9454
rect 5170 9415 5226 9424
rect 5276 9382 5304 10474
rect 5368 10266 5396 12718
rect 5460 10577 5488 18838
rect 5552 17921 5580 20567
rect 5908 20538 5960 20544
rect 6196 20262 6224 20946
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6184 20256 6236 20262
rect 6184 20198 6236 20204
rect 6196 20058 6224 20198
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6092 19984 6144 19990
rect 6092 19926 6144 19932
rect 6104 19378 6132 19926
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 5724 18760 5776 18766
rect 5724 18702 5776 18708
rect 5736 18154 5764 18702
rect 5724 18148 5776 18154
rect 5724 18090 5776 18096
rect 5538 17912 5594 17921
rect 5736 17882 5764 18090
rect 5538 17847 5594 17856
rect 5724 17876 5776 17882
rect 5724 17818 5776 17824
rect 5908 17740 5960 17746
rect 5908 17682 5960 17688
rect 5724 16176 5776 16182
rect 5724 16118 5776 16124
rect 5736 12986 5764 16118
rect 5920 14006 5948 17682
rect 6000 16652 6052 16658
rect 6000 16594 6052 16600
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5446 10568 5502 10577
rect 5446 10503 5502 10512
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5460 10266 5488 10406
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5448 10260 5500 10266
rect 5448 10202 5500 10208
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 5368 9761 5396 9862
rect 5354 9752 5410 9761
rect 5354 9687 5410 9696
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4436 9172 4488 9178
rect 5000 9166 5304 9194
rect 5368 9178 5396 9318
rect 4436 9114 4488 9120
rect 5276 8974 5304 9166
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 8974 5488 9998
rect 5552 9178 5580 12242
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 6012 12186 6040 16594
rect 6104 14618 6132 18770
rect 6196 17882 6224 19450
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 6196 15978 6224 16526
rect 6288 16114 6316 20878
rect 6644 20800 6696 20806
rect 6644 20742 6696 20748
rect 6656 20641 6684 20742
rect 6642 20632 6698 20641
rect 6642 20567 6698 20576
rect 6656 19961 6684 20567
rect 6840 20466 6868 21490
rect 6932 21010 6960 22766
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 7944 21078 7972 21490
rect 7932 21072 7984 21078
rect 7932 21014 7984 21020
rect 6920 21004 6972 21010
rect 6920 20946 6972 20952
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 6828 20460 6880 20466
rect 6828 20402 6880 20408
rect 7116 20398 7144 20946
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6642 19952 6698 19961
rect 6642 19887 6698 19896
rect 6552 19848 6604 19854
rect 6552 19790 6604 19796
rect 6736 19848 6788 19854
rect 7104 19848 7156 19854
rect 6788 19808 6868 19836
rect 6736 19790 6788 19796
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6380 17134 6408 19450
rect 6564 19394 6592 19790
rect 6734 19408 6790 19417
rect 6564 19366 6734 19394
rect 6734 19343 6790 19352
rect 6748 19281 6776 19343
rect 6840 19310 6868 19808
rect 7102 19816 7104 19825
rect 7156 19816 7158 19825
rect 7102 19751 7158 19760
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 6828 19304 6880 19310
rect 6734 19272 6790 19281
rect 6828 19246 6880 19252
rect 6734 19207 6790 19216
rect 6644 19168 6696 19174
rect 6644 19110 6696 19116
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6460 18896 6512 18902
rect 6460 18838 6512 18844
rect 6472 18426 6500 18838
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6564 18290 6592 18906
rect 6656 18737 6684 19110
rect 6748 18834 6776 19207
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6642 18728 6698 18737
rect 6698 18686 6776 18714
rect 6642 18663 6698 18672
rect 6748 18426 6776 18686
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6460 17740 6512 17746
rect 6460 17682 6512 17688
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 6472 17649 6500 17682
rect 6458 17640 6514 17649
rect 6458 17575 6514 17584
rect 6564 17241 6592 17682
rect 6550 17232 6606 17241
rect 6656 17202 6684 18294
rect 6736 18216 6788 18222
rect 6736 18158 6788 18164
rect 6550 17167 6606 17176
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6368 17128 6420 17134
rect 6552 17128 6604 17134
rect 6368 17070 6420 17076
rect 6458 17096 6514 17105
rect 6552 17070 6604 17076
rect 6458 17031 6514 17040
rect 6368 16652 6420 16658
rect 6368 16594 6420 16600
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6380 15994 6408 16594
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6288 15966 6408 15994
rect 6196 15706 6224 15914
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15484 6316 15966
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6196 15456 6316 15484
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 6104 12442 6132 14418
rect 6196 13818 6224 15456
rect 6380 14958 6408 15846
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6288 13938 6316 14214
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6196 13790 6316 13818
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6182 12336 6238 12345
rect 6182 12271 6238 12280
rect 5632 11620 5684 11626
rect 5632 11562 5684 11568
rect 5644 11529 5672 11562
rect 5630 11520 5686 11529
rect 5630 11455 5686 11464
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5644 9518 5672 10406
rect 5736 9994 5764 12174
rect 5816 12164 5868 12170
rect 6012 12158 6132 12186
rect 5816 12106 5868 12112
rect 5828 11898 5856 12106
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5828 11665 5856 11698
rect 5814 11656 5870 11665
rect 5814 11591 5870 11600
rect 5908 11552 5960 11558
rect 6012 11529 6040 12038
rect 5908 11494 5960 11500
rect 5998 11520 6054 11529
rect 5920 11218 5948 11494
rect 5998 11455 6054 11464
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5724 9988 5776 9994
rect 5724 9930 5776 9936
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 5080 8968 5132 8974
rect 5264 8968 5316 8974
rect 5132 8945 5212 8956
rect 5132 8936 5226 8945
rect 5132 8928 5170 8936
rect 5080 8910 5132 8916
rect 5264 8910 5316 8916
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5170 8871 5226 8880
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5080 8832 5132 8838
rect 5368 8786 5396 8842
rect 5132 8780 5396 8786
rect 5080 8774 5396 8780
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 5092 8758 5396 8774
rect 4588 8732 4884 8752
rect 4644 8730 4668 8732
rect 4724 8730 4748 8732
rect 4804 8730 4828 8732
rect 4666 8678 4668 8730
rect 4730 8678 4742 8730
rect 4804 8678 4806 8730
rect 4644 8676 4668 8678
rect 4724 8676 4748 8678
rect 4804 8676 4828 8678
rect 4588 8656 4884 8676
rect 5354 8664 5410 8673
rect 5354 8599 5410 8608
rect 5078 8528 5134 8537
rect 5368 8498 5396 8599
rect 5460 8566 5488 8774
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 5078 8463 5134 8472
rect 5356 8492 5408 8498
rect 5092 8430 5120 8463
rect 5356 8434 5408 8440
rect 5080 8424 5132 8430
rect 5080 8366 5132 8372
rect 5736 8294 5764 9454
rect 5828 9217 5856 10542
rect 5814 9208 5870 9217
rect 5920 9178 5948 11154
rect 6012 9178 6040 11455
rect 6104 10606 6132 12158
rect 6196 11898 6224 12271
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6182 11384 6238 11393
rect 6182 11319 6238 11328
rect 6196 11082 6224 11319
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 5814 9143 5870 9152
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6000 8968 6052 8974
rect 6000 8910 6052 8916
rect 6012 8566 6040 8910
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 6104 8430 6132 9862
rect 6196 9382 6224 10066
rect 6288 9518 6316 13790
rect 6276 9512 6328 9518
rect 6276 9454 6328 9460
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6196 8362 6224 9318
rect 6276 8832 6328 8838
rect 6380 8820 6408 13942
rect 6328 8792 6408 8820
rect 6276 8774 6328 8780
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 5724 8288 5776 8294
rect 5262 8256 5318 8265
rect 5724 8230 5776 8236
rect 5262 8191 5318 8200
rect 5276 8090 5304 8191
rect 5920 8090 5948 8298
rect 5264 8084 5316 8090
rect 5264 8026 5316 8032
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 4436 7880 4488 7886
rect 4434 7848 4436 7857
rect 4488 7848 4490 7857
rect 4434 7783 4490 7792
rect 4588 7644 4884 7664
rect 4644 7642 4668 7644
rect 4724 7642 4748 7644
rect 4804 7642 4828 7644
rect 4666 7590 4668 7642
rect 4730 7590 4742 7642
rect 4804 7590 4806 7642
rect 4644 7588 4668 7590
rect 4724 7588 4748 7590
rect 4804 7588 4828 7590
rect 4588 7568 4884 7588
rect 5276 7274 5304 8026
rect 5446 7984 5502 7993
rect 5446 7919 5502 7928
rect 6276 7948 6328 7954
rect 5460 7886 5488 7919
rect 6276 7890 6328 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6196 7410 6224 7686
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 7041 4752 7142
rect 4710 7032 4766 7041
rect 4710 6967 4766 6976
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4588 6556 4884 6576
rect 4644 6554 4668 6556
rect 4724 6554 4748 6556
rect 4804 6554 4828 6556
rect 4666 6502 4668 6554
rect 4730 6502 4742 6554
rect 4804 6502 4806 6554
rect 4644 6500 4668 6502
rect 4724 6500 4748 6502
rect 4804 6500 4828 6502
rect 4588 6480 4884 6500
rect 6288 5914 6316 7890
rect 6472 7886 6500 17031
rect 6564 16697 6592 17070
rect 6748 17066 6776 18158
rect 6840 17746 6868 19246
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17060 6788 17066
rect 6736 17002 6788 17008
rect 6840 16998 6868 17682
rect 6932 16998 6960 19314
rect 7380 19236 7432 19242
rect 7380 19178 7432 19184
rect 7012 18828 7064 18834
rect 7012 18770 7064 18776
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7024 17882 7052 18770
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7208 17678 7236 18770
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7208 17513 7236 17614
rect 7194 17504 7250 17513
rect 7194 17439 7250 17448
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6920 16992 6972 16998
rect 6920 16934 6972 16940
rect 6550 16688 6606 16697
rect 6550 16623 6552 16632
rect 6604 16623 6606 16632
rect 6736 16652 6788 16658
rect 6552 16594 6604 16600
rect 7024 16640 7052 17070
rect 6788 16612 7052 16640
rect 6736 16594 6788 16600
rect 6564 16563 6592 16594
rect 6552 16448 6604 16454
rect 6550 16416 6552 16425
rect 6644 16448 6696 16454
rect 6604 16416 6606 16425
rect 6644 16390 6696 16396
rect 6550 16351 6606 16360
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6564 10266 6592 13806
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6550 9616 6606 9625
rect 6550 9551 6606 9560
rect 6564 9178 6592 9551
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6550 9072 6606 9081
rect 6550 9007 6606 9016
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6366 7576 6422 7585
rect 6366 7511 6422 7520
rect 6380 7410 6408 7511
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6564 6730 6592 9007
rect 6656 8090 6684 16390
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6644 8084 6696 8090
rect 6644 8026 6696 8032
rect 6748 7546 6776 16186
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6840 15706 6868 16050
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6932 15162 6960 15914
rect 7196 15904 7248 15910
rect 7196 15846 7248 15852
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 7116 15026 7144 15438
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 14074 6868 14826
rect 7116 14498 7144 14962
rect 7208 14618 7236 15846
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7024 14470 7144 14498
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6840 13394 6868 14010
rect 7024 14006 7052 14470
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6932 13530 6960 13738
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6828 13388 6880 13394
rect 6828 13330 6880 13336
rect 7024 12986 7052 13670
rect 7116 13258 7144 14350
rect 7104 13252 7156 13258
rect 7104 13194 7156 13200
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 7208 12866 7236 14554
rect 7300 14414 7328 17818
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13394 7328 14214
rect 7288 13388 7340 13394
rect 7288 13330 7340 13336
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 7024 12838 7236 12866
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6840 11354 6868 12718
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6840 9042 6868 10406
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6840 6202 6868 8842
rect 6932 8634 6960 11154
rect 7024 10606 7052 12838
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11694 7144 12038
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 7116 9110 7144 11154
rect 7208 11150 7236 12174
rect 7300 11898 7328 13194
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7392 11370 7420 19178
rect 7576 18630 7604 19314
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7576 18222 7604 18566
rect 7564 18216 7616 18222
rect 7564 18158 7616 18164
rect 7760 18154 7788 20946
rect 8036 20602 8064 23520
rect 8668 21956 8720 21962
rect 8668 21898 8720 21904
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 8128 21350 8156 21626
rect 8576 21480 8628 21486
rect 8680 21457 8708 21898
rect 8576 21422 8628 21428
rect 8666 21448 8722 21457
rect 8116 21344 8168 21350
rect 8116 21286 8168 21292
rect 8128 20602 8156 21286
rect 8220 21244 8516 21264
rect 8276 21242 8300 21244
rect 8356 21242 8380 21244
rect 8436 21242 8460 21244
rect 8298 21190 8300 21242
rect 8362 21190 8374 21242
rect 8436 21190 8438 21242
rect 8276 21188 8300 21190
rect 8356 21188 8380 21190
rect 8436 21188 8460 21190
rect 8220 21168 8516 21188
rect 8588 21146 8616 21422
rect 8666 21383 8722 21392
rect 8680 21350 8708 21383
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8576 21140 8628 21146
rect 8576 21082 8628 21088
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8588 20398 8616 20742
rect 8576 20392 8628 20398
rect 8576 20334 8628 20340
rect 8668 20256 8720 20262
rect 8668 20198 8720 20204
rect 8220 20156 8516 20176
rect 8276 20154 8300 20156
rect 8356 20154 8380 20156
rect 8436 20154 8460 20156
rect 8298 20102 8300 20154
rect 8362 20102 8374 20154
rect 8436 20102 8438 20154
rect 8276 20100 8300 20102
rect 8356 20100 8380 20102
rect 8436 20100 8460 20102
rect 8220 20080 8516 20100
rect 8680 19922 8708 20198
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8668 19712 8720 19718
rect 8668 19654 8720 19660
rect 8680 19514 8708 19654
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8206 19408 8262 19417
rect 8206 19343 8262 19352
rect 8576 19372 8628 19378
rect 8220 19310 8248 19343
rect 8576 19314 8628 19320
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7852 18970 7880 19110
rect 8128 18970 8156 19178
rect 8220 19068 8516 19088
rect 8276 19066 8300 19068
rect 8356 19066 8380 19068
rect 8436 19066 8460 19068
rect 8298 19014 8300 19066
rect 8362 19014 8374 19066
rect 8436 19014 8438 19066
rect 8276 19012 8300 19014
rect 8356 19012 8380 19014
rect 8436 19012 8460 19014
rect 8220 18992 8516 19012
rect 8588 18970 8616 19314
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7484 17270 7512 17614
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7760 15688 7788 18090
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7840 17672 7892 17678
rect 7838 17640 7840 17649
rect 7892 17640 7894 17649
rect 7838 17575 7894 17584
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 7840 16720 7892 16726
rect 7840 16662 7892 16668
rect 7852 16250 7880 16662
rect 8036 16522 8064 17070
rect 8128 16590 8156 18022
rect 8220 17980 8516 18000
rect 8276 17978 8300 17980
rect 8356 17978 8380 17980
rect 8436 17978 8460 17980
rect 8298 17926 8300 17978
rect 8362 17926 8374 17978
rect 8436 17926 8438 17978
rect 8276 17924 8300 17926
rect 8356 17924 8380 17926
rect 8436 17924 8460 17926
rect 8220 17904 8516 17924
rect 8588 17542 8616 18770
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8220 16892 8516 16912
rect 8276 16890 8300 16892
rect 8356 16890 8380 16892
rect 8436 16890 8460 16892
rect 8298 16838 8300 16890
rect 8362 16838 8374 16890
rect 8436 16838 8438 16890
rect 8276 16836 8300 16838
rect 8356 16836 8380 16838
rect 8436 16836 8460 16838
rect 8220 16816 8516 16836
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8588 16522 8616 16934
rect 8680 16726 8708 19450
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7944 16250 7972 16390
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 8668 16108 8720 16114
rect 8668 16050 8720 16056
rect 8220 15804 8516 15824
rect 8276 15802 8300 15804
rect 8356 15802 8380 15804
rect 8436 15802 8460 15804
rect 8298 15750 8300 15802
rect 8362 15750 8374 15802
rect 8436 15750 8438 15802
rect 8276 15748 8300 15750
rect 8356 15748 8380 15750
rect 8436 15748 8460 15750
rect 8220 15728 8516 15748
rect 7760 15660 7880 15688
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14618 7512 14758
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7484 13530 7512 14418
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7576 13938 7604 14350
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7760 13870 7788 14214
rect 7748 13864 7800 13870
rect 7748 13806 7800 13812
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7760 12850 7788 13262
rect 7748 12844 7800 12850
rect 7668 12804 7748 12832
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7576 12345 7604 12718
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7300 11342 7420 11370
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7194 10976 7250 10985
rect 7194 10911 7250 10920
rect 7208 10810 7236 10911
rect 7196 10804 7248 10810
rect 7196 10746 7248 10752
rect 7104 9104 7156 9110
rect 7104 9046 7156 9052
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6920 8628 6972 8634
rect 6920 8570 6972 8576
rect 7024 7546 7052 8910
rect 7300 8106 7328 11342
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7392 9450 7420 11222
rect 7484 10713 7512 12174
rect 7668 11762 7696 12804
rect 7748 12786 7800 12792
rect 7852 12696 7880 15660
rect 8484 15632 8536 15638
rect 8312 15580 8484 15586
rect 8312 15574 8536 15580
rect 8312 15570 8524 15574
rect 8300 15564 8524 15570
rect 8352 15558 8524 15564
rect 8300 15506 8352 15512
rect 8312 15162 8340 15506
rect 8680 15366 8708 16050
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 13530 7972 13738
rect 8036 13569 8064 14418
rect 8128 14396 8156 14758
rect 8220 14716 8516 14736
rect 8276 14714 8300 14716
rect 8356 14714 8380 14716
rect 8436 14714 8460 14716
rect 8298 14662 8300 14714
rect 8362 14662 8374 14714
rect 8436 14662 8438 14714
rect 8276 14660 8300 14662
rect 8356 14660 8380 14662
rect 8436 14660 8460 14662
rect 8220 14640 8516 14660
rect 8772 14482 8800 23520
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8852 19916 8904 19922
rect 8852 19858 8904 19864
rect 8864 19689 8892 19858
rect 8850 19680 8906 19689
rect 8850 19615 8906 19624
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 8864 17746 8892 19450
rect 8956 18850 8984 21422
rect 9036 21344 9088 21350
rect 9036 21286 9088 21292
rect 9048 20058 9076 21286
rect 9312 21140 9364 21146
rect 9312 21082 9364 21088
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 8956 18822 9076 18850
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18154 8984 18566
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8208 14408 8260 14414
rect 8128 14368 8208 14396
rect 8022 13560 8078 13569
rect 7932 13524 7984 13530
rect 8022 13495 8078 13504
rect 7932 13466 7984 13472
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7944 12986 7972 13330
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7760 12668 7880 12696
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11218 7696 11698
rect 7656 11212 7708 11218
rect 7656 11154 7708 11160
rect 7470 10704 7526 10713
rect 7470 10639 7526 10648
rect 7564 10600 7616 10606
rect 7668 10588 7696 11154
rect 7616 10560 7696 10588
rect 7564 10542 7616 10548
rect 7576 10130 7604 10542
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7472 9920 7524 9926
rect 7470 9888 7472 9897
rect 7524 9888 7526 9897
rect 7470 9823 7526 9832
rect 7380 9444 7432 9450
rect 7380 9386 7432 9392
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7562 9072 7618 9081
rect 7380 9036 7432 9042
rect 7562 9007 7618 9016
rect 7380 8978 7432 8984
rect 7116 8078 7328 8106
rect 7392 8090 7420 8978
rect 7576 8906 7604 9007
rect 7668 8974 7696 9386
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7380 8084 7432 8090
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 6322 7144 8078
rect 7380 8026 7432 8032
rect 7196 8016 7248 8022
rect 7196 7958 7248 7964
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 6840 6174 6960 6202
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6276 5908 6328 5914
rect 6276 5850 6328 5856
rect 6840 5846 6868 6054
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 4588 5468 4884 5488
rect 4644 5466 4668 5468
rect 4724 5466 4748 5468
rect 4804 5466 4828 5468
rect 4666 5414 4668 5466
rect 4730 5414 4742 5466
rect 4804 5414 4806 5466
rect 4644 5412 4668 5414
rect 4724 5412 4748 5414
rect 4804 5412 4828 5414
rect 4588 5392 4884 5412
rect 4588 4380 4884 4400
rect 4644 4378 4668 4380
rect 4724 4378 4748 4380
rect 4804 4378 4828 4380
rect 4666 4326 4668 4378
rect 4730 4326 4742 4378
rect 4804 4326 4806 4378
rect 4644 4324 4668 4326
rect 4724 4324 4748 4326
rect 4804 4324 4828 4326
rect 4588 4304 4884 4324
rect 3606 4040 3662 4049
rect 3606 3975 3662 3984
rect 3516 3664 3568 3670
rect 3516 3606 3568 3612
rect 4588 3292 4884 3312
rect 4644 3290 4668 3292
rect 4724 3290 4748 3292
rect 4804 3290 4828 3292
rect 4666 3238 4668 3290
rect 4730 3238 4742 3290
rect 4804 3238 4806 3290
rect 4644 3236 4668 3238
rect 4724 3236 4748 3238
rect 4804 3236 4828 3238
rect 4588 3216 4884 3236
rect 6932 3058 6960 6174
rect 7208 5778 7236 7958
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7286 7440 7342 7449
rect 7286 7375 7342 7384
rect 7300 7002 7328 7375
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7392 6934 7420 7822
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5914 7328 6054
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 7484 3194 7512 8502
rect 7760 8378 7788 12668
rect 7840 11620 7892 11626
rect 7840 11562 7892 11568
rect 7852 10849 7880 11562
rect 7944 11540 7972 12922
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 8036 11898 8064 12650
rect 8128 12238 8156 14368
rect 8208 14350 8260 14356
rect 8864 13920 8892 15846
rect 8680 13892 8892 13920
rect 8220 13628 8516 13648
rect 8276 13626 8300 13628
rect 8356 13626 8380 13628
rect 8436 13626 8460 13628
rect 8298 13574 8300 13626
rect 8362 13574 8374 13626
rect 8436 13574 8438 13626
rect 8276 13572 8300 13574
rect 8356 13572 8380 13574
rect 8436 13572 8460 13574
rect 8220 13552 8516 13572
rect 8220 12540 8516 12560
rect 8276 12538 8300 12540
rect 8356 12538 8380 12540
rect 8436 12538 8460 12540
rect 8298 12486 8300 12538
rect 8362 12486 8374 12538
rect 8436 12486 8438 12538
rect 8276 12484 8300 12486
rect 8356 12484 8380 12486
rect 8436 12484 8460 12486
rect 8220 12464 8516 12484
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 8114 11792 8170 11801
rect 8114 11727 8170 11736
rect 8024 11552 8076 11558
rect 7944 11512 8024 11540
rect 8024 11494 8076 11500
rect 7838 10840 7894 10849
rect 8128 10810 8156 11727
rect 8220 11452 8516 11472
rect 8276 11450 8300 11452
rect 8356 11450 8380 11452
rect 8436 11450 8460 11452
rect 8298 11398 8300 11450
rect 8362 11398 8374 11450
rect 8436 11398 8438 11450
rect 8276 11396 8300 11398
rect 8356 11396 8380 11398
rect 8436 11396 8460 11398
rect 8220 11376 8516 11396
rect 8588 11354 8616 12038
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8208 11280 8260 11286
rect 8208 11222 8260 11228
rect 8220 10810 8248 11222
rect 7838 10775 7894 10784
rect 8116 10804 8168 10810
rect 7852 10266 7880 10775
rect 8116 10746 8168 10752
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 7930 10568 7986 10577
rect 7930 10503 7986 10512
rect 8024 10532 8076 10538
rect 7840 10260 7892 10266
rect 7840 10202 7892 10208
rect 7944 9568 7972 10503
rect 8024 10474 8076 10480
rect 8036 10305 8064 10474
rect 8220 10364 8516 10384
rect 8276 10362 8300 10364
rect 8356 10362 8380 10364
rect 8436 10362 8460 10364
rect 8298 10310 8300 10362
rect 8362 10310 8374 10362
rect 8436 10310 8438 10362
rect 8276 10308 8300 10310
rect 8356 10308 8380 10310
rect 8436 10308 8460 10310
rect 8022 10296 8078 10305
rect 8220 10288 8516 10308
rect 8022 10231 8078 10240
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 8022 9888 8078 9897
rect 8022 9823 8078 9832
rect 7852 9540 7972 9568
rect 7852 9217 7880 9540
rect 8036 9353 8064 9823
rect 8404 9518 8432 10066
rect 8588 9518 8616 10202
rect 8392 9512 8444 9518
rect 8114 9480 8170 9489
rect 8392 9454 8444 9460
rect 8576 9512 8628 9518
rect 8576 9454 8628 9460
rect 8114 9415 8170 9424
rect 8022 9344 8078 9353
rect 8022 9279 8078 9288
rect 7838 9208 7894 9217
rect 8128 9194 8156 9415
rect 8680 9364 8708 13892
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8772 12782 8800 13670
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8864 12374 8892 13738
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 9994 8800 10406
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8956 9761 8984 18090
rect 9048 16425 9076 18822
rect 9140 18222 9168 20334
rect 9218 19816 9274 19825
rect 9218 19751 9220 19760
rect 9272 19751 9274 19760
rect 9220 19722 9272 19728
rect 9324 19281 9352 21082
rect 9310 19272 9366 19281
rect 9310 19207 9366 19216
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9140 17066 9168 18158
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9140 16726 9168 17002
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9034 16416 9090 16425
rect 9034 16351 9090 16360
rect 9232 14346 9260 16594
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9324 13462 9352 19207
rect 9416 14890 9444 23520
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9588 21480 9640 21486
rect 9588 21422 9640 21428
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9508 20330 9536 20742
rect 9600 20398 9628 21422
rect 9692 20466 9720 21558
rect 9956 21412 10008 21418
rect 9956 21354 10008 21360
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9496 20324 9548 20330
rect 9496 20266 9548 20272
rect 9404 14884 9456 14890
rect 9404 14826 9456 14832
rect 9404 14476 9456 14482
rect 9404 14418 9456 14424
rect 9312 13456 9364 13462
rect 9312 13398 9364 13404
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9140 12238 9168 12718
rect 9416 12238 9444 14418
rect 9128 12232 9180 12238
rect 9048 12192 9128 12220
rect 8942 9752 8998 9761
rect 8942 9687 8998 9696
rect 9048 9518 9076 12192
rect 9128 12174 9180 12180
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9140 9926 9168 11630
rect 9324 11354 9352 12106
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9232 10538 9260 10950
rect 9310 10840 9366 10849
rect 9310 10775 9366 10784
rect 9220 10532 9272 10538
rect 9220 10474 9272 10480
rect 9324 10282 9352 10775
rect 9232 10254 9352 10282
rect 9232 10062 9260 10254
rect 9416 10130 9444 12174
rect 9508 11937 9536 20266
rect 9784 19718 9812 20878
rect 9968 20262 9996 21354
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9588 19168 9640 19174
rect 9586 19136 9588 19145
rect 9640 19136 9642 19145
rect 9586 19071 9642 19080
rect 9586 17096 9642 17105
rect 9586 17031 9588 17040
rect 9640 17031 9642 17040
rect 9588 17002 9640 17008
rect 9692 16794 9720 19246
rect 9784 17814 9812 19654
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9876 18057 9904 18362
rect 9862 18048 9918 18057
rect 9862 17983 9918 17992
rect 9772 17808 9824 17814
rect 9772 17750 9824 17756
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9586 16688 9642 16697
rect 9586 16623 9642 16632
rect 9600 16590 9628 16623
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9692 13870 9720 16730
rect 9772 15972 9824 15978
rect 9772 15914 9824 15920
rect 9784 15314 9812 15914
rect 9864 15360 9916 15366
rect 9784 15308 9864 15314
rect 9784 15302 9916 15308
rect 9784 15286 9904 15302
rect 9784 14890 9812 15286
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9784 14482 9812 14826
rect 9772 14476 9824 14482
rect 9772 14418 9824 14424
rect 9784 14074 9812 14418
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12850 9720 13194
rect 9784 12850 9812 13262
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9494 11928 9550 11937
rect 9494 11863 9550 11872
rect 9876 11762 9904 12718
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9692 11218 9720 11698
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9692 10690 9720 11154
rect 9784 10810 9812 11630
rect 9772 10804 9824 10810
rect 9772 10746 9824 10752
rect 9692 10662 9812 10690
rect 9784 10606 9812 10662
rect 9772 10600 9824 10606
rect 9772 10542 9824 10548
rect 9864 10600 9916 10606
rect 9864 10542 9916 10548
rect 9588 10464 9640 10470
rect 9494 10432 9550 10441
rect 9588 10406 9640 10412
rect 9494 10367 9550 10376
rect 9404 10124 9456 10130
rect 9404 10066 9456 10072
rect 9220 10056 9272 10062
rect 9508 10010 9536 10367
rect 9220 9998 9272 10004
rect 9416 9982 9536 10010
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 9140 9761 9168 9862
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 9128 9444 9180 9450
rect 9128 9386 9180 9392
rect 8680 9336 8800 9364
rect 8220 9276 8516 9296
rect 8276 9274 8300 9276
rect 8356 9274 8380 9276
rect 8436 9274 8460 9276
rect 8298 9222 8300 9274
rect 8362 9222 8374 9274
rect 8436 9222 8438 9274
rect 8276 9220 8300 9222
rect 8356 9220 8380 9222
rect 8436 9220 8460 9222
rect 8220 9200 8516 9220
rect 7838 9143 7894 9152
rect 8036 9166 8156 9194
rect 7668 8350 7788 8378
rect 7852 9042 7972 9058
rect 7852 9036 7984 9042
rect 7852 9030 7932 9036
rect 7562 7712 7618 7721
rect 7562 7647 7618 7656
rect 7576 7478 7604 7647
rect 7564 7472 7616 7478
rect 7564 7414 7616 7420
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 7002 7604 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7668 6866 7696 8350
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 7342 7788 8230
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7576 6118 7604 6734
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7760 4185 7788 6666
rect 7852 5370 7880 9030
rect 7932 8978 7984 8984
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7944 7886 7972 8434
rect 8036 8362 8064 9166
rect 8576 9104 8628 9110
rect 8576 9046 8628 9052
rect 8116 8560 8168 8566
rect 8116 8502 8168 8508
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7342 7972 7822
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 6798 7972 7278
rect 8128 7274 8156 8502
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 8362 8248 8434
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8496 8276 8524 8366
rect 8588 8344 8616 9046
rect 8668 8560 8720 8566
rect 8772 8548 8800 9336
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8944 8968 8996 8974
rect 8996 8928 9076 8956
rect 8944 8910 8996 8916
rect 8720 8520 8800 8548
rect 8668 8502 8720 8508
rect 8772 8362 8800 8427
rect 8760 8356 8812 8362
rect 8588 8316 8760 8344
rect 8760 8298 8812 8304
rect 8496 8248 8708 8276
rect 8220 8188 8516 8208
rect 8276 8186 8300 8188
rect 8356 8186 8380 8188
rect 8436 8186 8460 8188
rect 8298 8134 8300 8186
rect 8362 8134 8374 8186
rect 8436 8134 8438 8186
rect 8276 8132 8300 8134
rect 8356 8132 8380 8134
rect 8436 8132 8460 8134
rect 8220 8112 8516 8132
rect 8680 7834 8708 8248
rect 8772 8090 8800 8298
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8864 7993 8892 8910
rect 8850 7984 8906 7993
rect 9048 7954 9076 8928
rect 8850 7919 8906 7928
rect 9036 7948 9088 7954
rect 9036 7890 9088 7896
rect 9140 7886 9168 9386
rect 9310 9072 9366 9081
rect 9310 9007 9366 9016
rect 9416 9024 9444 9982
rect 9600 9654 9628 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9784 9722 9812 10066
rect 9876 9994 9904 10542
rect 9864 9988 9916 9994
rect 9864 9930 9916 9936
rect 9968 9897 9996 20198
rect 10152 19514 10180 23520
rect 10888 22794 10916 23520
rect 10704 22766 10916 22794
rect 10508 22364 10560 22370
rect 10508 22306 10560 22312
rect 10416 21004 10468 21010
rect 10416 20946 10468 20952
rect 10322 20088 10378 20097
rect 10322 20023 10378 20032
rect 10336 19854 10364 20023
rect 10324 19848 10376 19854
rect 10324 19790 10376 19796
rect 10140 19508 10192 19514
rect 10140 19450 10192 19456
rect 10428 19174 10456 20946
rect 10520 19786 10548 22306
rect 10600 20868 10652 20874
rect 10600 20810 10652 20816
rect 10612 20398 10640 20810
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10508 19780 10560 19786
rect 10508 19722 10560 19728
rect 10612 19417 10640 19790
rect 10598 19408 10654 19417
rect 10598 19343 10654 19352
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10060 18358 10088 19110
rect 10230 19000 10286 19009
rect 10230 18935 10286 18944
rect 10336 18986 10364 19110
rect 10612 18986 10640 19246
rect 10336 18958 10640 18986
rect 10048 18352 10100 18358
rect 10048 18294 10100 18300
rect 10060 10169 10088 18294
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10152 17134 10180 17614
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10244 15570 10272 18935
rect 10336 18222 10364 18958
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10428 16182 10456 18770
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10612 18290 10640 18702
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10600 18080 10652 18086
rect 10600 18022 10652 18028
rect 10612 17882 10640 18022
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10508 17740 10560 17746
rect 10508 17682 10560 17688
rect 10520 17338 10548 17682
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10520 16726 10548 17274
rect 10508 16720 10560 16726
rect 10508 16662 10560 16668
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10704 15994 10732 22766
rect 11532 22114 11560 23520
rect 12164 22296 12216 22302
rect 12164 22238 12216 22244
rect 11532 22086 11652 22114
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 10784 20800 10836 20806
rect 10784 20742 10836 20748
rect 10796 17134 10824 20742
rect 10980 20505 11008 20878
rect 10966 20496 11022 20505
rect 10966 20431 11022 20440
rect 10968 20324 11020 20330
rect 10888 20284 10968 20312
rect 10784 17128 10836 17134
rect 10784 17070 10836 17076
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16046 10824 16730
rect 10428 15966 10732 15994
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10428 15706 10456 15966
rect 10888 15858 10916 20284
rect 11072 20312 11100 21286
rect 11624 20602 11652 22086
rect 11852 21788 12148 21808
rect 11908 21786 11932 21788
rect 11988 21786 12012 21788
rect 12068 21786 12092 21788
rect 11930 21734 11932 21786
rect 11994 21734 12006 21786
rect 12068 21734 12070 21786
rect 11908 21732 11932 21734
rect 11988 21732 12012 21734
rect 12068 21732 12092 21734
rect 11852 21712 12148 21732
rect 12176 21350 12204 22238
rect 12268 22114 12296 23520
rect 12268 22086 12388 22114
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12268 21010 12296 21082
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 11852 20700 12148 20720
rect 11908 20698 11932 20700
rect 11988 20698 12012 20700
rect 12068 20698 12092 20700
rect 11930 20646 11932 20698
rect 11994 20646 12006 20698
rect 12068 20646 12070 20698
rect 11908 20644 11932 20646
rect 11988 20644 12012 20646
rect 12068 20644 12092 20646
rect 11852 20624 12148 20644
rect 12268 20602 12296 20946
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 11020 20284 11100 20312
rect 10968 20266 11020 20272
rect 11348 20262 11376 20538
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 11336 20256 11388 20262
rect 11336 20198 11388 20204
rect 12176 19990 12204 20334
rect 12164 19984 12216 19990
rect 11072 19910 11744 19938
rect 12164 19926 12216 19932
rect 11072 19854 11100 19910
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 10968 19168 11020 19174
rect 11072 19145 11100 19790
rect 10968 19110 11020 19116
rect 11058 19136 11114 19145
rect 10980 18986 11008 19110
rect 11058 19071 11114 19080
rect 10980 18958 11100 18986
rect 11072 18834 11100 18958
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11072 16402 11100 18634
rect 11256 18630 11284 19790
rect 11334 19408 11390 19417
rect 11334 19343 11390 19352
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11164 16658 11192 18090
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11072 16374 11192 16402
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 10520 15830 10916 15858
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10336 13326 10364 14962
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12442 10456 13262
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10140 12232 10192 12238
rect 10232 12232 10284 12238
rect 10140 12174 10192 12180
rect 10230 12200 10232 12209
rect 10284 12200 10286 12209
rect 10152 11626 10180 12174
rect 10230 12135 10286 12144
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 10138 10296 10194 10305
rect 10138 10231 10194 10240
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9954 9888 10010 9897
rect 9954 9823 10010 9832
rect 9772 9716 9824 9722
rect 9772 9658 9824 9664
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9692 9586 9904 9602
rect 9692 9580 9916 9586
rect 9692 9574 9864 9580
rect 9496 9512 9548 9518
rect 9692 9500 9720 9574
rect 9864 9522 9916 9528
rect 9548 9472 9720 9500
rect 9772 9512 9824 9518
rect 9496 9454 9548 9460
rect 10060 9466 10088 9930
rect 10152 9586 10180 10231
rect 10244 10062 10272 10678
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10336 10130 10364 10610
rect 10520 10418 10548 15830
rect 11072 15638 11100 16186
rect 11164 15706 11192 16374
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 14958 10824 15302
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10784 14952 10836 14958
rect 10784 14894 10836 14900
rect 11072 14550 11100 15098
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11060 14544 11112 14550
rect 11060 14486 11112 14492
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 10968 13932 11020 13938
rect 10968 13874 11020 13880
rect 10980 13530 11008 13874
rect 11072 13870 11100 14214
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11164 13530 11192 14758
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10704 12782 10732 13126
rect 11060 12844 11112 12850
rect 11060 12786 11112 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10692 12776 10744 12782
rect 11072 12730 11100 12786
rect 10692 12718 10744 12724
rect 10612 12594 10640 12718
rect 10796 12702 11100 12730
rect 10796 12594 10824 12702
rect 10612 12566 10824 12594
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10690 12472 10746 12481
rect 10690 12407 10692 12416
rect 10744 12407 10746 12416
rect 10692 12378 10744 12384
rect 10692 11212 10744 11218
rect 10692 11154 10744 11160
rect 10428 10390 10548 10418
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9824 9460 10088 9466
rect 9772 9454 10088 9460
rect 9784 9438 10088 9454
rect 9772 9172 9824 9178
rect 9824 9132 9996 9160
rect 9772 9114 9824 9120
rect 9968 9081 9996 9132
rect 9954 9072 10010 9081
rect 9496 9036 9548 9042
rect 9220 8424 9272 8430
rect 9220 8366 9272 8372
rect 9232 8294 9260 8366
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9128 7880 9180 7886
rect 8680 7818 8984 7834
rect 9128 7822 9180 7828
rect 9324 7818 9352 9007
rect 9416 8996 9496 9024
rect 8680 7812 8996 7818
rect 8680 7806 8944 7812
rect 8944 7754 8996 7760
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 8116 7268 8168 7274
rect 8116 7210 8168 7216
rect 8576 7268 8628 7274
rect 9416 7256 9444 8996
rect 9496 8978 9548 8984
rect 9680 9036 9732 9042
rect 9732 8996 9904 9024
rect 9954 9007 10010 9016
rect 9680 8978 9732 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9600 8894 9812 8922
rect 9508 8401 9536 8842
rect 9494 8392 9550 8401
rect 9494 8327 9550 8336
rect 9600 8276 9628 8894
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9784 8786 9812 8894
rect 9876 8888 9904 8996
rect 9876 8860 9996 8888
rect 9692 8650 9720 8774
rect 9784 8758 9904 8786
rect 9692 8622 9812 8650
rect 9508 8248 9628 8276
rect 9508 7886 9536 8248
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9600 7546 9628 7890
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9496 7268 9548 7274
rect 9416 7228 9496 7256
rect 8576 7210 8628 7216
rect 9496 7210 9548 7216
rect 8220 7100 8516 7120
rect 8276 7098 8300 7100
rect 8356 7098 8380 7100
rect 8436 7098 8460 7100
rect 8298 7046 8300 7098
rect 8362 7046 8374 7098
rect 8436 7046 8438 7098
rect 8276 7044 8300 7046
rect 8356 7044 8380 7046
rect 8436 7044 8460 7046
rect 8220 7024 8516 7044
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7944 6202 7972 6734
rect 8114 6488 8170 6497
rect 8588 6458 8616 7210
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 8114 6423 8170 6432
rect 8576 6452 8628 6458
rect 8024 6384 8076 6390
rect 8022 6352 8024 6361
rect 8076 6352 8078 6361
rect 8128 6322 8156 6423
rect 8576 6394 8628 6400
rect 8022 6287 8078 6296
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8300 6248 8352 6254
rect 7944 6196 8300 6202
rect 7944 6190 8352 6196
rect 7944 6174 8340 6190
rect 7944 5710 7972 6174
rect 8220 6012 8516 6032
rect 8276 6010 8300 6012
rect 8356 6010 8380 6012
rect 8436 6010 8460 6012
rect 8298 5958 8300 6010
rect 8362 5958 8374 6010
rect 8436 5958 8438 6010
rect 8276 5956 8300 5958
rect 8356 5956 8380 5958
rect 8436 5956 8460 5958
rect 8220 5936 8516 5956
rect 8024 5772 8076 5778
rect 8076 5732 8616 5760
rect 8024 5714 8076 5720
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 5166 7972 5646
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 8220 4924 8516 4944
rect 8276 4922 8300 4924
rect 8356 4922 8380 4924
rect 8436 4922 8460 4924
rect 8298 4870 8300 4922
rect 8362 4870 8374 4922
rect 8436 4870 8438 4922
rect 8276 4868 8300 4870
rect 8356 4868 8380 4870
rect 8436 4868 8460 4870
rect 8220 4848 8516 4868
rect 7746 4176 7802 4185
rect 7746 4111 7802 4120
rect 8588 4010 8616 5732
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 9140 3942 9168 5646
rect 9232 5574 9260 6802
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6254 9352 6598
rect 9508 6497 9536 7210
rect 9692 7002 9720 7482
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9784 6866 9812 8622
rect 9876 8378 9904 8758
rect 9968 8498 9996 8860
rect 10048 8832 10100 8838
rect 10048 8774 10100 8780
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10060 8378 10088 8774
rect 9876 8350 10088 8378
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 8022 10088 8230
rect 10048 8016 10100 8022
rect 10048 7958 10100 7964
rect 10060 7410 10088 7958
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10060 7002 10088 7142
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9494 6488 9550 6497
rect 9494 6423 9550 6432
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9232 4078 9260 5510
rect 9508 4214 9536 6423
rect 9876 5778 9904 6734
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 10060 6254 10088 6598
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9588 5772 9640 5778
rect 9588 5714 9640 5720
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9600 5370 9628 5714
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9600 4146 9628 5306
rect 10046 4856 10102 4865
rect 10046 4791 10048 4800
rect 10100 4791 10102 4800
rect 10048 4762 10100 4768
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 10244 4078 10272 9862
rect 10336 9518 10364 10066
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10336 8498 10364 9454
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10428 7546 10456 10390
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10520 9518 10548 10202
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 9512 10560 9518
rect 10508 9454 10560 9460
rect 10612 9382 10640 10066
rect 10600 9376 10652 9382
rect 10600 9318 10652 9324
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7206 10456 7346
rect 10416 7200 10468 7206
rect 10416 7142 10468 7148
rect 10520 6254 10548 7890
rect 10508 6248 10560 6254
rect 10508 6190 10560 6196
rect 10520 5710 10548 6190
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10520 5166 10548 5646
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10520 5030 10548 5102
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4622 10548 4966
rect 10508 4616 10560 4622
rect 10508 4558 10560 4564
rect 10704 4146 10732 11154
rect 10796 10674 10824 12566
rect 11072 12374 11100 12582
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11060 11620 11112 11626
rect 11060 11562 11112 11568
rect 11072 11354 11100 11562
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11256 11098 11284 18566
rect 11348 18170 11376 19343
rect 11440 18358 11468 19790
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11532 18358 11560 18770
rect 11624 18426 11652 19790
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11348 18142 11560 18170
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 11428 18080 11480 18086
rect 11428 18022 11480 18028
rect 11348 15994 11376 18022
rect 11440 17338 11468 18022
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11532 16454 11560 18142
rect 11716 17814 11744 19910
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12084 19825 12112 19858
rect 12070 19816 12126 19825
rect 12070 19751 12126 19760
rect 11852 19612 12148 19632
rect 11908 19610 11932 19612
rect 11988 19610 12012 19612
rect 12068 19610 12092 19612
rect 11930 19558 11932 19610
rect 11994 19558 12006 19610
rect 12068 19558 12070 19610
rect 11908 19556 11932 19558
rect 11988 19556 12012 19558
rect 12068 19556 12092 19558
rect 11852 19536 12148 19556
rect 12360 19446 12388 22086
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12532 21548 12584 21554
rect 12532 21490 12584 21496
rect 12544 20942 12572 21490
rect 12624 21480 12676 21486
rect 12624 21422 12676 21428
rect 12532 20936 12584 20942
rect 12532 20878 12584 20884
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12452 19310 12480 20742
rect 12544 20398 12572 20878
rect 12636 20641 12664 21422
rect 12622 20632 12678 20641
rect 12622 20567 12678 20576
rect 12532 20392 12584 20398
rect 12532 20334 12584 20340
rect 12544 19938 12572 20334
rect 12728 20330 12756 21830
rect 12808 21344 12860 21350
rect 12808 21286 12860 21292
rect 12716 20324 12768 20330
rect 12716 20266 12768 20272
rect 12728 20074 12756 20266
rect 12820 20262 12848 21286
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12728 20046 12848 20074
rect 12544 19910 12756 19938
rect 12532 19848 12584 19854
rect 12530 19816 12532 19825
rect 12584 19816 12586 19825
rect 12530 19751 12586 19760
rect 12532 19712 12584 19718
rect 12530 19680 12532 19689
rect 12624 19712 12676 19718
rect 12584 19680 12586 19689
rect 12624 19654 12676 19660
rect 12530 19615 12586 19624
rect 12636 19417 12664 19654
rect 12622 19408 12678 19417
rect 12622 19343 12678 19352
rect 12440 19304 12492 19310
rect 12254 19272 12310 19281
rect 12440 19246 12492 19252
rect 12530 19272 12586 19281
rect 12254 19207 12256 19216
rect 12308 19207 12310 19216
rect 12530 19207 12532 19216
rect 12256 19178 12308 19184
rect 12584 19207 12586 19216
rect 12728 19258 12756 19910
rect 12820 19378 12848 20046
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12808 19372 12860 19378
rect 12808 19314 12860 19320
rect 12912 19258 12940 19858
rect 12728 19230 12940 19258
rect 12532 19178 12584 19184
rect 12164 18896 12216 18902
rect 12162 18864 12164 18873
rect 12216 18864 12218 18873
rect 12728 18834 12756 19230
rect 12808 19168 12860 19174
rect 12808 19110 12860 19116
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12820 18970 12848 19110
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12162 18799 12218 18808
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12716 18828 12768 18834
rect 12716 18770 12768 18776
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 11852 18524 12148 18544
rect 11908 18522 11932 18524
rect 11988 18522 12012 18524
rect 12068 18522 12092 18524
rect 11930 18470 11932 18522
rect 11994 18470 12006 18522
rect 12068 18470 12070 18522
rect 11908 18468 11932 18470
rect 11988 18468 12012 18470
rect 12068 18468 12092 18470
rect 11852 18448 12148 18468
rect 12176 18442 12204 18702
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12254 18456 12310 18465
rect 12176 18414 12254 18442
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11716 17202 11744 17614
rect 11808 17610 11836 18294
rect 12176 18290 12204 18414
rect 12254 18391 12310 18400
rect 12164 18284 12216 18290
rect 12164 18226 12216 18232
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12268 17898 12296 18226
rect 12360 18154 12388 18566
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12176 17870 12296 17898
rect 12176 17678 12204 17870
rect 12452 17814 12480 18770
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12544 18154 12572 18566
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12256 17808 12308 17814
rect 12256 17750 12308 17756
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 11796 17604 11848 17610
rect 11796 17546 11848 17552
rect 11852 17436 12148 17456
rect 11908 17434 11932 17436
rect 11988 17434 12012 17436
rect 12068 17434 12092 17436
rect 11930 17382 11932 17434
rect 11994 17382 12006 17434
rect 12068 17382 12070 17434
rect 11908 17380 11932 17382
rect 11988 17380 12012 17382
rect 12068 17380 12092 17382
rect 11852 17360 12148 17380
rect 12176 17270 12204 17614
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11624 16114 11652 16526
rect 11716 16250 11744 16594
rect 11900 16590 11928 17138
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11852 16348 12148 16368
rect 11908 16346 11932 16348
rect 11988 16346 12012 16348
rect 12068 16346 12092 16348
rect 11930 16294 11932 16346
rect 11994 16294 12006 16346
rect 12068 16294 12070 16346
rect 11908 16292 11932 16294
rect 11988 16292 12012 16294
rect 12068 16292 12092 16294
rect 11852 16272 12148 16292
rect 12268 16289 12296 17750
rect 12346 17640 12402 17649
rect 12346 17575 12402 17584
rect 12360 17542 12388 17575
rect 12636 17542 12664 18634
rect 12728 18426 12756 18770
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12716 18148 12768 18154
rect 12716 18090 12768 18096
rect 12728 17882 12756 18090
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12438 17368 12494 17377
rect 12438 17303 12440 17312
rect 12492 17303 12494 17312
rect 12440 17274 12492 17280
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 16658 12480 17070
rect 12544 17066 12756 17082
rect 12532 17060 12756 17066
rect 12584 17054 12756 17060
rect 12532 17002 12584 17008
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12440 16652 12492 16658
rect 12440 16594 12492 16600
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12348 16448 12400 16454
rect 12348 16390 12400 16396
rect 12254 16280 12310 16289
rect 11704 16244 11756 16250
rect 12254 16215 12310 16224
rect 11704 16186 11756 16192
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11348 15966 11468 15994
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11348 14550 11376 15846
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11348 14074 11376 14486
rect 11336 14068 11388 14074
rect 11336 14010 11388 14016
rect 11440 13870 11468 15966
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 14278 11560 15846
rect 11624 15434 11652 16050
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11716 15162 11744 15506
rect 11852 15260 12148 15280
rect 11908 15258 11932 15260
rect 11988 15258 12012 15260
rect 12068 15258 12092 15260
rect 11930 15206 11932 15258
rect 11994 15206 12006 15258
rect 12068 15206 12070 15258
rect 11908 15204 11932 15206
rect 11988 15204 12012 15206
rect 12068 15204 12092 15206
rect 11852 15184 12148 15204
rect 12360 15162 12388 16390
rect 12440 16244 12492 16250
rect 12440 16186 12492 16192
rect 12452 16046 12480 16186
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12452 15502 12480 15982
rect 12440 15496 12492 15502
rect 12440 15438 12492 15444
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12452 14958 12480 15438
rect 11704 14952 11756 14958
rect 11704 14894 11756 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11428 13864 11480 13870
rect 11428 13806 11480 13812
rect 11624 13308 11652 14758
rect 11348 13280 11652 13308
rect 11348 12714 11376 13280
rect 11716 13190 11744 14894
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11852 14172 12148 14192
rect 11908 14170 11932 14172
rect 11988 14170 12012 14172
rect 12068 14170 12092 14172
rect 11930 14118 11932 14170
rect 11994 14118 12006 14170
rect 12068 14118 12070 14170
rect 11908 14116 11932 14118
rect 11988 14116 12012 14118
rect 12068 14116 12092 14118
rect 11852 14096 12148 14116
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13394 11836 13670
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 11348 11898 11376 12650
rect 11336 11892 11388 11898
rect 11336 11834 11388 11840
rect 11440 11762 11468 13126
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 12209 11560 12582
rect 11518 12200 11574 12209
rect 11518 12135 11574 12144
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11716 11694 11744 13126
rect 11852 13084 12148 13104
rect 11908 13082 11932 13084
rect 11988 13082 12012 13084
rect 12068 13082 12092 13084
rect 11930 13030 11932 13082
rect 11994 13030 12006 13082
rect 12068 13030 12070 13082
rect 11908 13028 11932 13030
rect 11988 13028 12012 13030
rect 12068 13028 12092 13030
rect 11852 13008 12148 13028
rect 11888 12912 11940 12918
rect 12176 12900 12204 14758
rect 12452 14414 12480 14894
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12544 13802 12572 16487
rect 12636 14618 12664 16934
rect 12728 14958 12756 17054
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12820 16726 12848 17002
rect 12808 16720 12860 16726
rect 12808 16662 12860 16668
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12728 14634 12756 14894
rect 12728 14618 12848 14634
rect 12624 14612 12676 14618
rect 12728 14612 12860 14618
rect 12728 14606 12808 14612
rect 12624 14554 12676 14560
rect 12808 14554 12860 14560
rect 12912 14006 12940 19110
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 13004 13870 13032 23520
rect 13082 20088 13138 20097
rect 13082 20023 13138 20032
rect 13096 19378 13124 20023
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13358 19680 13414 19689
rect 13358 19615 13414 19624
rect 13174 19544 13230 19553
rect 13174 19479 13176 19488
rect 13228 19479 13230 19488
rect 13176 19450 13228 19456
rect 13268 19440 13320 19446
rect 13268 19382 13320 19388
rect 13084 19372 13136 19378
rect 13084 19314 13136 19320
rect 13096 14074 13124 19314
rect 13280 18222 13308 19382
rect 13176 18216 13228 18222
rect 13176 18158 13228 18164
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13188 17134 13216 18158
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13188 14074 13216 14214
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13188 13870 13216 14010
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 13188 13326 13216 13806
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 11940 12872 12204 12900
rect 11888 12854 11940 12860
rect 12176 12714 12204 12872
rect 12360 12850 12388 13262
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11852 11996 12148 12016
rect 11908 11994 11932 11996
rect 11988 11994 12012 11996
rect 12068 11994 12092 11996
rect 11930 11942 11932 11994
rect 11994 11942 12006 11994
rect 12068 11942 12070 11994
rect 11908 11940 11932 11942
rect 11988 11940 12012 11942
rect 12068 11940 12092 11942
rect 11852 11920 12148 11940
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 12360 11218 12388 12786
rect 12532 12776 12584 12782
rect 12452 12736 12532 12764
rect 12452 11830 12480 12736
rect 12532 12718 12584 12724
rect 12636 12322 12664 13262
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12728 12986 12756 13194
rect 13280 13172 13308 18022
rect 13372 16017 13400 19615
rect 13464 16697 13492 19790
rect 13556 19446 13584 19790
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13648 19378 13676 23520
rect 14280 22840 14332 22846
rect 14280 22782 14332 22788
rect 13912 21412 13964 21418
rect 13912 21354 13964 21360
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13726 20632 13782 20641
rect 13832 20602 13860 21014
rect 13924 20806 13952 21354
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13726 20567 13782 20576
rect 13820 20596 13872 20602
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13648 18834 13676 19178
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 13648 18426 13676 18770
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13740 18086 13768 20567
rect 13820 20538 13872 20544
rect 14292 20262 14320 22782
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14188 19304 14240 19310
rect 14188 19246 14240 19252
rect 14200 18766 14228 19246
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14292 18834 14320 19110
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14278 18456 14334 18465
rect 14278 18391 14280 18400
rect 14332 18391 14334 18400
rect 14280 18362 14332 18368
rect 14188 18216 14240 18222
rect 14188 18158 14240 18164
rect 13728 18080 13780 18086
rect 13728 18022 13780 18028
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 14004 17740 14056 17746
rect 14004 17682 14056 17688
rect 13832 17338 13860 17682
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13450 16688 13506 16697
rect 13450 16623 13506 16632
rect 13358 16008 13414 16017
rect 13556 15978 13584 17070
rect 14016 16726 14044 17682
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13728 16652 13780 16658
rect 13912 16652 13964 16658
rect 13780 16612 13860 16640
rect 13728 16594 13780 16600
rect 13832 16250 13860 16612
rect 13912 16594 13964 16600
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13924 16046 13952 16594
rect 14004 16584 14056 16590
rect 14004 16526 14056 16532
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13358 15943 13414 15952
rect 13544 15972 13596 15978
rect 13188 13144 13308 13172
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12544 12294 12664 12322
rect 12544 12238 12572 12294
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12440 11688 12492 11694
rect 12544 11642 12572 12174
rect 12728 11694 12756 12922
rect 12492 11636 12572 11642
rect 12440 11630 12572 11636
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12452 11614 12572 11630
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11370 12480 11494
rect 12452 11342 12572 11370
rect 12544 11286 12572 11342
rect 12532 11280 12584 11286
rect 12532 11222 12584 11228
rect 11428 11212 11480 11218
rect 11612 11212 11664 11218
rect 11480 11172 11560 11200
rect 11428 11154 11480 11160
rect 11164 11070 11284 11098
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10796 9081 10824 9114
rect 10782 9072 10838 9081
rect 10888 9042 10916 10066
rect 11058 9752 11114 9761
rect 11058 9687 11114 9696
rect 10966 9072 11022 9081
rect 10782 9007 10838 9016
rect 10876 9036 10928 9042
rect 10966 9007 11022 9016
rect 10876 8978 10928 8984
rect 10980 8809 11008 9007
rect 10966 8800 11022 8809
rect 10966 8735 11022 8744
rect 11072 8362 11100 9687
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10888 7750 10916 8298
rect 10876 7744 10928 7750
rect 11164 7721 11192 11070
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11256 9722 11284 10950
rect 11348 10606 11376 10950
rect 11336 10600 11388 10606
rect 11336 10542 11388 10548
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10198 11468 10406
rect 11428 10192 11480 10198
rect 11428 10134 11480 10140
rect 11336 10056 11388 10062
rect 11336 9998 11388 10004
rect 11244 9716 11296 9722
rect 11244 9658 11296 9664
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 11256 9217 11284 9386
rect 11242 9208 11298 9217
rect 11242 9143 11298 9152
rect 11348 8906 11376 9998
rect 11532 9994 11560 11172
rect 11612 11154 11664 11160
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 11520 9988 11572 9994
rect 11520 9930 11572 9936
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11244 8832 11296 8838
rect 11440 8786 11468 9522
rect 11532 9042 11560 9930
rect 11624 9926 11652 11154
rect 11852 10908 12148 10928
rect 11908 10906 11932 10908
rect 11988 10906 12012 10908
rect 12068 10906 12092 10908
rect 11930 10854 11932 10906
rect 11994 10854 12006 10906
rect 12068 10854 12070 10906
rect 11908 10852 11932 10854
rect 11988 10852 12012 10854
rect 12068 10852 12092 10854
rect 11852 10832 12148 10852
rect 12360 10674 12388 11154
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12440 10804 12492 10810
rect 12440 10746 12492 10752
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12164 10600 12216 10606
rect 12164 10542 12216 10548
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11716 9194 11744 10406
rect 11852 9820 12148 9840
rect 11908 9818 11932 9820
rect 11988 9818 12012 9820
rect 12068 9818 12092 9820
rect 11930 9766 11932 9818
rect 11994 9766 12006 9818
rect 12068 9766 12070 9818
rect 11908 9764 11932 9766
rect 11988 9764 12012 9766
rect 12068 9764 12092 9766
rect 11852 9744 12148 9764
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11624 9166 11744 9194
rect 11520 9036 11572 9042
rect 11520 8978 11572 8984
rect 11244 8774 11296 8780
rect 11256 8634 11284 8774
rect 11348 8758 11468 8786
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11348 7954 11376 8758
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 10876 7686 10928 7692
rect 11150 7712 11206 7721
rect 10888 7274 10916 7686
rect 11150 7647 11206 7656
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10888 6458 10916 6598
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 11072 6118 11100 7142
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11256 5166 11284 6054
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 11256 4078 11284 5102
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 11244 4072 11296 4078
rect 11244 4014 11296 4020
rect 11348 3942 11376 6734
rect 11440 5370 11468 8502
rect 11532 7886 11560 8978
rect 11624 8106 11652 9166
rect 11704 9036 11756 9042
rect 11808 9024 11836 9386
rect 11756 8996 11836 9024
rect 11704 8978 11756 8984
rect 11716 8634 11744 8978
rect 11852 8732 12148 8752
rect 11908 8730 11932 8732
rect 11988 8730 12012 8732
rect 12068 8730 12092 8732
rect 11930 8678 11932 8730
rect 11994 8678 12006 8730
rect 12068 8678 12070 8730
rect 11908 8676 11932 8678
rect 11988 8676 12012 8678
rect 12068 8676 12092 8678
rect 11852 8656 12148 8676
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 12176 8566 12204 10542
rect 12452 10441 12480 10746
rect 13004 10606 13032 11086
rect 12992 10600 13044 10606
rect 12714 10568 12770 10577
rect 12992 10542 13044 10548
rect 12714 10503 12770 10512
rect 12438 10432 12494 10441
rect 12438 10367 12494 10376
rect 12268 9926 12296 9957
rect 12256 9920 12308 9926
rect 12254 9888 12256 9897
rect 12308 9888 12310 9897
rect 12254 9823 12310 9832
rect 12268 8956 12296 9823
rect 12346 9616 12402 9625
rect 12346 9551 12402 9560
rect 12360 9058 12388 9551
rect 12440 9512 12492 9518
rect 12492 9472 12664 9500
rect 12440 9454 12492 9460
rect 12636 9110 12664 9472
rect 12624 9104 12676 9110
rect 12360 9030 12572 9058
rect 12624 9046 12676 9052
rect 12440 8968 12492 8974
rect 12268 8928 12440 8956
rect 12440 8910 12492 8916
rect 12544 8809 12572 9030
rect 12622 8936 12678 8945
rect 12622 8871 12678 8880
rect 12636 8838 12664 8871
rect 12624 8832 12676 8838
rect 12530 8800 12586 8809
rect 12624 8774 12676 8780
rect 12530 8735 12586 8744
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11624 8078 11744 8106
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11716 7698 11744 8078
rect 11624 7670 11744 7698
rect 11624 7426 11652 7670
rect 11852 7644 12148 7664
rect 11908 7642 11932 7644
rect 11988 7642 12012 7644
rect 12068 7642 12092 7644
rect 11930 7590 11932 7642
rect 11994 7590 12006 7642
rect 12068 7590 12070 7642
rect 11908 7588 11932 7590
rect 11988 7588 12012 7590
rect 12068 7588 12092 7590
rect 11702 7576 11758 7585
rect 11852 7568 12148 7588
rect 12346 7576 12402 7585
rect 11702 7511 11758 7520
rect 12256 7540 12308 7546
rect 11532 7410 11652 7426
rect 11520 7404 11652 7410
rect 11572 7398 11652 7404
rect 11520 7346 11572 7352
rect 11624 6866 11652 7398
rect 11716 7342 11744 7511
rect 12728 7562 12756 10503
rect 12900 9920 12952 9926
rect 13004 9897 13032 10542
rect 12900 9862 12952 9868
rect 12990 9888 13046 9897
rect 12912 9722 12940 9862
rect 12990 9823 13046 9832
rect 12900 9716 12952 9722
rect 12900 9658 12952 9664
rect 12898 9480 12954 9489
rect 13004 9450 13032 9823
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 12898 9415 12954 9424
rect 12992 9444 13044 9450
rect 12912 9110 12940 9415
rect 12992 9386 13044 9392
rect 13096 9382 13124 9590
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13004 8498 13032 8774
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8022 13032 8434
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12992 8016 13044 8022
rect 12992 7958 13044 7964
rect 13096 7750 13124 8366
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 12346 7511 12402 7520
rect 12636 7534 12756 7562
rect 12256 7482 12308 7488
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 12164 7336 12216 7342
rect 12268 7313 12296 7482
rect 12360 7342 12388 7511
rect 12348 7336 12400 7342
rect 12164 7278 12216 7284
rect 12254 7304 12310 7313
rect 12176 7154 12204 7278
rect 12348 7278 12400 7284
rect 12254 7239 12310 7248
rect 12636 7206 12664 7534
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12728 7206 12756 7414
rect 13004 7410 13032 7686
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 12808 7336 12860 7342
rect 13188 7324 13216 13144
rect 13372 13002 13400 15943
rect 13544 15914 13596 15920
rect 13924 15706 13952 15982
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 14016 15638 14044 16526
rect 14108 16250 14136 17614
rect 14200 17270 14228 18158
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14280 17264 14332 17270
rect 14280 17206 14332 17212
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14200 16726 14228 17070
rect 14188 16720 14240 16726
rect 14188 16662 14240 16668
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14094 16144 14150 16153
rect 14094 16079 14150 16088
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13912 15564 13964 15570
rect 13912 15506 13964 15512
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 13740 13530 13768 13806
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13280 12974 13400 13002
rect 13280 8265 13308 12974
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 13726 12200 13782 12209
rect 13726 12135 13782 12144
rect 13740 11694 13768 12135
rect 13832 11898 13860 12310
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13542 9888 13598 9897
rect 13542 9823 13598 9832
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13372 9194 13400 9386
rect 13372 9178 13492 9194
rect 13372 9172 13504 9178
rect 13372 9166 13452 9172
rect 13266 8256 13322 8265
rect 13266 8191 13322 8200
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 12808 7278 12860 7284
rect 13096 7296 13216 7324
rect 12624 7200 12676 7206
rect 12176 7126 12572 7154
rect 12624 7142 12676 7148
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12268 7002 12388 7018
rect 12256 6996 12388 7002
rect 12308 6990 12388 6996
rect 12256 6938 12308 6944
rect 12164 6928 12216 6934
rect 12070 6896 12126 6905
rect 11612 6860 11664 6866
rect 12164 6870 12216 6876
rect 12070 6831 12126 6840
rect 11612 6802 11664 6808
rect 12084 6798 12112 6831
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 11852 6556 12148 6576
rect 11908 6554 11932 6556
rect 11988 6554 12012 6556
rect 12068 6554 12092 6556
rect 11930 6502 11932 6554
rect 11994 6502 12006 6554
rect 12068 6502 12070 6554
rect 11908 6500 11932 6502
rect 11988 6500 12012 6502
rect 12068 6500 12092 6502
rect 11852 6480 12148 6500
rect 11704 6452 11756 6458
rect 11704 6394 11756 6400
rect 11716 6254 11744 6394
rect 11794 6352 11850 6361
rect 11794 6287 11796 6296
rect 11848 6287 11850 6296
rect 11796 6258 11848 6264
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11520 6180 11572 6186
rect 11520 6122 11572 6128
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11532 4706 11560 6122
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11716 5370 11744 5714
rect 11852 5468 12148 5488
rect 11908 5466 11932 5468
rect 11988 5466 12012 5468
rect 12068 5466 12092 5468
rect 11930 5414 11932 5466
rect 11994 5414 12006 5466
rect 12068 5414 12070 5466
rect 11908 5412 11932 5414
rect 11988 5412 12012 5414
rect 12068 5412 12092 5414
rect 11852 5392 12148 5412
rect 11704 5364 11756 5370
rect 11704 5306 11756 5312
rect 11716 4826 11744 5306
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11532 4690 11652 4706
rect 11532 4684 11664 4690
rect 11532 4678 11612 4684
rect 11532 4146 11560 4678
rect 11612 4626 11664 4632
rect 12176 4570 12204 6870
rect 12256 6860 12308 6866
rect 12256 6802 12308 6808
rect 12268 6458 12296 6802
rect 12360 6769 12388 6990
rect 12544 6798 12572 7126
rect 12532 6792 12584 6798
rect 12346 6760 12402 6769
rect 12532 6734 12584 6740
rect 12346 6695 12402 6704
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12256 5840 12308 5846
rect 12254 5808 12256 5817
rect 12440 5840 12492 5846
rect 12308 5808 12310 5817
rect 12440 5782 12492 5788
rect 12254 5743 12310 5752
rect 12348 5568 12400 5574
rect 12348 5510 12400 5516
rect 12360 5098 12388 5510
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12360 4690 12388 5034
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12176 4542 12296 4570
rect 12268 4486 12296 4542
rect 12256 4480 12308 4486
rect 12256 4422 12308 4428
rect 11852 4380 12148 4400
rect 11908 4378 11932 4380
rect 11988 4378 12012 4380
rect 12068 4378 12092 4380
rect 11930 4326 11932 4378
rect 11994 4326 12006 4378
rect 12068 4326 12070 4378
rect 11908 4324 11932 4326
rect 11988 4324 12012 4326
rect 12068 4324 12092 4326
rect 11852 4304 12148 4324
rect 11520 4140 11572 4146
rect 11520 4082 11572 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 11336 3936 11388 3942
rect 11336 3878 11388 3884
rect 11428 3936 11480 3942
rect 11428 3878 11480 3884
rect 8220 3836 8516 3856
rect 8276 3834 8300 3836
rect 8356 3834 8380 3836
rect 8436 3834 8460 3836
rect 8298 3782 8300 3834
rect 8362 3782 8374 3834
rect 8436 3782 8438 3834
rect 8276 3780 8300 3782
rect 8356 3780 8380 3782
rect 8436 3780 8460 3782
rect 8220 3760 8516 3780
rect 11440 3670 11468 3878
rect 11900 3670 11928 4082
rect 12254 3904 12310 3913
rect 12254 3839 12310 3848
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 12268 3398 12296 3839
rect 12452 3602 12480 5782
rect 12636 5778 12664 7142
rect 12728 6934 12756 7142
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12820 5642 12848 7278
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12912 6458 12940 6802
rect 13096 6662 13124 7296
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13188 6730 13216 7142
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 13084 6384 13136 6390
rect 13082 6352 13084 6361
rect 13136 6352 13138 6361
rect 13082 6287 13138 6296
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 13004 5778 13032 6054
rect 12992 5772 13044 5778
rect 12912 5732 12992 5760
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12912 5574 12940 5732
rect 12992 5714 13044 5720
rect 13188 5574 13216 6666
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12636 4622 12664 5306
rect 12912 5234 12940 5510
rect 12900 5228 12952 5234
rect 12900 5170 12952 5176
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12530 4312 12586 4321
rect 12530 4247 12586 4256
rect 12544 3670 12572 4247
rect 12820 4214 12848 4558
rect 12808 4208 12860 4214
rect 12808 4150 12860 4156
rect 12716 4072 12768 4078
rect 12714 4040 12716 4049
rect 12768 4040 12770 4049
rect 12714 3975 12770 3984
rect 13004 3738 13032 5102
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 13096 4282 13124 4490
rect 13280 4282 13308 7346
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 13268 4276 13320 4282
rect 13268 4218 13320 4224
rect 13372 4214 13400 9166
rect 13452 9114 13504 9120
rect 13452 8424 13504 8430
rect 13556 8412 13584 9823
rect 13634 9616 13690 9625
rect 13634 9551 13690 9560
rect 13504 8384 13584 8412
rect 13452 8366 13504 8372
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13556 6848 13584 7822
rect 13648 7342 13676 9551
rect 13740 9217 13768 11154
rect 13924 9353 13952 15506
rect 14016 15162 14044 15574
rect 14004 15156 14056 15162
rect 14004 15098 14056 15104
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 11801 14044 14486
rect 14002 11792 14058 11801
rect 14002 11727 14058 11736
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 14016 11218 14044 11290
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14108 11098 14136 16079
rect 14200 15162 14228 16662
rect 14292 16454 14320 17206
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 14278 16280 14334 16289
rect 14278 16215 14334 16224
rect 14292 15910 14320 16215
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14384 15570 14412 23520
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 14832 21616 14884 21622
rect 14832 21558 14884 21564
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14476 21146 14504 21490
rect 14648 21412 14700 21418
rect 14648 21354 14700 21360
rect 14464 21140 14516 21146
rect 14464 21082 14516 21088
rect 14556 21004 14608 21010
rect 14556 20946 14608 20952
rect 14462 20496 14518 20505
rect 14462 20431 14518 20440
rect 14476 18698 14504 20431
rect 14464 18692 14516 18698
rect 14464 18634 14516 18640
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14200 11778 14228 14826
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14292 11898 14320 12582
rect 14384 12442 14412 13398
rect 14372 12436 14424 12442
rect 14372 12378 14424 12384
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14200 11750 14320 11778
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14016 11070 14136 11098
rect 14016 11014 14044 11070
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10538 14136 10950
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14108 10266 14136 10474
rect 14200 10305 14228 11290
rect 14186 10296 14242 10305
rect 14096 10260 14148 10266
rect 14186 10231 14242 10240
rect 14096 10202 14148 10208
rect 14200 10062 14228 10231
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 13910 9344 13966 9353
rect 13910 9279 13966 9288
rect 13726 9208 13782 9217
rect 13726 9143 13782 9152
rect 14186 9208 14242 9217
rect 14186 9143 14242 9152
rect 14096 8900 14148 8906
rect 14096 8842 14148 8848
rect 14108 8430 14136 8842
rect 14200 8838 14228 9143
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 13728 8288 13780 8294
rect 13726 8256 13728 8265
rect 13780 8256 13782 8265
rect 13726 8191 13782 8200
rect 13820 7744 13872 7750
rect 13726 7712 13782 7721
rect 13820 7686 13872 7692
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13726 7647 13782 7656
rect 13740 7449 13768 7647
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13636 6860 13688 6866
rect 13556 6820 13636 6848
rect 13688 6820 13768 6848
rect 13636 6802 13688 6808
rect 13740 6118 13768 6820
rect 13832 6746 13860 7686
rect 13924 7478 13952 7686
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 14002 7440 14058 7449
rect 14292 7392 14320 11750
rect 14476 11694 14504 18362
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14462 11520 14518 11529
rect 14462 11455 14518 11464
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14384 10198 14412 10406
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14384 8974 14412 9454
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14384 7449 14412 8910
rect 14002 7375 14058 7384
rect 14016 7342 14044 7375
rect 14200 7364 14320 7392
rect 14370 7440 14426 7449
rect 14370 7375 14426 7384
rect 14004 7336 14056 7342
rect 14004 7278 14056 7284
rect 13832 6718 13952 6746
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13832 6186 13860 6598
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 13464 4078 13492 4966
rect 13556 4826 13584 4966
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13740 4758 13768 6054
rect 13924 5914 13952 6718
rect 14096 6384 14148 6390
rect 14016 6332 14096 6338
rect 14200 6361 14228 7364
rect 14016 6326 14148 6332
rect 14186 6352 14242 6361
rect 14016 6310 14136 6326
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 13832 5794 13860 5850
rect 14016 5794 14044 6310
rect 14186 6287 14242 6296
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 14094 6216 14150 6225
rect 14094 6151 14150 6160
rect 14188 6180 14240 6186
rect 13832 5766 14044 5794
rect 13912 5296 13964 5302
rect 13912 5238 13964 5244
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13924 4570 13952 5238
rect 13740 4554 13952 4570
rect 13728 4548 13952 4554
rect 13780 4542 13952 4548
rect 13728 4490 13780 4496
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13556 4146 13584 4218
rect 13818 4176 13874 4185
rect 13544 4140 13596 4146
rect 13818 4111 13874 4120
rect 13544 4082 13596 4088
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13176 4004 13228 4010
rect 13176 3946 13228 3952
rect 13188 3738 13216 3946
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13176 3732 13228 3738
rect 13176 3674 13228 3680
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 13636 3528 13688 3534
rect 12438 3496 12494 3505
rect 13636 3470 13688 3476
rect 12438 3431 12440 3440
rect 12492 3431 12494 3440
rect 12440 3402 12492 3408
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 11852 3292 12148 3312
rect 11908 3290 11932 3292
rect 11988 3290 12012 3292
rect 12068 3290 12092 3292
rect 11930 3238 11932 3290
rect 11994 3238 12006 3290
rect 12068 3238 12070 3290
rect 11908 3236 11932 3238
rect 11988 3236 12012 3238
rect 12068 3236 12092 3238
rect 11852 3216 12148 3236
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 13648 3074 13676 3470
rect 13740 3194 13768 3878
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13648 3058 13768 3074
rect 6920 3052 6972 3058
rect 13648 3052 13780 3058
rect 13648 3046 13728 3052
rect 6920 2994 6972 3000
rect 13728 2994 13780 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3988 480 4016 2926
rect 12164 2848 12216 2854
rect 12164 2790 12216 2796
rect 8220 2748 8516 2768
rect 8276 2746 8300 2748
rect 8356 2746 8380 2748
rect 8436 2746 8460 2748
rect 8298 2694 8300 2746
rect 8362 2694 8374 2746
rect 8436 2694 8438 2746
rect 8276 2692 8300 2694
rect 8356 2692 8380 2694
rect 8436 2692 8460 2694
rect 8220 2672 8516 2692
rect 4588 2204 4884 2224
rect 4644 2202 4668 2204
rect 4724 2202 4748 2204
rect 4804 2202 4828 2204
rect 4666 2150 4668 2202
rect 4730 2150 4742 2202
rect 4804 2150 4806 2202
rect 4644 2148 4668 2150
rect 4724 2148 4748 2150
rect 4804 2148 4828 2150
rect 4588 2128 4884 2148
rect 11852 2204 12148 2224
rect 11908 2202 11932 2204
rect 11988 2202 12012 2204
rect 12068 2202 12092 2204
rect 11930 2150 11932 2202
rect 11994 2150 12006 2202
rect 12068 2150 12070 2202
rect 11908 2148 11932 2150
rect 11988 2148 12012 2150
rect 12068 2148 12092 2150
rect 11852 2128 12148 2148
rect 12176 1442 12204 2790
rect 13740 2428 13768 2994
rect 13832 2650 13860 4111
rect 13912 3664 13964 3670
rect 13912 3606 13964 3612
rect 13924 3233 13952 3606
rect 13910 3224 13966 3233
rect 13910 3159 13966 3168
rect 14108 2990 14136 6151
rect 14188 6122 14240 6128
rect 14200 4486 14228 6122
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14292 3466 14320 6258
rect 14476 6202 14504 11455
rect 14568 11234 14596 20946
rect 14660 20505 14688 21354
rect 14740 20528 14792 20534
rect 14646 20496 14702 20505
rect 14740 20470 14792 20476
rect 14646 20431 14702 20440
rect 14660 19854 14688 20431
rect 14648 19848 14700 19854
rect 14648 19790 14700 19796
rect 14752 19718 14780 20470
rect 14844 19922 14872 21558
rect 14936 21146 14964 21966
rect 14924 21140 14976 21146
rect 14924 21082 14976 21088
rect 14924 20392 14976 20398
rect 15016 20392 15068 20398
rect 14924 20334 14976 20340
rect 15014 20360 15016 20369
rect 15068 20360 15070 20369
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14660 18426 14688 19178
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14752 17678 14780 18770
rect 14936 18766 14964 20334
rect 15014 20295 15070 20304
rect 14924 18760 14976 18766
rect 14924 18702 14976 18708
rect 14936 18086 14964 18702
rect 14924 18080 14976 18086
rect 15016 18080 15068 18086
rect 14924 18022 14976 18028
rect 15014 18048 15016 18057
rect 15068 18048 15070 18057
rect 14740 17672 14792 17678
rect 14792 17632 14872 17660
rect 14740 17614 14792 17620
rect 14648 17536 14700 17542
rect 14648 17478 14700 17484
rect 14660 16561 14688 17478
rect 14844 17377 14872 17632
rect 14830 17368 14886 17377
rect 14830 17303 14886 17312
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14646 16552 14702 16561
rect 14646 16487 14702 16496
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14660 12238 14688 14418
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14752 11529 14780 17002
rect 14844 16590 14872 17303
rect 14936 17134 14964 18022
rect 15014 17983 15070 17992
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14936 15502 14964 17070
rect 15028 16153 15056 17614
rect 15014 16144 15070 16153
rect 15014 16079 15070 16088
rect 15016 16040 15068 16046
rect 15014 16008 15016 16017
rect 15068 16008 15070 16017
rect 15014 15943 15070 15952
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 15028 15434 15056 15846
rect 15016 15428 15068 15434
rect 15016 15370 15068 15376
rect 15016 14952 15068 14958
rect 14844 14912 15016 14940
rect 14844 12481 14872 14912
rect 15016 14894 15068 14900
rect 15120 14550 15148 23520
rect 15764 22794 15792 23520
rect 15304 22766 15792 22794
rect 15198 20768 15254 20777
rect 15198 20703 15254 20712
rect 15212 20398 15240 20703
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15212 20058 15240 20334
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15198 19544 15254 19553
rect 15198 19479 15254 19488
rect 15212 19446 15240 19479
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15212 16998 15240 18090
rect 15200 16992 15252 16998
rect 15200 16934 15252 16940
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15212 14074 15240 15506
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15304 13954 15332 22766
rect 15948 21542 16344 21570
rect 15948 21350 15976 21542
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 15396 20058 15424 21286
rect 15484 21244 15780 21264
rect 15540 21242 15564 21244
rect 15620 21242 15644 21244
rect 15700 21242 15724 21244
rect 15562 21190 15564 21242
rect 15626 21190 15638 21242
rect 15700 21190 15702 21242
rect 15540 21188 15564 21190
rect 15620 21188 15644 21190
rect 15700 21188 15724 21190
rect 15484 21168 15780 21188
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15488 20398 15516 20742
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15484 20156 15780 20176
rect 15540 20154 15564 20156
rect 15620 20154 15644 20156
rect 15700 20154 15724 20156
rect 15562 20102 15564 20154
rect 15626 20102 15638 20154
rect 15700 20102 15702 20154
rect 15540 20100 15564 20102
rect 15620 20100 15644 20102
rect 15700 20100 15724 20102
rect 15484 20080 15780 20100
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15568 19848 15620 19854
rect 15620 19808 15700 19836
rect 15568 19790 15620 19796
rect 15672 19281 15700 19808
rect 15658 19272 15714 19281
rect 15658 19207 15714 19216
rect 15384 19168 15436 19174
rect 15384 19110 15436 19116
rect 15396 17066 15424 19110
rect 15484 19068 15780 19088
rect 15540 19066 15564 19068
rect 15620 19066 15644 19068
rect 15700 19066 15724 19068
rect 15562 19014 15564 19066
rect 15626 19014 15638 19066
rect 15700 19014 15702 19066
rect 15540 19012 15564 19014
rect 15620 19012 15644 19014
rect 15700 19012 15724 19014
rect 15484 18992 15780 19012
rect 15484 17980 15780 18000
rect 15540 17978 15564 17980
rect 15620 17978 15644 17980
rect 15700 17978 15724 17980
rect 15562 17926 15564 17978
rect 15626 17926 15638 17978
rect 15700 17926 15702 17978
rect 15540 17924 15564 17926
rect 15620 17924 15644 17926
rect 15700 17924 15724 17926
rect 15484 17904 15780 17924
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15484 16892 15780 16912
rect 15540 16890 15564 16892
rect 15620 16890 15644 16892
rect 15700 16890 15724 16892
rect 15562 16838 15564 16890
rect 15626 16838 15638 16890
rect 15700 16838 15702 16890
rect 15540 16836 15564 16838
rect 15620 16836 15644 16838
rect 15700 16836 15724 16838
rect 15484 16816 15780 16836
rect 15474 16688 15530 16697
rect 15474 16623 15530 16632
rect 15488 16454 15516 16623
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15484 15804 15780 15824
rect 15540 15802 15564 15804
rect 15620 15802 15644 15804
rect 15700 15802 15724 15804
rect 15562 15750 15564 15802
rect 15626 15750 15638 15802
rect 15700 15750 15702 15802
rect 15540 15748 15564 15750
rect 15620 15748 15644 15750
rect 15700 15748 15724 15750
rect 15484 15728 15780 15748
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15580 15162 15608 15506
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15396 14822 15424 15098
rect 15750 15056 15806 15065
rect 15750 14991 15752 15000
rect 15804 14991 15806 15000
rect 15752 14962 15804 14968
rect 15384 14816 15436 14822
rect 15384 14758 15436 14764
rect 15212 13926 15332 13954
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14936 12646 14964 12786
rect 15016 12708 15068 12714
rect 15016 12650 15068 12656
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14830 12472 14886 12481
rect 14830 12407 14886 12416
rect 14738 11520 14794 11529
rect 14738 11455 14794 11464
rect 14568 11206 14780 11234
rect 14648 11076 14700 11082
rect 14648 11018 14700 11024
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14568 9518 14596 10950
rect 14660 9586 14688 11018
rect 14752 10554 14780 11206
rect 14844 10674 14872 12407
rect 14936 11762 14964 12582
rect 15028 12186 15056 12650
rect 15120 12374 15148 13806
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15212 12322 15240 13926
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12424 15332 13126
rect 15396 12753 15424 14758
rect 15484 14716 15780 14736
rect 15540 14714 15564 14716
rect 15620 14714 15644 14716
rect 15700 14714 15724 14716
rect 15562 14662 15564 14714
rect 15626 14662 15638 14714
rect 15700 14662 15702 14714
rect 15540 14660 15564 14662
rect 15620 14660 15644 14662
rect 15700 14660 15724 14662
rect 15484 14640 15780 14660
rect 15484 13628 15780 13648
rect 15540 13626 15564 13628
rect 15620 13626 15644 13628
rect 15700 13626 15724 13628
rect 15562 13574 15564 13626
rect 15626 13574 15638 13626
rect 15700 13574 15702 13626
rect 15540 13572 15564 13574
rect 15620 13572 15644 13574
rect 15700 13572 15724 13574
rect 15484 13552 15780 13572
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15476 12776 15528 12782
rect 15382 12744 15438 12753
rect 15764 12764 15792 13330
rect 15856 12889 15884 19926
rect 15948 18902 15976 19994
rect 15936 18896 15988 18902
rect 15936 18838 15988 18844
rect 15936 18624 15988 18630
rect 15936 18566 15988 18572
rect 15948 16658 15976 18566
rect 16040 17814 16068 21286
rect 16120 21004 16172 21010
rect 16120 20946 16172 20952
rect 16132 20534 16160 20946
rect 16120 20528 16172 20534
rect 16120 20470 16172 20476
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 18329 16160 19110
rect 16118 18320 16174 18329
rect 16118 18255 16174 18264
rect 16120 18080 16172 18086
rect 16120 18022 16172 18028
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16132 17066 16160 18022
rect 16120 17060 16172 17066
rect 16120 17002 16172 17008
rect 16224 16810 16252 21422
rect 16040 16782 16252 16810
rect 15936 16652 15988 16658
rect 15936 16594 15988 16600
rect 15936 15156 15988 15162
rect 15936 15098 15988 15104
rect 15948 14482 15976 15098
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15842 12880 15898 12889
rect 15842 12815 15898 12824
rect 15528 12736 15792 12764
rect 15476 12718 15528 12724
rect 15382 12679 15438 12688
rect 15764 12628 15792 12736
rect 15844 12640 15896 12646
rect 15764 12600 15844 12628
rect 15844 12582 15896 12588
rect 15484 12540 15780 12560
rect 15540 12538 15564 12540
rect 15620 12538 15644 12540
rect 15700 12538 15724 12540
rect 15562 12486 15564 12538
rect 15626 12486 15638 12538
rect 15700 12486 15702 12538
rect 15540 12484 15564 12486
rect 15620 12484 15644 12486
rect 15700 12484 15724 12486
rect 15484 12464 15780 12484
rect 15304 12396 15516 12424
rect 15212 12294 15332 12322
rect 15200 12232 15252 12238
rect 15028 12180 15200 12186
rect 15028 12174 15252 12180
rect 15028 12158 15240 12174
rect 15106 12064 15162 12073
rect 15106 11999 15162 12008
rect 15016 11824 15068 11830
rect 15014 11792 15016 11801
rect 15068 11792 15070 11801
rect 14924 11756 14976 11762
rect 15014 11727 15070 11736
rect 14924 11698 14976 11704
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14936 11082 14964 11562
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14752 10526 14872 10554
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14752 9518 14780 9862
rect 14844 9625 14872 10526
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9654 14964 9862
rect 14924 9648 14976 9654
rect 14830 9616 14886 9625
rect 14924 9590 14976 9596
rect 14830 9551 14886 9560
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14568 9110 14596 9318
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14568 8498 14596 8910
rect 14660 8566 14688 9114
rect 14648 8560 14700 8566
rect 14648 8502 14700 8508
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14648 8424 14700 8430
rect 14752 8401 14780 9318
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14648 8366 14700 8372
rect 14738 8392 14794 8401
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7206 14596 8230
rect 14660 7954 14688 8366
rect 14844 8362 14872 8910
rect 14738 8327 14794 8336
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14752 7818 14780 8026
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14384 6174 14504 6202
rect 14384 5817 14412 6174
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14370 5808 14426 5817
rect 14476 5778 14504 6054
rect 14370 5743 14426 5752
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 14384 5098 14412 5510
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 14384 4826 14412 5034
rect 14476 4826 14504 5714
rect 14660 4826 14688 6598
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4820 14516 4826
rect 14464 4762 14516 4768
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14384 4078 14412 4422
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14372 4072 14424 4078
rect 14372 4014 14424 4020
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14280 2984 14332 2990
rect 14384 2972 14412 4014
rect 14568 4010 14596 4218
rect 14556 4004 14608 4010
rect 14556 3946 14608 3952
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14646 3632 14702 3641
rect 14332 2944 14412 2972
rect 14280 2926 14332 2932
rect 14568 2650 14596 3606
rect 14646 3567 14648 3576
rect 14700 3567 14702 3576
rect 14648 3538 14700 3544
rect 13820 2644 13872 2650
rect 13820 2586 13872 2592
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14648 2576 14700 2582
rect 14752 2564 14780 7346
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14844 6322 14872 7142
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14844 3534 14872 5646
rect 14936 4865 14964 9046
rect 15028 5302 15056 11630
rect 15120 11218 15148 11999
rect 15304 11665 15332 12294
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15290 11656 15346 11665
rect 15290 11591 15346 11600
rect 15396 11558 15424 11834
rect 15488 11762 15516 12396
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 12102 15700 12242
rect 15948 12238 15976 14282
rect 16040 13025 16068 16782
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16132 16114 16160 16526
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16120 15972 16172 15978
rect 16120 15914 16172 15920
rect 16132 14657 16160 15914
rect 16118 14648 16174 14657
rect 16118 14583 16174 14592
rect 16120 14272 16172 14278
rect 16118 14240 16120 14249
rect 16172 14240 16174 14249
rect 16118 14175 16174 14184
rect 16224 13818 16252 16594
rect 16316 16130 16344 21542
rect 16396 21480 16448 21486
rect 16396 21422 16448 21428
rect 16408 20534 16436 21422
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 17882 16436 20198
rect 16500 20058 16528 23520
rect 17236 22302 17264 23520
rect 17880 22370 17908 23520
rect 17868 22364 17920 22370
rect 17868 22306 17920 22312
rect 17224 22296 17276 22302
rect 17224 22238 17276 22244
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16592 21146 16620 22170
rect 18616 21962 18644 23520
rect 19352 22658 19380 23520
rect 19430 23488 19486 23497
rect 19430 23423 19486 23432
rect 19444 22846 19472 23423
rect 19432 22840 19484 22846
rect 19432 22782 19484 22788
rect 19614 22808 19670 22817
rect 19996 22794 20024 23520
rect 19614 22743 19670 22752
rect 19904 22766 20024 22794
rect 19352 22630 19564 22658
rect 19340 22228 19392 22234
rect 19340 22170 19392 22176
rect 19352 22137 19380 22170
rect 19338 22128 19394 22137
rect 19338 22063 19394 22072
rect 18604 21956 18656 21962
rect 18604 21898 18656 21904
rect 19116 21788 19412 21808
rect 19172 21786 19196 21788
rect 19252 21786 19276 21788
rect 19332 21786 19356 21788
rect 19194 21734 19196 21786
rect 19258 21734 19270 21786
rect 19332 21734 19334 21786
rect 19172 21732 19196 21734
rect 19252 21732 19276 21734
rect 19332 21732 19356 21734
rect 19116 21712 19412 21732
rect 17316 21684 17368 21690
rect 17316 21626 17368 21632
rect 17224 21412 17276 21418
rect 17224 21354 17276 21360
rect 16856 21344 16908 21350
rect 16856 21286 16908 21292
rect 17132 21344 17184 21350
rect 17132 21286 17184 21292
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16764 21072 16816 21078
rect 16764 21014 16816 21020
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16580 19712 16632 19718
rect 16580 19654 16632 19660
rect 16488 18964 16540 18970
rect 16488 18906 16540 18912
rect 16500 17882 16528 18906
rect 16592 18834 16620 19654
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16672 18624 16724 18630
rect 16672 18566 16724 18572
rect 16684 18426 16712 18566
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16670 18184 16726 18193
rect 16670 18119 16726 18128
rect 16684 18086 16712 18119
rect 16672 18080 16724 18086
rect 16672 18022 16724 18028
rect 16396 17876 16448 17882
rect 16396 17818 16448 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16408 16289 16436 16526
rect 16394 16280 16450 16289
rect 16394 16215 16450 16224
rect 16316 16102 16436 16130
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16132 13790 16252 13818
rect 16026 13016 16082 13025
rect 16026 12951 16082 12960
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15764 11937 15792 12174
rect 15750 11928 15806 11937
rect 15750 11863 15806 11872
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15764 11626 15792 11863
rect 16026 11656 16082 11665
rect 15752 11620 15804 11626
rect 16026 11591 16082 11600
rect 15752 11562 15804 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15484 11452 15780 11472
rect 15540 11450 15564 11452
rect 15620 11450 15644 11452
rect 15700 11450 15724 11452
rect 15562 11398 15564 11450
rect 15626 11398 15638 11450
rect 15700 11398 15702 11450
rect 15540 11396 15564 11398
rect 15620 11396 15644 11398
rect 15700 11396 15724 11398
rect 15484 11376 15780 11396
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15384 11144 15436 11150
rect 15382 11112 15384 11121
rect 15436 11112 15438 11121
rect 15382 11047 15438 11056
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15290 10976 15346 10985
rect 15120 10742 15148 10950
rect 15290 10911 15346 10920
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15304 10606 15332 10911
rect 15856 10674 15884 11494
rect 15934 10704 15990 10713
rect 15844 10668 15896 10674
rect 15934 10639 15990 10648
rect 15844 10610 15896 10616
rect 15292 10600 15344 10606
rect 15292 10542 15344 10548
rect 15948 10470 15976 10639
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15108 9988 15160 9994
rect 15108 9930 15160 9936
rect 15120 6905 15148 9930
rect 15212 8922 15240 10406
rect 15484 10364 15780 10384
rect 15540 10362 15564 10364
rect 15620 10362 15644 10364
rect 15700 10362 15724 10364
rect 15562 10310 15564 10362
rect 15626 10310 15638 10362
rect 15700 10310 15702 10362
rect 15540 10308 15564 10310
rect 15620 10308 15644 10310
rect 15700 10308 15724 10310
rect 15484 10288 15780 10308
rect 15382 10160 15438 10169
rect 15292 10124 15344 10130
rect 15382 10095 15384 10104
rect 15292 10066 15344 10072
rect 15436 10095 15438 10104
rect 15384 10066 15436 10072
rect 15304 10033 15332 10066
rect 15290 10024 15346 10033
rect 15290 9959 15346 9968
rect 15948 9353 15976 10406
rect 15934 9344 15990 9353
rect 15484 9276 15780 9296
rect 15934 9279 15990 9288
rect 15540 9274 15564 9276
rect 15620 9274 15644 9276
rect 15700 9274 15724 9276
rect 15562 9222 15564 9274
rect 15626 9222 15638 9274
rect 15700 9222 15702 9274
rect 15540 9220 15564 9222
rect 15620 9220 15644 9222
rect 15700 9220 15724 9222
rect 15484 9200 15780 9220
rect 15476 9104 15528 9110
rect 15304 9052 15476 9058
rect 15304 9046 15528 9052
rect 15304 9042 15516 9046
rect 15292 9036 15516 9042
rect 15344 9030 15516 9036
rect 15292 8978 15344 8984
rect 15844 8968 15896 8974
rect 15212 8906 15516 8922
rect 15844 8910 15896 8916
rect 15212 8900 15528 8906
rect 15212 8894 15476 8900
rect 15476 8842 15528 8848
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15304 8634 15332 8774
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15396 8498 15424 8570
rect 15384 8492 15436 8498
rect 15212 8452 15384 8480
rect 15212 8294 15240 8452
rect 15384 8434 15436 8440
rect 15200 8288 15252 8294
rect 15488 8276 15516 8842
rect 15200 8230 15252 8236
rect 15396 8248 15516 8276
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15120 6322 15148 6831
rect 15212 6798 15240 7822
rect 15396 7585 15424 8248
rect 15484 8188 15780 8208
rect 15540 8186 15564 8188
rect 15620 8186 15644 8188
rect 15700 8186 15724 8188
rect 15562 8134 15564 8186
rect 15626 8134 15638 8186
rect 15700 8134 15702 8186
rect 15540 8132 15564 8134
rect 15620 8132 15644 8134
rect 15700 8132 15724 8134
rect 15484 8112 15780 8132
rect 15856 8022 15884 8910
rect 15948 8634 15976 9279
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15844 8016 15896 8022
rect 15844 7958 15896 7964
rect 15382 7576 15438 7585
rect 15382 7511 15438 7520
rect 15948 7478 15976 8366
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 15936 7472 15988 7478
rect 15936 7414 15988 7420
rect 15488 7313 15516 7414
rect 15474 7304 15530 7313
rect 15474 7239 15530 7248
rect 15484 7100 15780 7120
rect 15540 7098 15564 7100
rect 15620 7098 15644 7100
rect 15700 7098 15724 7100
rect 15562 7046 15564 7098
rect 15626 7046 15638 7098
rect 15700 7046 15702 7098
rect 15540 7044 15564 7046
rect 15620 7044 15644 7046
rect 15700 7044 15724 7046
rect 15484 7024 15780 7044
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15108 6316 15160 6322
rect 15108 6258 15160 6264
rect 15108 6112 15160 6118
rect 15108 6054 15160 6060
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 14922 4856 14978 4865
rect 14922 4791 14978 4800
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14936 4486 14964 4694
rect 15028 4554 15056 4966
rect 15120 4690 15148 6054
rect 15212 5166 15240 6734
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 15212 4758 15240 5102
rect 15200 4752 15252 4758
rect 15200 4694 15252 4700
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14936 3534 14964 4422
rect 15108 3936 15160 3942
rect 15212 3913 15240 4558
rect 15108 3878 15160 3884
rect 15198 3904 15254 3913
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14700 2536 14780 2564
rect 14648 2518 14700 2524
rect 15028 2514 15056 3538
rect 15120 2922 15148 3878
rect 15198 3839 15254 3848
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 13912 2440 13964 2446
rect 13740 2400 13912 2428
rect 13740 2106 13768 2400
rect 13912 2382 13964 2388
rect 15120 2378 15148 2858
rect 15304 2582 15332 6394
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15484 6012 15780 6032
rect 15540 6010 15564 6012
rect 15620 6010 15644 6012
rect 15700 6010 15724 6012
rect 15562 5958 15564 6010
rect 15626 5958 15638 6010
rect 15700 5958 15702 6010
rect 15540 5956 15564 5958
rect 15620 5956 15644 5958
rect 15700 5956 15724 5958
rect 15484 5936 15780 5956
rect 15948 5778 15976 6122
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 15568 5092 15620 5098
rect 15396 5052 15568 5080
rect 15396 3505 15424 5052
rect 15568 5034 15620 5040
rect 15484 4924 15780 4944
rect 15540 4922 15564 4924
rect 15620 4922 15644 4924
rect 15700 4922 15724 4924
rect 15562 4870 15564 4922
rect 15626 4870 15638 4922
rect 15700 4870 15702 4922
rect 15540 4868 15564 4870
rect 15620 4868 15644 4870
rect 15700 4868 15724 4870
rect 15484 4848 15780 4868
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15948 3924 15976 4082
rect 16040 4049 16068 11591
rect 16132 6458 16160 13790
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13326 16252 13670
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16224 12782 16252 13262
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12306 16252 12582
rect 16316 12442 16344 15982
rect 16408 13161 16436 16102
rect 16500 15978 16528 17002
rect 16776 16674 16804 21014
rect 16868 20777 16896 21286
rect 16948 20800 17000 20806
rect 16854 20768 16910 20777
rect 16948 20742 17000 20748
rect 16854 20703 16910 20712
rect 16854 20360 16910 20369
rect 16854 20295 16856 20304
rect 16908 20295 16910 20304
rect 16856 20266 16908 20272
rect 16960 19854 16988 20742
rect 17038 20632 17094 20641
rect 17038 20567 17094 20576
rect 17052 20369 17080 20567
rect 17038 20360 17094 20369
rect 17038 20295 17094 20304
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16960 19258 16988 19790
rect 16868 19230 16988 19258
rect 16868 19122 16896 19230
rect 16868 19094 16988 19122
rect 16854 18864 16910 18873
rect 16854 18799 16910 18808
rect 16868 18630 16896 18799
rect 16960 18698 16988 19094
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16856 18624 16908 18630
rect 16856 18566 16908 18572
rect 16856 17672 16908 17678
rect 16960 17660 16988 18634
rect 17144 18290 17172 21286
rect 17236 21146 17264 21354
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17236 19990 17264 21082
rect 17328 20466 17356 21626
rect 17684 21480 17736 21486
rect 17684 21422 17736 21428
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 17696 21146 17724 21422
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 19076 21078 19104 21422
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17224 19984 17276 19990
rect 17224 19926 17276 19932
rect 17512 19378 17540 20402
rect 17880 19446 17908 21014
rect 18328 21004 18380 21010
rect 18328 20946 18380 20952
rect 18340 20058 18368 20946
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18696 20868 18748 20874
rect 18696 20810 18748 20816
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 18052 19440 18104 19446
rect 18052 19382 18104 19388
rect 17500 19372 17552 19378
rect 17500 19314 17552 19320
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 17882 17264 18226
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17040 17808 17092 17814
rect 17040 17750 17092 17756
rect 16908 17632 16988 17660
rect 16856 17614 16908 17620
rect 16868 17134 16896 17614
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 17052 16998 17080 17750
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 16684 16646 16804 16674
rect 16856 16652 16908 16658
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 16500 14822 16528 15574
rect 16488 14816 16540 14822
rect 16488 14758 16540 14764
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 13870 16528 14418
rect 16488 13864 16540 13870
rect 16488 13806 16540 13812
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16500 13462 16528 13670
rect 16592 13530 16620 15846
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16488 13456 16540 13462
rect 16488 13398 16540 13404
rect 16394 13152 16450 13161
rect 16394 13087 16450 13096
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16408 12322 16436 12378
rect 16316 12306 16436 12322
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16304 12300 16436 12306
rect 16356 12294 16436 12300
rect 16304 12242 16356 12248
rect 16210 11656 16266 11665
rect 16210 11591 16266 11600
rect 16224 9450 16252 11591
rect 16592 11558 16620 12786
rect 16304 11552 16356 11558
rect 16488 11552 16540 11558
rect 16304 11494 16356 11500
rect 16408 11512 16488 11540
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16316 9178 16344 11494
rect 16408 9654 16436 11512
rect 16488 11494 16540 11500
rect 16580 11552 16632 11558
rect 16580 11494 16632 11500
rect 16592 11354 16620 11494
rect 16684 11370 16712 16646
rect 16856 16594 16908 16600
rect 16868 16250 16896 16594
rect 16856 16244 16908 16250
rect 16856 16186 16908 16192
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16776 12306 16804 12854
rect 16764 12300 16816 12306
rect 16764 12242 16816 12248
rect 16776 11830 16804 12242
rect 16868 12186 16896 15302
rect 16960 13530 16988 15370
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16868 12158 16988 12186
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16764 11824 16816 11830
rect 16764 11766 16816 11772
rect 16580 11348 16632 11354
rect 16684 11342 16804 11370
rect 16580 11290 16632 11296
rect 16672 11212 16724 11218
rect 16672 11154 16724 11160
rect 16488 11076 16540 11082
rect 16488 11018 16540 11024
rect 16500 10266 16528 11018
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 16488 10260 16540 10266
rect 16488 10202 16540 10208
rect 16396 9648 16448 9654
rect 16396 9590 16448 9596
rect 16500 9586 16528 10202
rect 16592 10033 16620 10406
rect 16578 10024 16634 10033
rect 16578 9959 16634 9968
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16592 9466 16620 9959
rect 16684 9654 16712 11154
rect 16776 10849 16804 11342
rect 16868 11234 16896 12038
rect 16960 11665 16988 12158
rect 16946 11656 17002 11665
rect 16946 11591 17002 11600
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16960 11354 16988 11494
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16868 11206 16988 11234
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16762 10840 16818 10849
rect 16762 10775 16818 10784
rect 16764 10600 16816 10606
rect 16764 10542 16816 10548
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16776 9602 16804 10542
rect 16868 10266 16896 10950
rect 16856 10260 16908 10266
rect 16856 10202 16908 10208
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16868 9722 16896 10066
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16776 9574 16896 9602
rect 16500 9438 16620 9466
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16408 9178 16436 9318
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16408 9058 16436 9114
rect 16224 9030 16436 9058
rect 16500 9042 16528 9438
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16488 9036 16540 9042
rect 16224 8430 16252 9030
rect 16488 8978 16540 8984
rect 16592 8922 16620 9318
rect 16868 9178 16896 9574
rect 16960 9518 16988 11206
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 16764 9104 16816 9110
rect 16764 9046 16816 9052
rect 16408 8906 16620 8922
rect 16396 8900 16620 8906
rect 16448 8894 16620 8900
rect 16396 8842 16448 8848
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16316 8498 16344 8570
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16212 8424 16264 8430
rect 16580 8424 16632 8430
rect 16212 8366 16264 8372
rect 16394 8392 16450 8401
rect 16224 6769 16252 8366
rect 16580 8366 16632 8372
rect 16394 8327 16450 8336
rect 16304 8016 16356 8022
rect 16304 7958 16356 7964
rect 16316 7478 16344 7958
rect 16408 7546 16436 8327
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16592 7002 16620 8366
rect 16776 8090 16804 9046
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16670 7440 16726 7449
rect 16670 7375 16726 7384
rect 16856 7404 16908 7410
rect 16580 6996 16632 7002
rect 16580 6938 16632 6944
rect 16684 6798 16712 7375
rect 16856 7346 16908 7352
rect 16672 6792 16724 6798
rect 16210 6760 16266 6769
rect 16672 6734 16724 6740
rect 16868 6730 16896 7346
rect 16948 7200 17000 7206
rect 16948 7142 17000 7148
rect 16960 6866 16988 7142
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16210 6695 16266 6704
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16120 6452 16172 6458
rect 16120 6394 16172 6400
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16316 6089 16344 6190
rect 16302 6080 16358 6089
rect 16302 6015 16358 6024
rect 16120 5704 16172 5710
rect 16316 5692 16344 6015
rect 16172 5664 16344 5692
rect 16120 5646 16172 5652
rect 16210 5400 16266 5409
rect 16210 5335 16266 5344
rect 16118 4312 16174 4321
rect 16118 4247 16174 4256
rect 16026 4040 16082 4049
rect 16132 4010 16160 4247
rect 16026 3975 16082 3984
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 15948 3896 16068 3924
rect 15484 3836 15780 3856
rect 15540 3834 15564 3836
rect 15620 3834 15644 3836
rect 15700 3834 15724 3836
rect 15562 3782 15564 3834
rect 15626 3782 15638 3834
rect 15700 3782 15702 3834
rect 15540 3780 15564 3782
rect 15620 3780 15644 3782
rect 15700 3780 15724 3782
rect 15484 3760 15780 3780
rect 15842 3632 15898 3641
rect 15568 3596 15620 3602
rect 15842 3567 15844 3576
rect 15568 3538 15620 3544
rect 15896 3567 15898 3576
rect 15844 3538 15896 3544
rect 15382 3496 15438 3505
rect 15382 3431 15438 3440
rect 15580 3126 15608 3538
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 15484 2748 15780 2768
rect 15540 2746 15564 2748
rect 15620 2746 15644 2748
rect 15700 2746 15724 2748
rect 15562 2694 15564 2746
rect 15626 2694 15638 2746
rect 15700 2694 15702 2746
rect 15540 2692 15564 2694
rect 15620 2692 15644 2694
rect 15700 2692 15724 2694
rect 15484 2672 15780 2692
rect 15948 2582 15976 3334
rect 16040 2972 16068 3896
rect 16224 3670 16252 5335
rect 16408 5098 16436 6598
rect 16868 5914 16896 6666
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 17052 5114 17080 16934
rect 17144 14958 17172 17478
rect 17500 17196 17552 17202
rect 17500 17138 17552 17144
rect 17316 15904 17368 15910
rect 17316 15846 17368 15852
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 17132 14952 17184 14958
rect 17132 14894 17184 14900
rect 17130 14784 17186 14793
rect 17130 14719 17186 14728
rect 17144 12374 17172 14719
rect 17236 13870 17264 15506
rect 17328 15366 17356 15846
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17314 15056 17370 15065
rect 17314 14991 17316 15000
rect 17368 14991 17370 15000
rect 17316 14962 17368 14968
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17328 14550 17356 14826
rect 17420 14618 17448 14894
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17316 14544 17368 14550
rect 17316 14486 17368 14492
rect 17224 13864 17276 13870
rect 17224 13806 17276 13812
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17328 12918 17356 13330
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17420 12782 17448 13466
rect 17512 12986 17540 17138
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17224 12368 17276 12374
rect 17224 12310 17276 12316
rect 17236 9489 17264 12310
rect 17328 12306 17356 12582
rect 17604 12458 17632 19314
rect 18064 18222 18092 19382
rect 18340 19378 18368 19994
rect 18328 19372 18380 19378
rect 18328 19314 18380 19320
rect 18432 19310 18460 20742
rect 18708 20466 18736 20810
rect 18984 20534 19012 20878
rect 19116 20700 19412 20720
rect 19172 20698 19196 20700
rect 19252 20698 19276 20700
rect 19332 20698 19356 20700
rect 19194 20646 19196 20698
rect 19258 20646 19270 20698
rect 19332 20646 19334 20698
rect 19172 20644 19196 20646
rect 19252 20644 19276 20646
rect 19332 20644 19356 20646
rect 19116 20624 19412 20644
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18248 18154 18276 19246
rect 18432 18902 18460 19246
rect 18420 18896 18472 18902
rect 18420 18838 18472 18844
rect 18418 18728 18474 18737
rect 18418 18663 18474 18672
rect 18432 18222 18460 18663
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 18236 18148 18288 18154
rect 18236 18090 18288 18096
rect 18432 17678 18460 18158
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17776 16516 17828 16522
rect 17776 16458 17828 16464
rect 17684 15564 17736 15570
rect 17684 15506 17736 15512
rect 17696 15162 17724 15506
rect 17684 15156 17736 15162
rect 17684 15098 17736 15104
rect 17696 14550 17724 15098
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17696 13530 17724 13670
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17696 12714 17724 13466
rect 17684 12708 17736 12714
rect 17684 12650 17736 12656
rect 17788 12594 17816 16458
rect 17880 16454 17908 17070
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17880 12850 17908 16390
rect 17972 15094 18000 17206
rect 18156 16998 18184 17614
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18144 16992 18196 16998
rect 18144 16934 18196 16940
rect 18156 16590 18184 16934
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18156 16028 18184 16526
rect 18248 16250 18276 17070
rect 18524 16402 18552 20334
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18432 16374 18552 16402
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18236 16040 18288 16046
rect 18156 16000 18236 16028
rect 18236 15982 18288 15988
rect 18052 15904 18104 15910
rect 18052 15846 18104 15852
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17972 14498 18000 15030
rect 18064 14618 18092 15846
rect 18248 15162 18276 15982
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18236 15156 18288 15162
rect 18236 15098 18288 15104
rect 18340 14958 18368 15642
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18156 14498 18184 14554
rect 17972 14470 18184 14498
rect 17960 14272 18012 14278
rect 17958 14240 17960 14249
rect 18012 14240 18014 14249
rect 17958 14175 18014 14184
rect 17960 13864 18012 13870
rect 17960 13806 18012 13812
rect 17972 13326 18000 13806
rect 18236 13796 18288 13802
rect 18236 13738 18288 13744
rect 18052 13524 18104 13530
rect 18052 13466 18104 13472
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17972 12782 18000 13262
rect 18064 12918 18092 13466
rect 18142 13424 18198 13433
rect 18248 13394 18276 13738
rect 18142 13359 18198 13368
rect 18236 13388 18288 13394
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17512 12430 17632 12458
rect 17696 12566 17816 12594
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17314 11792 17370 11801
rect 17314 11727 17370 11736
rect 17328 11694 17356 11727
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17328 11121 17356 11494
rect 17314 11112 17370 11121
rect 17314 11047 17370 11056
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10849 17356 10950
rect 17314 10840 17370 10849
rect 17314 10775 17370 10784
rect 17222 9480 17278 9489
rect 17222 9415 17278 9424
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 17144 6225 17172 8298
rect 17328 6361 17356 10775
rect 17420 10742 17448 11494
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17408 10600 17460 10606
rect 17406 10568 17408 10577
rect 17460 10568 17462 10577
rect 17406 10503 17462 10512
rect 17512 8945 17540 12430
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11762 17632 12038
rect 17592 11756 17644 11762
rect 17592 11698 17644 11704
rect 17590 11656 17646 11665
rect 17590 11591 17646 11600
rect 17498 8936 17554 8945
rect 17498 8871 17554 8880
rect 17408 6996 17460 7002
rect 17604 6984 17632 11591
rect 17460 6956 17632 6984
rect 17408 6938 17460 6944
rect 17696 6866 17724 12566
rect 17972 12306 18000 12718
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17788 11257 17816 11562
rect 18064 11558 18092 12242
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17774 11248 17830 11257
rect 17774 11183 17776 11192
rect 17828 11183 17830 11192
rect 17776 11154 17828 11160
rect 17788 11123 17816 11154
rect 18064 11150 18092 11494
rect 18156 11286 18184 13359
rect 18236 13330 18288 13336
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18144 11280 18196 11286
rect 18144 11222 18196 11228
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17776 11008 17828 11014
rect 17774 10976 17776 10985
rect 17828 10976 17830 10985
rect 17774 10911 17830 10920
rect 18052 10600 18104 10606
rect 18052 10542 18104 10548
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17788 7954 17816 8774
rect 17972 8498 18000 10202
rect 18064 8956 18092 10542
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 18156 9586 18184 9862
rect 18144 9580 18196 9586
rect 18144 9522 18196 9528
rect 18248 9178 18276 13126
rect 18326 11928 18382 11937
rect 18432 11898 18460 16374
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18524 15502 18552 15846
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18326 11863 18382 11872
rect 18420 11892 18472 11898
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18340 9042 18368 11863
rect 18420 11834 18472 11840
rect 18524 11626 18552 14554
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18418 11112 18474 11121
rect 18418 11047 18474 11056
rect 18432 10470 18460 11047
rect 18420 10464 18472 10470
rect 18420 10406 18472 10412
rect 18616 9466 18644 19858
rect 18708 18358 18736 20402
rect 18788 20256 18840 20262
rect 18788 20198 18840 20204
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18696 17536 18748 17542
rect 18696 17478 18748 17484
rect 18708 16658 18736 17478
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18800 12442 18828 20198
rect 19248 19916 19300 19922
rect 19352 19904 19380 20402
rect 19444 20398 19472 21286
rect 19536 20754 19564 22630
rect 19628 22098 19656 22743
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19536 20726 19656 20754
rect 19522 20632 19578 20641
rect 19522 20567 19578 20576
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19536 20058 19564 20567
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19628 19961 19656 20726
rect 19614 19952 19670 19961
rect 19300 19876 19472 19904
rect 19614 19887 19670 19896
rect 19248 19858 19300 19864
rect 19116 19612 19412 19632
rect 19172 19610 19196 19612
rect 19252 19610 19276 19612
rect 19332 19610 19356 19612
rect 19194 19558 19196 19610
rect 19258 19558 19270 19610
rect 19332 19558 19334 19610
rect 19172 19556 19196 19558
rect 19252 19556 19276 19558
rect 19332 19556 19356 19558
rect 19116 19536 19412 19556
rect 19444 19428 19472 19876
rect 19352 19400 19472 19428
rect 19352 19310 19380 19400
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 18880 19236 18932 19242
rect 18880 19178 18932 19184
rect 18892 18970 18920 19178
rect 19352 18970 19380 19246
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 18892 17814 18920 18906
rect 19168 18766 19196 18906
rect 19156 18760 19208 18766
rect 19154 18728 19156 18737
rect 19208 18728 19210 18737
rect 19154 18663 19210 18672
rect 19116 18524 19412 18544
rect 19172 18522 19196 18524
rect 19252 18522 19276 18524
rect 19332 18522 19356 18524
rect 19194 18470 19196 18522
rect 19258 18470 19270 18522
rect 19332 18470 19334 18522
rect 19172 18468 19196 18470
rect 19252 18468 19276 18470
rect 19332 18468 19356 18470
rect 19116 18448 19412 18468
rect 19614 18456 19670 18465
rect 19614 18391 19616 18400
rect 19668 18391 19670 18400
rect 19616 18362 19668 18368
rect 19248 18148 19300 18154
rect 19248 18090 19300 18096
rect 19260 17882 19288 18090
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 18880 17808 18932 17814
rect 18880 17750 18932 17756
rect 18972 17808 19024 17814
rect 18972 17750 19024 17756
rect 18984 17649 19012 17750
rect 18970 17640 19026 17649
rect 18970 17575 19026 17584
rect 19116 17436 19412 17456
rect 19172 17434 19196 17436
rect 19252 17434 19276 17436
rect 19332 17434 19356 17436
rect 19194 17382 19196 17434
rect 19258 17382 19270 17434
rect 19332 17382 19334 17434
rect 19172 17380 19196 17382
rect 19252 17380 19276 17382
rect 19332 17380 19356 17382
rect 19116 17360 19412 17380
rect 19720 17377 19748 21082
rect 19904 18086 19932 22766
rect 20732 21570 20760 23520
rect 21468 22386 21496 23520
rect 21468 22358 21588 22386
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20640 21542 20760 21570
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 19996 21321 20024 21354
rect 19982 21312 20038 21321
rect 19982 21247 20038 21256
rect 20548 20466 20576 21490
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19706 17368 19762 17377
rect 19706 17303 19762 17312
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18880 16788 18932 16794
rect 18880 16730 18932 16736
rect 18892 14958 18920 16730
rect 19076 16590 19104 17070
rect 19064 16584 19116 16590
rect 19064 16526 19116 16532
rect 19116 16348 19412 16368
rect 19172 16346 19196 16348
rect 19252 16346 19276 16348
rect 19332 16346 19356 16348
rect 19194 16294 19196 16346
rect 19258 16294 19270 16346
rect 19332 16294 19334 16346
rect 19172 16292 19196 16294
rect 19252 16292 19276 16294
rect 19332 16292 19356 16294
rect 19116 16272 19412 16292
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19444 15570 19472 15914
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18984 14550 19012 15438
rect 19116 15260 19412 15280
rect 19172 15258 19196 15260
rect 19252 15258 19276 15260
rect 19332 15258 19356 15260
rect 19194 15206 19196 15258
rect 19258 15206 19270 15258
rect 19332 15206 19334 15258
rect 19172 15204 19196 15206
rect 19252 15204 19276 15206
rect 19332 15204 19356 15206
rect 19116 15184 19412 15204
rect 19444 15162 19472 15506
rect 19720 15162 19748 17138
rect 19996 15910 20024 20266
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20074 17776 20130 17785
rect 20180 17746 20208 18022
rect 20074 17711 20130 17720
rect 20168 17740 20220 17746
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19904 15609 19932 15846
rect 19890 15600 19946 15609
rect 19890 15535 19946 15544
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 19076 14618 19104 14758
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 18984 14414 19012 14486
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 18984 14074 19012 14350
rect 19116 14172 19412 14192
rect 19172 14170 19196 14172
rect 19252 14170 19276 14172
rect 19332 14170 19356 14172
rect 19194 14118 19196 14170
rect 19258 14118 19270 14170
rect 19332 14118 19334 14170
rect 19172 14116 19196 14118
rect 19252 14116 19276 14118
rect 19332 14116 19356 14118
rect 19116 14096 19412 14116
rect 19444 14074 19472 14418
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19338 13968 19394 13977
rect 19260 13926 19338 13954
rect 19260 13530 19288 13926
rect 19338 13903 19394 13912
rect 19536 13870 19564 14350
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13530 19564 13806
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19432 13388 19484 13394
rect 19432 13330 19484 13336
rect 19116 13084 19412 13104
rect 19172 13082 19196 13084
rect 19252 13082 19276 13084
rect 19332 13082 19356 13084
rect 19194 13030 19196 13082
rect 19258 13030 19270 13082
rect 19332 13030 19334 13082
rect 19172 13028 19196 13030
rect 19252 13028 19276 13030
rect 19332 13028 19356 13030
rect 19116 13008 19412 13028
rect 19444 12986 19472 13330
rect 19720 13308 19748 14214
rect 19812 13530 19840 15302
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19800 13524 19852 13530
rect 19800 13466 19852 13472
rect 19720 13280 19840 13308
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12442 19380 12582
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 19340 12436 19392 12442
rect 19340 12378 19392 12384
rect 19616 12368 19668 12374
rect 19616 12310 19668 12316
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18696 11280 18748 11286
rect 18694 11248 18696 11257
rect 18748 11248 18750 11257
rect 18800 11218 18828 12242
rect 19116 11996 19412 12016
rect 19172 11994 19196 11996
rect 19252 11994 19276 11996
rect 19332 11994 19356 11996
rect 19194 11942 19196 11994
rect 19258 11942 19270 11994
rect 19332 11942 19334 11994
rect 19172 11940 19196 11942
rect 19252 11940 19276 11942
rect 19332 11940 19356 11942
rect 19116 11920 19412 11940
rect 19628 11937 19656 12310
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19720 11286 19748 12922
rect 19812 11694 19840 13280
rect 19904 12986 19932 14758
rect 19892 12980 19944 12986
rect 19892 12922 19944 12928
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 12442 19932 12582
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19892 12300 19944 12306
rect 19892 12242 19944 12248
rect 19904 11778 19932 12242
rect 19996 11898 20024 15438
rect 20088 14006 20116 17711
rect 20168 17682 20220 17688
rect 20272 16402 20300 19926
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 18970 20392 19790
rect 20536 19236 20588 19242
rect 20536 19178 20588 19184
rect 20548 18970 20576 19178
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20640 18630 20668 21542
rect 20720 21412 20772 21418
rect 20720 21354 20772 21360
rect 20732 20806 20760 21354
rect 20812 21344 20864 21350
rect 20812 21286 20864 21292
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 20824 21010 20852 21286
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 19990 20760 20742
rect 20824 20602 20852 20946
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20720 19984 20772 19990
rect 20720 19926 20772 19932
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20824 19514 20852 19858
rect 20812 19508 20864 19514
rect 20812 19450 20864 19456
rect 20916 19174 20944 20946
rect 20996 20800 21048 20806
rect 20994 20768 20996 20777
rect 21048 20768 21050 20777
rect 20994 20703 21050 20712
rect 21192 19446 21220 21286
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 20904 19168 20956 19174
rect 20904 19110 20956 19116
rect 21088 18828 21140 18834
rect 21088 18770 21140 18776
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20996 18624 21048 18630
rect 20996 18566 21048 18572
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20180 16374 20300 16402
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19904 11750 20024 11778
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11354 19932 11630
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 18694 11183 18750 11192
rect 18788 11212 18840 11218
rect 18788 11154 18840 11160
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 9489 18736 10406
rect 18800 9994 18828 11154
rect 19432 11008 19484 11014
rect 19432 10950 19484 10956
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19116 10908 19412 10928
rect 19172 10906 19196 10908
rect 19252 10906 19276 10908
rect 19332 10906 19356 10908
rect 19194 10854 19196 10906
rect 19258 10854 19270 10906
rect 19332 10854 19334 10906
rect 19172 10852 19196 10854
rect 19252 10852 19276 10854
rect 19332 10852 19356 10854
rect 19116 10832 19412 10852
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18878 10296 18934 10305
rect 18878 10231 18880 10240
rect 18932 10231 18934 10240
rect 18880 10202 18932 10208
rect 18984 10130 19012 10610
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19338 10432 19394 10441
rect 19076 10266 19104 10406
rect 19338 10367 19394 10376
rect 19154 10296 19210 10305
rect 19064 10260 19116 10266
rect 19154 10231 19156 10240
rect 19064 10202 19116 10208
rect 19208 10231 19210 10240
rect 19156 10202 19208 10208
rect 19352 10198 19380 10367
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 18972 10124 19024 10130
rect 18972 10066 19024 10072
rect 18788 9988 18840 9994
rect 18788 9930 18840 9936
rect 18984 9654 19012 10066
rect 19116 9820 19412 9840
rect 19172 9818 19196 9820
rect 19252 9818 19276 9820
rect 19332 9818 19356 9820
rect 19194 9766 19196 9818
rect 19258 9766 19270 9818
rect 19332 9766 19334 9818
rect 19172 9764 19196 9766
rect 19252 9764 19276 9766
rect 19332 9764 19356 9766
rect 19116 9744 19412 9764
rect 19444 9738 19472 10950
rect 19522 10024 19578 10033
rect 19522 9959 19578 9968
rect 19536 9926 19564 9959
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19522 9752 19578 9761
rect 19444 9710 19522 9738
rect 19628 9722 19656 10950
rect 19720 9994 19748 10950
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19522 9687 19578 9696
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 18972 9648 19024 9654
rect 18786 9616 18842 9625
rect 18972 9590 19024 9596
rect 18786 9551 18842 9560
rect 19338 9582 19394 9591
rect 18432 9438 18644 9466
rect 18694 9480 18750 9489
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18144 8968 18196 8974
rect 18064 8928 18144 8956
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17972 8362 18000 8434
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 18064 7449 18092 8928
rect 18144 8910 18196 8916
rect 18326 8800 18382 8809
rect 18432 8786 18460 9438
rect 18694 9415 18750 9424
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18382 8758 18460 8786
rect 18326 8735 18382 8744
rect 18050 7440 18106 7449
rect 18050 7375 18106 7384
rect 18064 7274 18092 7375
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 17684 6860 17736 6866
rect 17604 6820 17684 6848
rect 17314 6352 17370 6361
rect 17314 6287 17370 6296
rect 17130 6216 17186 6225
rect 17130 6151 17186 6160
rect 17408 5568 17460 5574
rect 17408 5510 17460 5516
rect 17420 5370 17448 5510
rect 17604 5409 17632 6820
rect 17684 6802 17736 6808
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5778 17724 6054
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17590 5400 17646 5409
rect 17408 5364 17460 5370
rect 17590 5335 17646 5344
rect 17408 5306 17460 5312
rect 16396 5092 16448 5098
rect 16396 5034 16448 5040
rect 16868 5086 17080 5114
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16316 3233 16344 3878
rect 16396 3460 16448 3466
rect 16396 3402 16448 3408
rect 16302 3224 16358 3233
rect 16302 3159 16358 3168
rect 16316 2990 16344 3159
rect 16120 2984 16172 2990
rect 16040 2944 16120 2972
rect 16120 2926 16172 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16132 2836 16160 2926
rect 16408 2836 16436 3402
rect 16500 2972 16528 4966
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16592 4078 16620 4626
rect 16684 4282 16712 4966
rect 16868 4570 16896 5086
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 17040 5024 17092 5030
rect 17040 4966 17092 4972
rect 16960 4758 16988 4966
rect 16948 4752 17000 4758
rect 16948 4694 17000 4700
rect 16868 4542 16988 4570
rect 16672 4276 16724 4282
rect 16672 4218 16724 4224
rect 16580 4072 16632 4078
rect 16580 4014 16632 4020
rect 16672 4072 16724 4078
rect 16672 4014 16724 4020
rect 16684 3194 16712 4014
rect 16856 4004 16908 4010
rect 16856 3946 16908 3952
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16580 2984 16632 2990
rect 16500 2944 16580 2972
rect 16580 2926 16632 2932
rect 16132 2808 16436 2836
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15936 2576 15988 2582
rect 15936 2518 15988 2524
rect 16132 2514 16160 2808
rect 16868 2650 16896 3946
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 15108 2372 15160 2378
rect 15108 2314 15160 2320
rect 16960 2310 16988 4542
rect 17052 2582 17080 4966
rect 17420 4622 17448 5306
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17604 4690 17632 5170
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17328 2990 17356 4422
rect 17604 4214 17632 4626
rect 17880 4486 17908 5714
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 4758 18092 5510
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18052 3936 18104 3942
rect 18052 3878 18104 3884
rect 18064 3670 18092 3878
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 18052 3664 18104 3670
rect 18052 3606 18104 3612
rect 17420 3194 17448 3606
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 18156 2650 18184 4082
rect 18248 3194 18276 4626
rect 18340 3942 18368 8735
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18432 7993 18460 8026
rect 18418 7984 18474 7993
rect 18418 7919 18474 7928
rect 18524 7886 18552 9114
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 6254 18460 7686
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18432 3602 18460 5510
rect 18616 4729 18644 9318
rect 18708 9042 18736 9415
rect 18800 9382 18828 9551
rect 18972 9512 19024 9518
rect 19156 9512 19208 9518
rect 19338 9517 19394 9526
rect 19616 9580 19668 9586
rect 19720 9568 19748 9930
rect 19668 9540 19748 9568
rect 19616 9522 19668 9528
rect 18972 9454 19024 9460
rect 19154 9480 19156 9489
rect 19432 9512 19484 9518
rect 19208 9480 19210 9489
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18708 8820 18736 8978
rect 18788 8968 18840 8974
rect 18984 8956 19012 9454
rect 19484 9472 19564 9500
rect 19432 9454 19484 9460
rect 19154 9415 19210 9424
rect 19536 9382 19564 9472
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19444 9194 19472 9318
rect 19812 9194 19840 11154
rect 19996 10130 20024 11750
rect 20088 10169 20116 12242
rect 20180 10606 20208 16374
rect 20258 16280 20314 16289
rect 20258 16215 20314 16224
rect 20272 16046 20300 16215
rect 20260 16040 20312 16046
rect 20260 15982 20312 15988
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 14634 20300 15846
rect 20364 15026 20392 17478
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20456 16658 20484 17070
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20456 16250 20484 16594
rect 20444 16244 20496 16250
rect 20444 16186 20496 16192
rect 20352 15020 20404 15026
rect 20352 14962 20404 14968
rect 20272 14606 20484 14634
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20272 14074 20300 14418
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20364 13954 20392 14486
rect 20272 13926 20392 13954
rect 20168 10600 20220 10606
rect 20168 10542 20220 10548
rect 20074 10160 20130 10169
rect 19984 10124 20036 10130
rect 20074 10095 20130 10104
rect 19984 10066 20036 10072
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19444 9166 19840 9194
rect 18840 8928 19012 8956
rect 18788 8910 18840 8916
rect 19432 8832 19484 8838
rect 18708 8792 18828 8820
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 18708 6866 18736 8230
rect 18800 7342 18828 8792
rect 19432 8774 19484 8780
rect 19116 8732 19412 8752
rect 19172 8730 19196 8732
rect 19252 8730 19276 8732
rect 19332 8730 19356 8732
rect 19194 8678 19196 8730
rect 19258 8678 19270 8730
rect 19332 8678 19334 8730
rect 19172 8676 19196 8678
rect 19252 8676 19276 8678
rect 19332 8676 19356 8678
rect 19116 8656 19412 8676
rect 19444 8090 19472 8774
rect 19628 8430 19656 9166
rect 19708 9036 19760 9042
rect 19708 8978 19760 8984
rect 19720 8634 19748 8978
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19616 8424 19668 8430
rect 19616 8366 19668 8372
rect 19524 8356 19576 8362
rect 19524 8298 19576 8304
rect 19432 8084 19484 8090
rect 19432 8026 19484 8032
rect 19536 7857 19564 8298
rect 19904 8276 19932 9862
rect 20180 9722 20208 9998
rect 20168 9716 20220 9722
rect 20168 9658 20220 9664
rect 20272 9602 20300 13926
rect 20456 13818 20484 14606
rect 20548 14550 20576 17478
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20456 13790 20576 13818
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 19706 8256 19762 8265
rect 19706 8191 19762 8200
rect 19812 8248 19932 8276
rect 19996 9574 20300 9602
rect 19616 7948 19668 7954
rect 19616 7890 19668 7896
rect 19522 7848 19578 7857
rect 19522 7783 19578 7792
rect 19628 7732 19656 7890
rect 19536 7704 19656 7732
rect 19116 7644 19412 7664
rect 19172 7642 19196 7644
rect 19252 7642 19276 7644
rect 19332 7642 19356 7644
rect 19194 7590 19196 7642
rect 19258 7590 19270 7642
rect 19332 7590 19334 7642
rect 19172 7588 19196 7590
rect 19252 7588 19276 7590
rect 19332 7588 19356 7590
rect 19116 7568 19412 7588
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 18788 7336 18840 7342
rect 18788 7278 18840 7284
rect 18800 7002 18828 7278
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18696 6860 18748 6866
rect 18696 6802 18748 6808
rect 18708 6089 18736 6802
rect 18694 6080 18750 6089
rect 18694 6015 18750 6024
rect 18708 5030 18736 6015
rect 18696 5024 18748 5030
rect 18696 4966 18748 4972
rect 18602 4720 18658 4729
rect 18602 4655 18658 4664
rect 18708 4570 18736 4966
rect 18616 4542 18736 4570
rect 18616 3602 18644 4542
rect 18800 3738 18828 6938
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18892 4826 18920 5646
rect 18984 4826 19012 7142
rect 19444 6662 19472 7346
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 19116 6556 19412 6576
rect 19172 6554 19196 6556
rect 19252 6554 19276 6556
rect 19332 6554 19356 6556
rect 19194 6502 19196 6554
rect 19258 6502 19270 6554
rect 19332 6502 19334 6554
rect 19172 6500 19196 6502
rect 19252 6500 19276 6502
rect 19332 6500 19356 6502
rect 19116 6480 19412 6500
rect 19536 6440 19564 7704
rect 19616 7540 19668 7546
rect 19616 7482 19668 7488
rect 19352 6412 19564 6440
rect 19352 5642 19380 6412
rect 19432 6180 19484 6186
rect 19432 6122 19484 6128
rect 19444 5710 19472 6122
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19340 5636 19392 5642
rect 19340 5578 19392 5584
rect 19116 5468 19412 5488
rect 19172 5466 19196 5468
rect 19252 5466 19276 5468
rect 19332 5466 19356 5468
rect 19194 5414 19196 5466
rect 19258 5414 19270 5466
rect 19332 5414 19334 5466
rect 19172 5412 19196 5414
rect 19252 5412 19276 5414
rect 19332 5412 19356 5414
rect 19116 5392 19412 5412
rect 19444 5370 19472 5646
rect 19432 5364 19484 5370
rect 19432 5306 19484 5312
rect 19536 5166 19564 5714
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18972 4820 19024 4826
rect 18972 4762 19024 4768
rect 19260 4758 19288 5034
rect 19628 4826 19656 7482
rect 19720 6254 19748 8191
rect 19812 7206 19840 8248
rect 19996 8090 20024 9574
rect 20260 9512 20312 9518
rect 20166 9480 20222 9489
rect 20364 9466 20392 12582
rect 20456 12442 20484 13262
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20456 11694 20484 12378
rect 20548 12102 20576 13790
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20444 11688 20496 11694
rect 20444 11630 20496 11636
rect 20548 10554 20576 12038
rect 20312 9460 20392 9466
rect 20260 9454 20392 9460
rect 20272 9438 20392 9454
rect 20166 9415 20222 9424
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 8498 20116 9318
rect 20180 9110 20208 9415
rect 20364 9178 20392 9438
rect 20456 10526 20576 10554
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20168 9104 20220 9110
rect 20456 9058 20484 10526
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20548 9450 20576 10406
rect 20536 9444 20588 9450
rect 20536 9386 20588 9392
rect 20168 9046 20220 9052
rect 20272 9030 20484 9058
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 20272 8378 20300 9030
rect 20548 8974 20576 9386
rect 20536 8968 20588 8974
rect 20536 8910 20588 8916
rect 20640 8514 20668 18158
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20812 18080 20864 18086
rect 20812 18022 20864 18028
rect 20732 15706 20760 18022
rect 20824 17338 20852 18022
rect 20916 17746 20944 18566
rect 20904 17740 20956 17746
rect 20904 17682 20956 17688
rect 21008 17626 21036 18566
rect 20916 17598 21036 17626
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20720 15428 20772 15434
rect 20720 15370 20772 15376
rect 20732 15162 20760 15370
rect 20824 15366 20852 17138
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20720 14952 20772 14958
rect 20720 14894 20772 14900
rect 20732 14482 20760 14894
rect 20812 14612 20864 14618
rect 20812 14554 20864 14560
rect 20720 14476 20772 14482
rect 20720 14418 20772 14424
rect 20732 14074 20760 14418
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20732 13394 20760 14010
rect 20824 13802 20852 14554
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20916 13546 20944 17598
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 21008 16658 21036 16934
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 21008 16250 21036 16594
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20996 15496 21048 15502
rect 20996 15438 21048 15444
rect 21008 13682 21036 15438
rect 21100 15162 21128 18770
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21192 17610 21220 18226
rect 21180 17604 21232 17610
rect 21180 17546 21232 17552
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 16658 21220 16934
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21192 15706 21220 16594
rect 21180 15700 21232 15706
rect 21180 15642 21232 15648
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21192 15366 21220 15438
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 21100 14550 21128 15098
rect 21088 14544 21140 14550
rect 21088 14486 21140 14492
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21008 13654 21128 13682
rect 20916 13518 21036 13546
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20720 12844 20772 12850
rect 20720 12786 20772 12792
rect 20732 11898 20760 12786
rect 20824 12714 20852 13126
rect 20916 12850 20944 13330
rect 20904 12844 20956 12850
rect 20904 12786 20956 12792
rect 20812 12708 20864 12714
rect 20812 12650 20864 12656
rect 20916 12306 20944 12786
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20732 11286 20760 11834
rect 20824 11354 20852 12174
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20720 11280 20772 11286
rect 20720 11222 20772 11228
rect 20824 10538 20852 11290
rect 20904 11212 20956 11218
rect 20904 11154 20956 11160
rect 20916 10674 20944 11154
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20812 10532 20864 10538
rect 20812 10474 20864 10480
rect 20916 10130 20944 10610
rect 20904 10124 20956 10130
rect 20904 10066 20956 10072
rect 20916 9042 20944 10066
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20088 8350 20300 8378
rect 20364 8486 20668 8514
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 20088 7970 20116 8350
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 19904 7942 20116 7970
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19800 6928 19852 6934
rect 19800 6870 19852 6876
rect 19812 6458 19840 6870
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19798 6352 19854 6361
rect 19798 6287 19854 6296
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19812 5250 19840 6287
rect 19904 5409 19932 7942
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19996 5914 20024 7686
rect 20088 7478 20116 7822
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 20076 7200 20128 7206
rect 20076 7142 20128 7148
rect 20088 6662 20116 7142
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20076 6248 20128 6254
rect 20076 6190 20128 6196
rect 19984 5908 20036 5914
rect 19984 5850 20036 5856
rect 19890 5400 19946 5409
rect 20088 5370 20116 6190
rect 20180 5642 20208 8026
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20272 7342 20300 7958
rect 20364 7546 20392 8486
rect 20628 8424 20680 8430
rect 20628 8366 20680 8372
rect 20444 7880 20496 7886
rect 20444 7822 20496 7828
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20352 7540 20404 7546
rect 20352 7482 20404 7488
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 20272 6458 20300 7278
rect 20364 6746 20392 7482
rect 20456 7410 20484 7822
rect 20444 7404 20496 7410
rect 20444 7346 20496 7352
rect 20548 6934 20576 7822
rect 20536 6928 20588 6934
rect 20640 6905 20668 8366
rect 20536 6870 20588 6876
rect 20626 6896 20682 6905
rect 20626 6831 20682 6840
rect 20720 6792 20772 6798
rect 20364 6718 20668 6746
rect 20720 6734 20772 6740
rect 20352 6656 20404 6662
rect 20352 6598 20404 6604
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20168 5636 20220 5642
rect 20168 5578 20220 5584
rect 19890 5335 19946 5344
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 19812 5222 19932 5250
rect 19616 4820 19668 4826
rect 19616 4762 19668 4768
rect 19248 4752 19300 4758
rect 19248 4694 19300 4700
rect 19708 4480 19760 4486
rect 19708 4422 19760 4428
rect 19116 4380 19412 4400
rect 19172 4378 19196 4380
rect 19252 4378 19276 4380
rect 19332 4378 19356 4380
rect 19194 4326 19196 4378
rect 19258 4326 19270 4378
rect 19332 4326 19334 4378
rect 19172 4324 19196 4326
rect 19252 4324 19276 4326
rect 19332 4324 19356 4326
rect 19116 4304 19412 4324
rect 19720 4146 19748 4422
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19800 4004 19852 4010
rect 19800 3946 19852 3952
rect 18880 3936 18932 3942
rect 18880 3878 18932 3884
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18616 3466 18644 3538
rect 18604 3460 18656 3466
rect 18604 3402 18656 3408
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 2922 18368 3334
rect 18616 3194 18644 3402
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18616 2990 18644 3130
rect 18604 2984 18656 2990
rect 18432 2944 18604 2972
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18340 2582 18368 2858
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18328 2440 18380 2446
rect 18432 2428 18460 2944
rect 18604 2926 18656 2932
rect 18708 2854 18736 3538
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18708 2650 18736 2790
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18892 2553 18920 3878
rect 19116 3292 19412 3312
rect 19172 3290 19196 3292
rect 19252 3290 19276 3292
rect 19332 3290 19356 3292
rect 19194 3238 19196 3290
rect 19258 3238 19270 3290
rect 19332 3238 19334 3290
rect 19172 3236 19196 3238
rect 19252 3236 19276 3238
rect 19332 3236 19356 3238
rect 19116 3216 19412 3236
rect 19812 3194 19840 3946
rect 19904 3913 19932 5222
rect 20088 4826 20116 5306
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20168 5024 20220 5030
rect 20168 4966 20220 4972
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19984 3936 20036 3942
rect 19890 3904 19946 3913
rect 19984 3878 20036 3884
rect 19890 3839 19946 3848
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19248 2848 19300 2854
rect 19904 2836 19932 3674
rect 19996 3398 20024 3878
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19996 2990 20024 3334
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19904 2808 20024 2836
rect 19248 2790 19300 2796
rect 19260 2582 19288 2790
rect 19248 2576 19300 2582
rect 18878 2544 18934 2553
rect 19248 2518 19300 2524
rect 18878 2479 18934 2488
rect 18380 2400 18460 2428
rect 18328 2382 18380 2388
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17788 2106 17816 2382
rect 19116 2204 19412 2224
rect 19172 2202 19196 2204
rect 19252 2202 19276 2204
rect 19332 2202 19356 2204
rect 19194 2150 19196 2202
rect 19258 2150 19270 2202
rect 19332 2150 19334 2202
rect 19172 2148 19196 2150
rect 19252 2148 19276 2150
rect 19332 2148 19356 2150
rect 19116 2128 19412 2148
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 17776 2100 17828 2106
rect 17776 2042 17828 2048
rect 11992 1414 12204 1442
rect 11992 480 12020 1414
rect 19996 480 20024 2808
rect 20088 2378 20116 4014
rect 20180 3738 20208 4966
rect 20272 4282 20300 5034
rect 20260 4276 20312 4282
rect 20260 4218 20312 4224
rect 20168 3732 20220 3738
rect 20168 3674 20220 3680
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20180 3126 20208 3470
rect 20364 3233 20392 6598
rect 20548 5710 20576 6598
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20456 4078 20484 4558
rect 20444 4072 20496 4078
rect 20444 4014 20496 4020
rect 20456 3534 20484 4014
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20350 3224 20406 3233
rect 20350 3159 20406 3168
rect 20168 3120 20220 3126
rect 20168 3062 20220 3068
rect 20076 2372 20128 2378
rect 20076 2314 20128 2320
rect 20548 1057 20576 5510
rect 20534 1048 20590 1057
rect 20534 983 20590 992
rect 3974 0 4030 480
rect 11978 0 12034 480
rect 19982 0 20038 480
rect 20640 377 20668 6718
rect 20732 6254 20760 6734
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20720 5092 20772 5098
rect 20720 5034 20772 5040
rect 20732 4486 20760 5034
rect 20824 4554 20852 8502
rect 20916 8498 20944 8978
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21008 7449 21036 13518
rect 21100 12986 21128 13654
rect 21192 13190 21220 13806
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21100 12374 21128 12922
rect 21192 12782 21220 13126
rect 21180 12776 21232 12782
rect 21180 12718 21232 12724
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21192 8634 21220 9318
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21284 8401 21312 20810
rect 21376 19310 21404 20878
rect 21560 20505 21588 22358
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21744 21554 21772 21830
rect 21732 21548 21784 21554
rect 21732 21490 21784 21496
rect 21732 21412 21784 21418
rect 21732 21354 21784 21360
rect 21546 20496 21602 20505
rect 21456 20460 21508 20466
rect 21546 20431 21602 20440
rect 21456 20402 21508 20408
rect 21468 19378 21496 20402
rect 21548 20256 21600 20262
rect 21548 20198 21600 20204
rect 21640 20256 21692 20262
rect 21640 20198 21692 20204
rect 21560 20058 21588 20198
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21652 19514 21680 20198
rect 21640 19508 21692 19514
rect 21640 19450 21692 19456
rect 21744 19394 21772 21354
rect 22112 20890 22140 23520
rect 22112 20862 22324 20890
rect 22100 20800 22152 20806
rect 22100 20742 22152 20748
rect 22112 19961 22140 20742
rect 22098 19952 22154 19961
rect 22098 19887 22154 19896
rect 21456 19372 21508 19378
rect 21456 19314 21508 19320
rect 21652 19366 21772 19394
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21376 18902 21404 19110
rect 21364 18896 21416 18902
rect 21364 18838 21416 18844
rect 21376 18426 21404 18838
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21364 18420 21416 18426
rect 21364 18362 21416 18368
rect 21456 18148 21508 18154
rect 21456 18090 21508 18096
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21376 17882 21404 18022
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21376 15978 21404 17546
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21364 15564 21416 15570
rect 21364 15506 21416 15512
rect 21376 11830 21404 15506
rect 21468 14618 21496 18090
rect 21560 15910 21588 18634
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21560 14958 21588 15846
rect 21548 14952 21600 14958
rect 21548 14894 21600 14900
rect 21456 14612 21508 14618
rect 21456 14554 21508 14560
rect 21652 13308 21680 19366
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 22098 19136 22154 19145
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 21836 18290 21864 18702
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21732 18080 21784 18086
rect 21732 18022 21784 18028
rect 21744 14074 21772 18022
rect 21836 17202 21864 18226
rect 21928 17762 21956 19110
rect 22098 19071 22154 19080
rect 22112 17882 22140 19071
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21928 17734 22140 17762
rect 21824 17196 21876 17202
rect 21824 17138 21876 17144
rect 21824 16992 21876 16998
rect 21824 16934 21876 16940
rect 21914 16960 21970 16969
rect 21836 16794 21864 16934
rect 21914 16895 21970 16904
rect 21824 16788 21876 16794
rect 21824 16730 21876 16736
rect 21928 15570 21956 16895
rect 21916 15564 21968 15570
rect 21916 15506 21968 15512
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21744 13462 21772 14010
rect 21732 13456 21784 13462
rect 21732 13398 21784 13404
rect 21652 13280 21772 13308
rect 21640 12708 21692 12714
rect 21640 12650 21692 12656
rect 21364 11824 21416 11830
rect 21364 11766 21416 11772
rect 21652 9586 21680 12650
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21744 9081 21772 13280
rect 21730 9072 21786 9081
rect 21730 9007 21786 9016
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 21270 8392 21326 8401
rect 21270 8327 21326 8336
rect 21916 7948 21968 7954
rect 21916 7890 21968 7896
rect 21548 7880 21600 7886
rect 21548 7822 21600 7828
rect 20994 7440 21050 7449
rect 20994 7375 21050 7384
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 6458 20944 7142
rect 21560 6882 21588 7822
rect 21640 7744 21692 7750
rect 21640 7686 21692 7692
rect 21652 7342 21680 7686
rect 21928 7585 21956 7890
rect 21914 7576 21970 7585
rect 21914 7511 21970 7520
rect 21732 7404 21784 7410
rect 21732 7346 21784 7352
rect 21640 7336 21692 7342
rect 21640 7278 21692 7284
rect 21560 6854 21680 6882
rect 21652 6662 21680 6854
rect 21640 6656 21692 6662
rect 21640 6598 21692 6604
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 21652 6254 21680 6598
rect 21640 6248 21692 6254
rect 21640 6190 21692 6196
rect 21744 6118 21772 7346
rect 21732 6112 21784 6118
rect 21732 6054 21784 6060
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20916 5166 20944 5646
rect 20904 5160 20956 5166
rect 20904 5102 20956 5108
rect 20916 4622 20944 5102
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20812 4548 20864 4554
rect 20812 4490 20864 4496
rect 20720 4480 20772 4486
rect 20720 4422 20772 4428
rect 20824 4434 20852 4490
rect 20732 2650 20760 4422
rect 20824 4406 20944 4434
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20720 2440 20772 2446
rect 20916 2428 20944 4406
rect 21284 3942 21312 4694
rect 21272 3936 21324 3942
rect 21272 3878 21324 3884
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 21192 2854 21220 3538
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21284 2514 21312 3878
rect 22020 2990 22048 9007
rect 22112 8537 22140 17734
rect 22296 16726 22324 20862
rect 22848 20369 22876 23520
rect 22834 20360 22890 20369
rect 22834 20295 22890 20304
rect 23584 17814 23612 23520
rect 23572 17808 23624 17814
rect 23572 17750 23624 17756
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22284 16448 22336 16454
rect 22284 16390 22336 16396
rect 22296 16046 22324 16390
rect 22284 16040 22336 16046
rect 22284 15982 22336 15988
rect 22296 15638 22324 15982
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 23386 11248 23442 11257
rect 23386 11183 23442 11192
rect 23400 11121 23428 11183
rect 23386 11112 23442 11121
rect 23386 11047 23442 11056
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22296 10198 22324 10406
rect 22284 10192 22336 10198
rect 22284 10134 22336 10140
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 22204 8906 22232 9522
rect 22296 9110 22324 9862
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22192 8900 22244 8906
rect 22192 8842 22244 8848
rect 22098 8528 22154 8537
rect 22098 8463 22154 8472
rect 22204 8430 22232 8842
rect 22284 8560 22336 8566
rect 22284 8502 22336 8508
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22296 8362 22324 8502
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 22296 6089 22324 8298
rect 22376 7744 22428 7750
rect 22376 7686 22428 7692
rect 22282 6080 22338 6089
rect 22282 6015 22338 6024
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22112 5030 22140 5714
rect 22284 5568 22336 5574
rect 22284 5510 22336 5516
rect 22100 5024 22152 5030
rect 22100 4966 22152 4972
rect 22112 2990 22140 4966
rect 22296 4826 22324 5510
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 22388 4282 22416 7686
rect 22376 4276 22428 4282
rect 22376 4218 22428 4224
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22296 3738 22324 3946
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22008 2984 22060 2990
rect 22008 2926 22060 2932
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22388 2802 22416 4218
rect 22112 2774 22416 2802
rect 21272 2508 21324 2514
rect 21272 2450 21324 2456
rect 22112 2446 22140 2774
rect 20772 2400 20944 2428
rect 22100 2440 22152 2446
rect 20720 2382 20772 2388
rect 22100 2382 22152 2388
rect 20732 2106 20760 2382
rect 20720 2100 20772 2106
rect 20720 2042 20772 2048
rect 20626 368 20682 377
rect 20626 303 20682 312
<< via2 >>
rect 1398 21428 1400 21448
rect 1400 21428 1452 21448
rect 1452 21428 1454 21448
rect 1398 21392 1454 21428
rect 1582 18672 1638 18728
rect 2778 19896 2834 19952
rect 1766 18128 1822 18184
rect 1674 13776 1730 13832
rect 1490 11872 1546 11928
rect 1858 9988 1914 10024
rect 1858 9968 1860 9988
rect 1860 9968 1912 9988
rect 1912 9968 1914 9988
rect 4066 19760 4122 19816
rect 3974 17856 4030 17912
rect 2778 14456 2834 14512
rect 3054 12300 3110 12336
rect 3054 12280 3056 12300
rect 3056 12280 3108 12300
rect 3108 12280 3110 12300
rect 3238 13812 3240 13832
rect 3240 13812 3292 13832
rect 3292 13812 3294 13832
rect 3238 13776 3294 13812
rect 2686 9580 2742 9616
rect 2686 9560 2688 9580
rect 2688 9560 2740 9580
rect 2740 9560 2742 9580
rect 1582 9460 1584 9480
rect 1584 9460 1636 9480
rect 1636 9460 1638 9480
rect 1582 9424 1638 9460
rect 3698 14048 3754 14104
rect 3606 12144 3662 12200
rect 2502 9172 2558 9208
rect 2502 9152 2504 9172
rect 2504 9152 2556 9172
rect 2556 9152 2558 9172
rect 4588 21786 4644 21788
rect 4668 21786 4724 21788
rect 4748 21786 4804 21788
rect 4828 21786 4884 21788
rect 4588 21734 4614 21786
rect 4614 21734 4644 21786
rect 4668 21734 4678 21786
rect 4678 21734 4724 21786
rect 4748 21734 4794 21786
rect 4794 21734 4804 21786
rect 4828 21734 4858 21786
rect 4858 21734 4884 21786
rect 4588 21732 4644 21734
rect 4668 21732 4724 21734
rect 4748 21732 4804 21734
rect 4828 21732 4884 21734
rect 4588 20698 4644 20700
rect 4668 20698 4724 20700
rect 4748 20698 4804 20700
rect 4828 20698 4884 20700
rect 4588 20646 4614 20698
rect 4614 20646 4644 20698
rect 4668 20646 4678 20698
rect 4678 20646 4724 20698
rect 4748 20646 4794 20698
rect 4794 20646 4804 20698
rect 4828 20646 4858 20698
rect 4858 20646 4884 20698
rect 4588 20644 4644 20646
rect 4668 20644 4724 20646
rect 4748 20644 4804 20646
rect 4828 20644 4884 20646
rect 4618 19796 4620 19816
rect 4620 19796 4672 19816
rect 4672 19796 4674 19816
rect 4618 19760 4674 19796
rect 4588 19610 4644 19612
rect 4668 19610 4724 19612
rect 4748 19610 4804 19612
rect 4828 19610 4884 19612
rect 4588 19558 4614 19610
rect 4614 19558 4644 19610
rect 4668 19558 4678 19610
rect 4678 19558 4724 19610
rect 4748 19558 4794 19610
rect 4794 19558 4804 19610
rect 4828 19558 4858 19610
rect 4858 19558 4884 19610
rect 4588 19556 4644 19558
rect 4668 19556 4724 19558
rect 4748 19556 4804 19558
rect 4828 19556 4884 19558
rect 4986 19508 5042 19544
rect 4986 19488 4988 19508
rect 4988 19488 5040 19508
rect 5040 19488 5042 19508
rect 5538 20576 5594 20632
rect 4526 19252 4528 19272
rect 4528 19252 4580 19272
rect 4580 19252 4582 19272
rect 4526 19216 4582 19252
rect 5354 19080 5410 19136
rect 4588 18522 4644 18524
rect 4668 18522 4724 18524
rect 4748 18522 4804 18524
rect 4828 18522 4884 18524
rect 4588 18470 4614 18522
rect 4614 18470 4644 18522
rect 4668 18470 4678 18522
rect 4678 18470 4724 18522
rect 4748 18470 4794 18522
rect 4794 18470 4804 18522
rect 4828 18470 4858 18522
rect 4858 18470 4884 18522
rect 4588 18468 4644 18470
rect 4668 18468 4724 18470
rect 4748 18468 4804 18470
rect 4828 18468 4884 18470
rect 4588 17434 4644 17436
rect 4668 17434 4724 17436
rect 4748 17434 4804 17436
rect 4828 17434 4884 17436
rect 4588 17382 4614 17434
rect 4614 17382 4644 17434
rect 4668 17382 4678 17434
rect 4678 17382 4724 17434
rect 4748 17382 4794 17434
rect 4794 17382 4804 17434
rect 4828 17382 4858 17434
rect 4858 17382 4884 17434
rect 4588 17380 4644 17382
rect 4668 17380 4724 17382
rect 4748 17380 4804 17382
rect 4828 17380 4884 17382
rect 4618 17176 4674 17232
rect 4588 16346 4644 16348
rect 4668 16346 4724 16348
rect 4748 16346 4804 16348
rect 4828 16346 4884 16348
rect 4588 16294 4614 16346
rect 4614 16294 4644 16346
rect 4668 16294 4678 16346
rect 4678 16294 4724 16346
rect 4748 16294 4794 16346
rect 4794 16294 4804 16346
rect 4828 16294 4858 16346
rect 4858 16294 4884 16346
rect 4588 16292 4644 16294
rect 4668 16292 4724 16294
rect 4748 16292 4804 16294
rect 4828 16292 4884 16294
rect 4588 15258 4644 15260
rect 4668 15258 4724 15260
rect 4748 15258 4804 15260
rect 4828 15258 4884 15260
rect 4588 15206 4614 15258
rect 4614 15206 4644 15258
rect 4668 15206 4678 15258
rect 4678 15206 4724 15258
rect 4748 15206 4794 15258
rect 4794 15206 4804 15258
rect 4828 15206 4858 15258
rect 4858 15206 4884 15258
rect 4588 15204 4644 15206
rect 4668 15204 4724 15206
rect 4748 15204 4804 15206
rect 4828 15204 4884 15206
rect 4066 14456 4122 14512
rect 4158 14068 4214 14104
rect 4158 14048 4160 14068
rect 4160 14048 4212 14068
rect 4212 14048 4214 14068
rect 4588 14170 4644 14172
rect 4668 14170 4724 14172
rect 4748 14170 4804 14172
rect 4828 14170 4884 14172
rect 4588 14118 4614 14170
rect 4614 14118 4644 14170
rect 4668 14118 4678 14170
rect 4678 14118 4724 14170
rect 4748 14118 4794 14170
rect 4794 14118 4804 14170
rect 4828 14118 4858 14170
rect 4858 14118 4884 14170
rect 4588 14116 4644 14118
rect 4668 14116 4724 14118
rect 4748 14116 4804 14118
rect 4828 14116 4884 14118
rect 4526 13524 4582 13560
rect 4526 13504 4528 13524
rect 4528 13504 4580 13524
rect 4580 13504 4582 13524
rect 4588 13082 4644 13084
rect 4668 13082 4724 13084
rect 4748 13082 4804 13084
rect 4828 13082 4884 13084
rect 4588 13030 4614 13082
rect 4614 13030 4644 13082
rect 4668 13030 4678 13082
rect 4678 13030 4724 13082
rect 4748 13030 4794 13082
rect 4794 13030 4804 13082
rect 4828 13030 4858 13082
rect 4858 13030 4884 13082
rect 4588 13028 4644 13030
rect 4668 13028 4724 13030
rect 4748 13028 4804 13030
rect 4828 13028 4884 13030
rect 4066 11756 4122 11792
rect 4066 11736 4068 11756
rect 4068 11736 4120 11756
rect 4120 11736 4122 11756
rect 4588 11994 4644 11996
rect 4668 11994 4724 11996
rect 4748 11994 4804 11996
rect 4828 11994 4884 11996
rect 4588 11942 4614 11994
rect 4614 11942 4644 11994
rect 4668 11942 4678 11994
rect 4678 11942 4724 11994
rect 4748 11942 4794 11994
rect 4794 11942 4804 11994
rect 4828 11942 4858 11994
rect 4858 11942 4884 11994
rect 4588 11940 4644 11942
rect 4668 11940 4724 11942
rect 4748 11940 4804 11942
rect 4828 11940 4884 11942
rect 3882 10104 3938 10160
rect 4342 11212 4398 11248
rect 4342 11192 4344 11212
rect 4344 11192 4396 11212
rect 4396 11192 4398 11212
rect 4802 11620 4858 11656
rect 4802 11600 4804 11620
rect 4804 11600 4856 11620
rect 4856 11600 4858 11620
rect 4894 11328 4950 11384
rect 4342 11056 4398 11112
rect 4588 10906 4644 10908
rect 4668 10906 4724 10908
rect 4748 10906 4804 10908
rect 4828 10906 4884 10908
rect 4588 10854 4614 10906
rect 4614 10854 4644 10906
rect 4668 10854 4678 10906
rect 4678 10854 4724 10906
rect 4748 10854 4794 10906
rect 4794 10854 4804 10906
rect 4828 10854 4858 10906
rect 4858 10854 4884 10906
rect 4588 10852 4644 10854
rect 4668 10852 4724 10854
rect 4748 10852 4804 10854
rect 4828 10852 4884 10854
rect 4526 10648 4582 10704
rect 4894 10240 4950 10296
rect 5078 11056 5134 11112
rect 3974 9288 4030 9344
rect 3698 9036 3754 9072
rect 3698 9016 3700 9036
rect 3700 9016 3752 9036
rect 3752 9016 3754 9036
rect 4066 8880 4122 8936
rect 4250 7268 4306 7304
rect 4250 7248 4252 7268
rect 4252 7248 4304 7268
rect 4304 7248 4306 7268
rect 4588 9818 4644 9820
rect 4668 9818 4724 9820
rect 4748 9818 4804 9820
rect 4828 9818 4884 9820
rect 4588 9766 4614 9818
rect 4614 9766 4644 9818
rect 4668 9766 4678 9818
rect 4678 9766 4724 9818
rect 4748 9766 4794 9818
rect 4794 9766 4804 9818
rect 4828 9766 4858 9818
rect 4858 9766 4884 9818
rect 4588 9764 4644 9766
rect 4668 9764 4724 9766
rect 4748 9764 4804 9766
rect 4828 9764 4884 9766
rect 5170 10376 5226 10432
rect 5170 9424 5226 9480
rect 5538 17856 5594 17912
rect 5446 10512 5502 10568
rect 5354 9696 5410 9752
rect 6642 20576 6698 20632
rect 6642 19896 6698 19952
rect 6734 19352 6790 19408
rect 7102 19796 7104 19816
rect 7104 19796 7156 19816
rect 7156 19796 7158 19816
rect 7102 19760 7158 19796
rect 6734 19216 6790 19272
rect 6642 18672 6698 18728
rect 6458 17584 6514 17640
rect 6550 17176 6606 17232
rect 6458 17040 6514 17096
rect 6182 12280 6238 12336
rect 5630 11464 5686 11520
rect 5814 11600 5870 11656
rect 5998 11464 6054 11520
rect 5170 8880 5226 8936
rect 4588 8730 4644 8732
rect 4668 8730 4724 8732
rect 4748 8730 4804 8732
rect 4828 8730 4884 8732
rect 4588 8678 4614 8730
rect 4614 8678 4644 8730
rect 4668 8678 4678 8730
rect 4678 8678 4724 8730
rect 4748 8678 4794 8730
rect 4794 8678 4804 8730
rect 4828 8678 4858 8730
rect 4858 8678 4884 8730
rect 4588 8676 4644 8678
rect 4668 8676 4724 8678
rect 4748 8676 4804 8678
rect 4828 8676 4884 8678
rect 5354 8608 5410 8664
rect 5078 8472 5134 8528
rect 5814 9152 5870 9208
rect 6182 11328 6238 11384
rect 5262 8200 5318 8256
rect 4434 7828 4436 7848
rect 4436 7828 4488 7848
rect 4488 7828 4490 7848
rect 4434 7792 4490 7828
rect 4588 7642 4644 7644
rect 4668 7642 4724 7644
rect 4748 7642 4804 7644
rect 4828 7642 4884 7644
rect 4588 7590 4614 7642
rect 4614 7590 4644 7642
rect 4668 7590 4678 7642
rect 4678 7590 4724 7642
rect 4748 7590 4794 7642
rect 4794 7590 4804 7642
rect 4828 7590 4858 7642
rect 4858 7590 4884 7642
rect 4588 7588 4644 7590
rect 4668 7588 4724 7590
rect 4748 7588 4804 7590
rect 4828 7588 4884 7590
rect 5446 7928 5502 7984
rect 4710 6976 4766 7032
rect 4588 6554 4644 6556
rect 4668 6554 4724 6556
rect 4748 6554 4804 6556
rect 4828 6554 4884 6556
rect 4588 6502 4614 6554
rect 4614 6502 4644 6554
rect 4668 6502 4678 6554
rect 4678 6502 4724 6554
rect 4748 6502 4794 6554
rect 4794 6502 4804 6554
rect 4828 6502 4858 6554
rect 4858 6502 4884 6554
rect 4588 6500 4644 6502
rect 4668 6500 4724 6502
rect 4748 6500 4804 6502
rect 4828 6500 4884 6502
rect 7194 17448 7250 17504
rect 6550 16652 6606 16688
rect 6550 16632 6552 16652
rect 6552 16632 6604 16652
rect 6604 16632 6606 16652
rect 6550 16396 6552 16416
rect 6552 16396 6604 16416
rect 6604 16396 6606 16416
rect 6550 16360 6606 16396
rect 6550 9560 6606 9616
rect 6550 9016 6606 9072
rect 6366 7520 6422 7576
rect 8220 21242 8276 21244
rect 8300 21242 8356 21244
rect 8380 21242 8436 21244
rect 8460 21242 8516 21244
rect 8220 21190 8246 21242
rect 8246 21190 8276 21242
rect 8300 21190 8310 21242
rect 8310 21190 8356 21242
rect 8380 21190 8426 21242
rect 8426 21190 8436 21242
rect 8460 21190 8490 21242
rect 8490 21190 8516 21242
rect 8220 21188 8276 21190
rect 8300 21188 8356 21190
rect 8380 21188 8436 21190
rect 8460 21188 8516 21190
rect 8666 21392 8722 21448
rect 8220 20154 8276 20156
rect 8300 20154 8356 20156
rect 8380 20154 8436 20156
rect 8460 20154 8516 20156
rect 8220 20102 8246 20154
rect 8246 20102 8276 20154
rect 8300 20102 8310 20154
rect 8310 20102 8356 20154
rect 8380 20102 8426 20154
rect 8426 20102 8436 20154
rect 8460 20102 8490 20154
rect 8490 20102 8516 20154
rect 8220 20100 8276 20102
rect 8300 20100 8356 20102
rect 8380 20100 8436 20102
rect 8460 20100 8516 20102
rect 8206 19352 8262 19408
rect 8220 19066 8276 19068
rect 8300 19066 8356 19068
rect 8380 19066 8436 19068
rect 8460 19066 8516 19068
rect 8220 19014 8246 19066
rect 8246 19014 8276 19066
rect 8300 19014 8310 19066
rect 8310 19014 8356 19066
rect 8380 19014 8426 19066
rect 8426 19014 8436 19066
rect 8460 19014 8490 19066
rect 8490 19014 8516 19066
rect 8220 19012 8276 19014
rect 8300 19012 8356 19014
rect 8380 19012 8436 19014
rect 8460 19012 8516 19014
rect 7838 17620 7840 17640
rect 7840 17620 7892 17640
rect 7892 17620 7894 17640
rect 7838 17584 7894 17620
rect 8220 17978 8276 17980
rect 8300 17978 8356 17980
rect 8380 17978 8436 17980
rect 8460 17978 8516 17980
rect 8220 17926 8246 17978
rect 8246 17926 8276 17978
rect 8300 17926 8310 17978
rect 8310 17926 8356 17978
rect 8380 17926 8426 17978
rect 8426 17926 8436 17978
rect 8460 17926 8490 17978
rect 8490 17926 8516 17978
rect 8220 17924 8276 17926
rect 8300 17924 8356 17926
rect 8380 17924 8436 17926
rect 8460 17924 8516 17926
rect 8220 16890 8276 16892
rect 8300 16890 8356 16892
rect 8380 16890 8436 16892
rect 8460 16890 8516 16892
rect 8220 16838 8246 16890
rect 8246 16838 8276 16890
rect 8300 16838 8310 16890
rect 8310 16838 8356 16890
rect 8380 16838 8426 16890
rect 8426 16838 8436 16890
rect 8460 16838 8490 16890
rect 8490 16838 8516 16890
rect 8220 16836 8276 16838
rect 8300 16836 8356 16838
rect 8380 16836 8436 16838
rect 8460 16836 8516 16838
rect 8220 15802 8276 15804
rect 8300 15802 8356 15804
rect 8380 15802 8436 15804
rect 8460 15802 8516 15804
rect 8220 15750 8246 15802
rect 8246 15750 8276 15802
rect 8300 15750 8310 15802
rect 8310 15750 8356 15802
rect 8380 15750 8426 15802
rect 8426 15750 8436 15802
rect 8460 15750 8490 15802
rect 8490 15750 8516 15802
rect 8220 15748 8276 15750
rect 8300 15748 8356 15750
rect 8380 15748 8436 15750
rect 8460 15748 8516 15750
rect 7562 12280 7618 12336
rect 7194 10920 7250 10976
rect 8220 14714 8276 14716
rect 8300 14714 8356 14716
rect 8380 14714 8436 14716
rect 8460 14714 8516 14716
rect 8220 14662 8246 14714
rect 8246 14662 8276 14714
rect 8300 14662 8310 14714
rect 8310 14662 8356 14714
rect 8380 14662 8426 14714
rect 8426 14662 8436 14714
rect 8460 14662 8490 14714
rect 8490 14662 8516 14714
rect 8220 14660 8276 14662
rect 8300 14660 8356 14662
rect 8380 14660 8436 14662
rect 8460 14660 8516 14662
rect 8850 19624 8906 19680
rect 8022 13504 8078 13560
rect 7470 10648 7526 10704
rect 7470 9868 7472 9888
rect 7472 9868 7524 9888
rect 7524 9868 7526 9888
rect 7470 9832 7526 9868
rect 7562 9016 7618 9072
rect 4588 5466 4644 5468
rect 4668 5466 4724 5468
rect 4748 5466 4804 5468
rect 4828 5466 4884 5468
rect 4588 5414 4614 5466
rect 4614 5414 4644 5466
rect 4668 5414 4678 5466
rect 4678 5414 4724 5466
rect 4748 5414 4794 5466
rect 4794 5414 4804 5466
rect 4828 5414 4858 5466
rect 4858 5414 4884 5466
rect 4588 5412 4644 5414
rect 4668 5412 4724 5414
rect 4748 5412 4804 5414
rect 4828 5412 4884 5414
rect 4588 4378 4644 4380
rect 4668 4378 4724 4380
rect 4748 4378 4804 4380
rect 4828 4378 4884 4380
rect 4588 4326 4614 4378
rect 4614 4326 4644 4378
rect 4668 4326 4678 4378
rect 4678 4326 4724 4378
rect 4748 4326 4794 4378
rect 4794 4326 4804 4378
rect 4828 4326 4858 4378
rect 4858 4326 4884 4378
rect 4588 4324 4644 4326
rect 4668 4324 4724 4326
rect 4748 4324 4804 4326
rect 4828 4324 4884 4326
rect 3606 3984 3662 4040
rect 4588 3290 4644 3292
rect 4668 3290 4724 3292
rect 4748 3290 4804 3292
rect 4828 3290 4884 3292
rect 4588 3238 4614 3290
rect 4614 3238 4644 3290
rect 4668 3238 4678 3290
rect 4678 3238 4724 3290
rect 4748 3238 4794 3290
rect 4794 3238 4804 3290
rect 4828 3238 4858 3290
rect 4858 3238 4884 3290
rect 4588 3236 4644 3238
rect 4668 3236 4724 3238
rect 4748 3236 4804 3238
rect 4828 3236 4884 3238
rect 7286 7384 7342 7440
rect 8220 13626 8276 13628
rect 8300 13626 8356 13628
rect 8380 13626 8436 13628
rect 8460 13626 8516 13628
rect 8220 13574 8246 13626
rect 8246 13574 8276 13626
rect 8300 13574 8310 13626
rect 8310 13574 8356 13626
rect 8380 13574 8426 13626
rect 8426 13574 8436 13626
rect 8460 13574 8490 13626
rect 8490 13574 8516 13626
rect 8220 13572 8276 13574
rect 8300 13572 8356 13574
rect 8380 13572 8436 13574
rect 8460 13572 8516 13574
rect 8220 12538 8276 12540
rect 8300 12538 8356 12540
rect 8380 12538 8436 12540
rect 8460 12538 8516 12540
rect 8220 12486 8246 12538
rect 8246 12486 8276 12538
rect 8300 12486 8310 12538
rect 8310 12486 8356 12538
rect 8380 12486 8426 12538
rect 8426 12486 8436 12538
rect 8460 12486 8490 12538
rect 8490 12486 8516 12538
rect 8220 12484 8276 12486
rect 8300 12484 8356 12486
rect 8380 12484 8436 12486
rect 8460 12484 8516 12486
rect 8114 11736 8170 11792
rect 7838 10784 7894 10840
rect 8220 11450 8276 11452
rect 8300 11450 8356 11452
rect 8380 11450 8436 11452
rect 8460 11450 8516 11452
rect 8220 11398 8246 11450
rect 8246 11398 8276 11450
rect 8300 11398 8310 11450
rect 8310 11398 8356 11450
rect 8380 11398 8426 11450
rect 8426 11398 8436 11450
rect 8460 11398 8490 11450
rect 8490 11398 8516 11450
rect 8220 11396 8276 11398
rect 8300 11396 8356 11398
rect 8380 11396 8436 11398
rect 8460 11396 8516 11398
rect 7930 10512 7986 10568
rect 8220 10362 8276 10364
rect 8300 10362 8356 10364
rect 8380 10362 8436 10364
rect 8460 10362 8516 10364
rect 8220 10310 8246 10362
rect 8246 10310 8276 10362
rect 8300 10310 8310 10362
rect 8310 10310 8356 10362
rect 8380 10310 8426 10362
rect 8426 10310 8436 10362
rect 8460 10310 8490 10362
rect 8490 10310 8516 10362
rect 8220 10308 8276 10310
rect 8300 10308 8356 10310
rect 8380 10308 8436 10310
rect 8460 10308 8516 10310
rect 8022 10240 8078 10296
rect 8022 9832 8078 9888
rect 8114 9424 8170 9480
rect 8022 9288 8078 9344
rect 7838 9152 7894 9208
rect 9218 19780 9274 19816
rect 9218 19760 9220 19780
rect 9220 19760 9272 19780
rect 9272 19760 9274 19780
rect 9310 19216 9366 19272
rect 9034 16360 9090 16416
rect 8942 9696 8998 9752
rect 9310 10784 9366 10840
rect 9586 19116 9588 19136
rect 9588 19116 9640 19136
rect 9640 19116 9642 19136
rect 9586 19080 9642 19116
rect 9586 17060 9642 17096
rect 9586 17040 9588 17060
rect 9588 17040 9640 17060
rect 9640 17040 9642 17060
rect 9862 17992 9918 18048
rect 9586 16632 9642 16688
rect 9494 11872 9550 11928
rect 9494 10376 9550 10432
rect 9126 9696 9182 9752
rect 8220 9274 8276 9276
rect 8300 9274 8356 9276
rect 8380 9274 8436 9276
rect 8460 9274 8516 9276
rect 8220 9222 8246 9274
rect 8246 9222 8276 9274
rect 8300 9222 8310 9274
rect 8310 9222 8356 9274
rect 8380 9222 8426 9274
rect 8426 9222 8436 9274
rect 8460 9222 8490 9274
rect 8490 9222 8516 9274
rect 8220 9220 8276 9222
rect 8300 9220 8356 9222
rect 8380 9220 8436 9222
rect 8460 9220 8516 9222
rect 7562 7656 7618 7712
rect 8220 8186 8276 8188
rect 8300 8186 8356 8188
rect 8380 8186 8436 8188
rect 8460 8186 8516 8188
rect 8220 8134 8246 8186
rect 8246 8134 8276 8186
rect 8300 8134 8310 8186
rect 8310 8134 8356 8186
rect 8380 8134 8426 8186
rect 8426 8134 8436 8186
rect 8460 8134 8490 8186
rect 8490 8134 8516 8186
rect 8220 8132 8276 8134
rect 8300 8132 8356 8134
rect 8380 8132 8436 8134
rect 8460 8132 8516 8134
rect 8850 7928 8906 7984
rect 9310 9016 9366 9072
rect 10322 20032 10378 20088
rect 10598 19352 10654 19408
rect 10230 18944 10286 19000
rect 10966 20440 11022 20496
rect 11852 21786 11908 21788
rect 11932 21786 11988 21788
rect 12012 21786 12068 21788
rect 12092 21786 12148 21788
rect 11852 21734 11878 21786
rect 11878 21734 11908 21786
rect 11932 21734 11942 21786
rect 11942 21734 11988 21786
rect 12012 21734 12058 21786
rect 12058 21734 12068 21786
rect 12092 21734 12122 21786
rect 12122 21734 12148 21786
rect 11852 21732 11908 21734
rect 11932 21732 11988 21734
rect 12012 21732 12068 21734
rect 12092 21732 12148 21734
rect 11852 20698 11908 20700
rect 11932 20698 11988 20700
rect 12012 20698 12068 20700
rect 12092 20698 12148 20700
rect 11852 20646 11878 20698
rect 11878 20646 11908 20698
rect 11932 20646 11942 20698
rect 11942 20646 11988 20698
rect 12012 20646 12058 20698
rect 12058 20646 12068 20698
rect 12092 20646 12122 20698
rect 12122 20646 12148 20698
rect 11852 20644 11908 20646
rect 11932 20644 11988 20646
rect 12012 20644 12068 20646
rect 12092 20644 12148 20646
rect 11058 19080 11114 19136
rect 11334 19352 11390 19408
rect 10230 12180 10232 12200
rect 10232 12180 10284 12200
rect 10284 12180 10286 12200
rect 10230 12144 10286 12180
rect 10138 10240 10194 10296
rect 10046 10104 10102 10160
rect 9954 9832 10010 9888
rect 10690 12436 10746 12472
rect 10690 12416 10692 12436
rect 10692 12416 10744 12436
rect 10744 12416 10746 12436
rect 9954 9016 10010 9072
rect 9494 8336 9550 8392
rect 8220 7098 8276 7100
rect 8300 7098 8356 7100
rect 8380 7098 8436 7100
rect 8460 7098 8516 7100
rect 8220 7046 8246 7098
rect 8246 7046 8276 7098
rect 8300 7046 8310 7098
rect 8310 7046 8356 7098
rect 8380 7046 8426 7098
rect 8426 7046 8436 7098
rect 8460 7046 8490 7098
rect 8490 7046 8516 7098
rect 8220 7044 8276 7046
rect 8300 7044 8356 7046
rect 8380 7044 8436 7046
rect 8460 7044 8516 7046
rect 8114 6432 8170 6488
rect 8022 6332 8024 6352
rect 8024 6332 8076 6352
rect 8076 6332 8078 6352
rect 8022 6296 8078 6332
rect 8220 6010 8276 6012
rect 8300 6010 8356 6012
rect 8380 6010 8436 6012
rect 8460 6010 8516 6012
rect 8220 5958 8246 6010
rect 8246 5958 8276 6010
rect 8300 5958 8310 6010
rect 8310 5958 8356 6010
rect 8380 5958 8426 6010
rect 8426 5958 8436 6010
rect 8460 5958 8490 6010
rect 8490 5958 8516 6010
rect 8220 5956 8276 5958
rect 8300 5956 8356 5958
rect 8380 5956 8436 5958
rect 8460 5956 8516 5958
rect 8220 4922 8276 4924
rect 8300 4922 8356 4924
rect 8380 4922 8436 4924
rect 8460 4922 8516 4924
rect 8220 4870 8246 4922
rect 8246 4870 8276 4922
rect 8300 4870 8310 4922
rect 8310 4870 8356 4922
rect 8380 4870 8426 4922
rect 8426 4870 8436 4922
rect 8460 4870 8490 4922
rect 8490 4870 8516 4922
rect 8220 4868 8276 4870
rect 8300 4868 8356 4870
rect 8380 4868 8436 4870
rect 8460 4868 8516 4870
rect 7746 4120 7802 4176
rect 9494 6432 9550 6488
rect 10046 4820 10102 4856
rect 10046 4800 10048 4820
rect 10048 4800 10100 4820
rect 10100 4800 10102 4820
rect 12070 19760 12126 19816
rect 11852 19610 11908 19612
rect 11932 19610 11988 19612
rect 12012 19610 12068 19612
rect 12092 19610 12148 19612
rect 11852 19558 11878 19610
rect 11878 19558 11908 19610
rect 11932 19558 11942 19610
rect 11942 19558 11988 19610
rect 12012 19558 12058 19610
rect 12058 19558 12068 19610
rect 12092 19558 12122 19610
rect 12122 19558 12148 19610
rect 11852 19556 11908 19558
rect 11932 19556 11988 19558
rect 12012 19556 12068 19558
rect 12092 19556 12148 19558
rect 12622 20576 12678 20632
rect 12530 19796 12532 19816
rect 12532 19796 12584 19816
rect 12584 19796 12586 19816
rect 12530 19760 12586 19796
rect 12530 19660 12532 19680
rect 12532 19660 12584 19680
rect 12584 19660 12586 19680
rect 12530 19624 12586 19660
rect 12622 19352 12678 19408
rect 12254 19236 12310 19272
rect 12254 19216 12256 19236
rect 12256 19216 12308 19236
rect 12308 19216 12310 19236
rect 12530 19236 12586 19272
rect 12530 19216 12532 19236
rect 12532 19216 12584 19236
rect 12584 19216 12586 19236
rect 12162 18844 12164 18864
rect 12164 18844 12216 18864
rect 12216 18844 12218 18864
rect 12162 18808 12218 18844
rect 11852 18522 11908 18524
rect 11932 18522 11988 18524
rect 12012 18522 12068 18524
rect 12092 18522 12148 18524
rect 11852 18470 11878 18522
rect 11878 18470 11908 18522
rect 11932 18470 11942 18522
rect 11942 18470 11988 18522
rect 12012 18470 12058 18522
rect 12058 18470 12068 18522
rect 12092 18470 12122 18522
rect 12122 18470 12148 18522
rect 11852 18468 11908 18470
rect 11932 18468 11988 18470
rect 12012 18468 12068 18470
rect 12092 18468 12148 18470
rect 12254 18400 12310 18456
rect 11852 17434 11908 17436
rect 11932 17434 11988 17436
rect 12012 17434 12068 17436
rect 12092 17434 12148 17436
rect 11852 17382 11878 17434
rect 11878 17382 11908 17434
rect 11932 17382 11942 17434
rect 11942 17382 11988 17434
rect 12012 17382 12058 17434
rect 12058 17382 12068 17434
rect 12092 17382 12122 17434
rect 12122 17382 12148 17434
rect 11852 17380 11908 17382
rect 11932 17380 11988 17382
rect 12012 17380 12068 17382
rect 12092 17380 12148 17382
rect 11852 16346 11908 16348
rect 11932 16346 11988 16348
rect 12012 16346 12068 16348
rect 12092 16346 12148 16348
rect 11852 16294 11878 16346
rect 11878 16294 11908 16346
rect 11932 16294 11942 16346
rect 11942 16294 11988 16346
rect 12012 16294 12058 16346
rect 12058 16294 12068 16346
rect 12092 16294 12122 16346
rect 12122 16294 12148 16346
rect 11852 16292 11908 16294
rect 11932 16292 11988 16294
rect 12012 16292 12068 16294
rect 12092 16292 12148 16294
rect 12346 17584 12402 17640
rect 12438 17332 12494 17368
rect 12438 17312 12440 17332
rect 12440 17312 12492 17332
rect 12492 17312 12494 17332
rect 12530 16496 12586 16552
rect 12254 16224 12310 16280
rect 11852 15258 11908 15260
rect 11932 15258 11988 15260
rect 12012 15258 12068 15260
rect 12092 15258 12148 15260
rect 11852 15206 11878 15258
rect 11878 15206 11908 15258
rect 11932 15206 11942 15258
rect 11942 15206 11988 15258
rect 12012 15206 12058 15258
rect 12058 15206 12068 15258
rect 12092 15206 12122 15258
rect 12122 15206 12148 15258
rect 11852 15204 11908 15206
rect 11932 15204 11988 15206
rect 12012 15204 12068 15206
rect 12092 15204 12148 15206
rect 11852 14170 11908 14172
rect 11932 14170 11988 14172
rect 12012 14170 12068 14172
rect 12092 14170 12148 14172
rect 11852 14118 11878 14170
rect 11878 14118 11908 14170
rect 11932 14118 11942 14170
rect 11942 14118 11988 14170
rect 12012 14118 12058 14170
rect 12058 14118 12068 14170
rect 12092 14118 12122 14170
rect 12122 14118 12148 14170
rect 11852 14116 11908 14118
rect 11932 14116 11988 14118
rect 12012 14116 12068 14118
rect 12092 14116 12148 14118
rect 11518 12144 11574 12200
rect 11852 13082 11908 13084
rect 11932 13082 11988 13084
rect 12012 13082 12068 13084
rect 12092 13082 12148 13084
rect 11852 13030 11878 13082
rect 11878 13030 11908 13082
rect 11932 13030 11942 13082
rect 11942 13030 11988 13082
rect 12012 13030 12058 13082
rect 12058 13030 12068 13082
rect 12092 13030 12122 13082
rect 12122 13030 12148 13082
rect 11852 13028 11908 13030
rect 11932 13028 11988 13030
rect 12012 13028 12068 13030
rect 12092 13028 12148 13030
rect 13082 20032 13138 20088
rect 13358 19624 13414 19680
rect 13174 19508 13230 19544
rect 13174 19488 13176 19508
rect 13176 19488 13228 19508
rect 13228 19488 13230 19508
rect 11852 11994 11908 11996
rect 11932 11994 11988 11996
rect 12012 11994 12068 11996
rect 12092 11994 12148 11996
rect 11852 11942 11878 11994
rect 11878 11942 11908 11994
rect 11932 11942 11942 11994
rect 11942 11942 11988 11994
rect 12012 11942 12058 11994
rect 12058 11942 12068 11994
rect 12092 11942 12122 11994
rect 12122 11942 12148 11994
rect 11852 11940 11908 11942
rect 11932 11940 11988 11942
rect 12012 11940 12068 11942
rect 12092 11940 12148 11942
rect 13726 20576 13782 20632
rect 14278 18420 14334 18456
rect 14278 18400 14280 18420
rect 14280 18400 14332 18420
rect 14332 18400 14334 18420
rect 13450 16632 13506 16688
rect 13358 15952 13414 16008
rect 10782 9016 10838 9072
rect 11058 9696 11114 9752
rect 10966 9016 11022 9072
rect 10966 8744 11022 8800
rect 11242 9152 11298 9208
rect 11852 10906 11908 10908
rect 11932 10906 11988 10908
rect 12012 10906 12068 10908
rect 12092 10906 12148 10908
rect 11852 10854 11878 10906
rect 11878 10854 11908 10906
rect 11932 10854 11942 10906
rect 11942 10854 11988 10906
rect 12012 10854 12058 10906
rect 12058 10854 12068 10906
rect 12092 10854 12122 10906
rect 12122 10854 12148 10906
rect 11852 10852 11908 10854
rect 11932 10852 11988 10854
rect 12012 10852 12068 10854
rect 12092 10852 12148 10854
rect 11852 9818 11908 9820
rect 11932 9818 11988 9820
rect 12012 9818 12068 9820
rect 12092 9818 12148 9820
rect 11852 9766 11878 9818
rect 11878 9766 11908 9818
rect 11932 9766 11942 9818
rect 11942 9766 11988 9818
rect 12012 9766 12058 9818
rect 12058 9766 12068 9818
rect 12092 9766 12122 9818
rect 12122 9766 12148 9818
rect 11852 9764 11908 9766
rect 11932 9764 11988 9766
rect 12012 9764 12068 9766
rect 12092 9764 12148 9766
rect 11150 7656 11206 7712
rect 11852 8730 11908 8732
rect 11932 8730 11988 8732
rect 12012 8730 12068 8732
rect 12092 8730 12148 8732
rect 11852 8678 11878 8730
rect 11878 8678 11908 8730
rect 11932 8678 11942 8730
rect 11942 8678 11988 8730
rect 12012 8678 12058 8730
rect 12058 8678 12068 8730
rect 12092 8678 12122 8730
rect 12122 8678 12148 8730
rect 11852 8676 11908 8678
rect 11932 8676 11988 8678
rect 12012 8676 12068 8678
rect 12092 8676 12148 8678
rect 12714 10512 12770 10568
rect 12438 10376 12494 10432
rect 12254 9868 12256 9888
rect 12256 9868 12308 9888
rect 12308 9868 12310 9888
rect 12254 9832 12310 9868
rect 12346 9560 12402 9616
rect 12622 8880 12678 8936
rect 12530 8744 12586 8800
rect 11852 7642 11908 7644
rect 11932 7642 11988 7644
rect 12012 7642 12068 7644
rect 12092 7642 12148 7644
rect 11852 7590 11878 7642
rect 11878 7590 11908 7642
rect 11932 7590 11942 7642
rect 11942 7590 11988 7642
rect 12012 7590 12058 7642
rect 12058 7590 12068 7642
rect 12092 7590 12122 7642
rect 12122 7590 12148 7642
rect 11852 7588 11908 7590
rect 11932 7588 11988 7590
rect 12012 7588 12068 7590
rect 12092 7588 12148 7590
rect 11702 7520 11758 7576
rect 12346 7520 12402 7576
rect 12990 9832 13046 9888
rect 12898 9424 12954 9480
rect 12254 7248 12310 7304
rect 14094 16088 14150 16144
rect 13726 12144 13782 12200
rect 13542 9832 13598 9888
rect 13266 8200 13322 8256
rect 12070 6840 12126 6896
rect 11852 6554 11908 6556
rect 11932 6554 11988 6556
rect 12012 6554 12068 6556
rect 12092 6554 12148 6556
rect 11852 6502 11878 6554
rect 11878 6502 11908 6554
rect 11932 6502 11942 6554
rect 11942 6502 11988 6554
rect 12012 6502 12058 6554
rect 12058 6502 12068 6554
rect 12092 6502 12122 6554
rect 12122 6502 12148 6554
rect 11852 6500 11908 6502
rect 11932 6500 11988 6502
rect 12012 6500 12068 6502
rect 12092 6500 12148 6502
rect 11794 6316 11850 6352
rect 11794 6296 11796 6316
rect 11796 6296 11848 6316
rect 11848 6296 11850 6316
rect 11852 5466 11908 5468
rect 11932 5466 11988 5468
rect 12012 5466 12068 5468
rect 12092 5466 12148 5468
rect 11852 5414 11878 5466
rect 11878 5414 11908 5466
rect 11932 5414 11942 5466
rect 11942 5414 11988 5466
rect 12012 5414 12058 5466
rect 12058 5414 12068 5466
rect 12092 5414 12122 5466
rect 12122 5414 12148 5466
rect 11852 5412 11908 5414
rect 11932 5412 11988 5414
rect 12012 5412 12068 5414
rect 12092 5412 12148 5414
rect 12346 6704 12402 6760
rect 12254 5788 12256 5808
rect 12256 5788 12308 5808
rect 12308 5788 12310 5808
rect 12254 5752 12310 5788
rect 11852 4378 11908 4380
rect 11932 4378 11988 4380
rect 12012 4378 12068 4380
rect 12092 4378 12148 4380
rect 11852 4326 11878 4378
rect 11878 4326 11908 4378
rect 11932 4326 11942 4378
rect 11942 4326 11988 4378
rect 12012 4326 12058 4378
rect 12058 4326 12068 4378
rect 12092 4326 12122 4378
rect 12122 4326 12148 4378
rect 11852 4324 11908 4326
rect 11932 4324 11988 4326
rect 12012 4324 12068 4326
rect 12092 4324 12148 4326
rect 8220 3834 8276 3836
rect 8300 3834 8356 3836
rect 8380 3834 8436 3836
rect 8460 3834 8516 3836
rect 8220 3782 8246 3834
rect 8246 3782 8276 3834
rect 8300 3782 8310 3834
rect 8310 3782 8356 3834
rect 8380 3782 8426 3834
rect 8426 3782 8436 3834
rect 8460 3782 8490 3834
rect 8490 3782 8516 3834
rect 8220 3780 8276 3782
rect 8300 3780 8356 3782
rect 8380 3780 8436 3782
rect 8460 3780 8516 3782
rect 12254 3848 12310 3904
rect 13082 6332 13084 6352
rect 13084 6332 13136 6352
rect 13136 6332 13138 6352
rect 13082 6296 13138 6332
rect 12530 4256 12586 4312
rect 12714 4020 12716 4040
rect 12716 4020 12768 4040
rect 12768 4020 12770 4040
rect 12714 3984 12770 4020
rect 13634 9560 13690 9616
rect 14002 11736 14058 11792
rect 14278 16224 14334 16280
rect 14462 20440 14518 20496
rect 14186 10240 14242 10296
rect 13910 9288 13966 9344
rect 13726 9152 13782 9208
rect 14186 9152 14242 9208
rect 13726 8236 13728 8256
rect 13728 8236 13780 8256
rect 13780 8236 13782 8256
rect 13726 8200 13782 8236
rect 13726 7656 13782 7712
rect 13726 7384 13782 7440
rect 14002 7384 14058 7440
rect 14462 11464 14518 11520
rect 14370 7384 14426 7440
rect 14186 6296 14242 6352
rect 14094 6160 14150 6216
rect 13818 4120 13874 4176
rect 12438 3460 12494 3496
rect 12438 3440 12440 3460
rect 12440 3440 12492 3460
rect 12492 3440 12494 3460
rect 11852 3290 11908 3292
rect 11932 3290 11988 3292
rect 12012 3290 12068 3292
rect 12092 3290 12148 3292
rect 11852 3238 11878 3290
rect 11878 3238 11908 3290
rect 11932 3238 11942 3290
rect 11942 3238 11988 3290
rect 12012 3238 12058 3290
rect 12058 3238 12068 3290
rect 12092 3238 12122 3290
rect 12122 3238 12148 3290
rect 11852 3236 11908 3238
rect 11932 3236 11988 3238
rect 12012 3236 12068 3238
rect 12092 3236 12148 3238
rect 8220 2746 8276 2748
rect 8300 2746 8356 2748
rect 8380 2746 8436 2748
rect 8460 2746 8516 2748
rect 8220 2694 8246 2746
rect 8246 2694 8276 2746
rect 8300 2694 8310 2746
rect 8310 2694 8356 2746
rect 8380 2694 8426 2746
rect 8426 2694 8436 2746
rect 8460 2694 8490 2746
rect 8490 2694 8516 2746
rect 8220 2692 8276 2694
rect 8300 2692 8356 2694
rect 8380 2692 8436 2694
rect 8460 2692 8516 2694
rect 4588 2202 4644 2204
rect 4668 2202 4724 2204
rect 4748 2202 4804 2204
rect 4828 2202 4884 2204
rect 4588 2150 4614 2202
rect 4614 2150 4644 2202
rect 4668 2150 4678 2202
rect 4678 2150 4724 2202
rect 4748 2150 4794 2202
rect 4794 2150 4804 2202
rect 4828 2150 4858 2202
rect 4858 2150 4884 2202
rect 4588 2148 4644 2150
rect 4668 2148 4724 2150
rect 4748 2148 4804 2150
rect 4828 2148 4884 2150
rect 11852 2202 11908 2204
rect 11932 2202 11988 2204
rect 12012 2202 12068 2204
rect 12092 2202 12148 2204
rect 11852 2150 11878 2202
rect 11878 2150 11908 2202
rect 11932 2150 11942 2202
rect 11942 2150 11988 2202
rect 12012 2150 12058 2202
rect 12058 2150 12068 2202
rect 12092 2150 12122 2202
rect 12122 2150 12148 2202
rect 11852 2148 11908 2150
rect 11932 2148 11988 2150
rect 12012 2148 12068 2150
rect 12092 2148 12148 2150
rect 13910 3168 13966 3224
rect 14646 20440 14702 20496
rect 15014 20340 15016 20360
rect 15016 20340 15068 20360
rect 15068 20340 15070 20360
rect 15014 20304 15070 20340
rect 15014 18028 15016 18048
rect 15016 18028 15068 18048
rect 15068 18028 15070 18048
rect 14830 17312 14886 17368
rect 14646 16496 14702 16552
rect 15014 17992 15070 18028
rect 15014 16088 15070 16144
rect 15014 15988 15016 16008
rect 15016 15988 15068 16008
rect 15068 15988 15070 16008
rect 15014 15952 15070 15988
rect 15198 20712 15254 20768
rect 15198 19488 15254 19544
rect 15484 21242 15540 21244
rect 15564 21242 15620 21244
rect 15644 21242 15700 21244
rect 15724 21242 15780 21244
rect 15484 21190 15510 21242
rect 15510 21190 15540 21242
rect 15564 21190 15574 21242
rect 15574 21190 15620 21242
rect 15644 21190 15690 21242
rect 15690 21190 15700 21242
rect 15724 21190 15754 21242
rect 15754 21190 15780 21242
rect 15484 21188 15540 21190
rect 15564 21188 15620 21190
rect 15644 21188 15700 21190
rect 15724 21188 15780 21190
rect 15484 20154 15540 20156
rect 15564 20154 15620 20156
rect 15644 20154 15700 20156
rect 15724 20154 15780 20156
rect 15484 20102 15510 20154
rect 15510 20102 15540 20154
rect 15564 20102 15574 20154
rect 15574 20102 15620 20154
rect 15644 20102 15690 20154
rect 15690 20102 15700 20154
rect 15724 20102 15754 20154
rect 15754 20102 15780 20154
rect 15484 20100 15540 20102
rect 15564 20100 15620 20102
rect 15644 20100 15700 20102
rect 15724 20100 15780 20102
rect 15658 19216 15714 19272
rect 15484 19066 15540 19068
rect 15564 19066 15620 19068
rect 15644 19066 15700 19068
rect 15724 19066 15780 19068
rect 15484 19014 15510 19066
rect 15510 19014 15540 19066
rect 15564 19014 15574 19066
rect 15574 19014 15620 19066
rect 15644 19014 15690 19066
rect 15690 19014 15700 19066
rect 15724 19014 15754 19066
rect 15754 19014 15780 19066
rect 15484 19012 15540 19014
rect 15564 19012 15620 19014
rect 15644 19012 15700 19014
rect 15724 19012 15780 19014
rect 15484 17978 15540 17980
rect 15564 17978 15620 17980
rect 15644 17978 15700 17980
rect 15724 17978 15780 17980
rect 15484 17926 15510 17978
rect 15510 17926 15540 17978
rect 15564 17926 15574 17978
rect 15574 17926 15620 17978
rect 15644 17926 15690 17978
rect 15690 17926 15700 17978
rect 15724 17926 15754 17978
rect 15754 17926 15780 17978
rect 15484 17924 15540 17926
rect 15564 17924 15620 17926
rect 15644 17924 15700 17926
rect 15724 17924 15780 17926
rect 15484 16890 15540 16892
rect 15564 16890 15620 16892
rect 15644 16890 15700 16892
rect 15724 16890 15780 16892
rect 15484 16838 15510 16890
rect 15510 16838 15540 16890
rect 15564 16838 15574 16890
rect 15574 16838 15620 16890
rect 15644 16838 15690 16890
rect 15690 16838 15700 16890
rect 15724 16838 15754 16890
rect 15754 16838 15780 16890
rect 15484 16836 15540 16838
rect 15564 16836 15620 16838
rect 15644 16836 15700 16838
rect 15724 16836 15780 16838
rect 15474 16632 15530 16688
rect 15484 15802 15540 15804
rect 15564 15802 15620 15804
rect 15644 15802 15700 15804
rect 15724 15802 15780 15804
rect 15484 15750 15510 15802
rect 15510 15750 15540 15802
rect 15564 15750 15574 15802
rect 15574 15750 15620 15802
rect 15644 15750 15690 15802
rect 15690 15750 15700 15802
rect 15724 15750 15754 15802
rect 15754 15750 15780 15802
rect 15484 15748 15540 15750
rect 15564 15748 15620 15750
rect 15644 15748 15700 15750
rect 15724 15748 15780 15750
rect 15750 15020 15806 15056
rect 15750 15000 15752 15020
rect 15752 15000 15804 15020
rect 15804 15000 15806 15020
rect 14830 12416 14886 12472
rect 14738 11464 14794 11520
rect 15484 14714 15540 14716
rect 15564 14714 15620 14716
rect 15644 14714 15700 14716
rect 15724 14714 15780 14716
rect 15484 14662 15510 14714
rect 15510 14662 15540 14714
rect 15564 14662 15574 14714
rect 15574 14662 15620 14714
rect 15644 14662 15690 14714
rect 15690 14662 15700 14714
rect 15724 14662 15754 14714
rect 15754 14662 15780 14714
rect 15484 14660 15540 14662
rect 15564 14660 15620 14662
rect 15644 14660 15700 14662
rect 15724 14660 15780 14662
rect 15484 13626 15540 13628
rect 15564 13626 15620 13628
rect 15644 13626 15700 13628
rect 15724 13626 15780 13628
rect 15484 13574 15510 13626
rect 15510 13574 15540 13626
rect 15564 13574 15574 13626
rect 15574 13574 15620 13626
rect 15644 13574 15690 13626
rect 15690 13574 15700 13626
rect 15724 13574 15754 13626
rect 15754 13574 15780 13626
rect 15484 13572 15540 13574
rect 15564 13572 15620 13574
rect 15644 13572 15700 13574
rect 15724 13572 15780 13574
rect 15382 12688 15438 12744
rect 16118 18264 16174 18320
rect 15842 12824 15898 12880
rect 15484 12538 15540 12540
rect 15564 12538 15620 12540
rect 15644 12538 15700 12540
rect 15724 12538 15780 12540
rect 15484 12486 15510 12538
rect 15510 12486 15540 12538
rect 15564 12486 15574 12538
rect 15574 12486 15620 12538
rect 15644 12486 15690 12538
rect 15690 12486 15700 12538
rect 15724 12486 15754 12538
rect 15754 12486 15780 12538
rect 15484 12484 15540 12486
rect 15564 12484 15620 12486
rect 15644 12484 15700 12486
rect 15724 12484 15780 12486
rect 15106 12008 15162 12064
rect 15014 11772 15016 11792
rect 15016 11772 15068 11792
rect 15068 11772 15070 11792
rect 15014 11736 15070 11772
rect 14830 9560 14886 9616
rect 14738 8336 14794 8392
rect 14370 5752 14426 5808
rect 14646 3596 14702 3632
rect 14646 3576 14648 3596
rect 14648 3576 14700 3596
rect 14700 3576 14702 3596
rect 15290 11600 15346 11656
rect 16118 14592 16174 14648
rect 16118 14220 16120 14240
rect 16120 14220 16172 14240
rect 16172 14220 16174 14240
rect 16118 14184 16174 14220
rect 19430 23432 19486 23488
rect 19614 22752 19670 22808
rect 19338 22072 19394 22128
rect 19116 21786 19172 21788
rect 19196 21786 19252 21788
rect 19276 21786 19332 21788
rect 19356 21786 19412 21788
rect 19116 21734 19142 21786
rect 19142 21734 19172 21786
rect 19196 21734 19206 21786
rect 19206 21734 19252 21786
rect 19276 21734 19322 21786
rect 19322 21734 19332 21786
rect 19356 21734 19386 21786
rect 19386 21734 19412 21786
rect 19116 21732 19172 21734
rect 19196 21732 19252 21734
rect 19276 21732 19332 21734
rect 19356 21732 19412 21734
rect 16670 18128 16726 18184
rect 16394 16224 16450 16280
rect 16026 12960 16082 13016
rect 15750 11872 15806 11928
rect 16026 11600 16082 11656
rect 15484 11450 15540 11452
rect 15564 11450 15620 11452
rect 15644 11450 15700 11452
rect 15724 11450 15780 11452
rect 15484 11398 15510 11450
rect 15510 11398 15540 11450
rect 15564 11398 15574 11450
rect 15574 11398 15620 11450
rect 15644 11398 15690 11450
rect 15690 11398 15700 11450
rect 15724 11398 15754 11450
rect 15754 11398 15780 11450
rect 15484 11396 15540 11398
rect 15564 11396 15620 11398
rect 15644 11396 15700 11398
rect 15724 11396 15780 11398
rect 15382 11092 15384 11112
rect 15384 11092 15436 11112
rect 15436 11092 15438 11112
rect 15382 11056 15438 11092
rect 15290 10920 15346 10976
rect 15934 10648 15990 10704
rect 15484 10362 15540 10364
rect 15564 10362 15620 10364
rect 15644 10362 15700 10364
rect 15724 10362 15780 10364
rect 15484 10310 15510 10362
rect 15510 10310 15540 10362
rect 15564 10310 15574 10362
rect 15574 10310 15620 10362
rect 15644 10310 15690 10362
rect 15690 10310 15700 10362
rect 15724 10310 15754 10362
rect 15754 10310 15780 10362
rect 15484 10308 15540 10310
rect 15564 10308 15620 10310
rect 15644 10308 15700 10310
rect 15724 10308 15780 10310
rect 15382 10124 15438 10160
rect 15382 10104 15384 10124
rect 15384 10104 15436 10124
rect 15436 10104 15438 10124
rect 15290 9968 15346 10024
rect 15934 9288 15990 9344
rect 15484 9274 15540 9276
rect 15564 9274 15620 9276
rect 15644 9274 15700 9276
rect 15724 9274 15780 9276
rect 15484 9222 15510 9274
rect 15510 9222 15540 9274
rect 15564 9222 15574 9274
rect 15574 9222 15620 9274
rect 15644 9222 15690 9274
rect 15690 9222 15700 9274
rect 15724 9222 15754 9274
rect 15754 9222 15780 9274
rect 15484 9220 15540 9222
rect 15564 9220 15620 9222
rect 15644 9220 15700 9222
rect 15724 9220 15780 9222
rect 15106 6840 15162 6896
rect 15484 8186 15540 8188
rect 15564 8186 15620 8188
rect 15644 8186 15700 8188
rect 15724 8186 15780 8188
rect 15484 8134 15510 8186
rect 15510 8134 15540 8186
rect 15564 8134 15574 8186
rect 15574 8134 15620 8186
rect 15644 8134 15690 8186
rect 15690 8134 15700 8186
rect 15724 8134 15754 8186
rect 15754 8134 15780 8186
rect 15484 8132 15540 8134
rect 15564 8132 15620 8134
rect 15644 8132 15700 8134
rect 15724 8132 15780 8134
rect 15382 7520 15438 7576
rect 15474 7248 15530 7304
rect 15484 7098 15540 7100
rect 15564 7098 15620 7100
rect 15644 7098 15700 7100
rect 15724 7098 15780 7100
rect 15484 7046 15510 7098
rect 15510 7046 15540 7098
rect 15564 7046 15574 7098
rect 15574 7046 15620 7098
rect 15644 7046 15690 7098
rect 15690 7046 15700 7098
rect 15724 7046 15754 7098
rect 15754 7046 15780 7098
rect 15484 7044 15540 7046
rect 15564 7044 15620 7046
rect 15644 7044 15700 7046
rect 15724 7044 15780 7046
rect 14922 4800 14978 4856
rect 15198 3848 15254 3904
rect 15484 6010 15540 6012
rect 15564 6010 15620 6012
rect 15644 6010 15700 6012
rect 15724 6010 15780 6012
rect 15484 5958 15510 6010
rect 15510 5958 15540 6010
rect 15564 5958 15574 6010
rect 15574 5958 15620 6010
rect 15644 5958 15690 6010
rect 15690 5958 15700 6010
rect 15724 5958 15754 6010
rect 15754 5958 15780 6010
rect 15484 5956 15540 5958
rect 15564 5956 15620 5958
rect 15644 5956 15700 5958
rect 15724 5956 15780 5958
rect 15484 4922 15540 4924
rect 15564 4922 15620 4924
rect 15644 4922 15700 4924
rect 15724 4922 15780 4924
rect 15484 4870 15510 4922
rect 15510 4870 15540 4922
rect 15564 4870 15574 4922
rect 15574 4870 15620 4922
rect 15644 4870 15690 4922
rect 15690 4870 15700 4922
rect 15724 4870 15754 4922
rect 15754 4870 15780 4922
rect 15484 4868 15540 4870
rect 15564 4868 15620 4870
rect 15644 4868 15700 4870
rect 15724 4868 15780 4870
rect 16854 20712 16910 20768
rect 16854 20324 16910 20360
rect 16854 20304 16856 20324
rect 16856 20304 16908 20324
rect 16908 20304 16910 20324
rect 17038 20576 17094 20632
rect 17038 20304 17094 20360
rect 16854 18808 16910 18864
rect 16394 13096 16450 13152
rect 16210 11600 16266 11656
rect 16578 9968 16634 10024
rect 16946 11600 17002 11656
rect 16762 10784 16818 10840
rect 16394 8336 16450 8392
rect 16670 7384 16726 7440
rect 16210 6704 16266 6760
rect 16302 6024 16358 6080
rect 16210 5344 16266 5400
rect 16118 4256 16174 4312
rect 16026 3984 16082 4040
rect 15484 3834 15540 3836
rect 15564 3834 15620 3836
rect 15644 3834 15700 3836
rect 15724 3834 15780 3836
rect 15484 3782 15510 3834
rect 15510 3782 15540 3834
rect 15564 3782 15574 3834
rect 15574 3782 15620 3834
rect 15644 3782 15690 3834
rect 15690 3782 15700 3834
rect 15724 3782 15754 3834
rect 15754 3782 15780 3834
rect 15484 3780 15540 3782
rect 15564 3780 15620 3782
rect 15644 3780 15700 3782
rect 15724 3780 15780 3782
rect 15842 3596 15898 3632
rect 15842 3576 15844 3596
rect 15844 3576 15896 3596
rect 15896 3576 15898 3596
rect 15382 3440 15438 3496
rect 15484 2746 15540 2748
rect 15564 2746 15620 2748
rect 15644 2746 15700 2748
rect 15724 2746 15780 2748
rect 15484 2694 15510 2746
rect 15510 2694 15540 2746
rect 15564 2694 15574 2746
rect 15574 2694 15620 2746
rect 15644 2694 15690 2746
rect 15690 2694 15700 2746
rect 15724 2694 15754 2746
rect 15754 2694 15780 2746
rect 15484 2692 15540 2694
rect 15564 2692 15620 2694
rect 15644 2692 15700 2694
rect 15724 2692 15780 2694
rect 17130 14728 17186 14784
rect 17314 15020 17370 15056
rect 17314 15000 17316 15020
rect 17316 15000 17368 15020
rect 17368 15000 17370 15020
rect 19116 20698 19172 20700
rect 19196 20698 19252 20700
rect 19276 20698 19332 20700
rect 19356 20698 19412 20700
rect 19116 20646 19142 20698
rect 19142 20646 19172 20698
rect 19196 20646 19206 20698
rect 19206 20646 19252 20698
rect 19276 20646 19322 20698
rect 19322 20646 19332 20698
rect 19356 20646 19386 20698
rect 19386 20646 19412 20698
rect 19116 20644 19172 20646
rect 19196 20644 19252 20646
rect 19276 20644 19332 20646
rect 19356 20644 19412 20646
rect 18418 18672 18474 18728
rect 17958 14220 17960 14240
rect 17960 14220 18012 14240
rect 18012 14220 18014 14240
rect 17958 14184 18014 14220
rect 18142 13368 18198 13424
rect 17314 11736 17370 11792
rect 17314 11056 17370 11112
rect 17314 10784 17370 10840
rect 17222 9424 17278 9480
rect 17406 10548 17408 10568
rect 17408 10548 17460 10568
rect 17460 10548 17462 10568
rect 17406 10512 17462 10548
rect 17590 11600 17646 11656
rect 17498 8880 17554 8936
rect 17774 11212 17830 11248
rect 17774 11192 17776 11212
rect 17776 11192 17828 11212
rect 17828 11192 17830 11212
rect 17774 10956 17776 10976
rect 17776 10956 17828 10976
rect 17828 10956 17830 10976
rect 17774 10920 17830 10956
rect 18326 11872 18382 11928
rect 18418 11056 18474 11112
rect 19522 20576 19578 20632
rect 19614 19896 19670 19952
rect 19116 19610 19172 19612
rect 19196 19610 19252 19612
rect 19276 19610 19332 19612
rect 19356 19610 19412 19612
rect 19116 19558 19142 19610
rect 19142 19558 19172 19610
rect 19196 19558 19206 19610
rect 19206 19558 19252 19610
rect 19276 19558 19322 19610
rect 19322 19558 19332 19610
rect 19356 19558 19386 19610
rect 19386 19558 19412 19610
rect 19116 19556 19172 19558
rect 19196 19556 19252 19558
rect 19276 19556 19332 19558
rect 19356 19556 19412 19558
rect 19154 18708 19156 18728
rect 19156 18708 19208 18728
rect 19208 18708 19210 18728
rect 19154 18672 19210 18708
rect 19116 18522 19172 18524
rect 19196 18522 19252 18524
rect 19276 18522 19332 18524
rect 19356 18522 19412 18524
rect 19116 18470 19142 18522
rect 19142 18470 19172 18522
rect 19196 18470 19206 18522
rect 19206 18470 19252 18522
rect 19276 18470 19322 18522
rect 19322 18470 19332 18522
rect 19356 18470 19386 18522
rect 19386 18470 19412 18522
rect 19116 18468 19172 18470
rect 19196 18468 19252 18470
rect 19276 18468 19332 18470
rect 19356 18468 19412 18470
rect 19614 18420 19670 18456
rect 19614 18400 19616 18420
rect 19616 18400 19668 18420
rect 19668 18400 19670 18420
rect 18970 17584 19026 17640
rect 19116 17434 19172 17436
rect 19196 17434 19252 17436
rect 19276 17434 19332 17436
rect 19356 17434 19412 17436
rect 19116 17382 19142 17434
rect 19142 17382 19172 17434
rect 19196 17382 19206 17434
rect 19206 17382 19252 17434
rect 19276 17382 19322 17434
rect 19322 17382 19332 17434
rect 19356 17382 19386 17434
rect 19386 17382 19412 17434
rect 19116 17380 19172 17382
rect 19196 17380 19252 17382
rect 19276 17380 19332 17382
rect 19356 17380 19412 17382
rect 19982 21256 20038 21312
rect 19706 17312 19762 17368
rect 19116 16346 19172 16348
rect 19196 16346 19252 16348
rect 19276 16346 19332 16348
rect 19356 16346 19412 16348
rect 19116 16294 19142 16346
rect 19142 16294 19172 16346
rect 19196 16294 19206 16346
rect 19206 16294 19252 16346
rect 19276 16294 19322 16346
rect 19322 16294 19332 16346
rect 19356 16294 19386 16346
rect 19386 16294 19412 16346
rect 19116 16292 19172 16294
rect 19196 16292 19252 16294
rect 19276 16292 19332 16294
rect 19356 16292 19412 16294
rect 19116 15258 19172 15260
rect 19196 15258 19252 15260
rect 19276 15258 19332 15260
rect 19356 15258 19412 15260
rect 19116 15206 19142 15258
rect 19142 15206 19172 15258
rect 19196 15206 19206 15258
rect 19206 15206 19252 15258
rect 19276 15206 19322 15258
rect 19322 15206 19332 15258
rect 19356 15206 19386 15258
rect 19386 15206 19412 15258
rect 19116 15204 19172 15206
rect 19196 15204 19252 15206
rect 19276 15204 19332 15206
rect 19356 15204 19412 15206
rect 20074 17720 20130 17776
rect 19890 15544 19946 15600
rect 19116 14170 19172 14172
rect 19196 14170 19252 14172
rect 19276 14170 19332 14172
rect 19356 14170 19412 14172
rect 19116 14118 19142 14170
rect 19142 14118 19172 14170
rect 19196 14118 19206 14170
rect 19206 14118 19252 14170
rect 19276 14118 19322 14170
rect 19322 14118 19332 14170
rect 19356 14118 19386 14170
rect 19386 14118 19412 14170
rect 19116 14116 19172 14118
rect 19196 14116 19252 14118
rect 19276 14116 19332 14118
rect 19356 14116 19412 14118
rect 19338 13912 19394 13968
rect 19116 13082 19172 13084
rect 19196 13082 19252 13084
rect 19276 13082 19332 13084
rect 19356 13082 19412 13084
rect 19116 13030 19142 13082
rect 19142 13030 19172 13082
rect 19196 13030 19206 13082
rect 19206 13030 19252 13082
rect 19276 13030 19322 13082
rect 19322 13030 19332 13082
rect 19356 13030 19386 13082
rect 19386 13030 19412 13082
rect 19116 13028 19172 13030
rect 19196 13028 19252 13030
rect 19276 13028 19332 13030
rect 19356 13028 19412 13030
rect 18694 11228 18696 11248
rect 18696 11228 18748 11248
rect 18748 11228 18750 11248
rect 18694 11192 18750 11228
rect 19116 11994 19172 11996
rect 19196 11994 19252 11996
rect 19276 11994 19332 11996
rect 19356 11994 19412 11996
rect 19116 11942 19142 11994
rect 19142 11942 19172 11994
rect 19196 11942 19206 11994
rect 19206 11942 19252 11994
rect 19276 11942 19322 11994
rect 19322 11942 19332 11994
rect 19356 11942 19386 11994
rect 19386 11942 19412 11994
rect 19116 11940 19172 11942
rect 19196 11940 19252 11942
rect 19276 11940 19332 11942
rect 19356 11940 19412 11942
rect 19614 11872 19670 11928
rect 20994 20748 20996 20768
rect 20996 20748 21048 20768
rect 21048 20748 21050 20768
rect 20994 20712 21050 20748
rect 19116 10906 19172 10908
rect 19196 10906 19252 10908
rect 19276 10906 19332 10908
rect 19356 10906 19412 10908
rect 19116 10854 19142 10906
rect 19142 10854 19172 10906
rect 19196 10854 19206 10906
rect 19206 10854 19252 10906
rect 19276 10854 19322 10906
rect 19322 10854 19332 10906
rect 19356 10854 19386 10906
rect 19386 10854 19412 10906
rect 19116 10852 19172 10854
rect 19196 10852 19252 10854
rect 19276 10852 19332 10854
rect 19356 10852 19412 10854
rect 18878 10260 18934 10296
rect 18878 10240 18880 10260
rect 18880 10240 18932 10260
rect 18932 10240 18934 10260
rect 19338 10376 19394 10432
rect 19154 10260 19210 10296
rect 19154 10240 19156 10260
rect 19156 10240 19208 10260
rect 19208 10240 19210 10260
rect 19116 9818 19172 9820
rect 19196 9818 19252 9820
rect 19276 9818 19332 9820
rect 19356 9818 19412 9820
rect 19116 9766 19142 9818
rect 19142 9766 19172 9818
rect 19196 9766 19206 9818
rect 19206 9766 19252 9818
rect 19276 9766 19322 9818
rect 19322 9766 19332 9818
rect 19356 9766 19386 9818
rect 19386 9766 19412 9818
rect 19116 9764 19172 9766
rect 19196 9764 19252 9766
rect 19276 9764 19332 9766
rect 19356 9764 19412 9766
rect 19522 9968 19578 10024
rect 19522 9696 19578 9752
rect 18786 9560 18842 9616
rect 19338 9580 19394 9582
rect 18326 8744 18382 8800
rect 18694 9424 18750 9480
rect 18050 7384 18106 7440
rect 17314 6296 17370 6352
rect 17130 6160 17186 6216
rect 17590 5344 17646 5400
rect 16302 3168 16358 3224
rect 18418 7928 18474 7984
rect 19338 9528 19340 9580
rect 19340 9528 19392 9580
rect 19392 9528 19394 9580
rect 19338 9526 19394 9528
rect 19154 9460 19156 9480
rect 19156 9460 19208 9480
rect 19208 9460 19210 9480
rect 19154 9424 19210 9460
rect 20258 16224 20314 16280
rect 20074 10104 20130 10160
rect 19116 8730 19172 8732
rect 19196 8730 19252 8732
rect 19276 8730 19332 8732
rect 19356 8730 19412 8732
rect 19116 8678 19142 8730
rect 19142 8678 19172 8730
rect 19196 8678 19206 8730
rect 19206 8678 19252 8730
rect 19276 8678 19322 8730
rect 19322 8678 19332 8730
rect 19356 8678 19386 8730
rect 19386 8678 19412 8730
rect 19116 8676 19172 8678
rect 19196 8676 19252 8678
rect 19276 8676 19332 8678
rect 19356 8676 19412 8678
rect 19706 8200 19762 8256
rect 19522 7792 19578 7848
rect 19116 7642 19172 7644
rect 19196 7642 19252 7644
rect 19276 7642 19332 7644
rect 19356 7642 19412 7644
rect 19116 7590 19142 7642
rect 19142 7590 19172 7642
rect 19196 7590 19206 7642
rect 19206 7590 19252 7642
rect 19276 7590 19322 7642
rect 19322 7590 19332 7642
rect 19356 7590 19386 7642
rect 19386 7590 19412 7642
rect 19116 7588 19172 7590
rect 19196 7588 19252 7590
rect 19276 7588 19332 7590
rect 19356 7588 19412 7590
rect 18694 6024 18750 6080
rect 18602 4664 18658 4720
rect 19116 6554 19172 6556
rect 19196 6554 19252 6556
rect 19276 6554 19332 6556
rect 19356 6554 19412 6556
rect 19116 6502 19142 6554
rect 19142 6502 19172 6554
rect 19196 6502 19206 6554
rect 19206 6502 19252 6554
rect 19276 6502 19322 6554
rect 19322 6502 19332 6554
rect 19356 6502 19386 6554
rect 19386 6502 19412 6554
rect 19116 6500 19172 6502
rect 19196 6500 19252 6502
rect 19276 6500 19332 6502
rect 19356 6500 19412 6502
rect 19116 5466 19172 5468
rect 19196 5466 19252 5468
rect 19276 5466 19332 5468
rect 19356 5466 19412 5468
rect 19116 5414 19142 5466
rect 19142 5414 19172 5466
rect 19196 5414 19206 5466
rect 19206 5414 19252 5466
rect 19276 5414 19322 5466
rect 19322 5414 19332 5466
rect 19356 5414 19386 5466
rect 19386 5414 19412 5466
rect 19116 5412 19172 5414
rect 19196 5412 19252 5414
rect 19276 5412 19332 5414
rect 19356 5412 19412 5414
rect 20166 9424 20222 9480
rect 19798 6296 19854 6352
rect 19890 5344 19946 5400
rect 20626 6840 20682 6896
rect 19116 4378 19172 4380
rect 19196 4378 19252 4380
rect 19276 4378 19332 4380
rect 19356 4378 19412 4380
rect 19116 4326 19142 4378
rect 19142 4326 19172 4378
rect 19196 4326 19206 4378
rect 19206 4326 19252 4378
rect 19276 4326 19322 4378
rect 19322 4326 19332 4378
rect 19356 4326 19386 4378
rect 19386 4326 19412 4378
rect 19116 4324 19172 4326
rect 19196 4324 19252 4326
rect 19276 4324 19332 4326
rect 19356 4324 19412 4326
rect 19116 3290 19172 3292
rect 19196 3290 19252 3292
rect 19276 3290 19332 3292
rect 19356 3290 19412 3292
rect 19116 3238 19142 3290
rect 19142 3238 19172 3290
rect 19196 3238 19206 3290
rect 19206 3238 19252 3290
rect 19276 3238 19322 3290
rect 19322 3238 19332 3290
rect 19356 3238 19386 3290
rect 19386 3238 19412 3290
rect 19116 3236 19172 3238
rect 19196 3236 19252 3238
rect 19276 3236 19332 3238
rect 19356 3236 19412 3238
rect 19890 3848 19946 3904
rect 18878 2488 18934 2544
rect 19116 2202 19172 2204
rect 19196 2202 19252 2204
rect 19276 2202 19332 2204
rect 19356 2202 19412 2204
rect 19116 2150 19142 2202
rect 19142 2150 19172 2202
rect 19196 2150 19206 2202
rect 19206 2150 19252 2202
rect 19276 2150 19322 2202
rect 19322 2150 19332 2202
rect 19356 2150 19386 2202
rect 19386 2150 19412 2202
rect 19116 2148 19172 2150
rect 19196 2148 19252 2150
rect 19276 2148 19332 2150
rect 19356 2148 19412 2150
rect 20350 3168 20406 3224
rect 20534 992 20590 1048
rect 21546 20440 21602 20496
rect 22098 19896 22154 19952
rect 22098 19080 22154 19136
rect 21914 16904 21970 16960
rect 21730 9016 21786 9072
rect 22006 9016 22062 9072
rect 21270 8336 21326 8392
rect 20994 7384 21050 7440
rect 21914 7520 21970 7576
rect 22834 20304 22890 20360
rect 23386 11192 23442 11248
rect 23386 11056 23442 11112
rect 22098 8472 22154 8528
rect 22282 6024 22338 6080
rect 20626 312 20682 368
<< metal3 >>
rect 19425 23490 19491 23493
rect 23520 23490 24000 23520
rect 19425 23488 24000 23490
rect 19425 23432 19430 23488
rect 19486 23432 24000 23488
rect 19425 23430 24000 23432
rect 19425 23427 19491 23430
rect 23520 23400 24000 23430
rect 19609 22810 19675 22813
rect 23520 22810 24000 22840
rect 19609 22808 24000 22810
rect 19609 22752 19614 22808
rect 19670 22752 24000 22808
rect 19609 22750 24000 22752
rect 19609 22747 19675 22750
rect 23520 22720 24000 22750
rect 19333 22130 19399 22133
rect 23520 22130 24000 22160
rect 19333 22128 24000 22130
rect 19333 22072 19338 22128
rect 19394 22072 24000 22128
rect 19333 22070 24000 22072
rect 19333 22067 19399 22070
rect 23520 22040 24000 22070
rect 4576 21792 4896 21793
rect 4576 21728 4584 21792
rect 4648 21728 4664 21792
rect 4728 21728 4744 21792
rect 4808 21728 4824 21792
rect 4888 21728 4896 21792
rect 4576 21727 4896 21728
rect 11840 21792 12160 21793
rect 11840 21728 11848 21792
rect 11912 21728 11928 21792
rect 11992 21728 12008 21792
rect 12072 21728 12088 21792
rect 12152 21728 12160 21792
rect 11840 21727 12160 21728
rect 19104 21792 19424 21793
rect 19104 21728 19112 21792
rect 19176 21728 19192 21792
rect 19256 21728 19272 21792
rect 19336 21728 19352 21792
rect 19416 21728 19424 21792
rect 19104 21727 19424 21728
rect 1393 21450 1459 21453
rect 8661 21450 8727 21453
rect 1393 21448 8727 21450
rect 1393 21392 1398 21448
rect 1454 21392 8666 21448
rect 8722 21392 8727 21448
rect 1393 21390 8727 21392
rect 1393 21387 1459 21390
rect 8661 21387 8727 21390
rect 19977 21314 20043 21317
rect 23520 21314 24000 21344
rect 19977 21312 24000 21314
rect 19977 21256 19982 21312
rect 20038 21256 24000 21312
rect 19977 21254 24000 21256
rect 19977 21251 20043 21254
rect 8208 21248 8528 21249
rect 8208 21184 8216 21248
rect 8280 21184 8296 21248
rect 8360 21184 8376 21248
rect 8440 21184 8456 21248
rect 8520 21184 8528 21248
rect 8208 21183 8528 21184
rect 15472 21248 15792 21249
rect 15472 21184 15480 21248
rect 15544 21184 15560 21248
rect 15624 21184 15640 21248
rect 15704 21184 15720 21248
rect 15784 21184 15792 21248
rect 23520 21224 24000 21254
rect 15472 21183 15792 21184
rect 15193 20770 15259 20773
rect 16849 20770 16915 20773
rect 15193 20768 16915 20770
rect 15193 20712 15198 20768
rect 15254 20712 16854 20768
rect 16910 20712 16915 20768
rect 15193 20710 16915 20712
rect 15193 20707 15259 20710
rect 16849 20707 16915 20710
rect 20989 20772 21055 20773
rect 20989 20768 21036 20772
rect 21100 20770 21106 20772
rect 20989 20712 20994 20768
rect 20989 20708 21036 20712
rect 21100 20710 21146 20770
rect 21100 20708 21106 20710
rect 20989 20707 21055 20708
rect 4576 20704 4896 20705
rect 4576 20640 4584 20704
rect 4648 20640 4664 20704
rect 4728 20640 4744 20704
rect 4808 20640 4824 20704
rect 4888 20640 4896 20704
rect 4576 20639 4896 20640
rect 11840 20704 12160 20705
rect 11840 20640 11848 20704
rect 11912 20640 11928 20704
rect 11992 20640 12008 20704
rect 12072 20640 12088 20704
rect 12152 20640 12160 20704
rect 11840 20639 12160 20640
rect 19104 20704 19424 20705
rect 19104 20640 19112 20704
rect 19176 20640 19192 20704
rect 19256 20640 19272 20704
rect 19336 20640 19352 20704
rect 19416 20640 19424 20704
rect 19104 20639 19424 20640
rect 5533 20634 5599 20637
rect 6637 20634 6703 20637
rect 5533 20632 6703 20634
rect 5533 20576 5538 20632
rect 5594 20576 6642 20632
rect 6698 20576 6703 20632
rect 5533 20574 6703 20576
rect 5533 20571 5599 20574
rect 6637 20571 6703 20574
rect 12617 20634 12683 20637
rect 13721 20634 13787 20637
rect 17033 20634 17099 20637
rect 12617 20632 17099 20634
rect 12617 20576 12622 20632
rect 12678 20576 13726 20632
rect 13782 20576 17038 20632
rect 17094 20576 17099 20632
rect 12617 20574 17099 20576
rect 12617 20571 12683 20574
rect 13721 20571 13787 20574
rect 17033 20571 17099 20574
rect 19517 20634 19583 20637
rect 23520 20634 24000 20664
rect 19517 20632 24000 20634
rect 19517 20576 19522 20632
rect 19578 20576 24000 20632
rect 19517 20574 24000 20576
rect 19517 20571 19583 20574
rect 23520 20544 24000 20574
rect 10961 20498 11027 20501
rect 14457 20498 14523 20501
rect 10961 20496 14523 20498
rect 10961 20440 10966 20496
rect 11022 20440 14462 20496
rect 14518 20440 14523 20496
rect 10961 20438 14523 20440
rect 10961 20435 11027 20438
rect 14457 20435 14523 20438
rect 14641 20498 14707 20501
rect 21541 20498 21607 20501
rect 14641 20496 21607 20498
rect 14641 20440 14646 20496
rect 14702 20440 21546 20496
rect 21602 20440 21607 20496
rect 14641 20438 21607 20440
rect 14641 20435 14707 20438
rect 21541 20435 21607 20438
rect 15009 20362 15075 20365
rect 16849 20362 16915 20365
rect 15009 20360 16915 20362
rect 15009 20304 15014 20360
rect 15070 20304 16854 20360
rect 16910 20304 16915 20360
rect 15009 20302 16915 20304
rect 15009 20299 15075 20302
rect 16849 20299 16915 20302
rect 17033 20362 17099 20365
rect 22829 20362 22895 20365
rect 17033 20360 22895 20362
rect 17033 20304 17038 20360
rect 17094 20304 22834 20360
rect 22890 20304 22895 20360
rect 17033 20302 22895 20304
rect 17033 20299 17099 20302
rect 22829 20299 22895 20302
rect 8208 20160 8528 20161
rect 8208 20096 8216 20160
rect 8280 20096 8296 20160
rect 8360 20096 8376 20160
rect 8440 20096 8456 20160
rect 8520 20096 8528 20160
rect 8208 20095 8528 20096
rect 15472 20160 15792 20161
rect 15472 20096 15480 20160
rect 15544 20096 15560 20160
rect 15624 20096 15640 20160
rect 15704 20096 15720 20160
rect 15784 20096 15792 20160
rect 15472 20095 15792 20096
rect 10317 20090 10383 20093
rect 13077 20090 13143 20093
rect 10317 20088 13143 20090
rect 10317 20032 10322 20088
rect 10378 20032 13082 20088
rect 13138 20032 13143 20088
rect 10317 20030 13143 20032
rect 10317 20027 10383 20030
rect 13077 20027 13143 20030
rect 0 19954 480 19984
rect 2773 19954 2839 19957
rect 0 19952 2839 19954
rect 0 19896 2778 19952
rect 2834 19896 2839 19952
rect 0 19894 2839 19896
rect 0 19864 480 19894
rect 2773 19891 2839 19894
rect 6637 19954 6703 19957
rect 19609 19954 19675 19957
rect 6637 19952 19675 19954
rect 6637 19896 6642 19952
rect 6698 19896 19614 19952
rect 19670 19896 19675 19952
rect 6637 19894 19675 19896
rect 6637 19891 6703 19894
rect 19609 19891 19675 19894
rect 22093 19954 22159 19957
rect 23520 19954 24000 19984
rect 22093 19952 24000 19954
rect 22093 19896 22098 19952
rect 22154 19896 24000 19952
rect 22093 19894 24000 19896
rect 22093 19891 22159 19894
rect 23520 19864 24000 19894
rect 4061 19818 4127 19821
rect 4613 19818 4679 19821
rect 4061 19816 4679 19818
rect 4061 19760 4066 19816
rect 4122 19760 4618 19816
rect 4674 19760 4679 19816
rect 4061 19758 4679 19760
rect 4061 19755 4127 19758
rect 4613 19755 4679 19758
rect 7097 19818 7163 19821
rect 9213 19818 9279 19821
rect 7097 19816 9279 19818
rect 7097 19760 7102 19816
rect 7158 19760 9218 19816
rect 9274 19760 9279 19816
rect 7097 19758 9279 19760
rect 7097 19755 7163 19758
rect 9213 19755 9279 19758
rect 12065 19818 12131 19821
rect 12525 19818 12591 19821
rect 12065 19816 12591 19818
rect 12065 19760 12070 19816
rect 12126 19760 12530 19816
rect 12586 19760 12591 19816
rect 12065 19758 12591 19760
rect 12065 19755 12131 19758
rect 12525 19755 12591 19758
rect 8845 19682 8911 19685
rect 4984 19680 8911 19682
rect 4984 19624 8850 19680
rect 8906 19624 8911 19680
rect 4984 19622 8911 19624
rect 4576 19616 4896 19617
rect 4576 19552 4584 19616
rect 4648 19552 4664 19616
rect 4728 19552 4744 19616
rect 4808 19552 4824 19616
rect 4888 19552 4896 19616
rect 4576 19551 4896 19552
rect 4984 19549 5044 19622
rect 8845 19619 8911 19622
rect 12525 19682 12591 19685
rect 13353 19682 13419 19685
rect 12525 19680 13419 19682
rect 12525 19624 12530 19680
rect 12586 19624 13358 19680
rect 13414 19624 13419 19680
rect 12525 19622 13419 19624
rect 12525 19619 12591 19622
rect 13353 19619 13419 19622
rect 11840 19616 12160 19617
rect 11840 19552 11848 19616
rect 11912 19552 11928 19616
rect 11992 19552 12008 19616
rect 12072 19552 12088 19616
rect 12152 19552 12160 19616
rect 11840 19551 12160 19552
rect 19104 19616 19424 19617
rect 19104 19552 19112 19616
rect 19176 19552 19192 19616
rect 19256 19552 19272 19616
rect 19336 19552 19352 19616
rect 19416 19552 19424 19616
rect 19104 19551 19424 19552
rect 4981 19544 5047 19549
rect 4981 19488 4986 19544
rect 5042 19488 5047 19544
rect 4981 19483 5047 19488
rect 13169 19546 13235 19549
rect 15193 19546 15259 19549
rect 13169 19544 15259 19546
rect 13169 19488 13174 19544
rect 13230 19488 15198 19544
rect 15254 19488 15259 19544
rect 13169 19486 15259 19488
rect 13169 19483 13235 19486
rect 15193 19483 15259 19486
rect 6729 19410 6795 19413
rect 8201 19410 8267 19413
rect 10593 19410 10659 19413
rect 11329 19410 11395 19413
rect 12617 19410 12683 19413
rect 6729 19408 11395 19410
rect 6729 19352 6734 19408
rect 6790 19352 8206 19408
rect 8262 19352 10598 19408
rect 10654 19352 11334 19408
rect 11390 19352 11395 19408
rect 6729 19350 11395 19352
rect 6729 19347 6795 19350
rect 8201 19347 8267 19350
rect 10593 19347 10659 19350
rect 11329 19347 11395 19350
rect 12022 19408 12683 19410
rect 12022 19352 12622 19408
rect 12678 19352 12683 19408
rect 12022 19350 12683 19352
rect 4521 19274 4587 19277
rect 6729 19274 6795 19277
rect 4521 19272 6795 19274
rect 4521 19216 4526 19272
rect 4582 19216 6734 19272
rect 6790 19216 6795 19272
rect 4521 19214 6795 19216
rect 4521 19211 4587 19214
rect 6729 19211 6795 19214
rect 9305 19274 9371 19277
rect 12022 19274 12082 19350
rect 12617 19347 12683 19350
rect 9305 19272 12082 19274
rect 9305 19216 9310 19272
rect 9366 19216 12082 19272
rect 9305 19214 12082 19216
rect 12249 19274 12315 19277
rect 12525 19274 12591 19277
rect 15653 19274 15719 19277
rect 12249 19272 12591 19274
rect 12249 19216 12254 19272
rect 12310 19216 12530 19272
rect 12586 19216 12591 19272
rect 12249 19214 12591 19216
rect 9305 19211 9371 19214
rect 12249 19211 12315 19214
rect 12525 19211 12591 19214
rect 12712 19272 15719 19274
rect 12712 19216 15658 19272
rect 15714 19216 15719 19272
rect 12712 19214 15719 19216
rect 4102 19076 4108 19140
rect 4172 19138 4178 19140
rect 5349 19138 5415 19141
rect 4172 19136 5415 19138
rect 4172 19080 5354 19136
rect 5410 19080 5415 19136
rect 4172 19078 5415 19080
rect 4172 19076 4178 19078
rect 5349 19075 5415 19078
rect 9581 19138 9647 19141
rect 11053 19138 11119 19141
rect 9581 19136 11119 19138
rect 9581 19080 9586 19136
rect 9642 19080 11058 19136
rect 11114 19080 11119 19136
rect 9581 19078 11119 19080
rect 9581 19075 9647 19078
rect 11053 19075 11119 19078
rect 8208 19072 8528 19073
rect 8208 19008 8216 19072
rect 8280 19008 8296 19072
rect 8360 19008 8376 19072
rect 8440 19008 8456 19072
rect 8520 19008 8528 19072
rect 8208 19007 8528 19008
rect 10225 19002 10291 19005
rect 12712 19002 12772 19214
rect 15653 19211 15719 19214
rect 22093 19138 22159 19141
rect 23520 19138 24000 19168
rect 22093 19136 24000 19138
rect 22093 19080 22098 19136
rect 22154 19080 24000 19136
rect 22093 19078 24000 19080
rect 22093 19075 22159 19078
rect 15472 19072 15792 19073
rect 15472 19008 15480 19072
rect 15544 19008 15560 19072
rect 15624 19008 15640 19072
rect 15704 19008 15720 19072
rect 15784 19008 15792 19072
rect 23520 19048 24000 19078
rect 15472 19007 15792 19008
rect 10225 19000 12772 19002
rect 10225 18944 10230 19000
rect 10286 18944 12772 19000
rect 10225 18942 12772 18944
rect 10225 18939 10291 18942
rect 12157 18866 12223 18869
rect 16849 18866 16915 18869
rect 12157 18864 16915 18866
rect 12157 18808 12162 18864
rect 12218 18808 16854 18864
rect 16910 18808 16915 18864
rect 12157 18806 16915 18808
rect 12157 18803 12223 18806
rect 16849 18803 16915 18806
rect 1577 18730 1643 18733
rect 6637 18730 6703 18733
rect 1577 18728 6703 18730
rect 1577 18672 1582 18728
rect 1638 18672 6642 18728
rect 6698 18672 6703 18728
rect 1577 18670 6703 18672
rect 1577 18667 1643 18670
rect 6637 18667 6703 18670
rect 18413 18730 18479 18733
rect 19149 18730 19215 18733
rect 18413 18728 19215 18730
rect 18413 18672 18418 18728
rect 18474 18672 19154 18728
rect 19210 18672 19215 18728
rect 18413 18670 19215 18672
rect 18413 18667 18479 18670
rect 19149 18667 19215 18670
rect 4576 18528 4896 18529
rect 4576 18464 4584 18528
rect 4648 18464 4664 18528
rect 4728 18464 4744 18528
rect 4808 18464 4824 18528
rect 4888 18464 4896 18528
rect 4576 18463 4896 18464
rect 11840 18528 12160 18529
rect 11840 18464 11848 18528
rect 11912 18464 11928 18528
rect 11992 18464 12008 18528
rect 12072 18464 12088 18528
rect 12152 18464 12160 18528
rect 11840 18463 12160 18464
rect 19104 18528 19424 18529
rect 19104 18464 19112 18528
rect 19176 18464 19192 18528
rect 19256 18464 19272 18528
rect 19336 18464 19352 18528
rect 19416 18464 19424 18528
rect 19104 18463 19424 18464
rect 12249 18458 12315 18461
rect 14273 18458 14339 18461
rect 12249 18456 14339 18458
rect 12249 18400 12254 18456
rect 12310 18400 14278 18456
rect 14334 18400 14339 18456
rect 12249 18398 14339 18400
rect 12249 18395 12315 18398
rect 14273 18395 14339 18398
rect 19609 18458 19675 18461
rect 23520 18458 24000 18488
rect 19609 18456 24000 18458
rect 19609 18400 19614 18456
rect 19670 18400 24000 18456
rect 19609 18398 24000 18400
rect 19609 18395 19675 18398
rect 23520 18368 24000 18398
rect 12566 18260 12572 18324
rect 12636 18322 12642 18324
rect 16113 18322 16179 18325
rect 12636 18320 16179 18322
rect 12636 18264 16118 18320
rect 16174 18264 16179 18320
rect 12636 18262 16179 18264
rect 12636 18260 12642 18262
rect 16113 18259 16179 18262
rect 1761 18186 1827 18189
rect 16665 18186 16731 18189
rect 1761 18184 16731 18186
rect 1761 18128 1766 18184
rect 1822 18128 16670 18184
rect 16726 18128 16731 18184
rect 1761 18126 16731 18128
rect 1761 18123 1827 18126
rect 16665 18123 16731 18126
rect 9857 18050 9923 18053
rect 15009 18050 15075 18053
rect 9857 18048 15075 18050
rect 9857 17992 9862 18048
rect 9918 17992 15014 18048
rect 15070 17992 15075 18048
rect 9857 17990 15075 17992
rect 9857 17987 9923 17990
rect 15009 17987 15075 17990
rect 8208 17984 8528 17985
rect 8208 17920 8216 17984
rect 8280 17920 8296 17984
rect 8360 17920 8376 17984
rect 8440 17920 8456 17984
rect 8520 17920 8528 17984
rect 8208 17919 8528 17920
rect 15472 17984 15792 17985
rect 15472 17920 15480 17984
rect 15544 17920 15560 17984
rect 15624 17920 15640 17984
rect 15704 17920 15720 17984
rect 15784 17920 15792 17984
rect 15472 17919 15792 17920
rect 3969 17914 4035 17917
rect 5533 17914 5599 17917
rect 3969 17912 5599 17914
rect 3969 17856 3974 17912
rect 4030 17856 5538 17912
rect 5594 17856 5599 17912
rect 3969 17854 5599 17856
rect 3969 17851 4035 17854
rect 5533 17851 5599 17854
rect 20069 17778 20135 17781
rect 23520 17778 24000 17808
rect 20069 17776 24000 17778
rect 20069 17720 20074 17776
rect 20130 17720 24000 17776
rect 20069 17718 24000 17720
rect 20069 17715 20135 17718
rect 23520 17688 24000 17718
rect 6453 17642 6519 17645
rect 7833 17642 7899 17645
rect 6453 17640 7899 17642
rect 6453 17584 6458 17640
rect 6514 17584 7838 17640
rect 7894 17584 7899 17640
rect 6453 17582 7899 17584
rect 6453 17579 6519 17582
rect 7833 17579 7899 17582
rect 12341 17642 12407 17645
rect 18965 17642 19031 17645
rect 12341 17640 19031 17642
rect 12341 17584 12346 17640
rect 12402 17584 18970 17640
rect 19026 17584 19031 17640
rect 12341 17582 19031 17584
rect 12341 17579 12407 17582
rect 18965 17579 19031 17582
rect 7189 17508 7255 17509
rect 7189 17506 7236 17508
rect 7144 17504 7236 17506
rect 7144 17448 7194 17504
rect 7144 17446 7236 17448
rect 7189 17444 7236 17446
rect 7300 17444 7306 17508
rect 7189 17443 7255 17444
rect 4576 17440 4896 17441
rect 4576 17376 4584 17440
rect 4648 17376 4664 17440
rect 4728 17376 4744 17440
rect 4808 17376 4824 17440
rect 4888 17376 4896 17440
rect 4576 17375 4896 17376
rect 11840 17440 12160 17441
rect 11840 17376 11848 17440
rect 11912 17376 11928 17440
rect 11992 17376 12008 17440
rect 12072 17376 12088 17440
rect 12152 17376 12160 17440
rect 11840 17375 12160 17376
rect 19104 17440 19424 17441
rect 19104 17376 19112 17440
rect 19176 17376 19192 17440
rect 19256 17376 19272 17440
rect 19336 17376 19352 17440
rect 19416 17376 19424 17440
rect 19104 17375 19424 17376
rect 12433 17370 12499 17373
rect 14825 17370 14891 17373
rect 12433 17368 14891 17370
rect 12433 17312 12438 17368
rect 12494 17312 14830 17368
rect 14886 17312 14891 17368
rect 12433 17310 14891 17312
rect 12433 17307 12499 17310
rect 14825 17307 14891 17310
rect 19558 17308 19564 17372
rect 19628 17370 19634 17372
rect 19701 17370 19767 17373
rect 19628 17368 19767 17370
rect 19628 17312 19706 17368
rect 19762 17312 19767 17368
rect 19628 17310 19767 17312
rect 19628 17308 19634 17310
rect 19701 17307 19767 17310
rect 4613 17234 4679 17237
rect 6545 17234 6611 17237
rect 4613 17232 6611 17234
rect 4613 17176 4618 17232
rect 4674 17176 6550 17232
rect 6606 17176 6611 17232
rect 4613 17174 6611 17176
rect 4613 17171 4679 17174
rect 6545 17171 6611 17174
rect 6453 17098 6519 17101
rect 9581 17098 9647 17101
rect 6453 17096 9647 17098
rect 6453 17040 6458 17096
rect 6514 17040 9586 17096
rect 9642 17040 9647 17096
rect 6453 17038 9647 17040
rect 6453 17035 6519 17038
rect 9581 17035 9647 17038
rect 21909 16962 21975 16965
rect 23520 16962 24000 16992
rect 21909 16960 24000 16962
rect 21909 16904 21914 16960
rect 21970 16904 24000 16960
rect 21909 16902 24000 16904
rect 21909 16899 21975 16902
rect 8208 16896 8528 16897
rect 8208 16832 8216 16896
rect 8280 16832 8296 16896
rect 8360 16832 8376 16896
rect 8440 16832 8456 16896
rect 8520 16832 8528 16896
rect 8208 16831 8528 16832
rect 15472 16896 15792 16897
rect 15472 16832 15480 16896
rect 15544 16832 15560 16896
rect 15624 16832 15640 16896
rect 15704 16832 15720 16896
rect 15784 16832 15792 16896
rect 23520 16872 24000 16902
rect 15472 16831 15792 16832
rect 6545 16690 6611 16693
rect 9581 16690 9647 16693
rect 6545 16688 9647 16690
rect 6545 16632 6550 16688
rect 6606 16632 9586 16688
rect 9642 16632 9647 16688
rect 6545 16630 9647 16632
rect 6545 16627 6611 16630
rect 9581 16627 9647 16630
rect 13445 16690 13511 16693
rect 15469 16690 15535 16693
rect 13445 16688 15535 16690
rect 13445 16632 13450 16688
rect 13506 16632 15474 16688
rect 15530 16632 15535 16688
rect 13445 16630 15535 16632
rect 13445 16627 13511 16630
rect 15469 16627 15535 16630
rect 12525 16554 12591 16557
rect 14641 16554 14707 16557
rect 12525 16552 14707 16554
rect 12525 16496 12530 16552
rect 12586 16496 14646 16552
rect 14702 16496 14707 16552
rect 12525 16494 14707 16496
rect 12525 16491 12591 16494
rect 14641 16491 14707 16494
rect 6545 16418 6611 16421
rect 9029 16418 9095 16421
rect 6545 16416 9095 16418
rect 6545 16360 6550 16416
rect 6606 16360 9034 16416
rect 9090 16360 9095 16416
rect 6545 16358 9095 16360
rect 6545 16355 6611 16358
rect 9029 16355 9095 16358
rect 4576 16352 4896 16353
rect 4576 16288 4584 16352
rect 4648 16288 4664 16352
rect 4728 16288 4744 16352
rect 4808 16288 4824 16352
rect 4888 16288 4896 16352
rect 4576 16287 4896 16288
rect 11840 16352 12160 16353
rect 11840 16288 11848 16352
rect 11912 16288 11928 16352
rect 11992 16288 12008 16352
rect 12072 16288 12088 16352
rect 12152 16288 12160 16352
rect 11840 16287 12160 16288
rect 19104 16352 19424 16353
rect 19104 16288 19112 16352
rect 19176 16288 19192 16352
rect 19256 16288 19272 16352
rect 19336 16288 19352 16352
rect 19416 16288 19424 16352
rect 19104 16287 19424 16288
rect 12249 16282 12315 16285
rect 14273 16282 14339 16285
rect 15878 16282 15884 16284
rect 12249 16280 15884 16282
rect 12249 16224 12254 16280
rect 12310 16224 14278 16280
rect 14334 16224 15884 16280
rect 12249 16222 15884 16224
rect 12249 16219 12315 16222
rect 14273 16219 14339 16222
rect 15878 16220 15884 16222
rect 15948 16282 15954 16284
rect 16389 16282 16455 16285
rect 15948 16280 16455 16282
rect 15948 16224 16394 16280
rect 16450 16224 16455 16280
rect 15948 16222 16455 16224
rect 15948 16220 15954 16222
rect 16389 16219 16455 16222
rect 20253 16282 20319 16285
rect 23520 16282 24000 16312
rect 20253 16280 24000 16282
rect 20253 16224 20258 16280
rect 20314 16224 24000 16280
rect 20253 16222 24000 16224
rect 20253 16219 20319 16222
rect 23520 16192 24000 16222
rect 14089 16146 14155 16149
rect 15009 16146 15075 16149
rect 14089 16144 15075 16146
rect 14089 16088 14094 16144
rect 14150 16088 15014 16144
rect 15070 16088 15075 16144
rect 14089 16086 15075 16088
rect 14089 16083 14155 16086
rect 15009 16083 15075 16086
rect 13353 16010 13419 16013
rect 15009 16010 15075 16013
rect 13353 16008 15075 16010
rect 13353 15952 13358 16008
rect 13414 15952 15014 16008
rect 15070 15952 15075 16008
rect 13353 15950 15075 15952
rect 13353 15947 13419 15950
rect 15009 15947 15075 15950
rect 8208 15808 8528 15809
rect 8208 15744 8216 15808
rect 8280 15744 8296 15808
rect 8360 15744 8376 15808
rect 8440 15744 8456 15808
rect 8520 15744 8528 15808
rect 8208 15743 8528 15744
rect 15472 15808 15792 15809
rect 15472 15744 15480 15808
rect 15544 15744 15560 15808
rect 15624 15744 15640 15808
rect 15704 15744 15720 15808
rect 15784 15744 15792 15808
rect 15472 15743 15792 15744
rect 19885 15602 19951 15605
rect 23520 15602 24000 15632
rect 19885 15600 24000 15602
rect 19885 15544 19890 15600
rect 19946 15544 24000 15600
rect 19885 15542 24000 15544
rect 19885 15539 19951 15542
rect 23520 15512 24000 15542
rect 4576 15264 4896 15265
rect 4576 15200 4584 15264
rect 4648 15200 4664 15264
rect 4728 15200 4744 15264
rect 4808 15200 4824 15264
rect 4888 15200 4896 15264
rect 4576 15199 4896 15200
rect 11840 15264 12160 15265
rect 11840 15200 11848 15264
rect 11912 15200 11928 15264
rect 11992 15200 12008 15264
rect 12072 15200 12088 15264
rect 12152 15200 12160 15264
rect 11840 15199 12160 15200
rect 19104 15264 19424 15265
rect 19104 15200 19112 15264
rect 19176 15200 19192 15264
rect 19256 15200 19272 15264
rect 19336 15200 19352 15264
rect 19416 15200 19424 15264
rect 19104 15199 19424 15200
rect 15745 15058 15811 15061
rect 17309 15058 17375 15061
rect 15745 15056 17375 15058
rect 15745 15000 15750 15056
rect 15806 15000 17314 15056
rect 17370 15000 17375 15056
rect 15745 14998 17375 15000
rect 15745 14995 15811 14998
rect 17309 14995 17375 14998
rect 17125 14786 17191 14789
rect 23520 14786 24000 14816
rect 17125 14784 24000 14786
rect 17125 14728 17130 14784
rect 17186 14728 24000 14784
rect 17125 14726 24000 14728
rect 17125 14723 17191 14726
rect 8208 14720 8528 14721
rect 8208 14656 8216 14720
rect 8280 14656 8296 14720
rect 8360 14656 8376 14720
rect 8440 14656 8456 14720
rect 8520 14656 8528 14720
rect 8208 14655 8528 14656
rect 15472 14720 15792 14721
rect 15472 14656 15480 14720
rect 15544 14656 15560 14720
rect 15624 14656 15640 14720
rect 15704 14656 15720 14720
rect 15784 14656 15792 14720
rect 23520 14696 24000 14726
rect 15472 14655 15792 14656
rect 16113 14650 16179 14653
rect 16070 14648 16179 14650
rect 16070 14592 16118 14648
rect 16174 14592 16179 14648
rect 16070 14587 16179 14592
rect 2773 14514 2839 14517
rect 4061 14514 4127 14517
rect 2773 14512 4127 14514
rect 2773 14456 2778 14512
rect 2834 14456 4066 14512
rect 4122 14456 4127 14512
rect 2773 14454 4127 14456
rect 2773 14451 2839 14454
rect 4061 14451 4127 14454
rect 11462 14452 11468 14516
rect 11532 14514 11538 14516
rect 16070 14514 16130 14587
rect 11532 14454 16130 14514
rect 11532 14452 11538 14454
rect 16113 14242 16179 14245
rect 17953 14242 18019 14245
rect 16113 14240 18019 14242
rect 16113 14184 16118 14240
rect 16174 14184 17958 14240
rect 18014 14184 18019 14240
rect 16113 14182 18019 14184
rect 16113 14179 16179 14182
rect 17953 14179 18019 14182
rect 4576 14176 4896 14177
rect 4576 14112 4584 14176
rect 4648 14112 4664 14176
rect 4728 14112 4744 14176
rect 4808 14112 4824 14176
rect 4888 14112 4896 14176
rect 4576 14111 4896 14112
rect 11840 14176 12160 14177
rect 11840 14112 11848 14176
rect 11912 14112 11928 14176
rect 11992 14112 12008 14176
rect 12072 14112 12088 14176
rect 12152 14112 12160 14176
rect 11840 14111 12160 14112
rect 19104 14176 19424 14177
rect 19104 14112 19112 14176
rect 19176 14112 19192 14176
rect 19256 14112 19272 14176
rect 19336 14112 19352 14176
rect 19416 14112 19424 14176
rect 19104 14111 19424 14112
rect 3693 14106 3759 14109
rect 4153 14106 4219 14109
rect 23520 14106 24000 14136
rect 3693 14104 4219 14106
rect 3693 14048 3698 14104
rect 3754 14048 4158 14104
rect 4214 14048 4219 14104
rect 3693 14046 4219 14048
rect 3693 14043 3759 14046
rect 4153 14043 4219 14046
rect 19612 14046 24000 14106
rect 1669 13834 1735 13837
rect 3233 13834 3299 13837
rect 3696 13834 3756 14043
rect 19333 13970 19399 13973
rect 19612 13970 19672 14046
rect 23520 14016 24000 14046
rect 19333 13968 19672 13970
rect 19333 13912 19338 13968
rect 19394 13912 19672 13968
rect 19333 13910 19672 13912
rect 19333 13907 19399 13910
rect 1669 13832 3756 13834
rect 1669 13776 1674 13832
rect 1730 13776 3238 13832
rect 3294 13776 3756 13832
rect 1669 13774 3756 13776
rect 1669 13771 1735 13774
rect 3233 13771 3299 13774
rect 8208 13632 8528 13633
rect 8208 13568 8216 13632
rect 8280 13568 8296 13632
rect 8360 13568 8376 13632
rect 8440 13568 8456 13632
rect 8520 13568 8528 13632
rect 8208 13567 8528 13568
rect 15472 13632 15792 13633
rect 15472 13568 15480 13632
rect 15544 13568 15560 13632
rect 15624 13568 15640 13632
rect 15704 13568 15720 13632
rect 15784 13568 15792 13632
rect 15472 13567 15792 13568
rect 4521 13562 4587 13565
rect 8017 13562 8083 13565
rect 4521 13560 8083 13562
rect 4521 13504 4526 13560
rect 4582 13504 8022 13560
rect 8078 13504 8083 13560
rect 4521 13502 8083 13504
rect 4521 13499 4587 13502
rect 8017 13499 8083 13502
rect 18137 13426 18203 13429
rect 23520 13426 24000 13456
rect 18137 13424 24000 13426
rect 18137 13368 18142 13424
rect 18198 13368 24000 13424
rect 18137 13366 24000 13368
rect 18137 13363 18203 13366
rect 23520 13336 24000 13366
rect 14774 13092 14780 13156
rect 14844 13154 14850 13156
rect 16389 13154 16455 13157
rect 14844 13152 16455 13154
rect 14844 13096 16394 13152
rect 16450 13096 16455 13152
rect 14844 13094 16455 13096
rect 14844 13092 14850 13094
rect 16389 13091 16455 13094
rect 4576 13088 4896 13089
rect 4576 13024 4584 13088
rect 4648 13024 4664 13088
rect 4728 13024 4744 13088
rect 4808 13024 4824 13088
rect 4888 13024 4896 13088
rect 4576 13023 4896 13024
rect 11840 13088 12160 13089
rect 11840 13024 11848 13088
rect 11912 13024 11928 13088
rect 11992 13024 12008 13088
rect 12072 13024 12088 13088
rect 12152 13024 12160 13088
rect 11840 13023 12160 13024
rect 19104 13088 19424 13089
rect 19104 13024 19112 13088
rect 19176 13024 19192 13088
rect 19256 13024 19272 13088
rect 19336 13024 19352 13088
rect 19416 13024 19424 13088
rect 19104 13023 19424 13024
rect 14958 12956 14964 13020
rect 15028 13018 15034 13020
rect 16021 13018 16087 13021
rect 15028 13016 16087 13018
rect 15028 12960 16026 13016
rect 16082 12960 16087 13016
rect 15028 12958 16087 12960
rect 15028 12956 15034 12958
rect 16021 12955 16087 12958
rect 15142 12820 15148 12884
rect 15212 12882 15218 12884
rect 15837 12882 15903 12885
rect 15212 12880 15903 12882
rect 15212 12824 15842 12880
rect 15898 12824 15903 12880
rect 15212 12822 15903 12824
rect 15212 12820 15218 12822
rect 15837 12819 15903 12822
rect 15377 12748 15443 12749
rect 9254 12684 9260 12748
rect 9324 12746 9330 12748
rect 12566 12746 12572 12748
rect 9324 12686 12572 12746
rect 9324 12684 9330 12686
rect 12566 12684 12572 12686
rect 12636 12684 12642 12748
rect 15326 12684 15332 12748
rect 15396 12746 15443 12748
rect 15396 12744 15488 12746
rect 15438 12688 15488 12744
rect 15396 12686 15488 12688
rect 15396 12684 15443 12686
rect 15377 12683 15443 12684
rect 23520 12610 24000 12640
rect 16990 12550 24000 12610
rect 8208 12544 8528 12545
rect 8208 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8528 12544
rect 8208 12479 8528 12480
rect 15472 12544 15792 12545
rect 15472 12480 15480 12544
rect 15544 12480 15560 12544
rect 15624 12480 15640 12544
rect 15704 12480 15720 12544
rect 15784 12480 15792 12544
rect 15472 12479 15792 12480
rect 10685 12474 10751 12477
rect 14825 12474 14891 12477
rect 10685 12472 14891 12474
rect 10685 12416 10690 12472
rect 10746 12416 14830 12472
rect 14886 12416 14891 12472
rect 10685 12414 14891 12416
rect 10685 12411 10751 12414
rect 14825 12411 14891 12414
rect 3049 12338 3115 12341
rect 6177 12338 6243 12341
rect 7557 12338 7623 12341
rect 3049 12336 7623 12338
rect 3049 12280 3054 12336
rect 3110 12280 6182 12336
rect 6238 12280 7562 12336
rect 7618 12280 7623 12336
rect 3049 12278 7623 12280
rect 3049 12275 3115 12278
rect 6177 12275 6243 12278
rect 7557 12275 7623 12278
rect 3601 12202 3667 12205
rect 10225 12202 10291 12205
rect 3601 12200 10291 12202
rect 3601 12144 3606 12200
rect 3662 12144 10230 12200
rect 10286 12144 10291 12200
rect 3601 12142 10291 12144
rect 3601 12139 3667 12142
rect 10225 12139 10291 12142
rect 11513 12202 11579 12205
rect 13721 12202 13787 12205
rect 11513 12200 13787 12202
rect 11513 12144 11518 12200
rect 11574 12144 13726 12200
rect 13782 12144 13787 12200
rect 11513 12142 13787 12144
rect 11513 12139 11579 12142
rect 13721 12139 13787 12142
rect 15101 12066 15167 12069
rect 16990 12066 17050 12550
rect 23520 12520 24000 12550
rect 15101 12064 17050 12066
rect 15101 12008 15106 12064
rect 15162 12008 17050 12064
rect 15101 12006 17050 12008
rect 15101 12003 15167 12006
rect 4576 12000 4896 12001
rect 0 11930 480 11960
rect 4576 11936 4584 12000
rect 4648 11936 4664 12000
rect 4728 11936 4744 12000
rect 4808 11936 4824 12000
rect 4888 11936 4896 12000
rect 4576 11935 4896 11936
rect 11840 12000 12160 12001
rect 11840 11936 11848 12000
rect 11912 11936 11928 12000
rect 11992 11936 12008 12000
rect 12072 11936 12088 12000
rect 12152 11936 12160 12000
rect 11840 11935 12160 11936
rect 19104 12000 19424 12001
rect 19104 11936 19112 12000
rect 19176 11936 19192 12000
rect 19256 11936 19272 12000
rect 19336 11936 19352 12000
rect 19416 11936 19424 12000
rect 19104 11935 19424 11936
rect 1485 11930 1551 11933
rect 0 11928 1551 11930
rect 0 11872 1490 11928
rect 1546 11872 1551 11928
rect 0 11870 1551 11872
rect 0 11840 480 11870
rect 1485 11867 1551 11870
rect 8702 11868 8708 11932
rect 8772 11930 8778 11932
rect 9489 11930 9555 11933
rect 8772 11928 9555 11930
rect 8772 11872 9494 11928
rect 9550 11872 9555 11928
rect 8772 11870 9555 11872
rect 8772 11868 8778 11870
rect 9489 11867 9555 11870
rect 15745 11930 15811 11933
rect 18321 11930 18387 11933
rect 15745 11928 18387 11930
rect 15745 11872 15750 11928
rect 15806 11872 18326 11928
rect 18382 11872 18387 11928
rect 15745 11870 18387 11872
rect 15745 11867 15811 11870
rect 18321 11867 18387 11870
rect 19609 11930 19675 11933
rect 23520 11930 24000 11960
rect 19609 11928 24000 11930
rect 19609 11872 19614 11928
rect 19670 11872 24000 11928
rect 19609 11870 24000 11872
rect 19609 11867 19675 11870
rect 23520 11840 24000 11870
rect 4061 11796 4127 11797
rect 4061 11794 4108 11796
rect 4016 11792 4108 11794
rect 4016 11736 4066 11792
rect 4016 11734 4108 11736
rect 4061 11732 4108 11734
rect 4172 11732 4178 11796
rect 8109 11794 8175 11797
rect 13997 11794 14063 11797
rect 8109 11792 14063 11794
rect 8109 11736 8114 11792
rect 8170 11736 14002 11792
rect 14058 11736 14063 11792
rect 8109 11734 14063 11736
rect 4061 11731 4127 11732
rect 8109 11731 8175 11734
rect 13997 11731 14063 11734
rect 15009 11794 15075 11797
rect 17309 11794 17375 11797
rect 15009 11792 17375 11794
rect 15009 11736 15014 11792
rect 15070 11736 17314 11792
rect 17370 11736 17375 11792
rect 15009 11734 17375 11736
rect 15009 11731 15075 11734
rect 16254 11661 16314 11734
rect 17309 11731 17375 11734
rect 4797 11658 4863 11661
rect 5809 11658 5875 11661
rect 4797 11656 5875 11658
rect 4797 11600 4802 11656
rect 4858 11600 5814 11656
rect 5870 11600 5875 11656
rect 4797 11598 5875 11600
rect 4797 11595 4863 11598
rect 5809 11595 5875 11598
rect 15285 11658 15351 11661
rect 16021 11658 16087 11661
rect 15285 11656 16087 11658
rect 15285 11600 15290 11656
rect 15346 11600 16026 11656
rect 16082 11600 16087 11656
rect 15285 11598 16087 11600
rect 15285 11595 15351 11598
rect 16021 11595 16087 11598
rect 16205 11656 16314 11661
rect 16205 11600 16210 11656
rect 16266 11600 16314 11656
rect 16205 11598 16314 11600
rect 16941 11658 17007 11661
rect 17585 11658 17651 11661
rect 16941 11656 17651 11658
rect 16941 11600 16946 11656
rect 17002 11600 17590 11656
rect 17646 11600 17651 11656
rect 16941 11598 17651 11600
rect 16205 11595 16271 11598
rect 16941 11595 17007 11598
rect 17585 11595 17651 11598
rect 5625 11522 5691 11525
rect 5993 11522 6059 11525
rect 5625 11520 6059 11522
rect 5625 11464 5630 11520
rect 5686 11464 5998 11520
rect 6054 11464 6059 11520
rect 5625 11462 6059 11464
rect 5625 11459 5691 11462
rect 5993 11459 6059 11462
rect 14457 11522 14523 11525
rect 14733 11522 14799 11525
rect 14457 11520 14799 11522
rect 14457 11464 14462 11520
rect 14518 11464 14738 11520
rect 14794 11464 14799 11520
rect 14457 11462 14799 11464
rect 14457 11459 14523 11462
rect 14733 11459 14799 11462
rect 8208 11456 8528 11457
rect 8208 11392 8216 11456
rect 8280 11392 8296 11456
rect 8360 11392 8376 11456
rect 8440 11392 8456 11456
rect 8520 11392 8528 11456
rect 8208 11391 8528 11392
rect 15472 11456 15792 11457
rect 15472 11392 15480 11456
rect 15544 11392 15560 11456
rect 15624 11392 15640 11456
rect 15704 11392 15720 11456
rect 15784 11392 15792 11456
rect 15472 11391 15792 11392
rect 4889 11386 4955 11389
rect 6177 11386 6243 11389
rect 21030 11386 21036 11388
rect 4889 11384 6243 11386
rect 4889 11328 4894 11384
rect 4950 11328 6182 11384
rect 6238 11328 6243 11384
rect 4889 11326 6243 11328
rect 4889 11323 4955 11326
rect 6177 11323 6243 11326
rect 16622 11326 21036 11386
rect 4337 11250 4403 11253
rect 16622 11250 16682 11326
rect 21030 11324 21036 11326
rect 21100 11324 21106 11388
rect 4337 11248 16682 11250
rect 4337 11192 4342 11248
rect 4398 11192 16682 11248
rect 4337 11190 16682 11192
rect 17769 11250 17835 11253
rect 18689 11250 18755 11253
rect 17769 11248 18755 11250
rect 17769 11192 17774 11248
rect 17830 11192 18694 11248
rect 18750 11192 18755 11248
rect 17769 11190 18755 11192
rect 4337 11187 4403 11190
rect 17769 11187 17835 11190
rect 18689 11187 18755 11190
rect 23381 11250 23447 11253
rect 23520 11250 24000 11280
rect 23381 11248 24000 11250
rect 23381 11192 23386 11248
rect 23442 11192 24000 11248
rect 23381 11190 24000 11192
rect 23381 11187 23447 11190
rect 23520 11160 24000 11190
rect 4337 11114 4403 11117
rect 5073 11114 5139 11117
rect 4337 11112 5139 11114
rect 4337 11056 4342 11112
rect 4398 11056 5078 11112
rect 5134 11056 5139 11112
rect 4337 11054 5139 11056
rect 4337 11051 4403 11054
rect 5073 11051 5139 11054
rect 15377 11114 15443 11117
rect 17309 11114 17375 11117
rect 15377 11112 17375 11114
rect 15377 11056 15382 11112
rect 15438 11056 17314 11112
rect 17370 11056 17375 11112
rect 15377 11054 17375 11056
rect 15377 11051 15443 11054
rect 17309 11051 17375 11054
rect 18413 11114 18479 11117
rect 23381 11114 23447 11117
rect 18413 11112 23447 11114
rect 18413 11056 18418 11112
rect 18474 11056 23386 11112
rect 23442 11056 23447 11112
rect 18413 11054 23447 11056
rect 18413 11051 18479 11054
rect 23381 11051 23447 11054
rect 7189 10980 7255 10981
rect 7189 10976 7236 10980
rect 7300 10978 7306 10980
rect 15285 10978 15351 10981
rect 17769 10978 17835 10981
rect 7189 10920 7194 10976
rect 7189 10916 7236 10920
rect 7300 10918 7346 10978
rect 15285 10976 17835 10978
rect 15285 10920 15290 10976
rect 15346 10920 17774 10976
rect 17830 10920 17835 10976
rect 15285 10918 17835 10920
rect 7300 10916 7306 10918
rect 7189 10915 7255 10916
rect 15285 10915 15351 10918
rect 17769 10915 17835 10918
rect 4576 10912 4896 10913
rect 4576 10848 4584 10912
rect 4648 10848 4664 10912
rect 4728 10848 4744 10912
rect 4808 10848 4824 10912
rect 4888 10848 4896 10912
rect 4576 10847 4896 10848
rect 11840 10912 12160 10913
rect 11840 10848 11848 10912
rect 11912 10848 11928 10912
rect 11992 10848 12008 10912
rect 12072 10848 12088 10912
rect 12152 10848 12160 10912
rect 11840 10847 12160 10848
rect 19104 10912 19424 10913
rect 19104 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19272 10912
rect 19336 10848 19352 10912
rect 19416 10848 19424 10912
rect 19104 10847 19424 10848
rect 7833 10842 7899 10845
rect 9305 10842 9371 10845
rect 7833 10840 9371 10842
rect 7833 10784 7838 10840
rect 7894 10784 9310 10840
rect 9366 10784 9371 10840
rect 7833 10782 9371 10784
rect 7833 10779 7899 10782
rect 9305 10779 9371 10782
rect 16757 10842 16823 10845
rect 17309 10842 17375 10845
rect 16757 10840 17375 10842
rect 16757 10784 16762 10840
rect 16818 10784 17314 10840
rect 17370 10784 17375 10840
rect 16757 10782 17375 10784
rect 16757 10779 16823 10782
rect 17309 10779 17375 10782
rect 4521 10706 4587 10709
rect 7465 10706 7531 10709
rect 15929 10708 15995 10709
rect 4521 10704 7531 10706
rect 4521 10648 4526 10704
rect 4582 10648 7470 10704
rect 7526 10648 7531 10704
rect 4521 10646 7531 10648
rect 4521 10643 4587 10646
rect 7465 10643 7531 10646
rect 15878 10644 15884 10708
rect 15948 10706 15995 10708
rect 15948 10704 16040 10706
rect 15990 10648 16040 10704
rect 15948 10646 16040 10648
rect 15948 10644 15995 10646
rect 15929 10643 15995 10644
rect 5441 10570 5507 10573
rect 5168 10568 5507 10570
rect 5168 10512 5446 10568
rect 5502 10512 5507 10568
rect 5168 10510 5507 10512
rect 5168 10437 5228 10510
rect 5441 10507 5507 10510
rect 7925 10570 7991 10573
rect 9254 10570 9260 10572
rect 7925 10568 9260 10570
rect 7925 10512 7930 10568
rect 7986 10512 9260 10568
rect 7925 10510 9260 10512
rect 7925 10507 7991 10510
rect 9254 10508 9260 10510
rect 9324 10508 9330 10572
rect 12709 10570 12775 10573
rect 17401 10570 17467 10573
rect 12709 10568 17467 10570
rect 12709 10512 12714 10568
rect 12770 10512 17406 10568
rect 17462 10512 17467 10568
rect 12709 10510 17467 10512
rect 12709 10507 12775 10510
rect 17401 10507 17467 10510
rect 5165 10432 5231 10437
rect 5165 10376 5170 10432
rect 5226 10376 5231 10432
rect 5165 10371 5231 10376
rect 9489 10434 9555 10437
rect 12433 10434 12499 10437
rect 9489 10432 12499 10434
rect 9489 10376 9494 10432
rect 9550 10376 12438 10432
rect 12494 10376 12499 10432
rect 9489 10374 12499 10376
rect 9489 10371 9555 10374
rect 12433 10371 12499 10374
rect 19333 10434 19399 10437
rect 23520 10434 24000 10464
rect 19333 10432 24000 10434
rect 19333 10376 19338 10432
rect 19394 10376 24000 10432
rect 19333 10374 24000 10376
rect 19333 10371 19399 10374
rect 8208 10368 8528 10369
rect 8208 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8528 10368
rect 8208 10303 8528 10304
rect 15472 10368 15792 10369
rect 15472 10304 15480 10368
rect 15544 10304 15560 10368
rect 15624 10304 15640 10368
rect 15704 10304 15720 10368
rect 15784 10304 15792 10368
rect 23520 10344 24000 10374
rect 15472 10303 15792 10304
rect 4889 10298 4955 10301
rect 8017 10298 8083 10301
rect 4889 10296 8083 10298
rect 4889 10240 4894 10296
rect 4950 10240 8022 10296
rect 8078 10240 8083 10296
rect 4889 10238 8083 10240
rect 4889 10235 4955 10238
rect 8017 10235 8083 10238
rect 10133 10298 10199 10301
rect 14181 10298 14247 10301
rect 10133 10296 14247 10298
rect 10133 10240 10138 10296
rect 10194 10240 14186 10296
rect 14242 10240 14247 10296
rect 10133 10238 14247 10240
rect 10133 10235 10199 10238
rect 14181 10235 14247 10238
rect 18873 10298 18939 10301
rect 19149 10298 19215 10301
rect 18873 10296 19215 10298
rect 18873 10240 18878 10296
rect 18934 10240 19154 10296
rect 19210 10240 19215 10296
rect 18873 10238 19215 10240
rect 18873 10235 18939 10238
rect 19149 10235 19215 10238
rect 3877 10162 3943 10165
rect 10041 10162 10107 10165
rect 3877 10160 10107 10162
rect 3877 10104 3882 10160
rect 3938 10104 10046 10160
rect 10102 10104 10107 10160
rect 3877 10102 10107 10104
rect 3877 10099 3943 10102
rect 10041 10099 10107 10102
rect 15377 10162 15443 10165
rect 20069 10162 20135 10165
rect 15377 10160 20135 10162
rect 15377 10104 15382 10160
rect 15438 10104 20074 10160
rect 20130 10104 20135 10160
rect 15377 10102 20135 10104
rect 15377 10099 15443 10102
rect 20069 10099 20135 10102
rect 1853 10026 1919 10029
rect 15142 10026 15148 10028
rect 1853 10024 15148 10026
rect 1853 9968 1858 10024
rect 1914 9968 15148 10024
rect 1853 9966 15148 9968
rect 1853 9963 1919 9966
rect 15142 9964 15148 9966
rect 15212 9964 15218 10028
rect 15285 10026 15351 10029
rect 16573 10026 16639 10029
rect 19517 10028 19583 10029
rect 19517 10026 19564 10028
rect 15285 10024 16639 10026
rect 15285 9968 15290 10024
rect 15346 9968 16578 10024
rect 16634 9968 16639 10024
rect 15285 9966 16639 9968
rect 19472 10024 19564 10026
rect 19472 9968 19522 10024
rect 19472 9966 19564 9968
rect 15285 9963 15351 9966
rect 16573 9963 16639 9966
rect 19517 9964 19564 9966
rect 19628 9964 19634 10028
rect 19517 9963 19583 9964
rect 7465 9890 7531 9893
rect 5996 9888 7531 9890
rect 5996 9832 7470 9888
rect 7526 9832 7531 9888
rect 5996 9830 7531 9832
rect 4576 9824 4896 9825
rect 4576 9760 4584 9824
rect 4648 9760 4664 9824
rect 4728 9760 4744 9824
rect 4808 9760 4824 9824
rect 4888 9760 4896 9824
rect 4576 9759 4896 9760
rect 5349 9754 5415 9757
rect 5996 9754 6056 9830
rect 7465 9827 7531 9830
rect 8017 9890 8083 9893
rect 9949 9890 10015 9893
rect 8017 9888 10015 9890
rect 8017 9832 8022 9888
rect 8078 9832 9954 9888
rect 10010 9832 10015 9888
rect 8017 9830 10015 9832
rect 8017 9827 8083 9830
rect 9949 9827 10015 9830
rect 12249 9890 12315 9893
rect 12985 9890 13051 9893
rect 13537 9890 13603 9893
rect 15288 9890 15348 9963
rect 12249 9888 15348 9890
rect 12249 9832 12254 9888
rect 12310 9832 12990 9888
rect 13046 9832 13542 9888
rect 13598 9832 15348 9888
rect 12249 9830 15348 9832
rect 12249 9827 12315 9830
rect 12985 9827 13051 9830
rect 13537 9827 13603 9830
rect 11840 9824 12160 9825
rect 11840 9760 11848 9824
rect 11912 9760 11928 9824
rect 11992 9760 12008 9824
rect 12072 9760 12088 9824
rect 12152 9760 12160 9824
rect 11840 9759 12160 9760
rect 19104 9824 19424 9825
rect 19104 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19272 9824
rect 19336 9760 19352 9824
rect 19416 9760 19424 9824
rect 19104 9759 19424 9760
rect 8937 9754 9003 9757
rect 5349 9752 6056 9754
rect 5349 9696 5354 9752
rect 5410 9696 6056 9752
rect 5349 9694 6056 9696
rect 6134 9752 9003 9754
rect 6134 9696 8942 9752
rect 8998 9696 9003 9752
rect 6134 9694 9003 9696
rect 5349 9691 5415 9694
rect 2681 9618 2747 9621
rect 6134 9618 6194 9694
rect 8937 9691 9003 9694
rect 9121 9754 9187 9757
rect 11053 9754 11119 9757
rect 9121 9752 11119 9754
rect 9121 9696 9126 9752
rect 9182 9696 11058 9752
rect 11114 9696 11119 9752
rect 9121 9694 11119 9696
rect 9121 9691 9187 9694
rect 11053 9691 11119 9694
rect 19517 9754 19583 9757
rect 23520 9754 24000 9784
rect 19517 9752 24000 9754
rect 19517 9696 19522 9752
rect 19578 9696 24000 9752
rect 19517 9694 24000 9696
rect 19517 9691 19583 9694
rect 23520 9664 24000 9694
rect 2681 9616 6194 9618
rect 2681 9560 2686 9616
rect 2742 9560 6194 9616
rect 2681 9558 6194 9560
rect 6545 9618 6611 9621
rect 12341 9618 12407 9621
rect 13629 9618 13695 9621
rect 6545 9616 12407 9618
rect 6545 9560 6550 9616
rect 6606 9560 12346 9616
rect 12402 9560 12407 9616
rect 6545 9558 12407 9560
rect 2681 9555 2747 9558
rect 6545 9555 6611 9558
rect 12341 9555 12407 9558
rect 12758 9616 13695 9618
rect 12758 9560 13634 9616
rect 13690 9560 13695 9616
rect 12758 9558 13695 9560
rect 1577 9482 1643 9485
rect 5165 9482 5231 9485
rect 1577 9480 5231 9482
rect 1577 9424 1582 9480
rect 1638 9424 5170 9480
rect 5226 9424 5231 9480
rect 1577 9422 5231 9424
rect 1577 9419 1643 9422
rect 5165 9419 5231 9422
rect 8109 9482 8175 9485
rect 12758 9482 12818 9558
rect 13629 9555 13695 9558
rect 14825 9618 14891 9621
rect 18781 9618 18847 9621
rect 14825 9616 18847 9618
rect 14825 9560 14830 9616
rect 14886 9560 18786 9616
rect 18842 9560 18847 9616
rect 14825 9558 18847 9560
rect 14825 9555 14891 9558
rect 18781 9555 18847 9558
rect 19333 9584 19399 9587
rect 19333 9582 19442 9584
rect 19333 9526 19338 9582
rect 19394 9526 19442 9582
rect 19333 9521 19442 9526
rect 8109 9480 12818 9482
rect 8109 9424 8114 9480
rect 8170 9424 12818 9480
rect 8109 9422 12818 9424
rect 12893 9482 12959 9485
rect 17217 9482 17283 9485
rect 18689 9482 18755 9485
rect 19149 9482 19215 9485
rect 12893 9480 17283 9482
rect 12893 9424 12898 9480
rect 12954 9424 17222 9480
rect 17278 9424 17283 9480
rect 12893 9422 17283 9424
rect 8109 9419 8175 9422
rect 12893 9419 12959 9422
rect 17217 9419 17283 9422
rect 17358 9480 19215 9482
rect 17358 9424 18694 9480
rect 18750 9424 19154 9480
rect 19210 9424 19215 9480
rect 17358 9422 19215 9424
rect 19382 9482 19442 9521
rect 20161 9482 20227 9485
rect 19382 9480 20227 9482
rect 19382 9424 20166 9480
rect 20222 9424 20227 9480
rect 19382 9422 20227 9424
rect 3969 9346 4035 9349
rect 8017 9346 8083 9349
rect 13905 9346 13971 9349
rect 3969 9344 8083 9346
rect 3969 9288 3974 9344
rect 4030 9288 8022 9344
rect 8078 9288 8083 9344
rect 3969 9286 8083 9288
rect 3969 9283 4035 9286
rect 8017 9283 8083 9286
rect 9814 9344 13971 9346
rect 9814 9288 13910 9344
rect 13966 9288 13971 9344
rect 9814 9286 13971 9288
rect 8208 9280 8528 9281
rect 8208 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8528 9280
rect 8208 9215 8528 9216
rect 2497 9210 2563 9213
rect 5809 9210 5875 9213
rect 7833 9210 7899 9213
rect 2497 9208 5875 9210
rect 2497 9152 2502 9208
rect 2558 9152 5814 9208
rect 5870 9152 5875 9208
rect 2497 9150 5875 9152
rect 2497 9147 2563 9150
rect 5809 9147 5875 9150
rect 6686 9208 7899 9210
rect 6686 9152 7838 9208
rect 7894 9152 7899 9208
rect 6686 9150 7899 9152
rect 3693 9074 3759 9077
rect 6545 9074 6611 9077
rect 6686 9074 6746 9150
rect 7833 9147 7899 9150
rect 3693 9072 6746 9074
rect 3693 9016 3698 9072
rect 3754 9016 6550 9072
rect 6606 9016 6746 9072
rect 3693 9014 6746 9016
rect 7557 9074 7623 9077
rect 9305 9074 9371 9077
rect 9814 9074 9874 9286
rect 13905 9283 13971 9286
rect 15929 9346 15995 9349
rect 17358 9346 17418 9422
rect 18689 9419 18755 9422
rect 19149 9419 19215 9422
rect 20161 9419 20227 9422
rect 15929 9344 17418 9346
rect 15929 9288 15934 9344
rect 15990 9288 17418 9344
rect 15929 9286 17418 9288
rect 15929 9283 15995 9286
rect 15472 9280 15792 9281
rect 15472 9216 15480 9280
rect 15544 9216 15560 9280
rect 15624 9216 15640 9280
rect 15704 9216 15720 9280
rect 15784 9216 15792 9280
rect 15472 9215 15792 9216
rect 11237 9210 11303 9213
rect 13721 9210 13787 9213
rect 14181 9210 14247 9213
rect 11237 9208 14247 9210
rect 11237 9152 11242 9208
rect 11298 9152 13726 9208
rect 13782 9152 14186 9208
rect 14242 9152 14247 9208
rect 11237 9150 14247 9152
rect 11237 9147 11303 9150
rect 13721 9147 13787 9150
rect 14181 9147 14247 9150
rect 7557 9072 8954 9074
rect 7557 9016 7562 9072
rect 7618 9016 8954 9072
rect 7557 9014 8954 9016
rect 3693 9011 3759 9014
rect 6545 9011 6611 9014
rect 7557 9011 7623 9014
rect 4061 8938 4127 8941
rect 5165 8938 5231 8941
rect 8702 8938 8708 8940
rect 4061 8936 5090 8938
rect 4061 8880 4066 8936
rect 4122 8880 5090 8936
rect 4061 8878 5090 8880
rect 4061 8875 4127 8878
rect 5030 8802 5090 8878
rect 5165 8936 8708 8938
rect 5165 8880 5170 8936
rect 5226 8880 8708 8936
rect 5165 8878 8708 8880
rect 5165 8875 5231 8878
rect 8702 8876 8708 8878
rect 8772 8876 8778 8940
rect 8894 8938 8954 9014
rect 9305 9072 9874 9074
rect 9305 9016 9310 9072
rect 9366 9016 9874 9072
rect 9305 9014 9874 9016
rect 9949 9074 10015 9077
rect 10777 9074 10843 9077
rect 9949 9072 10843 9074
rect 9949 9016 9954 9072
rect 10010 9016 10782 9072
rect 10838 9016 10843 9072
rect 9949 9014 10843 9016
rect 9305 9011 9371 9014
rect 9949 9011 10015 9014
rect 10777 9011 10843 9014
rect 10961 9074 11027 9077
rect 21725 9074 21791 9077
rect 10961 9072 21791 9074
rect 10961 9016 10966 9072
rect 11022 9016 21730 9072
rect 21786 9016 21791 9072
rect 10961 9014 21791 9016
rect 10961 9011 11027 9014
rect 21725 9011 21791 9014
rect 22001 9074 22067 9077
rect 23520 9074 24000 9104
rect 22001 9072 24000 9074
rect 22001 9016 22006 9072
rect 22062 9016 24000 9072
rect 22001 9014 24000 9016
rect 22001 9011 22067 9014
rect 23520 8984 24000 9014
rect 12617 8938 12683 8941
rect 17493 8938 17559 8941
rect 20478 8938 20484 8940
rect 8894 8878 12450 8938
rect 10961 8802 11027 8805
rect 5030 8800 11027 8802
rect 5030 8744 10966 8800
rect 11022 8744 11027 8800
rect 5030 8742 11027 8744
rect 10961 8739 11027 8742
rect 4576 8736 4896 8737
rect 4576 8672 4584 8736
rect 4648 8672 4664 8736
rect 4728 8672 4744 8736
rect 4808 8672 4824 8736
rect 4888 8672 4896 8736
rect 4576 8671 4896 8672
rect 11840 8736 12160 8737
rect 11840 8672 11848 8736
rect 11912 8672 11928 8736
rect 11992 8672 12008 8736
rect 12072 8672 12088 8736
rect 12152 8672 12160 8736
rect 11840 8671 12160 8672
rect 5349 8666 5415 8669
rect 11462 8666 11468 8668
rect 5349 8664 11468 8666
rect 5349 8608 5354 8664
rect 5410 8608 11468 8664
rect 5349 8606 11468 8608
rect 5349 8603 5415 8606
rect 11462 8604 11468 8606
rect 11532 8604 11538 8668
rect 12390 8666 12450 8878
rect 12617 8936 17559 8938
rect 12617 8880 12622 8936
rect 12678 8880 17498 8936
rect 17554 8880 17559 8936
rect 12617 8878 17559 8880
rect 12617 8875 12683 8878
rect 17493 8875 17559 8878
rect 18462 8878 20484 8938
rect 12525 8802 12591 8805
rect 18321 8802 18387 8805
rect 12525 8800 18387 8802
rect 12525 8744 12530 8800
rect 12586 8744 18326 8800
rect 18382 8744 18387 8800
rect 12525 8742 18387 8744
rect 12525 8739 12591 8742
rect 18321 8739 18387 8742
rect 18462 8666 18522 8878
rect 20478 8876 20484 8878
rect 20548 8876 20554 8940
rect 19104 8736 19424 8737
rect 19104 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19272 8736
rect 19336 8672 19352 8736
rect 19416 8672 19424 8736
rect 19104 8671 19424 8672
rect 12390 8606 18522 8666
rect 5073 8530 5139 8533
rect 22093 8530 22159 8533
rect 5073 8528 22159 8530
rect 5073 8472 5078 8528
rect 5134 8472 22098 8528
rect 22154 8472 22159 8528
rect 5073 8470 22159 8472
rect 5073 8467 5139 8470
rect 22093 8467 22159 8470
rect 9489 8394 9555 8397
rect 14733 8394 14799 8397
rect 16389 8394 16455 8397
rect 7974 8334 8770 8394
rect 5257 8258 5323 8261
rect 7974 8258 8034 8334
rect 5257 8256 8034 8258
rect 5257 8200 5262 8256
rect 5318 8200 8034 8256
rect 5257 8198 8034 8200
rect 8710 8258 8770 8334
rect 9489 8392 14799 8394
rect 9489 8336 9494 8392
rect 9550 8336 14738 8392
rect 14794 8336 14799 8392
rect 9489 8334 14799 8336
rect 9489 8331 9555 8334
rect 14733 8331 14799 8334
rect 15334 8392 16455 8394
rect 15334 8336 16394 8392
rect 16450 8336 16455 8392
rect 15334 8334 16455 8336
rect 13261 8258 13327 8261
rect 8710 8256 13327 8258
rect 8710 8200 13266 8256
rect 13322 8200 13327 8256
rect 8710 8198 13327 8200
rect 5257 8195 5323 8198
rect 13261 8195 13327 8198
rect 13721 8258 13787 8261
rect 15334 8258 15394 8334
rect 16389 8331 16455 8334
rect 20478 8332 20484 8396
rect 20548 8394 20554 8396
rect 21265 8394 21331 8397
rect 20548 8392 21331 8394
rect 20548 8336 21270 8392
rect 21326 8336 21331 8392
rect 20548 8334 21331 8336
rect 20548 8332 20554 8334
rect 21265 8331 21331 8334
rect 13721 8256 15394 8258
rect 13721 8200 13726 8256
rect 13782 8200 15394 8256
rect 13721 8198 15394 8200
rect 19701 8258 19767 8261
rect 23520 8258 24000 8288
rect 19701 8256 24000 8258
rect 19701 8200 19706 8256
rect 19762 8200 24000 8256
rect 19701 8198 24000 8200
rect 13721 8195 13787 8198
rect 19701 8195 19767 8198
rect 8208 8192 8528 8193
rect 8208 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8528 8192
rect 8208 8127 8528 8128
rect 15472 8192 15792 8193
rect 15472 8128 15480 8192
rect 15544 8128 15560 8192
rect 15624 8128 15640 8192
rect 15704 8128 15720 8192
rect 15784 8128 15792 8192
rect 23520 8168 24000 8198
rect 15472 8127 15792 8128
rect 15326 8122 15332 8124
rect 8710 8062 15332 8122
rect 5441 7986 5507 7989
rect 8710 7986 8770 8062
rect 15326 8060 15332 8062
rect 15396 8060 15402 8124
rect 5441 7984 8770 7986
rect 5441 7928 5446 7984
rect 5502 7928 8770 7984
rect 5441 7926 8770 7928
rect 8845 7986 8911 7989
rect 18413 7986 18479 7989
rect 8845 7984 18479 7986
rect 8845 7928 8850 7984
rect 8906 7928 18418 7984
rect 18474 7928 18479 7984
rect 8845 7926 18479 7928
rect 5441 7923 5507 7926
rect 8845 7923 8911 7926
rect 18413 7923 18479 7926
rect 4429 7850 4495 7853
rect 19517 7850 19583 7853
rect 4429 7848 19583 7850
rect 4429 7792 4434 7848
rect 4490 7792 19522 7848
rect 19578 7792 19583 7848
rect 4429 7790 19583 7792
rect 4429 7787 4495 7790
rect 19517 7787 19583 7790
rect 7557 7714 7623 7717
rect 11145 7714 11211 7717
rect 7557 7712 11211 7714
rect 7557 7656 7562 7712
rect 7618 7656 11150 7712
rect 11206 7656 11211 7712
rect 7557 7654 11211 7656
rect 7557 7651 7623 7654
rect 11145 7651 11211 7654
rect 13721 7714 13787 7717
rect 13721 7712 15578 7714
rect 13721 7656 13726 7712
rect 13782 7656 15578 7712
rect 13721 7654 15578 7656
rect 13721 7651 13787 7654
rect 4576 7648 4896 7649
rect 4576 7584 4584 7648
rect 4648 7584 4664 7648
rect 4728 7584 4744 7648
rect 4808 7584 4824 7648
rect 4888 7584 4896 7648
rect 4576 7583 4896 7584
rect 11840 7648 12160 7649
rect 11840 7584 11848 7648
rect 11912 7584 11928 7648
rect 11992 7584 12008 7648
rect 12072 7584 12088 7648
rect 12152 7584 12160 7648
rect 11840 7583 12160 7584
rect 6361 7578 6427 7581
rect 11697 7578 11763 7581
rect 6361 7576 11763 7578
rect 6361 7520 6366 7576
rect 6422 7520 11702 7576
rect 11758 7520 11763 7576
rect 6361 7518 11763 7520
rect 6361 7515 6427 7518
rect 11697 7515 11763 7518
rect 12341 7578 12407 7581
rect 15377 7578 15443 7581
rect 12341 7576 15443 7578
rect 12341 7520 12346 7576
rect 12402 7520 15382 7576
rect 15438 7520 15443 7576
rect 12341 7518 15443 7520
rect 15518 7578 15578 7654
rect 19104 7648 19424 7649
rect 19104 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19272 7648
rect 19336 7584 19352 7648
rect 19416 7584 19424 7648
rect 19104 7583 19424 7584
rect 21909 7578 21975 7581
rect 23520 7578 24000 7608
rect 15518 7518 18338 7578
rect 12341 7515 12407 7518
rect 15377 7515 15443 7518
rect 7281 7442 7347 7445
rect 13721 7442 13787 7445
rect 7281 7440 13787 7442
rect 7281 7384 7286 7440
rect 7342 7384 13726 7440
rect 13782 7384 13787 7440
rect 7281 7382 13787 7384
rect 7281 7379 7347 7382
rect 13721 7379 13787 7382
rect 13997 7442 14063 7445
rect 14365 7442 14431 7445
rect 16665 7442 16731 7445
rect 18045 7442 18111 7445
rect 13997 7440 18111 7442
rect 13997 7384 14002 7440
rect 14058 7384 14370 7440
rect 14426 7384 16670 7440
rect 16726 7384 18050 7440
rect 18106 7384 18111 7440
rect 13997 7382 18111 7384
rect 18278 7442 18338 7518
rect 21909 7576 24000 7578
rect 21909 7520 21914 7576
rect 21970 7520 24000 7576
rect 21909 7518 24000 7520
rect 21909 7515 21975 7518
rect 23520 7488 24000 7518
rect 20989 7442 21055 7445
rect 18278 7440 21055 7442
rect 18278 7384 20994 7440
rect 21050 7384 21055 7440
rect 18278 7382 21055 7384
rect 13997 7379 14063 7382
rect 14365 7379 14431 7382
rect 16665 7379 16731 7382
rect 18045 7379 18111 7382
rect 20989 7379 21055 7382
rect 4245 7306 4311 7309
rect 12249 7306 12315 7309
rect 15469 7306 15535 7309
rect 4245 7304 8770 7306
rect 4245 7248 4250 7304
rect 4306 7248 8770 7304
rect 4245 7246 8770 7248
rect 4245 7243 4311 7246
rect 8710 7170 8770 7246
rect 12249 7304 15535 7306
rect 12249 7248 12254 7304
rect 12310 7248 15474 7304
rect 15530 7248 15535 7304
rect 12249 7246 15535 7248
rect 12249 7243 12315 7246
rect 15469 7243 15535 7246
rect 14958 7170 14964 7172
rect 8710 7110 14964 7170
rect 14958 7108 14964 7110
rect 15028 7108 15034 7172
rect 8208 7104 8528 7105
rect 8208 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8528 7104
rect 8208 7039 8528 7040
rect 15472 7104 15792 7105
rect 15472 7040 15480 7104
rect 15544 7040 15560 7104
rect 15624 7040 15640 7104
rect 15704 7040 15720 7104
rect 15784 7040 15792 7104
rect 15472 7039 15792 7040
rect 4705 7034 4771 7037
rect 14774 7034 14780 7036
rect 4705 7032 8034 7034
rect 4705 6976 4710 7032
rect 4766 6976 8034 7032
rect 4705 6974 8034 6976
rect 4705 6971 4771 6974
rect 7974 6898 8034 6974
rect 8710 6974 14780 7034
rect 8710 6898 8770 6974
rect 14774 6972 14780 6974
rect 14844 6972 14850 7036
rect 7974 6838 8770 6898
rect 12065 6898 12131 6901
rect 15101 6898 15167 6901
rect 12065 6896 15167 6898
rect 12065 6840 12070 6896
rect 12126 6840 15106 6896
rect 15162 6840 15167 6896
rect 12065 6838 15167 6840
rect 12065 6835 12131 6838
rect 15101 6835 15167 6838
rect 20621 6898 20687 6901
rect 23520 6898 24000 6928
rect 20621 6896 24000 6898
rect 20621 6840 20626 6896
rect 20682 6840 24000 6896
rect 20621 6838 24000 6840
rect 20621 6835 20687 6838
rect 23520 6808 24000 6838
rect 12341 6762 12407 6765
rect 16205 6762 16271 6765
rect 12341 6760 16271 6762
rect 12341 6704 12346 6760
rect 12402 6704 16210 6760
rect 16266 6704 16271 6760
rect 12341 6702 16271 6704
rect 12341 6699 12407 6702
rect 16205 6699 16271 6702
rect 4576 6560 4896 6561
rect 4576 6496 4584 6560
rect 4648 6496 4664 6560
rect 4728 6496 4744 6560
rect 4808 6496 4824 6560
rect 4888 6496 4896 6560
rect 4576 6495 4896 6496
rect 11840 6560 12160 6561
rect 11840 6496 11848 6560
rect 11912 6496 11928 6560
rect 11992 6496 12008 6560
rect 12072 6496 12088 6560
rect 12152 6496 12160 6560
rect 11840 6495 12160 6496
rect 19104 6560 19424 6561
rect 19104 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19272 6560
rect 19336 6496 19352 6560
rect 19416 6496 19424 6560
rect 19104 6495 19424 6496
rect 8109 6490 8175 6493
rect 9489 6490 9555 6493
rect 8109 6488 9555 6490
rect 8109 6432 8114 6488
rect 8170 6432 9494 6488
rect 9550 6432 9555 6488
rect 8109 6430 9555 6432
rect 8109 6427 8175 6430
rect 9489 6427 9555 6430
rect 8017 6354 8083 6357
rect 11789 6354 11855 6357
rect 8017 6352 11855 6354
rect 8017 6296 8022 6352
rect 8078 6296 11794 6352
rect 11850 6296 11855 6352
rect 8017 6294 11855 6296
rect 8017 6291 8083 6294
rect 11789 6291 11855 6294
rect 13077 6354 13143 6357
rect 14181 6354 14247 6357
rect 13077 6352 14247 6354
rect 13077 6296 13082 6352
rect 13138 6296 14186 6352
rect 14242 6296 14247 6352
rect 13077 6294 14247 6296
rect 13077 6291 13143 6294
rect 14181 6291 14247 6294
rect 17309 6354 17375 6357
rect 19793 6354 19859 6357
rect 17309 6352 19859 6354
rect 17309 6296 17314 6352
rect 17370 6296 19798 6352
rect 19854 6296 19859 6352
rect 17309 6294 19859 6296
rect 17309 6291 17375 6294
rect 19793 6291 19859 6294
rect 14089 6218 14155 6221
rect 17125 6218 17191 6221
rect 14089 6216 17191 6218
rect 14089 6160 14094 6216
rect 14150 6160 17130 6216
rect 17186 6160 17191 6216
rect 14089 6158 17191 6160
rect 14089 6155 14155 6158
rect 17125 6155 17191 6158
rect 16297 6082 16363 6085
rect 18689 6082 18755 6085
rect 16297 6080 18755 6082
rect 16297 6024 16302 6080
rect 16358 6024 18694 6080
rect 18750 6024 18755 6080
rect 16297 6022 18755 6024
rect 16297 6019 16363 6022
rect 18689 6019 18755 6022
rect 22277 6082 22343 6085
rect 23520 6082 24000 6112
rect 22277 6080 24000 6082
rect 22277 6024 22282 6080
rect 22338 6024 24000 6080
rect 22277 6022 24000 6024
rect 22277 6019 22343 6022
rect 8208 6016 8528 6017
rect 8208 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8528 6016
rect 8208 5951 8528 5952
rect 15472 6016 15792 6017
rect 15472 5952 15480 6016
rect 15544 5952 15560 6016
rect 15624 5952 15640 6016
rect 15704 5952 15720 6016
rect 15784 5952 15792 6016
rect 23520 5992 24000 6022
rect 15472 5951 15792 5952
rect 12249 5810 12315 5813
rect 14365 5810 14431 5813
rect 12249 5808 14431 5810
rect 12249 5752 12254 5808
rect 12310 5752 14370 5808
rect 14426 5752 14431 5808
rect 12249 5750 14431 5752
rect 12249 5747 12315 5750
rect 14365 5747 14431 5750
rect 4576 5472 4896 5473
rect 4576 5408 4584 5472
rect 4648 5408 4664 5472
rect 4728 5408 4744 5472
rect 4808 5408 4824 5472
rect 4888 5408 4896 5472
rect 4576 5407 4896 5408
rect 11840 5472 12160 5473
rect 11840 5408 11848 5472
rect 11912 5408 11928 5472
rect 11992 5408 12008 5472
rect 12072 5408 12088 5472
rect 12152 5408 12160 5472
rect 11840 5407 12160 5408
rect 19104 5472 19424 5473
rect 19104 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19272 5472
rect 19336 5408 19352 5472
rect 19416 5408 19424 5472
rect 19104 5407 19424 5408
rect 16205 5402 16271 5405
rect 17585 5402 17651 5405
rect 16205 5400 17651 5402
rect 16205 5344 16210 5400
rect 16266 5344 17590 5400
rect 17646 5344 17651 5400
rect 16205 5342 17651 5344
rect 16205 5339 16271 5342
rect 17585 5339 17651 5342
rect 19885 5402 19951 5405
rect 23520 5402 24000 5432
rect 19885 5400 24000 5402
rect 19885 5344 19890 5400
rect 19946 5344 24000 5400
rect 19885 5342 24000 5344
rect 19885 5339 19951 5342
rect 23520 5312 24000 5342
rect 8208 4928 8528 4929
rect 8208 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8528 4928
rect 8208 4863 8528 4864
rect 15472 4928 15792 4929
rect 15472 4864 15480 4928
rect 15544 4864 15560 4928
rect 15624 4864 15640 4928
rect 15704 4864 15720 4928
rect 15784 4864 15792 4928
rect 15472 4863 15792 4864
rect 10041 4858 10107 4861
rect 14917 4858 14983 4861
rect 10041 4856 14983 4858
rect 10041 4800 10046 4856
rect 10102 4800 14922 4856
rect 14978 4800 14983 4856
rect 10041 4798 14983 4800
rect 10041 4795 10107 4798
rect 14917 4795 14983 4798
rect 18597 4722 18663 4725
rect 23520 4722 24000 4752
rect 18597 4720 24000 4722
rect 18597 4664 18602 4720
rect 18658 4664 24000 4720
rect 18597 4662 24000 4664
rect 18597 4659 18663 4662
rect 23520 4632 24000 4662
rect 4576 4384 4896 4385
rect 4576 4320 4584 4384
rect 4648 4320 4664 4384
rect 4728 4320 4744 4384
rect 4808 4320 4824 4384
rect 4888 4320 4896 4384
rect 4576 4319 4896 4320
rect 11840 4384 12160 4385
rect 11840 4320 11848 4384
rect 11912 4320 11928 4384
rect 11992 4320 12008 4384
rect 12072 4320 12088 4384
rect 12152 4320 12160 4384
rect 11840 4319 12160 4320
rect 19104 4384 19424 4385
rect 19104 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19272 4384
rect 19336 4320 19352 4384
rect 19416 4320 19424 4384
rect 19104 4319 19424 4320
rect 12525 4314 12591 4317
rect 16113 4314 16179 4317
rect 12525 4312 16179 4314
rect 12525 4256 12530 4312
rect 12586 4256 16118 4312
rect 16174 4256 16179 4312
rect 12525 4254 16179 4256
rect 12525 4251 12591 4254
rect 16113 4251 16179 4254
rect 7741 4178 7807 4181
rect 13813 4178 13879 4181
rect 7741 4176 13879 4178
rect 7741 4120 7746 4176
rect 7802 4120 13818 4176
rect 13874 4120 13879 4176
rect 7741 4118 13879 4120
rect 7741 4115 7807 4118
rect 13813 4115 13879 4118
rect 0 4042 480 4072
rect 3601 4042 3667 4045
rect 0 4040 3667 4042
rect 0 3984 3606 4040
rect 3662 3984 3667 4040
rect 0 3982 3667 3984
rect 0 3952 480 3982
rect 3601 3979 3667 3982
rect 12709 4042 12775 4045
rect 16021 4042 16087 4045
rect 12709 4040 16087 4042
rect 12709 3984 12714 4040
rect 12770 3984 16026 4040
rect 16082 3984 16087 4040
rect 12709 3982 16087 3984
rect 12709 3979 12775 3982
rect 16021 3979 16087 3982
rect 12249 3906 12315 3909
rect 15193 3906 15259 3909
rect 12249 3904 15259 3906
rect 12249 3848 12254 3904
rect 12310 3848 15198 3904
rect 15254 3848 15259 3904
rect 12249 3846 15259 3848
rect 12249 3843 12315 3846
rect 15193 3843 15259 3846
rect 19885 3906 19951 3909
rect 23520 3906 24000 3936
rect 19885 3904 24000 3906
rect 19885 3848 19890 3904
rect 19946 3848 24000 3904
rect 19885 3846 24000 3848
rect 19885 3843 19951 3846
rect 8208 3840 8528 3841
rect 8208 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8528 3840
rect 8208 3775 8528 3776
rect 15472 3840 15792 3841
rect 15472 3776 15480 3840
rect 15544 3776 15560 3840
rect 15624 3776 15640 3840
rect 15704 3776 15720 3840
rect 15784 3776 15792 3840
rect 23520 3816 24000 3846
rect 15472 3775 15792 3776
rect 14641 3634 14707 3637
rect 15837 3634 15903 3637
rect 14641 3632 15903 3634
rect 14641 3576 14646 3632
rect 14702 3576 15842 3632
rect 15898 3576 15903 3632
rect 14641 3574 15903 3576
rect 14641 3571 14707 3574
rect 15837 3571 15903 3574
rect 12433 3498 12499 3501
rect 15377 3498 15443 3501
rect 12433 3496 15443 3498
rect 12433 3440 12438 3496
rect 12494 3440 15382 3496
rect 15438 3440 15443 3496
rect 12433 3438 15443 3440
rect 12433 3435 12499 3438
rect 15377 3435 15443 3438
rect 4576 3296 4896 3297
rect 4576 3232 4584 3296
rect 4648 3232 4664 3296
rect 4728 3232 4744 3296
rect 4808 3232 4824 3296
rect 4888 3232 4896 3296
rect 4576 3231 4896 3232
rect 11840 3296 12160 3297
rect 11840 3232 11848 3296
rect 11912 3232 11928 3296
rect 11992 3232 12008 3296
rect 12072 3232 12088 3296
rect 12152 3232 12160 3296
rect 11840 3231 12160 3232
rect 19104 3296 19424 3297
rect 19104 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19272 3296
rect 19336 3232 19352 3296
rect 19416 3232 19424 3296
rect 19104 3231 19424 3232
rect 13905 3226 13971 3229
rect 16297 3226 16363 3229
rect 13905 3224 16363 3226
rect 13905 3168 13910 3224
rect 13966 3168 16302 3224
rect 16358 3168 16363 3224
rect 13905 3166 16363 3168
rect 13905 3163 13971 3166
rect 16297 3163 16363 3166
rect 20345 3226 20411 3229
rect 23520 3226 24000 3256
rect 20345 3224 24000 3226
rect 20345 3168 20350 3224
rect 20406 3168 24000 3224
rect 20345 3166 24000 3168
rect 20345 3163 20411 3166
rect 23520 3136 24000 3166
rect 8208 2752 8528 2753
rect 8208 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8528 2752
rect 8208 2687 8528 2688
rect 15472 2752 15792 2753
rect 15472 2688 15480 2752
rect 15544 2688 15560 2752
rect 15624 2688 15640 2752
rect 15704 2688 15720 2752
rect 15784 2688 15792 2752
rect 15472 2687 15792 2688
rect 18873 2546 18939 2549
rect 23520 2546 24000 2576
rect 18873 2544 24000 2546
rect 18873 2488 18878 2544
rect 18934 2488 24000 2544
rect 18873 2486 24000 2488
rect 18873 2483 18939 2486
rect 23520 2456 24000 2486
rect 4576 2208 4896 2209
rect 4576 2144 4584 2208
rect 4648 2144 4664 2208
rect 4728 2144 4744 2208
rect 4808 2144 4824 2208
rect 4888 2144 4896 2208
rect 4576 2143 4896 2144
rect 11840 2208 12160 2209
rect 11840 2144 11848 2208
rect 11912 2144 11928 2208
rect 11992 2144 12008 2208
rect 12072 2144 12088 2208
rect 12152 2144 12160 2208
rect 11840 2143 12160 2144
rect 19104 2208 19424 2209
rect 19104 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19272 2208
rect 19336 2144 19352 2208
rect 19416 2144 19424 2208
rect 19104 2143 19424 2144
rect 20478 1668 20484 1732
rect 20548 1730 20554 1732
rect 23520 1730 24000 1760
rect 20548 1670 24000 1730
rect 20548 1668 20554 1670
rect 23520 1640 24000 1670
rect 20529 1050 20595 1053
rect 23520 1050 24000 1080
rect 20529 1048 24000 1050
rect 20529 992 20534 1048
rect 20590 992 24000 1048
rect 20529 990 24000 992
rect 20529 987 20595 990
rect 23520 960 24000 990
rect 20621 370 20687 373
rect 23520 370 24000 400
rect 20621 368 24000 370
rect 20621 312 20626 368
rect 20682 312 24000 368
rect 20621 310 24000 312
rect 20621 307 20687 310
rect 23520 280 24000 310
<< via3 >>
rect 4584 21788 4648 21792
rect 4584 21732 4588 21788
rect 4588 21732 4644 21788
rect 4644 21732 4648 21788
rect 4584 21728 4648 21732
rect 4664 21788 4728 21792
rect 4664 21732 4668 21788
rect 4668 21732 4724 21788
rect 4724 21732 4728 21788
rect 4664 21728 4728 21732
rect 4744 21788 4808 21792
rect 4744 21732 4748 21788
rect 4748 21732 4804 21788
rect 4804 21732 4808 21788
rect 4744 21728 4808 21732
rect 4824 21788 4888 21792
rect 4824 21732 4828 21788
rect 4828 21732 4884 21788
rect 4884 21732 4888 21788
rect 4824 21728 4888 21732
rect 11848 21788 11912 21792
rect 11848 21732 11852 21788
rect 11852 21732 11908 21788
rect 11908 21732 11912 21788
rect 11848 21728 11912 21732
rect 11928 21788 11992 21792
rect 11928 21732 11932 21788
rect 11932 21732 11988 21788
rect 11988 21732 11992 21788
rect 11928 21728 11992 21732
rect 12008 21788 12072 21792
rect 12008 21732 12012 21788
rect 12012 21732 12068 21788
rect 12068 21732 12072 21788
rect 12008 21728 12072 21732
rect 12088 21788 12152 21792
rect 12088 21732 12092 21788
rect 12092 21732 12148 21788
rect 12148 21732 12152 21788
rect 12088 21728 12152 21732
rect 19112 21788 19176 21792
rect 19112 21732 19116 21788
rect 19116 21732 19172 21788
rect 19172 21732 19176 21788
rect 19112 21728 19176 21732
rect 19192 21788 19256 21792
rect 19192 21732 19196 21788
rect 19196 21732 19252 21788
rect 19252 21732 19256 21788
rect 19192 21728 19256 21732
rect 19272 21788 19336 21792
rect 19272 21732 19276 21788
rect 19276 21732 19332 21788
rect 19332 21732 19336 21788
rect 19272 21728 19336 21732
rect 19352 21788 19416 21792
rect 19352 21732 19356 21788
rect 19356 21732 19412 21788
rect 19412 21732 19416 21788
rect 19352 21728 19416 21732
rect 8216 21244 8280 21248
rect 8216 21188 8220 21244
rect 8220 21188 8276 21244
rect 8276 21188 8280 21244
rect 8216 21184 8280 21188
rect 8296 21244 8360 21248
rect 8296 21188 8300 21244
rect 8300 21188 8356 21244
rect 8356 21188 8360 21244
rect 8296 21184 8360 21188
rect 8376 21244 8440 21248
rect 8376 21188 8380 21244
rect 8380 21188 8436 21244
rect 8436 21188 8440 21244
rect 8376 21184 8440 21188
rect 8456 21244 8520 21248
rect 8456 21188 8460 21244
rect 8460 21188 8516 21244
rect 8516 21188 8520 21244
rect 8456 21184 8520 21188
rect 15480 21244 15544 21248
rect 15480 21188 15484 21244
rect 15484 21188 15540 21244
rect 15540 21188 15544 21244
rect 15480 21184 15544 21188
rect 15560 21244 15624 21248
rect 15560 21188 15564 21244
rect 15564 21188 15620 21244
rect 15620 21188 15624 21244
rect 15560 21184 15624 21188
rect 15640 21244 15704 21248
rect 15640 21188 15644 21244
rect 15644 21188 15700 21244
rect 15700 21188 15704 21244
rect 15640 21184 15704 21188
rect 15720 21244 15784 21248
rect 15720 21188 15724 21244
rect 15724 21188 15780 21244
rect 15780 21188 15784 21244
rect 15720 21184 15784 21188
rect 21036 20768 21100 20772
rect 21036 20712 21050 20768
rect 21050 20712 21100 20768
rect 21036 20708 21100 20712
rect 4584 20700 4648 20704
rect 4584 20644 4588 20700
rect 4588 20644 4644 20700
rect 4644 20644 4648 20700
rect 4584 20640 4648 20644
rect 4664 20700 4728 20704
rect 4664 20644 4668 20700
rect 4668 20644 4724 20700
rect 4724 20644 4728 20700
rect 4664 20640 4728 20644
rect 4744 20700 4808 20704
rect 4744 20644 4748 20700
rect 4748 20644 4804 20700
rect 4804 20644 4808 20700
rect 4744 20640 4808 20644
rect 4824 20700 4888 20704
rect 4824 20644 4828 20700
rect 4828 20644 4884 20700
rect 4884 20644 4888 20700
rect 4824 20640 4888 20644
rect 11848 20700 11912 20704
rect 11848 20644 11852 20700
rect 11852 20644 11908 20700
rect 11908 20644 11912 20700
rect 11848 20640 11912 20644
rect 11928 20700 11992 20704
rect 11928 20644 11932 20700
rect 11932 20644 11988 20700
rect 11988 20644 11992 20700
rect 11928 20640 11992 20644
rect 12008 20700 12072 20704
rect 12008 20644 12012 20700
rect 12012 20644 12068 20700
rect 12068 20644 12072 20700
rect 12008 20640 12072 20644
rect 12088 20700 12152 20704
rect 12088 20644 12092 20700
rect 12092 20644 12148 20700
rect 12148 20644 12152 20700
rect 12088 20640 12152 20644
rect 19112 20700 19176 20704
rect 19112 20644 19116 20700
rect 19116 20644 19172 20700
rect 19172 20644 19176 20700
rect 19112 20640 19176 20644
rect 19192 20700 19256 20704
rect 19192 20644 19196 20700
rect 19196 20644 19252 20700
rect 19252 20644 19256 20700
rect 19192 20640 19256 20644
rect 19272 20700 19336 20704
rect 19272 20644 19276 20700
rect 19276 20644 19332 20700
rect 19332 20644 19336 20700
rect 19272 20640 19336 20644
rect 19352 20700 19416 20704
rect 19352 20644 19356 20700
rect 19356 20644 19412 20700
rect 19412 20644 19416 20700
rect 19352 20640 19416 20644
rect 8216 20156 8280 20160
rect 8216 20100 8220 20156
rect 8220 20100 8276 20156
rect 8276 20100 8280 20156
rect 8216 20096 8280 20100
rect 8296 20156 8360 20160
rect 8296 20100 8300 20156
rect 8300 20100 8356 20156
rect 8356 20100 8360 20156
rect 8296 20096 8360 20100
rect 8376 20156 8440 20160
rect 8376 20100 8380 20156
rect 8380 20100 8436 20156
rect 8436 20100 8440 20156
rect 8376 20096 8440 20100
rect 8456 20156 8520 20160
rect 8456 20100 8460 20156
rect 8460 20100 8516 20156
rect 8516 20100 8520 20156
rect 8456 20096 8520 20100
rect 15480 20156 15544 20160
rect 15480 20100 15484 20156
rect 15484 20100 15540 20156
rect 15540 20100 15544 20156
rect 15480 20096 15544 20100
rect 15560 20156 15624 20160
rect 15560 20100 15564 20156
rect 15564 20100 15620 20156
rect 15620 20100 15624 20156
rect 15560 20096 15624 20100
rect 15640 20156 15704 20160
rect 15640 20100 15644 20156
rect 15644 20100 15700 20156
rect 15700 20100 15704 20156
rect 15640 20096 15704 20100
rect 15720 20156 15784 20160
rect 15720 20100 15724 20156
rect 15724 20100 15780 20156
rect 15780 20100 15784 20156
rect 15720 20096 15784 20100
rect 4584 19612 4648 19616
rect 4584 19556 4588 19612
rect 4588 19556 4644 19612
rect 4644 19556 4648 19612
rect 4584 19552 4648 19556
rect 4664 19612 4728 19616
rect 4664 19556 4668 19612
rect 4668 19556 4724 19612
rect 4724 19556 4728 19612
rect 4664 19552 4728 19556
rect 4744 19612 4808 19616
rect 4744 19556 4748 19612
rect 4748 19556 4804 19612
rect 4804 19556 4808 19612
rect 4744 19552 4808 19556
rect 4824 19612 4888 19616
rect 4824 19556 4828 19612
rect 4828 19556 4884 19612
rect 4884 19556 4888 19612
rect 4824 19552 4888 19556
rect 11848 19612 11912 19616
rect 11848 19556 11852 19612
rect 11852 19556 11908 19612
rect 11908 19556 11912 19612
rect 11848 19552 11912 19556
rect 11928 19612 11992 19616
rect 11928 19556 11932 19612
rect 11932 19556 11988 19612
rect 11988 19556 11992 19612
rect 11928 19552 11992 19556
rect 12008 19612 12072 19616
rect 12008 19556 12012 19612
rect 12012 19556 12068 19612
rect 12068 19556 12072 19612
rect 12008 19552 12072 19556
rect 12088 19612 12152 19616
rect 12088 19556 12092 19612
rect 12092 19556 12148 19612
rect 12148 19556 12152 19612
rect 12088 19552 12152 19556
rect 19112 19612 19176 19616
rect 19112 19556 19116 19612
rect 19116 19556 19172 19612
rect 19172 19556 19176 19612
rect 19112 19552 19176 19556
rect 19192 19612 19256 19616
rect 19192 19556 19196 19612
rect 19196 19556 19252 19612
rect 19252 19556 19256 19612
rect 19192 19552 19256 19556
rect 19272 19612 19336 19616
rect 19272 19556 19276 19612
rect 19276 19556 19332 19612
rect 19332 19556 19336 19612
rect 19272 19552 19336 19556
rect 19352 19612 19416 19616
rect 19352 19556 19356 19612
rect 19356 19556 19412 19612
rect 19412 19556 19416 19612
rect 19352 19552 19416 19556
rect 4108 19076 4172 19140
rect 8216 19068 8280 19072
rect 8216 19012 8220 19068
rect 8220 19012 8276 19068
rect 8276 19012 8280 19068
rect 8216 19008 8280 19012
rect 8296 19068 8360 19072
rect 8296 19012 8300 19068
rect 8300 19012 8356 19068
rect 8356 19012 8360 19068
rect 8296 19008 8360 19012
rect 8376 19068 8440 19072
rect 8376 19012 8380 19068
rect 8380 19012 8436 19068
rect 8436 19012 8440 19068
rect 8376 19008 8440 19012
rect 8456 19068 8520 19072
rect 8456 19012 8460 19068
rect 8460 19012 8516 19068
rect 8516 19012 8520 19068
rect 8456 19008 8520 19012
rect 15480 19068 15544 19072
rect 15480 19012 15484 19068
rect 15484 19012 15540 19068
rect 15540 19012 15544 19068
rect 15480 19008 15544 19012
rect 15560 19068 15624 19072
rect 15560 19012 15564 19068
rect 15564 19012 15620 19068
rect 15620 19012 15624 19068
rect 15560 19008 15624 19012
rect 15640 19068 15704 19072
rect 15640 19012 15644 19068
rect 15644 19012 15700 19068
rect 15700 19012 15704 19068
rect 15640 19008 15704 19012
rect 15720 19068 15784 19072
rect 15720 19012 15724 19068
rect 15724 19012 15780 19068
rect 15780 19012 15784 19068
rect 15720 19008 15784 19012
rect 4584 18524 4648 18528
rect 4584 18468 4588 18524
rect 4588 18468 4644 18524
rect 4644 18468 4648 18524
rect 4584 18464 4648 18468
rect 4664 18524 4728 18528
rect 4664 18468 4668 18524
rect 4668 18468 4724 18524
rect 4724 18468 4728 18524
rect 4664 18464 4728 18468
rect 4744 18524 4808 18528
rect 4744 18468 4748 18524
rect 4748 18468 4804 18524
rect 4804 18468 4808 18524
rect 4744 18464 4808 18468
rect 4824 18524 4888 18528
rect 4824 18468 4828 18524
rect 4828 18468 4884 18524
rect 4884 18468 4888 18524
rect 4824 18464 4888 18468
rect 11848 18524 11912 18528
rect 11848 18468 11852 18524
rect 11852 18468 11908 18524
rect 11908 18468 11912 18524
rect 11848 18464 11912 18468
rect 11928 18524 11992 18528
rect 11928 18468 11932 18524
rect 11932 18468 11988 18524
rect 11988 18468 11992 18524
rect 11928 18464 11992 18468
rect 12008 18524 12072 18528
rect 12008 18468 12012 18524
rect 12012 18468 12068 18524
rect 12068 18468 12072 18524
rect 12008 18464 12072 18468
rect 12088 18524 12152 18528
rect 12088 18468 12092 18524
rect 12092 18468 12148 18524
rect 12148 18468 12152 18524
rect 12088 18464 12152 18468
rect 19112 18524 19176 18528
rect 19112 18468 19116 18524
rect 19116 18468 19172 18524
rect 19172 18468 19176 18524
rect 19112 18464 19176 18468
rect 19192 18524 19256 18528
rect 19192 18468 19196 18524
rect 19196 18468 19252 18524
rect 19252 18468 19256 18524
rect 19192 18464 19256 18468
rect 19272 18524 19336 18528
rect 19272 18468 19276 18524
rect 19276 18468 19332 18524
rect 19332 18468 19336 18524
rect 19272 18464 19336 18468
rect 19352 18524 19416 18528
rect 19352 18468 19356 18524
rect 19356 18468 19412 18524
rect 19412 18468 19416 18524
rect 19352 18464 19416 18468
rect 12572 18260 12636 18324
rect 8216 17980 8280 17984
rect 8216 17924 8220 17980
rect 8220 17924 8276 17980
rect 8276 17924 8280 17980
rect 8216 17920 8280 17924
rect 8296 17980 8360 17984
rect 8296 17924 8300 17980
rect 8300 17924 8356 17980
rect 8356 17924 8360 17980
rect 8296 17920 8360 17924
rect 8376 17980 8440 17984
rect 8376 17924 8380 17980
rect 8380 17924 8436 17980
rect 8436 17924 8440 17980
rect 8376 17920 8440 17924
rect 8456 17980 8520 17984
rect 8456 17924 8460 17980
rect 8460 17924 8516 17980
rect 8516 17924 8520 17980
rect 8456 17920 8520 17924
rect 15480 17980 15544 17984
rect 15480 17924 15484 17980
rect 15484 17924 15540 17980
rect 15540 17924 15544 17980
rect 15480 17920 15544 17924
rect 15560 17980 15624 17984
rect 15560 17924 15564 17980
rect 15564 17924 15620 17980
rect 15620 17924 15624 17980
rect 15560 17920 15624 17924
rect 15640 17980 15704 17984
rect 15640 17924 15644 17980
rect 15644 17924 15700 17980
rect 15700 17924 15704 17980
rect 15640 17920 15704 17924
rect 15720 17980 15784 17984
rect 15720 17924 15724 17980
rect 15724 17924 15780 17980
rect 15780 17924 15784 17980
rect 15720 17920 15784 17924
rect 7236 17504 7300 17508
rect 7236 17448 7250 17504
rect 7250 17448 7300 17504
rect 7236 17444 7300 17448
rect 4584 17436 4648 17440
rect 4584 17380 4588 17436
rect 4588 17380 4644 17436
rect 4644 17380 4648 17436
rect 4584 17376 4648 17380
rect 4664 17436 4728 17440
rect 4664 17380 4668 17436
rect 4668 17380 4724 17436
rect 4724 17380 4728 17436
rect 4664 17376 4728 17380
rect 4744 17436 4808 17440
rect 4744 17380 4748 17436
rect 4748 17380 4804 17436
rect 4804 17380 4808 17436
rect 4744 17376 4808 17380
rect 4824 17436 4888 17440
rect 4824 17380 4828 17436
rect 4828 17380 4884 17436
rect 4884 17380 4888 17436
rect 4824 17376 4888 17380
rect 11848 17436 11912 17440
rect 11848 17380 11852 17436
rect 11852 17380 11908 17436
rect 11908 17380 11912 17436
rect 11848 17376 11912 17380
rect 11928 17436 11992 17440
rect 11928 17380 11932 17436
rect 11932 17380 11988 17436
rect 11988 17380 11992 17436
rect 11928 17376 11992 17380
rect 12008 17436 12072 17440
rect 12008 17380 12012 17436
rect 12012 17380 12068 17436
rect 12068 17380 12072 17436
rect 12008 17376 12072 17380
rect 12088 17436 12152 17440
rect 12088 17380 12092 17436
rect 12092 17380 12148 17436
rect 12148 17380 12152 17436
rect 12088 17376 12152 17380
rect 19112 17436 19176 17440
rect 19112 17380 19116 17436
rect 19116 17380 19172 17436
rect 19172 17380 19176 17436
rect 19112 17376 19176 17380
rect 19192 17436 19256 17440
rect 19192 17380 19196 17436
rect 19196 17380 19252 17436
rect 19252 17380 19256 17436
rect 19192 17376 19256 17380
rect 19272 17436 19336 17440
rect 19272 17380 19276 17436
rect 19276 17380 19332 17436
rect 19332 17380 19336 17436
rect 19272 17376 19336 17380
rect 19352 17436 19416 17440
rect 19352 17380 19356 17436
rect 19356 17380 19412 17436
rect 19412 17380 19416 17436
rect 19352 17376 19416 17380
rect 19564 17308 19628 17372
rect 8216 16892 8280 16896
rect 8216 16836 8220 16892
rect 8220 16836 8276 16892
rect 8276 16836 8280 16892
rect 8216 16832 8280 16836
rect 8296 16892 8360 16896
rect 8296 16836 8300 16892
rect 8300 16836 8356 16892
rect 8356 16836 8360 16892
rect 8296 16832 8360 16836
rect 8376 16892 8440 16896
rect 8376 16836 8380 16892
rect 8380 16836 8436 16892
rect 8436 16836 8440 16892
rect 8376 16832 8440 16836
rect 8456 16892 8520 16896
rect 8456 16836 8460 16892
rect 8460 16836 8516 16892
rect 8516 16836 8520 16892
rect 8456 16832 8520 16836
rect 15480 16892 15544 16896
rect 15480 16836 15484 16892
rect 15484 16836 15540 16892
rect 15540 16836 15544 16892
rect 15480 16832 15544 16836
rect 15560 16892 15624 16896
rect 15560 16836 15564 16892
rect 15564 16836 15620 16892
rect 15620 16836 15624 16892
rect 15560 16832 15624 16836
rect 15640 16892 15704 16896
rect 15640 16836 15644 16892
rect 15644 16836 15700 16892
rect 15700 16836 15704 16892
rect 15640 16832 15704 16836
rect 15720 16892 15784 16896
rect 15720 16836 15724 16892
rect 15724 16836 15780 16892
rect 15780 16836 15784 16892
rect 15720 16832 15784 16836
rect 4584 16348 4648 16352
rect 4584 16292 4588 16348
rect 4588 16292 4644 16348
rect 4644 16292 4648 16348
rect 4584 16288 4648 16292
rect 4664 16348 4728 16352
rect 4664 16292 4668 16348
rect 4668 16292 4724 16348
rect 4724 16292 4728 16348
rect 4664 16288 4728 16292
rect 4744 16348 4808 16352
rect 4744 16292 4748 16348
rect 4748 16292 4804 16348
rect 4804 16292 4808 16348
rect 4744 16288 4808 16292
rect 4824 16348 4888 16352
rect 4824 16292 4828 16348
rect 4828 16292 4884 16348
rect 4884 16292 4888 16348
rect 4824 16288 4888 16292
rect 11848 16348 11912 16352
rect 11848 16292 11852 16348
rect 11852 16292 11908 16348
rect 11908 16292 11912 16348
rect 11848 16288 11912 16292
rect 11928 16348 11992 16352
rect 11928 16292 11932 16348
rect 11932 16292 11988 16348
rect 11988 16292 11992 16348
rect 11928 16288 11992 16292
rect 12008 16348 12072 16352
rect 12008 16292 12012 16348
rect 12012 16292 12068 16348
rect 12068 16292 12072 16348
rect 12008 16288 12072 16292
rect 12088 16348 12152 16352
rect 12088 16292 12092 16348
rect 12092 16292 12148 16348
rect 12148 16292 12152 16348
rect 12088 16288 12152 16292
rect 19112 16348 19176 16352
rect 19112 16292 19116 16348
rect 19116 16292 19172 16348
rect 19172 16292 19176 16348
rect 19112 16288 19176 16292
rect 19192 16348 19256 16352
rect 19192 16292 19196 16348
rect 19196 16292 19252 16348
rect 19252 16292 19256 16348
rect 19192 16288 19256 16292
rect 19272 16348 19336 16352
rect 19272 16292 19276 16348
rect 19276 16292 19332 16348
rect 19332 16292 19336 16348
rect 19272 16288 19336 16292
rect 19352 16348 19416 16352
rect 19352 16292 19356 16348
rect 19356 16292 19412 16348
rect 19412 16292 19416 16348
rect 19352 16288 19416 16292
rect 15884 16220 15948 16284
rect 8216 15804 8280 15808
rect 8216 15748 8220 15804
rect 8220 15748 8276 15804
rect 8276 15748 8280 15804
rect 8216 15744 8280 15748
rect 8296 15804 8360 15808
rect 8296 15748 8300 15804
rect 8300 15748 8356 15804
rect 8356 15748 8360 15804
rect 8296 15744 8360 15748
rect 8376 15804 8440 15808
rect 8376 15748 8380 15804
rect 8380 15748 8436 15804
rect 8436 15748 8440 15804
rect 8376 15744 8440 15748
rect 8456 15804 8520 15808
rect 8456 15748 8460 15804
rect 8460 15748 8516 15804
rect 8516 15748 8520 15804
rect 8456 15744 8520 15748
rect 15480 15804 15544 15808
rect 15480 15748 15484 15804
rect 15484 15748 15540 15804
rect 15540 15748 15544 15804
rect 15480 15744 15544 15748
rect 15560 15804 15624 15808
rect 15560 15748 15564 15804
rect 15564 15748 15620 15804
rect 15620 15748 15624 15804
rect 15560 15744 15624 15748
rect 15640 15804 15704 15808
rect 15640 15748 15644 15804
rect 15644 15748 15700 15804
rect 15700 15748 15704 15804
rect 15640 15744 15704 15748
rect 15720 15804 15784 15808
rect 15720 15748 15724 15804
rect 15724 15748 15780 15804
rect 15780 15748 15784 15804
rect 15720 15744 15784 15748
rect 4584 15260 4648 15264
rect 4584 15204 4588 15260
rect 4588 15204 4644 15260
rect 4644 15204 4648 15260
rect 4584 15200 4648 15204
rect 4664 15260 4728 15264
rect 4664 15204 4668 15260
rect 4668 15204 4724 15260
rect 4724 15204 4728 15260
rect 4664 15200 4728 15204
rect 4744 15260 4808 15264
rect 4744 15204 4748 15260
rect 4748 15204 4804 15260
rect 4804 15204 4808 15260
rect 4744 15200 4808 15204
rect 4824 15260 4888 15264
rect 4824 15204 4828 15260
rect 4828 15204 4884 15260
rect 4884 15204 4888 15260
rect 4824 15200 4888 15204
rect 11848 15260 11912 15264
rect 11848 15204 11852 15260
rect 11852 15204 11908 15260
rect 11908 15204 11912 15260
rect 11848 15200 11912 15204
rect 11928 15260 11992 15264
rect 11928 15204 11932 15260
rect 11932 15204 11988 15260
rect 11988 15204 11992 15260
rect 11928 15200 11992 15204
rect 12008 15260 12072 15264
rect 12008 15204 12012 15260
rect 12012 15204 12068 15260
rect 12068 15204 12072 15260
rect 12008 15200 12072 15204
rect 12088 15260 12152 15264
rect 12088 15204 12092 15260
rect 12092 15204 12148 15260
rect 12148 15204 12152 15260
rect 12088 15200 12152 15204
rect 19112 15260 19176 15264
rect 19112 15204 19116 15260
rect 19116 15204 19172 15260
rect 19172 15204 19176 15260
rect 19112 15200 19176 15204
rect 19192 15260 19256 15264
rect 19192 15204 19196 15260
rect 19196 15204 19252 15260
rect 19252 15204 19256 15260
rect 19192 15200 19256 15204
rect 19272 15260 19336 15264
rect 19272 15204 19276 15260
rect 19276 15204 19332 15260
rect 19332 15204 19336 15260
rect 19272 15200 19336 15204
rect 19352 15260 19416 15264
rect 19352 15204 19356 15260
rect 19356 15204 19412 15260
rect 19412 15204 19416 15260
rect 19352 15200 19416 15204
rect 8216 14716 8280 14720
rect 8216 14660 8220 14716
rect 8220 14660 8276 14716
rect 8276 14660 8280 14716
rect 8216 14656 8280 14660
rect 8296 14716 8360 14720
rect 8296 14660 8300 14716
rect 8300 14660 8356 14716
rect 8356 14660 8360 14716
rect 8296 14656 8360 14660
rect 8376 14716 8440 14720
rect 8376 14660 8380 14716
rect 8380 14660 8436 14716
rect 8436 14660 8440 14716
rect 8376 14656 8440 14660
rect 8456 14716 8520 14720
rect 8456 14660 8460 14716
rect 8460 14660 8516 14716
rect 8516 14660 8520 14716
rect 8456 14656 8520 14660
rect 15480 14716 15544 14720
rect 15480 14660 15484 14716
rect 15484 14660 15540 14716
rect 15540 14660 15544 14716
rect 15480 14656 15544 14660
rect 15560 14716 15624 14720
rect 15560 14660 15564 14716
rect 15564 14660 15620 14716
rect 15620 14660 15624 14716
rect 15560 14656 15624 14660
rect 15640 14716 15704 14720
rect 15640 14660 15644 14716
rect 15644 14660 15700 14716
rect 15700 14660 15704 14716
rect 15640 14656 15704 14660
rect 15720 14716 15784 14720
rect 15720 14660 15724 14716
rect 15724 14660 15780 14716
rect 15780 14660 15784 14716
rect 15720 14656 15784 14660
rect 11468 14452 11532 14516
rect 4584 14172 4648 14176
rect 4584 14116 4588 14172
rect 4588 14116 4644 14172
rect 4644 14116 4648 14172
rect 4584 14112 4648 14116
rect 4664 14172 4728 14176
rect 4664 14116 4668 14172
rect 4668 14116 4724 14172
rect 4724 14116 4728 14172
rect 4664 14112 4728 14116
rect 4744 14172 4808 14176
rect 4744 14116 4748 14172
rect 4748 14116 4804 14172
rect 4804 14116 4808 14172
rect 4744 14112 4808 14116
rect 4824 14172 4888 14176
rect 4824 14116 4828 14172
rect 4828 14116 4884 14172
rect 4884 14116 4888 14172
rect 4824 14112 4888 14116
rect 11848 14172 11912 14176
rect 11848 14116 11852 14172
rect 11852 14116 11908 14172
rect 11908 14116 11912 14172
rect 11848 14112 11912 14116
rect 11928 14172 11992 14176
rect 11928 14116 11932 14172
rect 11932 14116 11988 14172
rect 11988 14116 11992 14172
rect 11928 14112 11992 14116
rect 12008 14172 12072 14176
rect 12008 14116 12012 14172
rect 12012 14116 12068 14172
rect 12068 14116 12072 14172
rect 12008 14112 12072 14116
rect 12088 14172 12152 14176
rect 12088 14116 12092 14172
rect 12092 14116 12148 14172
rect 12148 14116 12152 14172
rect 12088 14112 12152 14116
rect 19112 14172 19176 14176
rect 19112 14116 19116 14172
rect 19116 14116 19172 14172
rect 19172 14116 19176 14172
rect 19112 14112 19176 14116
rect 19192 14172 19256 14176
rect 19192 14116 19196 14172
rect 19196 14116 19252 14172
rect 19252 14116 19256 14172
rect 19192 14112 19256 14116
rect 19272 14172 19336 14176
rect 19272 14116 19276 14172
rect 19276 14116 19332 14172
rect 19332 14116 19336 14172
rect 19272 14112 19336 14116
rect 19352 14172 19416 14176
rect 19352 14116 19356 14172
rect 19356 14116 19412 14172
rect 19412 14116 19416 14172
rect 19352 14112 19416 14116
rect 8216 13628 8280 13632
rect 8216 13572 8220 13628
rect 8220 13572 8276 13628
rect 8276 13572 8280 13628
rect 8216 13568 8280 13572
rect 8296 13628 8360 13632
rect 8296 13572 8300 13628
rect 8300 13572 8356 13628
rect 8356 13572 8360 13628
rect 8296 13568 8360 13572
rect 8376 13628 8440 13632
rect 8376 13572 8380 13628
rect 8380 13572 8436 13628
rect 8436 13572 8440 13628
rect 8376 13568 8440 13572
rect 8456 13628 8520 13632
rect 8456 13572 8460 13628
rect 8460 13572 8516 13628
rect 8516 13572 8520 13628
rect 8456 13568 8520 13572
rect 15480 13628 15544 13632
rect 15480 13572 15484 13628
rect 15484 13572 15540 13628
rect 15540 13572 15544 13628
rect 15480 13568 15544 13572
rect 15560 13628 15624 13632
rect 15560 13572 15564 13628
rect 15564 13572 15620 13628
rect 15620 13572 15624 13628
rect 15560 13568 15624 13572
rect 15640 13628 15704 13632
rect 15640 13572 15644 13628
rect 15644 13572 15700 13628
rect 15700 13572 15704 13628
rect 15640 13568 15704 13572
rect 15720 13628 15784 13632
rect 15720 13572 15724 13628
rect 15724 13572 15780 13628
rect 15780 13572 15784 13628
rect 15720 13568 15784 13572
rect 14780 13092 14844 13156
rect 4584 13084 4648 13088
rect 4584 13028 4588 13084
rect 4588 13028 4644 13084
rect 4644 13028 4648 13084
rect 4584 13024 4648 13028
rect 4664 13084 4728 13088
rect 4664 13028 4668 13084
rect 4668 13028 4724 13084
rect 4724 13028 4728 13084
rect 4664 13024 4728 13028
rect 4744 13084 4808 13088
rect 4744 13028 4748 13084
rect 4748 13028 4804 13084
rect 4804 13028 4808 13084
rect 4744 13024 4808 13028
rect 4824 13084 4888 13088
rect 4824 13028 4828 13084
rect 4828 13028 4884 13084
rect 4884 13028 4888 13084
rect 4824 13024 4888 13028
rect 11848 13084 11912 13088
rect 11848 13028 11852 13084
rect 11852 13028 11908 13084
rect 11908 13028 11912 13084
rect 11848 13024 11912 13028
rect 11928 13084 11992 13088
rect 11928 13028 11932 13084
rect 11932 13028 11988 13084
rect 11988 13028 11992 13084
rect 11928 13024 11992 13028
rect 12008 13084 12072 13088
rect 12008 13028 12012 13084
rect 12012 13028 12068 13084
rect 12068 13028 12072 13084
rect 12008 13024 12072 13028
rect 12088 13084 12152 13088
rect 12088 13028 12092 13084
rect 12092 13028 12148 13084
rect 12148 13028 12152 13084
rect 12088 13024 12152 13028
rect 19112 13084 19176 13088
rect 19112 13028 19116 13084
rect 19116 13028 19172 13084
rect 19172 13028 19176 13084
rect 19112 13024 19176 13028
rect 19192 13084 19256 13088
rect 19192 13028 19196 13084
rect 19196 13028 19252 13084
rect 19252 13028 19256 13084
rect 19192 13024 19256 13028
rect 19272 13084 19336 13088
rect 19272 13028 19276 13084
rect 19276 13028 19332 13084
rect 19332 13028 19336 13084
rect 19272 13024 19336 13028
rect 19352 13084 19416 13088
rect 19352 13028 19356 13084
rect 19356 13028 19412 13084
rect 19412 13028 19416 13084
rect 19352 13024 19416 13028
rect 14964 12956 15028 13020
rect 15148 12820 15212 12884
rect 9260 12684 9324 12748
rect 12572 12684 12636 12748
rect 15332 12744 15396 12748
rect 15332 12688 15382 12744
rect 15382 12688 15396 12744
rect 15332 12684 15396 12688
rect 8216 12540 8280 12544
rect 8216 12484 8220 12540
rect 8220 12484 8276 12540
rect 8276 12484 8280 12540
rect 8216 12480 8280 12484
rect 8296 12540 8360 12544
rect 8296 12484 8300 12540
rect 8300 12484 8356 12540
rect 8356 12484 8360 12540
rect 8296 12480 8360 12484
rect 8376 12540 8440 12544
rect 8376 12484 8380 12540
rect 8380 12484 8436 12540
rect 8436 12484 8440 12540
rect 8376 12480 8440 12484
rect 8456 12540 8520 12544
rect 8456 12484 8460 12540
rect 8460 12484 8516 12540
rect 8516 12484 8520 12540
rect 8456 12480 8520 12484
rect 15480 12540 15544 12544
rect 15480 12484 15484 12540
rect 15484 12484 15540 12540
rect 15540 12484 15544 12540
rect 15480 12480 15544 12484
rect 15560 12540 15624 12544
rect 15560 12484 15564 12540
rect 15564 12484 15620 12540
rect 15620 12484 15624 12540
rect 15560 12480 15624 12484
rect 15640 12540 15704 12544
rect 15640 12484 15644 12540
rect 15644 12484 15700 12540
rect 15700 12484 15704 12540
rect 15640 12480 15704 12484
rect 15720 12540 15784 12544
rect 15720 12484 15724 12540
rect 15724 12484 15780 12540
rect 15780 12484 15784 12540
rect 15720 12480 15784 12484
rect 4584 11996 4648 12000
rect 4584 11940 4588 11996
rect 4588 11940 4644 11996
rect 4644 11940 4648 11996
rect 4584 11936 4648 11940
rect 4664 11996 4728 12000
rect 4664 11940 4668 11996
rect 4668 11940 4724 11996
rect 4724 11940 4728 11996
rect 4664 11936 4728 11940
rect 4744 11996 4808 12000
rect 4744 11940 4748 11996
rect 4748 11940 4804 11996
rect 4804 11940 4808 11996
rect 4744 11936 4808 11940
rect 4824 11996 4888 12000
rect 4824 11940 4828 11996
rect 4828 11940 4884 11996
rect 4884 11940 4888 11996
rect 4824 11936 4888 11940
rect 11848 11996 11912 12000
rect 11848 11940 11852 11996
rect 11852 11940 11908 11996
rect 11908 11940 11912 11996
rect 11848 11936 11912 11940
rect 11928 11996 11992 12000
rect 11928 11940 11932 11996
rect 11932 11940 11988 11996
rect 11988 11940 11992 11996
rect 11928 11936 11992 11940
rect 12008 11996 12072 12000
rect 12008 11940 12012 11996
rect 12012 11940 12068 11996
rect 12068 11940 12072 11996
rect 12008 11936 12072 11940
rect 12088 11996 12152 12000
rect 12088 11940 12092 11996
rect 12092 11940 12148 11996
rect 12148 11940 12152 11996
rect 12088 11936 12152 11940
rect 19112 11996 19176 12000
rect 19112 11940 19116 11996
rect 19116 11940 19172 11996
rect 19172 11940 19176 11996
rect 19112 11936 19176 11940
rect 19192 11996 19256 12000
rect 19192 11940 19196 11996
rect 19196 11940 19252 11996
rect 19252 11940 19256 11996
rect 19192 11936 19256 11940
rect 19272 11996 19336 12000
rect 19272 11940 19276 11996
rect 19276 11940 19332 11996
rect 19332 11940 19336 11996
rect 19272 11936 19336 11940
rect 19352 11996 19416 12000
rect 19352 11940 19356 11996
rect 19356 11940 19412 11996
rect 19412 11940 19416 11996
rect 19352 11936 19416 11940
rect 8708 11868 8772 11932
rect 4108 11792 4172 11796
rect 4108 11736 4122 11792
rect 4122 11736 4172 11792
rect 4108 11732 4172 11736
rect 8216 11452 8280 11456
rect 8216 11396 8220 11452
rect 8220 11396 8276 11452
rect 8276 11396 8280 11452
rect 8216 11392 8280 11396
rect 8296 11452 8360 11456
rect 8296 11396 8300 11452
rect 8300 11396 8356 11452
rect 8356 11396 8360 11452
rect 8296 11392 8360 11396
rect 8376 11452 8440 11456
rect 8376 11396 8380 11452
rect 8380 11396 8436 11452
rect 8436 11396 8440 11452
rect 8376 11392 8440 11396
rect 8456 11452 8520 11456
rect 8456 11396 8460 11452
rect 8460 11396 8516 11452
rect 8516 11396 8520 11452
rect 8456 11392 8520 11396
rect 15480 11452 15544 11456
rect 15480 11396 15484 11452
rect 15484 11396 15540 11452
rect 15540 11396 15544 11452
rect 15480 11392 15544 11396
rect 15560 11452 15624 11456
rect 15560 11396 15564 11452
rect 15564 11396 15620 11452
rect 15620 11396 15624 11452
rect 15560 11392 15624 11396
rect 15640 11452 15704 11456
rect 15640 11396 15644 11452
rect 15644 11396 15700 11452
rect 15700 11396 15704 11452
rect 15640 11392 15704 11396
rect 15720 11452 15784 11456
rect 15720 11396 15724 11452
rect 15724 11396 15780 11452
rect 15780 11396 15784 11452
rect 15720 11392 15784 11396
rect 21036 11324 21100 11388
rect 7236 10976 7300 10980
rect 7236 10920 7250 10976
rect 7250 10920 7300 10976
rect 7236 10916 7300 10920
rect 4584 10908 4648 10912
rect 4584 10852 4588 10908
rect 4588 10852 4644 10908
rect 4644 10852 4648 10908
rect 4584 10848 4648 10852
rect 4664 10908 4728 10912
rect 4664 10852 4668 10908
rect 4668 10852 4724 10908
rect 4724 10852 4728 10908
rect 4664 10848 4728 10852
rect 4744 10908 4808 10912
rect 4744 10852 4748 10908
rect 4748 10852 4804 10908
rect 4804 10852 4808 10908
rect 4744 10848 4808 10852
rect 4824 10908 4888 10912
rect 4824 10852 4828 10908
rect 4828 10852 4884 10908
rect 4884 10852 4888 10908
rect 4824 10848 4888 10852
rect 11848 10908 11912 10912
rect 11848 10852 11852 10908
rect 11852 10852 11908 10908
rect 11908 10852 11912 10908
rect 11848 10848 11912 10852
rect 11928 10908 11992 10912
rect 11928 10852 11932 10908
rect 11932 10852 11988 10908
rect 11988 10852 11992 10908
rect 11928 10848 11992 10852
rect 12008 10908 12072 10912
rect 12008 10852 12012 10908
rect 12012 10852 12068 10908
rect 12068 10852 12072 10908
rect 12008 10848 12072 10852
rect 12088 10908 12152 10912
rect 12088 10852 12092 10908
rect 12092 10852 12148 10908
rect 12148 10852 12152 10908
rect 12088 10848 12152 10852
rect 19112 10908 19176 10912
rect 19112 10852 19116 10908
rect 19116 10852 19172 10908
rect 19172 10852 19176 10908
rect 19112 10848 19176 10852
rect 19192 10908 19256 10912
rect 19192 10852 19196 10908
rect 19196 10852 19252 10908
rect 19252 10852 19256 10908
rect 19192 10848 19256 10852
rect 19272 10908 19336 10912
rect 19272 10852 19276 10908
rect 19276 10852 19332 10908
rect 19332 10852 19336 10908
rect 19272 10848 19336 10852
rect 19352 10908 19416 10912
rect 19352 10852 19356 10908
rect 19356 10852 19412 10908
rect 19412 10852 19416 10908
rect 19352 10848 19416 10852
rect 15884 10704 15948 10708
rect 15884 10648 15934 10704
rect 15934 10648 15948 10704
rect 15884 10644 15948 10648
rect 9260 10508 9324 10572
rect 8216 10364 8280 10368
rect 8216 10308 8220 10364
rect 8220 10308 8276 10364
rect 8276 10308 8280 10364
rect 8216 10304 8280 10308
rect 8296 10364 8360 10368
rect 8296 10308 8300 10364
rect 8300 10308 8356 10364
rect 8356 10308 8360 10364
rect 8296 10304 8360 10308
rect 8376 10364 8440 10368
rect 8376 10308 8380 10364
rect 8380 10308 8436 10364
rect 8436 10308 8440 10364
rect 8376 10304 8440 10308
rect 8456 10364 8520 10368
rect 8456 10308 8460 10364
rect 8460 10308 8516 10364
rect 8516 10308 8520 10364
rect 8456 10304 8520 10308
rect 15480 10364 15544 10368
rect 15480 10308 15484 10364
rect 15484 10308 15540 10364
rect 15540 10308 15544 10364
rect 15480 10304 15544 10308
rect 15560 10364 15624 10368
rect 15560 10308 15564 10364
rect 15564 10308 15620 10364
rect 15620 10308 15624 10364
rect 15560 10304 15624 10308
rect 15640 10364 15704 10368
rect 15640 10308 15644 10364
rect 15644 10308 15700 10364
rect 15700 10308 15704 10364
rect 15640 10304 15704 10308
rect 15720 10364 15784 10368
rect 15720 10308 15724 10364
rect 15724 10308 15780 10364
rect 15780 10308 15784 10364
rect 15720 10304 15784 10308
rect 15148 9964 15212 10028
rect 19564 10024 19628 10028
rect 19564 9968 19578 10024
rect 19578 9968 19628 10024
rect 19564 9964 19628 9968
rect 4584 9820 4648 9824
rect 4584 9764 4588 9820
rect 4588 9764 4644 9820
rect 4644 9764 4648 9820
rect 4584 9760 4648 9764
rect 4664 9820 4728 9824
rect 4664 9764 4668 9820
rect 4668 9764 4724 9820
rect 4724 9764 4728 9820
rect 4664 9760 4728 9764
rect 4744 9820 4808 9824
rect 4744 9764 4748 9820
rect 4748 9764 4804 9820
rect 4804 9764 4808 9820
rect 4744 9760 4808 9764
rect 4824 9820 4888 9824
rect 4824 9764 4828 9820
rect 4828 9764 4884 9820
rect 4884 9764 4888 9820
rect 4824 9760 4888 9764
rect 11848 9820 11912 9824
rect 11848 9764 11852 9820
rect 11852 9764 11908 9820
rect 11908 9764 11912 9820
rect 11848 9760 11912 9764
rect 11928 9820 11992 9824
rect 11928 9764 11932 9820
rect 11932 9764 11988 9820
rect 11988 9764 11992 9820
rect 11928 9760 11992 9764
rect 12008 9820 12072 9824
rect 12008 9764 12012 9820
rect 12012 9764 12068 9820
rect 12068 9764 12072 9820
rect 12008 9760 12072 9764
rect 12088 9820 12152 9824
rect 12088 9764 12092 9820
rect 12092 9764 12148 9820
rect 12148 9764 12152 9820
rect 12088 9760 12152 9764
rect 19112 9820 19176 9824
rect 19112 9764 19116 9820
rect 19116 9764 19172 9820
rect 19172 9764 19176 9820
rect 19112 9760 19176 9764
rect 19192 9820 19256 9824
rect 19192 9764 19196 9820
rect 19196 9764 19252 9820
rect 19252 9764 19256 9820
rect 19192 9760 19256 9764
rect 19272 9820 19336 9824
rect 19272 9764 19276 9820
rect 19276 9764 19332 9820
rect 19332 9764 19336 9820
rect 19272 9760 19336 9764
rect 19352 9820 19416 9824
rect 19352 9764 19356 9820
rect 19356 9764 19412 9820
rect 19412 9764 19416 9820
rect 19352 9760 19416 9764
rect 8216 9276 8280 9280
rect 8216 9220 8220 9276
rect 8220 9220 8276 9276
rect 8276 9220 8280 9276
rect 8216 9216 8280 9220
rect 8296 9276 8360 9280
rect 8296 9220 8300 9276
rect 8300 9220 8356 9276
rect 8356 9220 8360 9276
rect 8296 9216 8360 9220
rect 8376 9276 8440 9280
rect 8376 9220 8380 9276
rect 8380 9220 8436 9276
rect 8436 9220 8440 9276
rect 8376 9216 8440 9220
rect 8456 9276 8520 9280
rect 8456 9220 8460 9276
rect 8460 9220 8516 9276
rect 8516 9220 8520 9276
rect 8456 9216 8520 9220
rect 15480 9276 15544 9280
rect 15480 9220 15484 9276
rect 15484 9220 15540 9276
rect 15540 9220 15544 9276
rect 15480 9216 15544 9220
rect 15560 9276 15624 9280
rect 15560 9220 15564 9276
rect 15564 9220 15620 9276
rect 15620 9220 15624 9276
rect 15560 9216 15624 9220
rect 15640 9276 15704 9280
rect 15640 9220 15644 9276
rect 15644 9220 15700 9276
rect 15700 9220 15704 9276
rect 15640 9216 15704 9220
rect 15720 9276 15784 9280
rect 15720 9220 15724 9276
rect 15724 9220 15780 9276
rect 15780 9220 15784 9276
rect 15720 9216 15784 9220
rect 8708 8876 8772 8940
rect 4584 8732 4648 8736
rect 4584 8676 4588 8732
rect 4588 8676 4644 8732
rect 4644 8676 4648 8732
rect 4584 8672 4648 8676
rect 4664 8732 4728 8736
rect 4664 8676 4668 8732
rect 4668 8676 4724 8732
rect 4724 8676 4728 8732
rect 4664 8672 4728 8676
rect 4744 8732 4808 8736
rect 4744 8676 4748 8732
rect 4748 8676 4804 8732
rect 4804 8676 4808 8732
rect 4744 8672 4808 8676
rect 4824 8732 4888 8736
rect 4824 8676 4828 8732
rect 4828 8676 4884 8732
rect 4884 8676 4888 8732
rect 4824 8672 4888 8676
rect 11848 8732 11912 8736
rect 11848 8676 11852 8732
rect 11852 8676 11908 8732
rect 11908 8676 11912 8732
rect 11848 8672 11912 8676
rect 11928 8732 11992 8736
rect 11928 8676 11932 8732
rect 11932 8676 11988 8732
rect 11988 8676 11992 8732
rect 11928 8672 11992 8676
rect 12008 8732 12072 8736
rect 12008 8676 12012 8732
rect 12012 8676 12068 8732
rect 12068 8676 12072 8732
rect 12008 8672 12072 8676
rect 12088 8732 12152 8736
rect 12088 8676 12092 8732
rect 12092 8676 12148 8732
rect 12148 8676 12152 8732
rect 12088 8672 12152 8676
rect 11468 8604 11532 8668
rect 20484 8876 20548 8940
rect 19112 8732 19176 8736
rect 19112 8676 19116 8732
rect 19116 8676 19172 8732
rect 19172 8676 19176 8732
rect 19112 8672 19176 8676
rect 19192 8732 19256 8736
rect 19192 8676 19196 8732
rect 19196 8676 19252 8732
rect 19252 8676 19256 8732
rect 19192 8672 19256 8676
rect 19272 8732 19336 8736
rect 19272 8676 19276 8732
rect 19276 8676 19332 8732
rect 19332 8676 19336 8732
rect 19272 8672 19336 8676
rect 19352 8732 19416 8736
rect 19352 8676 19356 8732
rect 19356 8676 19412 8732
rect 19412 8676 19416 8732
rect 19352 8672 19416 8676
rect 20484 8332 20548 8396
rect 8216 8188 8280 8192
rect 8216 8132 8220 8188
rect 8220 8132 8276 8188
rect 8276 8132 8280 8188
rect 8216 8128 8280 8132
rect 8296 8188 8360 8192
rect 8296 8132 8300 8188
rect 8300 8132 8356 8188
rect 8356 8132 8360 8188
rect 8296 8128 8360 8132
rect 8376 8188 8440 8192
rect 8376 8132 8380 8188
rect 8380 8132 8436 8188
rect 8436 8132 8440 8188
rect 8376 8128 8440 8132
rect 8456 8188 8520 8192
rect 8456 8132 8460 8188
rect 8460 8132 8516 8188
rect 8516 8132 8520 8188
rect 8456 8128 8520 8132
rect 15480 8188 15544 8192
rect 15480 8132 15484 8188
rect 15484 8132 15540 8188
rect 15540 8132 15544 8188
rect 15480 8128 15544 8132
rect 15560 8188 15624 8192
rect 15560 8132 15564 8188
rect 15564 8132 15620 8188
rect 15620 8132 15624 8188
rect 15560 8128 15624 8132
rect 15640 8188 15704 8192
rect 15640 8132 15644 8188
rect 15644 8132 15700 8188
rect 15700 8132 15704 8188
rect 15640 8128 15704 8132
rect 15720 8188 15784 8192
rect 15720 8132 15724 8188
rect 15724 8132 15780 8188
rect 15780 8132 15784 8188
rect 15720 8128 15784 8132
rect 15332 8060 15396 8124
rect 4584 7644 4648 7648
rect 4584 7588 4588 7644
rect 4588 7588 4644 7644
rect 4644 7588 4648 7644
rect 4584 7584 4648 7588
rect 4664 7644 4728 7648
rect 4664 7588 4668 7644
rect 4668 7588 4724 7644
rect 4724 7588 4728 7644
rect 4664 7584 4728 7588
rect 4744 7644 4808 7648
rect 4744 7588 4748 7644
rect 4748 7588 4804 7644
rect 4804 7588 4808 7644
rect 4744 7584 4808 7588
rect 4824 7644 4888 7648
rect 4824 7588 4828 7644
rect 4828 7588 4884 7644
rect 4884 7588 4888 7644
rect 4824 7584 4888 7588
rect 11848 7644 11912 7648
rect 11848 7588 11852 7644
rect 11852 7588 11908 7644
rect 11908 7588 11912 7644
rect 11848 7584 11912 7588
rect 11928 7644 11992 7648
rect 11928 7588 11932 7644
rect 11932 7588 11988 7644
rect 11988 7588 11992 7644
rect 11928 7584 11992 7588
rect 12008 7644 12072 7648
rect 12008 7588 12012 7644
rect 12012 7588 12068 7644
rect 12068 7588 12072 7644
rect 12008 7584 12072 7588
rect 12088 7644 12152 7648
rect 12088 7588 12092 7644
rect 12092 7588 12148 7644
rect 12148 7588 12152 7644
rect 12088 7584 12152 7588
rect 19112 7644 19176 7648
rect 19112 7588 19116 7644
rect 19116 7588 19172 7644
rect 19172 7588 19176 7644
rect 19112 7584 19176 7588
rect 19192 7644 19256 7648
rect 19192 7588 19196 7644
rect 19196 7588 19252 7644
rect 19252 7588 19256 7644
rect 19192 7584 19256 7588
rect 19272 7644 19336 7648
rect 19272 7588 19276 7644
rect 19276 7588 19332 7644
rect 19332 7588 19336 7644
rect 19272 7584 19336 7588
rect 19352 7644 19416 7648
rect 19352 7588 19356 7644
rect 19356 7588 19412 7644
rect 19412 7588 19416 7644
rect 19352 7584 19416 7588
rect 14964 7108 15028 7172
rect 8216 7100 8280 7104
rect 8216 7044 8220 7100
rect 8220 7044 8276 7100
rect 8276 7044 8280 7100
rect 8216 7040 8280 7044
rect 8296 7100 8360 7104
rect 8296 7044 8300 7100
rect 8300 7044 8356 7100
rect 8356 7044 8360 7100
rect 8296 7040 8360 7044
rect 8376 7100 8440 7104
rect 8376 7044 8380 7100
rect 8380 7044 8436 7100
rect 8436 7044 8440 7100
rect 8376 7040 8440 7044
rect 8456 7100 8520 7104
rect 8456 7044 8460 7100
rect 8460 7044 8516 7100
rect 8516 7044 8520 7100
rect 8456 7040 8520 7044
rect 15480 7100 15544 7104
rect 15480 7044 15484 7100
rect 15484 7044 15540 7100
rect 15540 7044 15544 7100
rect 15480 7040 15544 7044
rect 15560 7100 15624 7104
rect 15560 7044 15564 7100
rect 15564 7044 15620 7100
rect 15620 7044 15624 7100
rect 15560 7040 15624 7044
rect 15640 7100 15704 7104
rect 15640 7044 15644 7100
rect 15644 7044 15700 7100
rect 15700 7044 15704 7100
rect 15640 7040 15704 7044
rect 15720 7100 15784 7104
rect 15720 7044 15724 7100
rect 15724 7044 15780 7100
rect 15780 7044 15784 7100
rect 15720 7040 15784 7044
rect 14780 6972 14844 7036
rect 4584 6556 4648 6560
rect 4584 6500 4588 6556
rect 4588 6500 4644 6556
rect 4644 6500 4648 6556
rect 4584 6496 4648 6500
rect 4664 6556 4728 6560
rect 4664 6500 4668 6556
rect 4668 6500 4724 6556
rect 4724 6500 4728 6556
rect 4664 6496 4728 6500
rect 4744 6556 4808 6560
rect 4744 6500 4748 6556
rect 4748 6500 4804 6556
rect 4804 6500 4808 6556
rect 4744 6496 4808 6500
rect 4824 6556 4888 6560
rect 4824 6500 4828 6556
rect 4828 6500 4884 6556
rect 4884 6500 4888 6556
rect 4824 6496 4888 6500
rect 11848 6556 11912 6560
rect 11848 6500 11852 6556
rect 11852 6500 11908 6556
rect 11908 6500 11912 6556
rect 11848 6496 11912 6500
rect 11928 6556 11992 6560
rect 11928 6500 11932 6556
rect 11932 6500 11988 6556
rect 11988 6500 11992 6556
rect 11928 6496 11992 6500
rect 12008 6556 12072 6560
rect 12008 6500 12012 6556
rect 12012 6500 12068 6556
rect 12068 6500 12072 6556
rect 12008 6496 12072 6500
rect 12088 6556 12152 6560
rect 12088 6500 12092 6556
rect 12092 6500 12148 6556
rect 12148 6500 12152 6556
rect 12088 6496 12152 6500
rect 19112 6556 19176 6560
rect 19112 6500 19116 6556
rect 19116 6500 19172 6556
rect 19172 6500 19176 6556
rect 19112 6496 19176 6500
rect 19192 6556 19256 6560
rect 19192 6500 19196 6556
rect 19196 6500 19252 6556
rect 19252 6500 19256 6556
rect 19192 6496 19256 6500
rect 19272 6556 19336 6560
rect 19272 6500 19276 6556
rect 19276 6500 19332 6556
rect 19332 6500 19336 6556
rect 19272 6496 19336 6500
rect 19352 6556 19416 6560
rect 19352 6500 19356 6556
rect 19356 6500 19412 6556
rect 19412 6500 19416 6556
rect 19352 6496 19416 6500
rect 8216 6012 8280 6016
rect 8216 5956 8220 6012
rect 8220 5956 8276 6012
rect 8276 5956 8280 6012
rect 8216 5952 8280 5956
rect 8296 6012 8360 6016
rect 8296 5956 8300 6012
rect 8300 5956 8356 6012
rect 8356 5956 8360 6012
rect 8296 5952 8360 5956
rect 8376 6012 8440 6016
rect 8376 5956 8380 6012
rect 8380 5956 8436 6012
rect 8436 5956 8440 6012
rect 8376 5952 8440 5956
rect 8456 6012 8520 6016
rect 8456 5956 8460 6012
rect 8460 5956 8516 6012
rect 8516 5956 8520 6012
rect 8456 5952 8520 5956
rect 15480 6012 15544 6016
rect 15480 5956 15484 6012
rect 15484 5956 15540 6012
rect 15540 5956 15544 6012
rect 15480 5952 15544 5956
rect 15560 6012 15624 6016
rect 15560 5956 15564 6012
rect 15564 5956 15620 6012
rect 15620 5956 15624 6012
rect 15560 5952 15624 5956
rect 15640 6012 15704 6016
rect 15640 5956 15644 6012
rect 15644 5956 15700 6012
rect 15700 5956 15704 6012
rect 15640 5952 15704 5956
rect 15720 6012 15784 6016
rect 15720 5956 15724 6012
rect 15724 5956 15780 6012
rect 15780 5956 15784 6012
rect 15720 5952 15784 5956
rect 4584 5468 4648 5472
rect 4584 5412 4588 5468
rect 4588 5412 4644 5468
rect 4644 5412 4648 5468
rect 4584 5408 4648 5412
rect 4664 5468 4728 5472
rect 4664 5412 4668 5468
rect 4668 5412 4724 5468
rect 4724 5412 4728 5468
rect 4664 5408 4728 5412
rect 4744 5468 4808 5472
rect 4744 5412 4748 5468
rect 4748 5412 4804 5468
rect 4804 5412 4808 5468
rect 4744 5408 4808 5412
rect 4824 5468 4888 5472
rect 4824 5412 4828 5468
rect 4828 5412 4884 5468
rect 4884 5412 4888 5468
rect 4824 5408 4888 5412
rect 11848 5468 11912 5472
rect 11848 5412 11852 5468
rect 11852 5412 11908 5468
rect 11908 5412 11912 5468
rect 11848 5408 11912 5412
rect 11928 5468 11992 5472
rect 11928 5412 11932 5468
rect 11932 5412 11988 5468
rect 11988 5412 11992 5468
rect 11928 5408 11992 5412
rect 12008 5468 12072 5472
rect 12008 5412 12012 5468
rect 12012 5412 12068 5468
rect 12068 5412 12072 5468
rect 12008 5408 12072 5412
rect 12088 5468 12152 5472
rect 12088 5412 12092 5468
rect 12092 5412 12148 5468
rect 12148 5412 12152 5468
rect 12088 5408 12152 5412
rect 19112 5468 19176 5472
rect 19112 5412 19116 5468
rect 19116 5412 19172 5468
rect 19172 5412 19176 5468
rect 19112 5408 19176 5412
rect 19192 5468 19256 5472
rect 19192 5412 19196 5468
rect 19196 5412 19252 5468
rect 19252 5412 19256 5468
rect 19192 5408 19256 5412
rect 19272 5468 19336 5472
rect 19272 5412 19276 5468
rect 19276 5412 19332 5468
rect 19332 5412 19336 5468
rect 19272 5408 19336 5412
rect 19352 5468 19416 5472
rect 19352 5412 19356 5468
rect 19356 5412 19412 5468
rect 19412 5412 19416 5468
rect 19352 5408 19416 5412
rect 8216 4924 8280 4928
rect 8216 4868 8220 4924
rect 8220 4868 8276 4924
rect 8276 4868 8280 4924
rect 8216 4864 8280 4868
rect 8296 4924 8360 4928
rect 8296 4868 8300 4924
rect 8300 4868 8356 4924
rect 8356 4868 8360 4924
rect 8296 4864 8360 4868
rect 8376 4924 8440 4928
rect 8376 4868 8380 4924
rect 8380 4868 8436 4924
rect 8436 4868 8440 4924
rect 8376 4864 8440 4868
rect 8456 4924 8520 4928
rect 8456 4868 8460 4924
rect 8460 4868 8516 4924
rect 8516 4868 8520 4924
rect 8456 4864 8520 4868
rect 15480 4924 15544 4928
rect 15480 4868 15484 4924
rect 15484 4868 15540 4924
rect 15540 4868 15544 4924
rect 15480 4864 15544 4868
rect 15560 4924 15624 4928
rect 15560 4868 15564 4924
rect 15564 4868 15620 4924
rect 15620 4868 15624 4924
rect 15560 4864 15624 4868
rect 15640 4924 15704 4928
rect 15640 4868 15644 4924
rect 15644 4868 15700 4924
rect 15700 4868 15704 4924
rect 15640 4864 15704 4868
rect 15720 4924 15784 4928
rect 15720 4868 15724 4924
rect 15724 4868 15780 4924
rect 15780 4868 15784 4924
rect 15720 4864 15784 4868
rect 4584 4380 4648 4384
rect 4584 4324 4588 4380
rect 4588 4324 4644 4380
rect 4644 4324 4648 4380
rect 4584 4320 4648 4324
rect 4664 4380 4728 4384
rect 4664 4324 4668 4380
rect 4668 4324 4724 4380
rect 4724 4324 4728 4380
rect 4664 4320 4728 4324
rect 4744 4380 4808 4384
rect 4744 4324 4748 4380
rect 4748 4324 4804 4380
rect 4804 4324 4808 4380
rect 4744 4320 4808 4324
rect 4824 4380 4888 4384
rect 4824 4324 4828 4380
rect 4828 4324 4884 4380
rect 4884 4324 4888 4380
rect 4824 4320 4888 4324
rect 11848 4380 11912 4384
rect 11848 4324 11852 4380
rect 11852 4324 11908 4380
rect 11908 4324 11912 4380
rect 11848 4320 11912 4324
rect 11928 4380 11992 4384
rect 11928 4324 11932 4380
rect 11932 4324 11988 4380
rect 11988 4324 11992 4380
rect 11928 4320 11992 4324
rect 12008 4380 12072 4384
rect 12008 4324 12012 4380
rect 12012 4324 12068 4380
rect 12068 4324 12072 4380
rect 12008 4320 12072 4324
rect 12088 4380 12152 4384
rect 12088 4324 12092 4380
rect 12092 4324 12148 4380
rect 12148 4324 12152 4380
rect 12088 4320 12152 4324
rect 19112 4380 19176 4384
rect 19112 4324 19116 4380
rect 19116 4324 19172 4380
rect 19172 4324 19176 4380
rect 19112 4320 19176 4324
rect 19192 4380 19256 4384
rect 19192 4324 19196 4380
rect 19196 4324 19252 4380
rect 19252 4324 19256 4380
rect 19192 4320 19256 4324
rect 19272 4380 19336 4384
rect 19272 4324 19276 4380
rect 19276 4324 19332 4380
rect 19332 4324 19336 4380
rect 19272 4320 19336 4324
rect 19352 4380 19416 4384
rect 19352 4324 19356 4380
rect 19356 4324 19412 4380
rect 19412 4324 19416 4380
rect 19352 4320 19416 4324
rect 8216 3836 8280 3840
rect 8216 3780 8220 3836
rect 8220 3780 8276 3836
rect 8276 3780 8280 3836
rect 8216 3776 8280 3780
rect 8296 3836 8360 3840
rect 8296 3780 8300 3836
rect 8300 3780 8356 3836
rect 8356 3780 8360 3836
rect 8296 3776 8360 3780
rect 8376 3836 8440 3840
rect 8376 3780 8380 3836
rect 8380 3780 8436 3836
rect 8436 3780 8440 3836
rect 8376 3776 8440 3780
rect 8456 3836 8520 3840
rect 8456 3780 8460 3836
rect 8460 3780 8516 3836
rect 8516 3780 8520 3836
rect 8456 3776 8520 3780
rect 15480 3836 15544 3840
rect 15480 3780 15484 3836
rect 15484 3780 15540 3836
rect 15540 3780 15544 3836
rect 15480 3776 15544 3780
rect 15560 3836 15624 3840
rect 15560 3780 15564 3836
rect 15564 3780 15620 3836
rect 15620 3780 15624 3836
rect 15560 3776 15624 3780
rect 15640 3836 15704 3840
rect 15640 3780 15644 3836
rect 15644 3780 15700 3836
rect 15700 3780 15704 3836
rect 15640 3776 15704 3780
rect 15720 3836 15784 3840
rect 15720 3780 15724 3836
rect 15724 3780 15780 3836
rect 15780 3780 15784 3836
rect 15720 3776 15784 3780
rect 4584 3292 4648 3296
rect 4584 3236 4588 3292
rect 4588 3236 4644 3292
rect 4644 3236 4648 3292
rect 4584 3232 4648 3236
rect 4664 3292 4728 3296
rect 4664 3236 4668 3292
rect 4668 3236 4724 3292
rect 4724 3236 4728 3292
rect 4664 3232 4728 3236
rect 4744 3292 4808 3296
rect 4744 3236 4748 3292
rect 4748 3236 4804 3292
rect 4804 3236 4808 3292
rect 4744 3232 4808 3236
rect 4824 3292 4888 3296
rect 4824 3236 4828 3292
rect 4828 3236 4884 3292
rect 4884 3236 4888 3292
rect 4824 3232 4888 3236
rect 11848 3292 11912 3296
rect 11848 3236 11852 3292
rect 11852 3236 11908 3292
rect 11908 3236 11912 3292
rect 11848 3232 11912 3236
rect 11928 3292 11992 3296
rect 11928 3236 11932 3292
rect 11932 3236 11988 3292
rect 11988 3236 11992 3292
rect 11928 3232 11992 3236
rect 12008 3292 12072 3296
rect 12008 3236 12012 3292
rect 12012 3236 12068 3292
rect 12068 3236 12072 3292
rect 12008 3232 12072 3236
rect 12088 3292 12152 3296
rect 12088 3236 12092 3292
rect 12092 3236 12148 3292
rect 12148 3236 12152 3292
rect 12088 3232 12152 3236
rect 19112 3292 19176 3296
rect 19112 3236 19116 3292
rect 19116 3236 19172 3292
rect 19172 3236 19176 3292
rect 19112 3232 19176 3236
rect 19192 3292 19256 3296
rect 19192 3236 19196 3292
rect 19196 3236 19252 3292
rect 19252 3236 19256 3292
rect 19192 3232 19256 3236
rect 19272 3292 19336 3296
rect 19272 3236 19276 3292
rect 19276 3236 19332 3292
rect 19332 3236 19336 3292
rect 19272 3232 19336 3236
rect 19352 3292 19416 3296
rect 19352 3236 19356 3292
rect 19356 3236 19412 3292
rect 19412 3236 19416 3292
rect 19352 3232 19416 3236
rect 8216 2748 8280 2752
rect 8216 2692 8220 2748
rect 8220 2692 8276 2748
rect 8276 2692 8280 2748
rect 8216 2688 8280 2692
rect 8296 2748 8360 2752
rect 8296 2692 8300 2748
rect 8300 2692 8356 2748
rect 8356 2692 8360 2748
rect 8296 2688 8360 2692
rect 8376 2748 8440 2752
rect 8376 2692 8380 2748
rect 8380 2692 8436 2748
rect 8436 2692 8440 2748
rect 8376 2688 8440 2692
rect 8456 2748 8520 2752
rect 8456 2692 8460 2748
rect 8460 2692 8516 2748
rect 8516 2692 8520 2748
rect 8456 2688 8520 2692
rect 15480 2748 15544 2752
rect 15480 2692 15484 2748
rect 15484 2692 15540 2748
rect 15540 2692 15544 2748
rect 15480 2688 15544 2692
rect 15560 2748 15624 2752
rect 15560 2692 15564 2748
rect 15564 2692 15620 2748
rect 15620 2692 15624 2748
rect 15560 2688 15624 2692
rect 15640 2748 15704 2752
rect 15640 2692 15644 2748
rect 15644 2692 15700 2748
rect 15700 2692 15704 2748
rect 15640 2688 15704 2692
rect 15720 2748 15784 2752
rect 15720 2692 15724 2748
rect 15724 2692 15780 2748
rect 15780 2692 15784 2748
rect 15720 2688 15784 2692
rect 4584 2204 4648 2208
rect 4584 2148 4588 2204
rect 4588 2148 4644 2204
rect 4644 2148 4648 2204
rect 4584 2144 4648 2148
rect 4664 2204 4728 2208
rect 4664 2148 4668 2204
rect 4668 2148 4724 2204
rect 4724 2148 4728 2204
rect 4664 2144 4728 2148
rect 4744 2204 4808 2208
rect 4744 2148 4748 2204
rect 4748 2148 4804 2204
rect 4804 2148 4808 2204
rect 4744 2144 4808 2148
rect 4824 2204 4888 2208
rect 4824 2148 4828 2204
rect 4828 2148 4884 2204
rect 4884 2148 4888 2204
rect 4824 2144 4888 2148
rect 11848 2204 11912 2208
rect 11848 2148 11852 2204
rect 11852 2148 11908 2204
rect 11908 2148 11912 2204
rect 11848 2144 11912 2148
rect 11928 2204 11992 2208
rect 11928 2148 11932 2204
rect 11932 2148 11988 2204
rect 11988 2148 11992 2204
rect 11928 2144 11992 2148
rect 12008 2204 12072 2208
rect 12008 2148 12012 2204
rect 12012 2148 12068 2204
rect 12068 2148 12072 2204
rect 12008 2144 12072 2148
rect 12088 2204 12152 2208
rect 12088 2148 12092 2204
rect 12092 2148 12148 2204
rect 12148 2148 12152 2204
rect 12088 2144 12152 2148
rect 19112 2204 19176 2208
rect 19112 2148 19116 2204
rect 19116 2148 19172 2204
rect 19172 2148 19176 2204
rect 19112 2144 19176 2148
rect 19192 2204 19256 2208
rect 19192 2148 19196 2204
rect 19196 2148 19252 2204
rect 19252 2148 19256 2204
rect 19192 2144 19256 2148
rect 19272 2204 19336 2208
rect 19272 2148 19276 2204
rect 19276 2148 19332 2204
rect 19332 2148 19336 2204
rect 19272 2144 19336 2148
rect 19352 2204 19416 2208
rect 19352 2148 19356 2204
rect 19356 2148 19412 2204
rect 19412 2148 19416 2204
rect 19352 2144 19416 2148
rect 20484 1668 20548 1732
<< metal4 >>
rect 4576 21792 4896 21808
rect 4576 21728 4584 21792
rect 4648 21728 4664 21792
rect 4728 21728 4744 21792
rect 4808 21728 4824 21792
rect 4888 21728 4896 21792
rect 4576 20704 4896 21728
rect 4576 20640 4584 20704
rect 4648 20640 4664 20704
rect 4728 20640 4744 20704
rect 4808 20640 4824 20704
rect 4888 20640 4896 20704
rect 4576 19616 4896 20640
rect 4576 19552 4584 19616
rect 4648 19552 4664 19616
rect 4728 19552 4744 19616
rect 4808 19552 4824 19616
rect 4888 19552 4896 19616
rect 4107 19140 4173 19141
rect 4107 19076 4108 19140
rect 4172 19076 4173 19140
rect 4107 19075 4173 19076
rect 4110 11797 4170 19075
rect 4576 18528 4896 19552
rect 4576 18464 4584 18528
rect 4648 18464 4664 18528
rect 4728 18464 4744 18528
rect 4808 18464 4824 18528
rect 4888 18464 4896 18528
rect 4576 17440 4896 18464
rect 8208 21248 8528 21808
rect 8208 21184 8216 21248
rect 8280 21184 8296 21248
rect 8360 21184 8376 21248
rect 8440 21184 8456 21248
rect 8520 21184 8528 21248
rect 8208 20160 8528 21184
rect 8208 20096 8216 20160
rect 8280 20096 8296 20160
rect 8360 20096 8376 20160
rect 8440 20096 8456 20160
rect 8520 20096 8528 20160
rect 8208 19072 8528 20096
rect 8208 19008 8216 19072
rect 8280 19008 8296 19072
rect 8360 19008 8376 19072
rect 8440 19008 8456 19072
rect 8520 19008 8528 19072
rect 8208 17984 8528 19008
rect 8208 17920 8216 17984
rect 8280 17920 8296 17984
rect 8360 17920 8376 17984
rect 8440 17920 8456 17984
rect 8520 17920 8528 17984
rect 7235 17508 7301 17509
rect 7235 17444 7236 17508
rect 7300 17444 7301 17508
rect 7235 17443 7301 17444
rect 4576 17376 4584 17440
rect 4648 17376 4664 17440
rect 4728 17376 4744 17440
rect 4808 17376 4824 17440
rect 4888 17376 4896 17440
rect 4576 16352 4896 17376
rect 4576 16288 4584 16352
rect 4648 16288 4664 16352
rect 4728 16288 4744 16352
rect 4808 16288 4824 16352
rect 4888 16288 4896 16352
rect 4576 15264 4896 16288
rect 4576 15200 4584 15264
rect 4648 15200 4664 15264
rect 4728 15200 4744 15264
rect 4808 15200 4824 15264
rect 4888 15200 4896 15264
rect 4576 14176 4896 15200
rect 4576 14112 4584 14176
rect 4648 14112 4664 14176
rect 4728 14112 4744 14176
rect 4808 14112 4824 14176
rect 4888 14112 4896 14176
rect 4576 13088 4896 14112
rect 4576 13024 4584 13088
rect 4648 13024 4664 13088
rect 4728 13024 4744 13088
rect 4808 13024 4824 13088
rect 4888 13024 4896 13088
rect 4576 12000 4896 13024
rect 4576 11936 4584 12000
rect 4648 11936 4664 12000
rect 4728 11936 4744 12000
rect 4808 11936 4824 12000
rect 4888 11936 4896 12000
rect 4107 11796 4173 11797
rect 4107 11732 4108 11796
rect 4172 11732 4173 11796
rect 4107 11731 4173 11732
rect 4576 10912 4896 11936
rect 7238 10981 7298 17443
rect 8208 16896 8528 17920
rect 8208 16832 8216 16896
rect 8280 16832 8296 16896
rect 8360 16832 8376 16896
rect 8440 16832 8456 16896
rect 8520 16832 8528 16896
rect 8208 15808 8528 16832
rect 8208 15744 8216 15808
rect 8280 15744 8296 15808
rect 8360 15744 8376 15808
rect 8440 15744 8456 15808
rect 8520 15744 8528 15808
rect 8208 14720 8528 15744
rect 8208 14656 8216 14720
rect 8280 14656 8296 14720
rect 8360 14656 8376 14720
rect 8440 14656 8456 14720
rect 8520 14656 8528 14720
rect 8208 13632 8528 14656
rect 11840 21792 12160 21808
rect 11840 21728 11848 21792
rect 11912 21728 11928 21792
rect 11992 21728 12008 21792
rect 12072 21728 12088 21792
rect 12152 21728 12160 21792
rect 11840 20704 12160 21728
rect 11840 20640 11848 20704
rect 11912 20640 11928 20704
rect 11992 20640 12008 20704
rect 12072 20640 12088 20704
rect 12152 20640 12160 20704
rect 11840 19616 12160 20640
rect 11840 19552 11848 19616
rect 11912 19552 11928 19616
rect 11992 19552 12008 19616
rect 12072 19552 12088 19616
rect 12152 19552 12160 19616
rect 11840 18528 12160 19552
rect 11840 18464 11848 18528
rect 11912 18464 11928 18528
rect 11992 18464 12008 18528
rect 12072 18464 12088 18528
rect 12152 18464 12160 18528
rect 11840 17440 12160 18464
rect 15472 21248 15792 21808
rect 15472 21184 15480 21248
rect 15544 21184 15560 21248
rect 15624 21184 15640 21248
rect 15704 21184 15720 21248
rect 15784 21184 15792 21248
rect 15472 20160 15792 21184
rect 15472 20096 15480 20160
rect 15544 20096 15560 20160
rect 15624 20096 15640 20160
rect 15704 20096 15720 20160
rect 15784 20096 15792 20160
rect 15472 19072 15792 20096
rect 15472 19008 15480 19072
rect 15544 19008 15560 19072
rect 15624 19008 15640 19072
rect 15704 19008 15720 19072
rect 15784 19008 15792 19072
rect 12571 18324 12637 18325
rect 12571 18260 12572 18324
rect 12636 18260 12637 18324
rect 12571 18259 12637 18260
rect 11840 17376 11848 17440
rect 11912 17376 11928 17440
rect 11992 17376 12008 17440
rect 12072 17376 12088 17440
rect 12152 17376 12160 17440
rect 11840 16352 12160 17376
rect 11840 16288 11848 16352
rect 11912 16288 11928 16352
rect 11992 16288 12008 16352
rect 12072 16288 12088 16352
rect 12152 16288 12160 16352
rect 11840 15264 12160 16288
rect 11840 15200 11848 15264
rect 11912 15200 11928 15264
rect 11992 15200 12008 15264
rect 12072 15200 12088 15264
rect 12152 15200 12160 15264
rect 11467 14516 11533 14517
rect 11467 14452 11468 14516
rect 11532 14452 11533 14516
rect 11467 14451 11533 14452
rect 8208 13568 8216 13632
rect 8280 13568 8296 13632
rect 8360 13568 8376 13632
rect 8440 13568 8456 13632
rect 8520 13568 8528 13632
rect 8208 12544 8528 13568
rect 9259 12748 9325 12749
rect 9259 12684 9260 12748
rect 9324 12684 9325 12748
rect 9259 12683 9325 12684
rect 8208 12480 8216 12544
rect 8280 12480 8296 12544
rect 8360 12480 8376 12544
rect 8440 12480 8456 12544
rect 8520 12480 8528 12544
rect 8208 11456 8528 12480
rect 8707 11932 8773 11933
rect 8707 11868 8708 11932
rect 8772 11868 8773 11932
rect 8707 11867 8773 11868
rect 8208 11392 8216 11456
rect 8280 11392 8296 11456
rect 8360 11392 8376 11456
rect 8440 11392 8456 11456
rect 8520 11392 8528 11456
rect 7235 10980 7301 10981
rect 7235 10916 7236 10980
rect 7300 10916 7301 10980
rect 7235 10915 7301 10916
rect 4576 10848 4584 10912
rect 4648 10848 4664 10912
rect 4728 10848 4744 10912
rect 4808 10848 4824 10912
rect 4888 10848 4896 10912
rect 4576 9824 4896 10848
rect 4576 9760 4584 9824
rect 4648 9760 4664 9824
rect 4728 9760 4744 9824
rect 4808 9760 4824 9824
rect 4888 9760 4896 9824
rect 4576 8736 4896 9760
rect 4576 8672 4584 8736
rect 4648 8672 4664 8736
rect 4728 8672 4744 8736
rect 4808 8672 4824 8736
rect 4888 8672 4896 8736
rect 4576 7648 4896 8672
rect 4576 7584 4584 7648
rect 4648 7584 4664 7648
rect 4728 7584 4744 7648
rect 4808 7584 4824 7648
rect 4888 7584 4896 7648
rect 4576 6560 4896 7584
rect 4576 6496 4584 6560
rect 4648 6496 4664 6560
rect 4728 6496 4744 6560
rect 4808 6496 4824 6560
rect 4888 6496 4896 6560
rect 4576 5472 4896 6496
rect 4576 5408 4584 5472
rect 4648 5408 4664 5472
rect 4728 5408 4744 5472
rect 4808 5408 4824 5472
rect 4888 5408 4896 5472
rect 4576 4384 4896 5408
rect 4576 4320 4584 4384
rect 4648 4320 4664 4384
rect 4728 4320 4744 4384
rect 4808 4320 4824 4384
rect 4888 4320 4896 4384
rect 4576 3296 4896 4320
rect 4576 3232 4584 3296
rect 4648 3232 4664 3296
rect 4728 3232 4744 3296
rect 4808 3232 4824 3296
rect 4888 3232 4896 3296
rect 4576 2208 4896 3232
rect 4576 2144 4584 2208
rect 4648 2144 4664 2208
rect 4728 2144 4744 2208
rect 4808 2144 4824 2208
rect 4888 2144 4896 2208
rect 4576 2128 4896 2144
rect 8208 10368 8528 11392
rect 8208 10304 8216 10368
rect 8280 10304 8296 10368
rect 8360 10304 8376 10368
rect 8440 10304 8456 10368
rect 8520 10304 8528 10368
rect 8208 9280 8528 10304
rect 8208 9216 8216 9280
rect 8280 9216 8296 9280
rect 8360 9216 8376 9280
rect 8440 9216 8456 9280
rect 8520 9216 8528 9280
rect 8208 8192 8528 9216
rect 8710 8941 8770 11867
rect 9262 10573 9322 12683
rect 9259 10572 9325 10573
rect 9259 10508 9260 10572
rect 9324 10508 9325 10572
rect 9259 10507 9325 10508
rect 8707 8940 8773 8941
rect 8707 8876 8708 8940
rect 8772 8876 8773 8940
rect 8707 8875 8773 8876
rect 11470 8669 11530 14451
rect 11840 14176 12160 15200
rect 11840 14112 11848 14176
rect 11912 14112 11928 14176
rect 11992 14112 12008 14176
rect 12072 14112 12088 14176
rect 12152 14112 12160 14176
rect 11840 13088 12160 14112
rect 11840 13024 11848 13088
rect 11912 13024 11928 13088
rect 11992 13024 12008 13088
rect 12072 13024 12088 13088
rect 12152 13024 12160 13088
rect 11840 12000 12160 13024
rect 12574 12749 12634 18259
rect 15472 17984 15792 19008
rect 15472 17920 15480 17984
rect 15544 17920 15560 17984
rect 15624 17920 15640 17984
rect 15704 17920 15720 17984
rect 15784 17920 15792 17984
rect 15472 16896 15792 17920
rect 15472 16832 15480 16896
rect 15544 16832 15560 16896
rect 15624 16832 15640 16896
rect 15704 16832 15720 16896
rect 15784 16832 15792 16896
rect 15472 15808 15792 16832
rect 19104 21792 19424 21808
rect 19104 21728 19112 21792
rect 19176 21728 19192 21792
rect 19256 21728 19272 21792
rect 19336 21728 19352 21792
rect 19416 21728 19424 21792
rect 19104 20704 19424 21728
rect 21035 20772 21101 20773
rect 21035 20708 21036 20772
rect 21100 20708 21101 20772
rect 21035 20707 21101 20708
rect 19104 20640 19112 20704
rect 19176 20640 19192 20704
rect 19256 20640 19272 20704
rect 19336 20640 19352 20704
rect 19416 20640 19424 20704
rect 19104 19616 19424 20640
rect 19104 19552 19112 19616
rect 19176 19552 19192 19616
rect 19256 19552 19272 19616
rect 19336 19552 19352 19616
rect 19416 19552 19424 19616
rect 19104 18528 19424 19552
rect 19104 18464 19112 18528
rect 19176 18464 19192 18528
rect 19256 18464 19272 18528
rect 19336 18464 19352 18528
rect 19416 18464 19424 18528
rect 19104 17440 19424 18464
rect 19104 17376 19112 17440
rect 19176 17376 19192 17440
rect 19256 17376 19272 17440
rect 19336 17376 19352 17440
rect 19416 17376 19424 17440
rect 19104 16352 19424 17376
rect 19563 17372 19629 17373
rect 19563 17308 19564 17372
rect 19628 17308 19629 17372
rect 19563 17307 19629 17308
rect 19104 16288 19112 16352
rect 19176 16288 19192 16352
rect 19256 16288 19272 16352
rect 19336 16288 19352 16352
rect 19416 16288 19424 16352
rect 15883 16284 15949 16285
rect 15883 16220 15884 16284
rect 15948 16220 15949 16284
rect 15883 16219 15949 16220
rect 15472 15744 15480 15808
rect 15544 15744 15560 15808
rect 15624 15744 15640 15808
rect 15704 15744 15720 15808
rect 15784 15744 15792 15808
rect 15472 14720 15792 15744
rect 15472 14656 15480 14720
rect 15544 14656 15560 14720
rect 15624 14656 15640 14720
rect 15704 14656 15720 14720
rect 15784 14656 15792 14720
rect 15472 13632 15792 14656
rect 15472 13568 15480 13632
rect 15544 13568 15560 13632
rect 15624 13568 15640 13632
rect 15704 13568 15720 13632
rect 15784 13568 15792 13632
rect 14779 13156 14845 13157
rect 14779 13092 14780 13156
rect 14844 13092 14845 13156
rect 14779 13091 14845 13092
rect 12571 12748 12637 12749
rect 12571 12684 12572 12748
rect 12636 12684 12637 12748
rect 12571 12683 12637 12684
rect 11840 11936 11848 12000
rect 11912 11936 11928 12000
rect 11992 11936 12008 12000
rect 12072 11936 12088 12000
rect 12152 11936 12160 12000
rect 11840 10912 12160 11936
rect 11840 10848 11848 10912
rect 11912 10848 11928 10912
rect 11992 10848 12008 10912
rect 12072 10848 12088 10912
rect 12152 10848 12160 10912
rect 11840 9824 12160 10848
rect 11840 9760 11848 9824
rect 11912 9760 11928 9824
rect 11992 9760 12008 9824
rect 12072 9760 12088 9824
rect 12152 9760 12160 9824
rect 11840 8736 12160 9760
rect 11840 8672 11848 8736
rect 11912 8672 11928 8736
rect 11992 8672 12008 8736
rect 12072 8672 12088 8736
rect 12152 8672 12160 8736
rect 11467 8668 11533 8669
rect 11467 8604 11468 8668
rect 11532 8604 11533 8668
rect 11467 8603 11533 8604
rect 8208 8128 8216 8192
rect 8280 8128 8296 8192
rect 8360 8128 8376 8192
rect 8440 8128 8456 8192
rect 8520 8128 8528 8192
rect 8208 7104 8528 8128
rect 8208 7040 8216 7104
rect 8280 7040 8296 7104
rect 8360 7040 8376 7104
rect 8440 7040 8456 7104
rect 8520 7040 8528 7104
rect 8208 6016 8528 7040
rect 8208 5952 8216 6016
rect 8280 5952 8296 6016
rect 8360 5952 8376 6016
rect 8440 5952 8456 6016
rect 8520 5952 8528 6016
rect 8208 4928 8528 5952
rect 8208 4864 8216 4928
rect 8280 4864 8296 4928
rect 8360 4864 8376 4928
rect 8440 4864 8456 4928
rect 8520 4864 8528 4928
rect 8208 3840 8528 4864
rect 8208 3776 8216 3840
rect 8280 3776 8296 3840
rect 8360 3776 8376 3840
rect 8440 3776 8456 3840
rect 8520 3776 8528 3840
rect 8208 2752 8528 3776
rect 8208 2688 8216 2752
rect 8280 2688 8296 2752
rect 8360 2688 8376 2752
rect 8440 2688 8456 2752
rect 8520 2688 8528 2752
rect 8208 2128 8528 2688
rect 11840 7648 12160 8672
rect 11840 7584 11848 7648
rect 11912 7584 11928 7648
rect 11992 7584 12008 7648
rect 12072 7584 12088 7648
rect 12152 7584 12160 7648
rect 11840 6560 12160 7584
rect 14782 7037 14842 13091
rect 14963 13020 15029 13021
rect 14963 12956 14964 13020
rect 15028 12956 15029 13020
rect 14963 12955 15029 12956
rect 14966 7173 15026 12955
rect 15147 12884 15213 12885
rect 15147 12820 15148 12884
rect 15212 12820 15213 12884
rect 15147 12819 15213 12820
rect 15150 10029 15210 12819
rect 15331 12748 15397 12749
rect 15331 12684 15332 12748
rect 15396 12684 15397 12748
rect 15331 12683 15397 12684
rect 15147 10028 15213 10029
rect 15147 9964 15148 10028
rect 15212 9964 15213 10028
rect 15147 9963 15213 9964
rect 15334 8125 15394 12683
rect 15472 12544 15792 13568
rect 15472 12480 15480 12544
rect 15544 12480 15560 12544
rect 15624 12480 15640 12544
rect 15704 12480 15720 12544
rect 15784 12480 15792 12544
rect 15472 11456 15792 12480
rect 15472 11392 15480 11456
rect 15544 11392 15560 11456
rect 15624 11392 15640 11456
rect 15704 11392 15720 11456
rect 15784 11392 15792 11456
rect 15472 10368 15792 11392
rect 15886 10709 15946 16219
rect 19104 15264 19424 16288
rect 19104 15200 19112 15264
rect 19176 15200 19192 15264
rect 19256 15200 19272 15264
rect 19336 15200 19352 15264
rect 19416 15200 19424 15264
rect 19104 14176 19424 15200
rect 19104 14112 19112 14176
rect 19176 14112 19192 14176
rect 19256 14112 19272 14176
rect 19336 14112 19352 14176
rect 19416 14112 19424 14176
rect 19104 13088 19424 14112
rect 19104 13024 19112 13088
rect 19176 13024 19192 13088
rect 19256 13024 19272 13088
rect 19336 13024 19352 13088
rect 19416 13024 19424 13088
rect 19104 12000 19424 13024
rect 19104 11936 19112 12000
rect 19176 11936 19192 12000
rect 19256 11936 19272 12000
rect 19336 11936 19352 12000
rect 19416 11936 19424 12000
rect 19104 10912 19424 11936
rect 19104 10848 19112 10912
rect 19176 10848 19192 10912
rect 19256 10848 19272 10912
rect 19336 10848 19352 10912
rect 19416 10848 19424 10912
rect 15883 10708 15949 10709
rect 15883 10644 15884 10708
rect 15948 10644 15949 10708
rect 15883 10643 15949 10644
rect 15472 10304 15480 10368
rect 15544 10304 15560 10368
rect 15624 10304 15640 10368
rect 15704 10304 15720 10368
rect 15784 10304 15792 10368
rect 15472 9280 15792 10304
rect 15472 9216 15480 9280
rect 15544 9216 15560 9280
rect 15624 9216 15640 9280
rect 15704 9216 15720 9280
rect 15784 9216 15792 9280
rect 15472 8192 15792 9216
rect 15472 8128 15480 8192
rect 15544 8128 15560 8192
rect 15624 8128 15640 8192
rect 15704 8128 15720 8192
rect 15784 8128 15792 8192
rect 15331 8124 15397 8125
rect 15331 8060 15332 8124
rect 15396 8060 15397 8124
rect 15331 8059 15397 8060
rect 14963 7172 15029 7173
rect 14963 7108 14964 7172
rect 15028 7108 15029 7172
rect 14963 7107 15029 7108
rect 15472 7104 15792 8128
rect 15472 7040 15480 7104
rect 15544 7040 15560 7104
rect 15624 7040 15640 7104
rect 15704 7040 15720 7104
rect 15784 7040 15792 7104
rect 14779 7036 14845 7037
rect 14779 6972 14780 7036
rect 14844 6972 14845 7036
rect 14779 6971 14845 6972
rect 11840 6496 11848 6560
rect 11912 6496 11928 6560
rect 11992 6496 12008 6560
rect 12072 6496 12088 6560
rect 12152 6496 12160 6560
rect 11840 5472 12160 6496
rect 11840 5408 11848 5472
rect 11912 5408 11928 5472
rect 11992 5408 12008 5472
rect 12072 5408 12088 5472
rect 12152 5408 12160 5472
rect 11840 4384 12160 5408
rect 11840 4320 11848 4384
rect 11912 4320 11928 4384
rect 11992 4320 12008 4384
rect 12072 4320 12088 4384
rect 12152 4320 12160 4384
rect 11840 3296 12160 4320
rect 11840 3232 11848 3296
rect 11912 3232 11928 3296
rect 11992 3232 12008 3296
rect 12072 3232 12088 3296
rect 12152 3232 12160 3296
rect 11840 2208 12160 3232
rect 11840 2144 11848 2208
rect 11912 2144 11928 2208
rect 11992 2144 12008 2208
rect 12072 2144 12088 2208
rect 12152 2144 12160 2208
rect 11840 2128 12160 2144
rect 15472 6016 15792 7040
rect 15472 5952 15480 6016
rect 15544 5952 15560 6016
rect 15624 5952 15640 6016
rect 15704 5952 15720 6016
rect 15784 5952 15792 6016
rect 15472 4928 15792 5952
rect 15472 4864 15480 4928
rect 15544 4864 15560 4928
rect 15624 4864 15640 4928
rect 15704 4864 15720 4928
rect 15784 4864 15792 4928
rect 15472 3840 15792 4864
rect 15472 3776 15480 3840
rect 15544 3776 15560 3840
rect 15624 3776 15640 3840
rect 15704 3776 15720 3840
rect 15784 3776 15792 3840
rect 15472 2752 15792 3776
rect 15472 2688 15480 2752
rect 15544 2688 15560 2752
rect 15624 2688 15640 2752
rect 15704 2688 15720 2752
rect 15784 2688 15792 2752
rect 15472 2128 15792 2688
rect 19104 9824 19424 10848
rect 19566 10029 19626 17307
rect 21038 11389 21098 20707
rect 21035 11388 21101 11389
rect 21035 11324 21036 11388
rect 21100 11324 21101 11388
rect 21035 11323 21101 11324
rect 19563 10028 19629 10029
rect 19563 9964 19564 10028
rect 19628 9964 19629 10028
rect 19563 9963 19629 9964
rect 19104 9760 19112 9824
rect 19176 9760 19192 9824
rect 19256 9760 19272 9824
rect 19336 9760 19352 9824
rect 19416 9760 19424 9824
rect 19104 8736 19424 9760
rect 20483 8940 20549 8941
rect 20483 8876 20484 8940
rect 20548 8876 20549 8940
rect 20483 8875 20549 8876
rect 19104 8672 19112 8736
rect 19176 8672 19192 8736
rect 19256 8672 19272 8736
rect 19336 8672 19352 8736
rect 19416 8672 19424 8736
rect 19104 7648 19424 8672
rect 20486 8397 20546 8875
rect 20483 8396 20549 8397
rect 20483 8332 20484 8396
rect 20548 8332 20549 8396
rect 20483 8331 20549 8332
rect 19104 7584 19112 7648
rect 19176 7584 19192 7648
rect 19256 7584 19272 7648
rect 19336 7584 19352 7648
rect 19416 7584 19424 7648
rect 19104 6560 19424 7584
rect 19104 6496 19112 6560
rect 19176 6496 19192 6560
rect 19256 6496 19272 6560
rect 19336 6496 19352 6560
rect 19416 6496 19424 6560
rect 19104 5472 19424 6496
rect 19104 5408 19112 5472
rect 19176 5408 19192 5472
rect 19256 5408 19272 5472
rect 19336 5408 19352 5472
rect 19416 5408 19424 5472
rect 19104 4384 19424 5408
rect 19104 4320 19112 4384
rect 19176 4320 19192 4384
rect 19256 4320 19272 4384
rect 19336 4320 19352 4384
rect 19416 4320 19424 4384
rect 19104 3296 19424 4320
rect 19104 3232 19112 3296
rect 19176 3232 19192 3296
rect 19256 3232 19272 3296
rect 19336 3232 19352 3296
rect 19416 3232 19424 3296
rect 19104 2208 19424 3232
rect 19104 2144 19112 2208
rect 19176 2144 19192 2208
rect 19256 2144 19272 2208
rect 19336 2144 19352 2208
rect 19416 2144 19424 2208
rect 19104 2128 19424 2144
rect 20486 1733 20546 8331
rect 20483 1732 20549 1733
rect 20483 1668 20484 1732
rect 20548 1668 20549 1732
rect 20483 1667 20549 1668
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1605641404
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1605641404
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1605641404
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1605641404
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1605641404
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1605641404
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1605641404
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1605641404
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1605641404
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1605641404
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1605641404
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1605641404
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1605641404
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1605641404
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1605641404
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1605641404
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1605641404
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1605641404
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1605641404
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1605641404
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_119
timestamp 1605641404
transform 1 0 12052 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_114 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_110
timestamp 1605641404
transform 1 0 11224 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1605641404
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _64_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1605641404
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_125
timestamp 1605641404
transform 1 0 12604 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1605641404
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1605641404
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _40_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 12696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _38_
timestamp 1605641404
transform 1 0 12880 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1605641404
transform 1 0 12972 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1605641404
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 13156 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14352 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13340 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 14168 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_0_142
timestamp 1605641404
transform 1 0 14168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1605641404
transform 1 0 13984 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 15456 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 16008 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1605641404
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_153
timestamp 1605641404
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp 1605641404
transform 1 0 16928 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1605641404
transform 1 0 15640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1605641404
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1605641404
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1605641404
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1605641404
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 17204 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1605641404
transform 1 0 18400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1605641404
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 18308 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 18584 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 20056 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 21160 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 20240 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1605641404
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp 1605641404
transform 1 0 19780 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1605641404
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 1605641404
transform 1 0 20056 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 21896 0 1 2720
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1605641404
transform -1 0 22816 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1605641404
transform -1 0 22816 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_227
timestamp 1605641404
transform 1 0 21988 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_224
timestamp 1605641404
transform 1 0 21712 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_231
timestamp 1605641404
transform 1 0 22356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1605641404
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1605641404
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1605641404
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1605641404
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1605641404
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1605641404
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1605641404
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1605641404
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1605641404
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1605641404
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _35_
timestamp 1605641404
transform 1 0 10672 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11132 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1605641404
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_93
timestamp 1605641404
transform 1 0 9660 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_101
timestamp 1605641404
transform 1 0 10396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1605641404
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 12144 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 13156 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1605641404
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_129
timestamp 1605641404
transform 1 0 12972 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_2_140
timestamp 1605641404
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_151
timestamp 1605641404
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 15272 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 16928 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1605641404
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_170
timestamp 1605641404
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 18584 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1605641404
transform 1 0 18400 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 20240 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 20884 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1605641404
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_206
timestamp 1605641404
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_212
timestamp 1605641404
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1605641404
transform -1 0 22816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_231
timestamp 1605641404
transform 1 0 22356 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1605641404
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1605641404
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1605641404
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1605641404
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1605641404
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1605641404
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1605641404
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1605641404
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1605641404
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 9108 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1605641404
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp 1605641404
transform 1 0 9016 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 10212 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_3_96
timestamp 1605641404
transform 1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_108
timestamp 1605641404
transform 1 0 11040 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 12696 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11224 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1605641404
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_119
timestamp 1605641404
transform 1 0 12052 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_123
timestamp 1605641404
transform 1 0 12420 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1605641404
transform 1 0 13064 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 14260 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 13248 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_141
timestamp 1605641404
transform 1 0 14076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 15916 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_159
timestamp 1605641404
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 19044 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 18032 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1605641404
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1605641404
transform 1 0 17388 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_3_193
timestamp 1605641404
transform 1 0 18860 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 20056 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 20700 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_3_204
timestamp 1605641404
transform 1 0 19872 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_210
timestamp 1605641404
transform 1 0 20424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1605641404
transform -1 0 22816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_229
timestamp 1605641404
transform 1 0 22172 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1605641404
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1605641404
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1605641404
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1605641404
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1605641404
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1605641404
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1605641404
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1605641404
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _36_
timestamp 1605641404
transform 1 0 9108 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1605641404
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_80
timestamp 1605641404
transform 1 0 8464 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_86
timestamp 1605641404
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _39_
timestamp 1605641404
transform 1 0 10028 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 10488 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1605641404
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 1605641404
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1605641404
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_100
timestamp 1605641404
transform 1 0 10304 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13156 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 12144 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp 1605641404
transform 1 0 11960 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1605641404
transform 1 0 12972 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_4_140
timestamp 1605641404
transform 1 0 13984 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 1605641404
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16192 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 15640 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1605641404
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_154
timestamp 1605641404
transform 1 0 15272 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_162
timestamp 1605641404
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_173
timestamp 1605641404
transform 1 0 17020 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 17388 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18676 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_4_186
timestamp 1605641404
transform 1 0 18216 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_190
timestamp 1605641404
transform 1 0 18584 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 19688 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 20884 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1605641404
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_200
timestamp 1605641404
transform 1 0 19504 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1605641404
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1605641404
transform -1 0 22816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_231
timestamp 1605641404
transform 1 0 22356 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1605641404
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1605641404
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1605641404
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1605641404
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1605641404
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1605641404
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1605641404
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1605641404
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1605641404
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 8188 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_5_74
timestamp 1605641404
transform 1 0 7912 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _41_
timestamp 1605641404
transform 1 0 10212 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 10672 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1605641404
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_98
timestamp 1605641404
transform 1 0 10120 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_102
timestamp 1605641404
transform 1 0 10488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _42_
timestamp 1605641404
transform 1 0 12420 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12880 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1605641404
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1605641404
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_126
timestamp 1605641404
transform 1 0 12696 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 14720 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_144
timestamp 1605641404
transform 1 0 14352 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1605641404
transform 1 0 15088 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_170
timestamp 1605641404
transform 1 0 16744 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1605641404
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_181
timestamp 1605641404
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19688 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 20884 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 1605641404
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_211
timestamp 1605641404
transform 1 0 20516 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1605641404
transform -1 0 22816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 1605641404
transform 1 0 22356 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1605641404
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1605641404
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1605641404
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1605641404
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1605641404
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1605641404
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1605641404
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1605641404
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1605641404
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1605641404
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1605641404
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1605641404
transform 1 0 5796 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1605641404
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1605641404
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1605641404
transform 1 0 6164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_62
timestamp 1605641404
transform 1 0 6808 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_56
timestamp 1605641404
transform 1 0 6256 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1605641404
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _57_
timestamp 1605641404
transform 1 0 6256 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _37_
timestamp 1605641404
transform 1 0 6808 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1605641404
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 7268 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 8280 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 7912 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_6_72
timestamp 1605641404
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1605641404
transform 1 0 8096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp 1605641404
transform 1 0 9752 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1605641404
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1605641404
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 10028 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 9660 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_101
timestamp 1605641404
transform 1 0 10396 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_106
timestamp 1605641404
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1605641404
transform 1 0 10488 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 10948 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 10580 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 12420 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13064 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12972 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1605641404
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_prog_clk
timestamp 1605641404
transform 1 0 12696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_123
timestamp 1605641404
transform 1 0 12420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1605641404
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_127
timestamp 1605641404
transform 1 0 12788 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14720 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 14628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_145
timestamp 1605641404
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1605641404
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1605641404
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 15732 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 15548 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16284 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16100 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1605641404
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_154
timestamp 1605641404
transform 1 0 15272 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1605641404
transform 1 0 15916 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1605641404
transform 1 0 15548 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_163
timestamp 1605641404
transform 1 0 16100 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 17848 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18400 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18400 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1605641404
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_179
timestamp 1605641404
transform 1 0 17572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_186
timestamp 1605641404
transform 1 0 18216 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_181
timestamp 1605641404
transform 1 0 17756 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_184
timestamp 1605641404
transform 1 0 18032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 20056 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20884 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 20608 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1605641404
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_197
timestamp 1605641404
transform 1 0 19228 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1605641404
transform 1 0 20608 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1605641404
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1605641404
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1605641404
transform -1 0 22816 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1605641404
transform -1 0 22816 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_231
timestamp 1605641404
transform 1 0 22356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_228
timestamp 1605641404
transform 1 0 22080 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_232
timestamp 1605641404
transform 1 0 22448 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1605641404
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1605641404
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1605641404
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1605641404
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1605641404
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1605641404
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _59_
timestamp 1605641404
transform 1 0 5428 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp 1605641404
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_59
timestamp 1605641404
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 7912 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_72
timestamp 1605641404
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10856 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 9660 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1605641404
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1605641404
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_102
timestamp 1605641404
transform 1 0 10488 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 11868 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 12880 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_115
timestamp 1605641404
transform 1 0 11684 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_126
timestamp 1605641404
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13524 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_8_132
timestamp 1605641404
transform 1 0 13248 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1605641404
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 17020 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1605641404
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp 1605641404
transform 1 0 16744 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 19136 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1605641404
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20884 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1605641404
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1605641404
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1605641404
transform -1 0 22816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_231
timestamp 1605641404
transform 1 0 22356 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1605641404
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1605641404
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1605641404
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _61_
timestamp 1605641404
transform 1 0 4232 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_27
timestamp 1605641404
transform 1 0 3588 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1605641404
transform 1 0 4140 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_37
timestamp 1605641404
transform 1 0 4508 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5704 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1605641404
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_48
timestamp 1605641404
transform 1 0 5520 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1605641404
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_62
timestamp 1605641404
transform 1 0 6808 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 8188 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7176 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1605641404
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 9844 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 10948 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_93
timestamp 1605641404
transform 1 0 9660 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_104
timestamp 1605641404
transform 1 0 10672 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1605641404
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_116
timestamp 1605641404
transform 1 0 11776 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 14076 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 13432 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp 1605641404
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp 1605641404
transform 1 0 13800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 16192 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1605641404
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_168
timestamp 1605641404
transform 1 0 16560 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 18676 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 18124 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1605641404
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1605641404
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_184
timestamp 1605641404
transform 1 0 18032 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_189
timestamp 1605641404
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 21160 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_212
timestamp 1605641404
transform 1 0 20608 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1605641404
transform -1 0 22816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_227
timestamp 1605641404
transform 1 0 21988 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1605641404
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1605641404
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_15
timestamp 1605641404
transform 1 0 2484 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _50_
timestamp 1605641404
transform 1 0 4416 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _63_
timestamp 1605641404
transform 1 0 3496 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4876 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1605641404
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1605641404
transform 1 0 4232 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_23
timestamp 1605641404
transform 1 0 3220 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp 1605641404
transform 1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1605641404
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_39
timestamp 1605641404
transform 1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5888 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 6900 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_50
timestamp 1605641404
transform 1 0 5704 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_61
timestamp 1605641404
transform 1 0 6716 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 7912 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1605641404
transform 1 0 7728 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 9660 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1605641404
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 1605641404
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1605641404
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 11316 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 11868 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_115
timestamp 1605641404
transform 1 0 11684 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13524 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_10_133
timestamp 1605641404
transform 1 0 13340 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1605641404
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15364 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 17020 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1605641404
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_154
timestamp 1605641404
transform 1 0 15272 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_171
timestamp 1605641404
transform 1 0 16836 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 18492 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19964 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1605641404
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 21896 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1605641404
transform -1 0 22816 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_224
timestamp 1605641404
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp 1605641404
transform 1 0 22264 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _62_
timestamp 1605641404
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1605641404
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1605641404
transform 1 0 2576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1605641404
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp 1605641404
transform 1 0 2484 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_21
timestamp 1605641404
transform 1 0 3036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _58_
timestamp 1605641404
transform 1 0 3220 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3496 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4692 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1605641404
transform 1 0 4508 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1605641404
transform 1 0 4324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 5704 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 7084 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1605641404
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_48
timestamp 1605641404
transform 1 0 5520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1605641404
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 1605641404
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 8648 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7636 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_69
timestamp 1605641404
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1605641404
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 10304 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_98
timestamp 1605641404
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 12420 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1605641404
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_prog_clk
timestamp 1605641404
transform 1 0 11960 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_116
timestamp 1605641404
transform 1 0 11776 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1605641404
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 15088 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13432 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 1605641404
transform 1 0 13248 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_150
timestamp 1605641404
transform 1 0 14904 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1605641404
transform 1 0 17020 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 17204 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1605641404
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_prog_clk
timestamp 1605641404
transform 1 0 18676 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_179
timestamp 1605641404
transform 1 0 17572 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1605641404
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1605641404
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_194
timestamp 1605641404
transform 1 0 18952 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 20516 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 20884 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19688 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1605641404
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1605641404
transform -1 0 22816 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 1605641404
transform 1 0 22356 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _55_
timestamp 1605641404
transform 1 0 2484 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _60_
timestamp 1605641404
transform 1 0 2024 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2944 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1605641404
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_3
timestamp 1605641404
transform 1 0 1380 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_9
timestamp 1605641404
transform 1 0 1932 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1605641404
transform 1 0 2300 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_18
timestamp 1605641404
transform 1 0 2760 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _49_
timestamp 1605641404
transform 1 0 4048 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 4508 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1605641404
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1605641404
transform 1 0 4324 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1605641404
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 5520 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6532 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_46
timestamp 1605641404
transform 1 0 5336 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1605641404
transform 1 0 6348 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 7544 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1605641404
transform 1 0 7360 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1605641404
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1605641404
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 1605641404
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_109
timestamp 1605641404
transform 1 0 11132 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11408 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 13064 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_12_128
timestamp 1605641404
transform 1 0 12880 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _46_
timestamp 1605641404
transform 1 0 14720 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_146
timestamp 1605641404
transform 1 0 14536 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_151
timestamp 1605641404
transform 1 0 14996 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16376 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1605641404
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_163
timestamp 1605641404
transform 1 0 16100 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 18032 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 18584 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1605641404
transform 1 0 17848 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 1605641404
transform 1 0 18400 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20884 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1605641404
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1605641404
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1605641404
transform -1 0 22816 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_231
timestamp 1605641404
transform 1 0 22356 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1605641404
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1605641404
transform 1 0 1840 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1605641404
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1605641404
transform 1 0 1748 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1605641404
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1605641404
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _56_
timestamp 1605641404
transform 1 0 1564 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _54_
timestamp 1605641404
transform 1 0 1472 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_18
timestamp 1605641404
transform 1 0 2760 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_19
timestamp 1605641404
transform 1 0 2852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2024 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 3036 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 2944 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1605641404
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1605641404
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 1605641404
transform 1 0 3864 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1605641404
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 4048 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_39
timestamp 1605641404
transform 1 0 4692 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_41
timestamp 1605641404
transform 1 0 4876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 4324 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4876 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 5060 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 5888 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1605641404
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1605641404
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1605641404
transform 1 0 6808 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_50
timestamp 1605641404
transform 1 0 5704 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 7544 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7176 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 8188 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_75
timestamp 1605641404
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_86
timestamp 1605641404
transform 1 0 9016 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1605641404
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_86
timestamp 1605641404
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_98
timestamp 1605641404
transform 1 0 10120 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1605641404
transform 1 0 9660 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1605641404
transform 1 0 9476 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 1605641404
transform 1 0 10028 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_prog_clk
timestamp 1605641404
transform 1 0 9200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1605641404
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 9200 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 9752 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 10304 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 10212 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _44_
timestamp 1605641404
transform 1 0 11868 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 13156 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 11960 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1605641404
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1605641404
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1605641404
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_128
timestamp 1605641404
transform 1 0 12880 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_116
timestamp 1605641404
transform 1 0 11776 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 14628 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 13616 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1605641404
transform 1 0 14628 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1605641404
transform 1 0 13432 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_145
timestamp 1605641404
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_151
timestamp 1605641404
transform 1 0 14996 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 17020 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 16928 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16008 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1605641404
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_158
timestamp 1605641404
transform 1 0 15640 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_171
timestamp 1605641404
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_170
timestamp 1605641404
transform 1 0 16744 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_176
timestamp 1605641404
transform 1 0 17296 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_182
timestamp 1605641404
transform 1 0 17848 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_177
timestamp 1605641404
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_prog_clk
timestamp 1605641404
transform 1 0 17572 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1605641404
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 18032 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 17572 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp 1605641404
transform 1 0 18400 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1605641404
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 18584 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 19044 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19596 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 20884 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 21160 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1605641404
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_216
timestamp 1605641404
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_199
timestamp 1605641404
transform 1 0 19412 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_210
timestamp 1605641404
transform 1 0 20424 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1605641404
transform -1 0 22816 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1605641404
transform -1 0 22816 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_227
timestamp 1605641404
transform 1 0 21988 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_231
timestamp 1605641404
transform 1 0 22356 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 2576 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 1564 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1605641404
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1605641404
transform 1 0 1380 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_14
timestamp 1605641404
transform 1 0 2392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _48_
timestamp 1605641404
transform 1 0 4600 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 5060 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_25
timestamp 1605641404
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1605641404
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_41
timestamp 1605641404
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 6900 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1605641404
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1605641404
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_62
timestamp 1605641404
transform 1 0 6808 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 9108 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 7452 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_67
timestamp 1605641404
transform 1 0 7268 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1605641404
transform 1 0 8924 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10948 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_15_103
timestamp 1605641404
transform 1 0 10580 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 12420 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 12972 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1605641404
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_prog_clk
timestamp 1605641404
transform 1 0 11960 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_116
timestamp 1605641404
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_121
timestamp 1605641404
transform 1 0 12236 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1605641404
transform 1 0 12788 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1605641404
transform 1 0 14444 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 1605641404
transform 1 0 14996 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 15548 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_prog_clk
timestamp 1605641404
transform 1 0 15180 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_156
timestamp 1605641404
transform 1 0 15456 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 18032 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1605641404
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_prog_clk
timestamp 1605641404
transform 1 0 17664 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_178
timestamp 1605641404
transform 1 0 17480 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 20148 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20884 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_205
timestamp 1605641404
transform 1 0 19964 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_211
timestamp 1605641404
transform 1 0 20516 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1605641404
transform -1 0 22816 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 1605641404
transform 1 0 22356 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 1380 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1605641404
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1605641404
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 4876 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 4324 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 3404 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1605641404
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1605641404
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1605641404
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_32
timestamp 1605641404
transform 1 0 4048 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_39
timestamp 1605641404
transform 1 0 4692 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 6532 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_57
timestamp 1605641404
transform 1 0 6348 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 7728 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1605641404
transform 1 0 7360 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 9660 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1605641404
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1605641404
transform 1 0 9200 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1605641404
transform 1 0 11132 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 12972 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 11316 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1605641404
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 14812 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 14444 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15364 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1605641404
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1605641404
transform 1 0 15272 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_171
timestamp 1605641404
transform 1 0 16836 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18216 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 17204 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_184
timestamp 1605641404
transform 1 0 18032 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 20148 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 20884 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1605641404
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_prog_clk
timestamp 1605641404
transform 1 0 19872 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_202
timestamp 1605641404
transform 1 0 19688 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_211
timestamp 1605641404
transform 1 0 20516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1605641404
transform -1 0 22816 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_231
timestamp 1605641404
transform 1 0 22356 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 3036 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1380 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1605641404
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_19
timestamp 1605641404
transform 1 0 2852 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 4692 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 4140 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_17_30
timestamp 1605641404
transform 1 0 3864 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_37
timestamp 1605641404
transform 1 0 4508 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 7084 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1605641404
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_prog_clk
timestamp 1605641404
transform 1 0 6348 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_55
timestamp 1605641404
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp 1605641404
transform 1 0 6624 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_62
timestamp 1605641404
transform 1 0 6808 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 7636 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1605641404
transform 1 0 7452 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1605641404
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 9292 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 9844 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_93
timestamp 1605641404
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 11776 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 12420 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1605641404
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_left_width_0_height_0__pin_52_
timestamp 1605641404
transform 1 0 11500 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_111
timestamp 1605641404
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_120
timestamp 1605641404
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 14260 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 13892 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15088 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15916 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1605641404
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1605641404
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1605641404
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 19780 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20332 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_17_200
timestamp 1605641404
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1605641404
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 21988 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1605641404
transform -1 0 22816 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_225
timestamp 1605641404
transform 1 0 21804 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 1605641404
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1380 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1605641404
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_19
timestamp 1605641404
transform 1 0 2852 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 4140 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 4692 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 3404 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1605641404
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_prog_clk
timestamp 1605641404
transform 1 0 3128 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 1605641404
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_32
timestamp 1605641404
transform 1 0 4048 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1605641404
transform 1 0 4508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6348 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_55
timestamp 1605641404
transform 1 0 6164 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 7544 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 8556 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_18_66
timestamp 1605641404
transform 1 0 7176 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1605641404
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1605641404
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1605641404
transform 1 0 11132 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_prog_clk
timestamp 1605641404
transform 1 0 9844 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_prog_clk
timestamp 1605641404
transform 1 0 10672 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1605641404
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_93
timestamp 1605641404
transform 1 0 9660 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_98
timestamp 1605641404
transform 1 0 10120 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_18_107
timestamp 1605641404
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 12972 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 14720 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__decap_3  FILLER_18_145
timestamp 1605641404
transform 1 0 14444 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16192 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1605641404
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_163
timestamp 1605641404
transform 1 0 16100 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 17940 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_18_180
timestamp 1605641404
transform 1 0 17664 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 20884 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1605641404
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_199
timestamp 1605641404
transform 1 0 19412 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1605641404
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1605641404
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 1605641404
transform 1 0 22356 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 1656 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 2116 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 1564 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1605641404
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1605641404
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1605641404
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1605641404
transform 1 0 1380 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_9
timestamp 1605641404
transform 1 0 1932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 3312 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 4324 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 5060 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1605641404
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1605641404
transform 1 0 3128 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_40
timestamp 1605641404
transform 1 0 4784 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1605641404
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_32
timestamp 1605641404
transform 1 0 4048 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 6808 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5336 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1605641404
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1605641404
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_44
timestamp 1605641404
transform 1 0 5152 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_62
timestamp 1605641404
transform 1 0 6808 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 7268 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 7728 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 7820 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_prog_clk
timestamp 1605641404
transform 1 0 7452 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_66
timestamp 1605641404
transform 1 0 7176 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_66
timestamp 1605641404
transform 1 0 7176 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_71
timestamp 1605641404
transform 1 0 7636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 9200 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 9752 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 10764 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 10028 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1605641404
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_89
timestamp 1605641404
transform 1 0 9292 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_93
timestamp 1605641404
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1605641404
transform 1 0 10580 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11500 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 12420 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1605641404
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_left_width_0_height_0__pin_52_
timestamp 1605641404
transform 1 0 11776 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1605641404
transform 1 0 11592 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _45_
timestamp 1605641404
transform 1 0 15088 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 13892 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 14720 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 13616 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1605641404
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15364 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16284 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1605641404
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_prog_clk
timestamp 1605641404
transform 1 0 17112 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_171
timestamp 1605641404
transform 1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1605641404
transform 1 0 16100 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 17388 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 18032 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 17940 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1605641404
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_181
timestamp 1605641404
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_181
timestamp 1605641404
transform 1 0 17756 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 20884 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 20884 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19872 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1605641404
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_200
timestamp 1605641404
transform 1 0 19504 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 1605641404
transform 1 0 20700 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_199
timestamp 1605641404
transform 1 0 19412 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1605641404
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1605641404
transform -1 0 22816 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1605641404
transform -1 0 22816 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_231
timestamp 1605641404
transform 1 0 22356 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_231
timestamp 1605641404
transform 1 0 22356 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2208 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 1656 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1605641404
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1605641404
transform 1 0 1380 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1605641404
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1605641404
transform 1 0 3036 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 3220 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 4876 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_39
timestamp 1605641404
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1605641404
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1605641404
transform 1 0 6348 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 7820 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1605641404
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 9844 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_prog_clk
timestamp 1605641404
transform 1 0 9476 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1605641404
transform 1 0 9292 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_94
timestamp 1605641404
transform 1 0 9752 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 11684 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 12420 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 13156 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1605641404
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_111
timestamp 1605641404
transform 1 0 11316 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_119
timestamp 1605641404
transform 1 0 12052 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_127
timestamp 1605641404
transform 1 0 12788 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14812 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_21_147
timestamp 1605641404
transform 1 0 14628 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _47_
timestamp 1605641404
transform 1 0 16468 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16928 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_165
timestamp 1605641404
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_170
timestamp 1605641404
transform 1 0 16744 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 18032 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1605641404
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1605641404
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 19872 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 20516 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1605641404
transform 1 0 19504 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1605641404
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1605641404
transform -1 0 22816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_227
timestamp 1605641404
transform 1 0 21988 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 2576 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 1564 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1605641404
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1605641404
transform 1 0 1380 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_14
timestamp 1605641404
transform 1 0 2392 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 4048 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1605641404
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_prog_clk
timestamp 1605641404
transform 1 0 3680 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1605641404
transform 1 0 3404 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 6624 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 6072 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_prog_clk
timestamp 1605641404
transform 1 0 5796 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_48
timestamp 1605641404
transform 1 0 5520 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_58
timestamp 1605641404
transform 1 0 6440 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 7636 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 8648 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_69
timestamp 1605641404
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_80
timestamp 1605641404
transform 1 0 8464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_86
timestamp 1605641404
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 9660 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1605641404
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_prog_clk
timestamp 1605641404
transform 1 0 9200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_91
timestamp 1605641404
transform 1 0 9476 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_109
timestamp 1605641404
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 11316 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 12972 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_127
timestamp 1605641404
transform 1 0 12788 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 14628 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1605641404
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1605641404
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 15364 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 16376 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1605641404
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1605641404
transform 1 0 15272 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_164
timestamp 1605641404
transform 1 0 16192 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 19044 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 18032 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_182
timestamp 1605641404
transform 1 0 17848 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1605641404
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 20240 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 20884 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1605641404
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_204
timestamp 1605641404
transform 1 0 19872 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_212
timestamp 1605641404
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1605641404
transform -1 0 22816 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_231
timestamp 1605641404
transform 1 0 22356 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 1472 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1605641404
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 1605641404
transform 1 0 1380 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_20
timestamp 1605641404
transform 1 0 2944 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 3312 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 4324 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_33
timestamp 1605641404
transform 1 0 4140 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 6164 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 7084 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1605641404
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1605641404
transform 1 0 5796 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1605641404
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_62
timestamp 1605641404
transform 1 0 6808 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 8740 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_81
timestamp 1605641404
transform 1 0 8556 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_87
timestamp 1605641404
transform 1 0 9108 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 9292 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 10948 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_23_105
timestamp 1605641404
transform 1 0 10764 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 12420 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1605641404
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_left_width_0_height_0__pin_52_
timestamp 1605641404
transform 1 0 11960 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_116
timestamp 1605641404
transform 1 0 11776 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_121
timestamp 1605641404
transform 1 0 12236 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14444 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_prog_clk
timestamp 1605641404
transform 1 0 14168 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_139
timestamp 1605641404
transform 1 0 13892 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 16284 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_161
timestamp 1605641404
transform 1 0 15916 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 18032 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1605641404
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1605641404
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 19872 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 20884 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1605641404
transform 1 0 19504 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1605641404
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1605641404
transform -1 0 22816 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_231
timestamp 1605641404
transform 1 0 22356 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 1656 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1605641404
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_3
timestamp 1605641404
transform 1 0 1380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _77_
timestamp 1605641404
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 3404 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4784 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1605641404
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_22
timestamp 1605641404
transform 1 0 3128 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1605641404
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_36
timestamp 1605641404
transform 1 0 4416 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 6624 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1605641404
transform 1 0 6256 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_64
timestamp 1605641404
transform 1 0 6992 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 8832 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7176 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1605641404
transform 1 0 8648 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 9660 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1605641404
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_89
timestamp 1605641404
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1605641404
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 11316 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 12512 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_24_120
timestamp 1605641404
transform 1 0 12144 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 14168 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_140
timestamp 1605641404
transform 1 0 13984 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1605641404
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 15272 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 17112 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1605641404
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_170
timestamp 1605641404
transform 1 0 16744 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 18768 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1605641404
transform 1 0 18584 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 20884 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 19780 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1605641404
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1605641404
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_212
timestamp 1605641404
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 21896 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1605641404
transform -1 0 22816 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_224
timestamp 1605641404
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_230
timestamp 1605641404
transform 1 0 22264 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _53_
timestamp 1605641404
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 1840 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1605641404
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_6
timestamp 1605641404
transform 1 0 1656 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 3588 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4600 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_25_24
timestamp 1605641404
transform 1 0 3312 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1605641404
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _52_
timestamp 1605641404
transform 1 0 6256 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1605641404
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1605641404
transform 1 0 6072 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1605641404
transform 1 0 6532 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _34_
timestamp 1605641404
transform 1 0 8832 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1605641404
transform 1 0 7636 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_82
timestamp 1605641404
transform 1 0 8648 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_87
timestamp 1605641404
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 10948 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 9292 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_105
timestamp 1605641404
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 12512 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1605641404
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_prog_clk
timestamp 1605641404
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_116
timestamp 1605641404
transform 1 0 11776 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_123
timestamp 1605641404
transform 1 0 12420 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 14260 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  FILLER_25_140
timestamp 1605641404
transform 1 0 13984 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 16376 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16928 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1605641404
transform 1 0 16192 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_170
timestamp 1605641404
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 18032 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 18584 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1605641404
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_181
timestamp 1605641404
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_188
timestamp 1605641404
transform 1 0 18400 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 20240 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 20792 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_25_206
timestamp 1605641404
transform 1 0 20056 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1605641404
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1605641404
transform -1 0 22816 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_230
timestamp 1605641404
transform 1 0 22264 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_10
timestamp 1605641404
transform 1 0 2024 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp 1605641404
transform 1 0 1380 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_9
timestamp 1605641404
transform 1 0 1932 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1605641404
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1605641404
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1605641404
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1605641404
transform 1 0 1564 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1605641404
transform 1 0 1656 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 2208 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 2116 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 4048 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 4600 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 4600 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1605641404
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1605641404
transform 1 0 3588 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_36
timestamp 1605641404
transform 1 0 4416 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_28
timestamp 1605641404
transform 1 0 3680 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1605641404
transform 1 0 4416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _78_
timestamp 1605641404
transform 1 0 6808 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 5612 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6624 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1605641404
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1605641404
transform 1 0 5428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_58
timestamp 1605641404
transform 1 0 6440 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1605641404
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8280 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7452 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 9108 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_26_76
timestamp 1605641404
transform 1 0 8096 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_87
timestamp 1605641404
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_66
timestamp 1605641404
transform 1 0 7176 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_85
timestamp 1605641404
transform 1 0 8924 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 10764 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 9660 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1605641404
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_prog_clk
timestamp 1605641404
transform 1 0 9292 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_109
timestamp 1605641404
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1605641404
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_109
timestamp 1605641404
transform 1 0 11132 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 11316 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 11316 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 12420 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 12420 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1605641404
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_120
timestamp 1605641404
transform 1 0 12144 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1605641404
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 14076 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 14352 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_prog_clk
timestamp 1605641404
transform 1 0 14076 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_139
timestamp 1605641404
transform 1 0 13892 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1605641404
transform 1 0 14904 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_139
timestamp 1605641404
transform 1 0 13892 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 16100 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 16008 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1605641404
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_prog_clk
timestamp 1605641404
transform 1 0 15824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_158
timestamp 1605641404
transform 1 0 15640 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_160
timestamp 1605641404
transform 1 0 15824 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1605641404
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_178
timestamp 1605641404
transform 1 0 17480 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_184
timestamp 1605641404
transform 1 0 18032 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_prog_clk
timestamp 1605641404
transform 1 0 17664 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1605641404
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_190
timestamp 1605641404
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1605641404
transform 1 0 18952 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1605641404
transform 1 0 18216 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 18768 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 19136 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 19780 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 20884 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1605641404
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_212
timestamp 1605641404
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1605641404
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 21436 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1605641404
transform -1 0 22816 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1605641404
transform -1 0 22816 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_231
timestamp 1605641404
transform 1 0 22356 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_219
timestamp 1605641404
transform 1 0 21252 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_230
timestamp 1605641404
transform 1 0 22264 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 1564 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1605641404
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1605641404
transform 1 0 1380 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_21
timestamp 1605641404
transform 1 0 3036 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 3220 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4324 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1605641404
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1605641404
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1605641404
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _80_
timestamp 1605641404
transform 1 0 5980 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 6716 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1605641404
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_57
timestamp 1605641404
transform 1 0 6348 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 8832 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1605641404
transform 1 0 8648 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 10672 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1605641404
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1605641404
transform 1 0 9200 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_102
timestamp 1605641404
transform 1 0 10488 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_108
timestamp 1605641404
transform 1 0 11040 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 12420 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1605641404
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 14076 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_28_139
timestamp 1605641404
transform 1 0 13892 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_150
timestamp 1605641404
transform 1 0 14904 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1605641404
transform 1 0 16284 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 16836 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1605641404
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_163
timestamp 1605641404
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1605641404
transform 1 0 16652 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1605641404
transform 1 0 18492 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1605641404
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 20884 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1605641404
transform 1 0 20148 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1605641404
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1605641404
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1605641404
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1605641404
transform 1 0 21896 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1605641404
transform -1 0 22816 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_224
timestamp 1605641404
transform 1 0 21712 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_230
timestamp 1605641404
transform 1 0 22264 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 1564 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1605641404
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1605641404
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1605641404
transform 1 0 3036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 3220 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 5060 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_28
timestamp 1605641404
transform 1 0 3680 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_41
timestamp 1605641404
transform 1 0 4876 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1605641404
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1605641404
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8464 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 1605641404
transform 1 0 8280 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1605641404
transform 1 0 10120 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_96
timestamp 1605641404
transform 1 0 9936 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1605641404
transform 1 0 10948 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 11316 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 12420 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1605641404
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1605641404
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 14076 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14904 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_prog_clk
timestamp 1605641404
transform 1 0 14628 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1605641404
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 1605641404
transform 1 0 14444 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 16652 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_166
timestamp 1605641404
transform 1 0 16376 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1605641404
transform 1 0 18124 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1605641404
transform 1 0 18676 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1605641404
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_178
timestamp 1605641404
transform 1 0 17480 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1605641404
transform 1 0 17848 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_184
timestamp 1605641404
transform 1 0 18032 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_189
timestamp 1605641404
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 20332 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 1605641404
transform 1 0 20148 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_218
timestamp 1605641404
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 21344 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1605641404
transform -1 0 22816 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_229
timestamp 1605641404
transform 1 0 22172 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 1932 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1605641404
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1605641404
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 4048 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4876 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1605641404
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_25
timestamp 1605641404
transform 1 0 3404 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_36
timestamp 1605641404
transform 1 0 4416 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_40
timestamp 1605641404
transform 1 0 4784 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6164 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_prog_clk
timestamp 1605641404
transform 1 0 5888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_50
timestamp 1605641404
transform 1 0 5704 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1605641404
transform 1 0 8832 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 7820 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_71
timestamp 1605641404
transform 1 0 7636 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1605641404
transform 1 0 8648 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1605641404
transform 1 0 10028 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 11040 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1605641404
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1605641404
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_93
timestamp 1605641404
transform 1 0 9660 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_106
timestamp 1605641404
transform 1 0 10856 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 11592 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12604 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_112
timestamp 1605641404
transform 1 0 11408 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_123
timestamp 1605641404
transform 1 0 12420 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 14260 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1605641404
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1605641404
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 15272 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1605641404
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_170
timestamp 1605641404
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1605641404
transform 1 0 19136 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1605641404
transform 1 0 17480 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1605641404
transform 1 0 17296 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1605641404
transform 1 0 18952 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 20884 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1605641404
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1605641404
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1605641404
transform 1 0 22080 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1605641404
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1605641404
transform 1 0 21896 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 1605641404
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_231
timestamp 1605641404
transform 1 0 22356 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 3036 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 1380 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1605641404
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1605641404
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 4416 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_31_30
timestamp 1605641404
transform 1 0 3864 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6808 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1605641404
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_57
timestamp 1605641404
transform 1 0 6348 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 8188 0 1 19040
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_6  FILLER_31_71
timestamp 1605641404
transform 1 0 7636 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10672 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_prog_clk
timestamp 1605641404
transform 1 0 10304 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1605641404
transform 1 0 10120 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1605641404
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 12420 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1605641404
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1605641404
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 13432 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 14168 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_132
timestamp 1605641404
transform 1 0 13248 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_139
timestamp 1605641404
transform 1 0 13892 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 15824 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1605641404
transform 1 0 16928 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_158
timestamp 1605641404
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1605641404
transform 1 0 16652 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1605641404
transform 1 0 18032 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1605641404
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1605641404
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_193
timestamp 1605641404
transform 1 0 18860 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1605641404
transform 1 0 20884 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1605641404
transform 1 0 19412 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1605641404
transform 1 0 22080 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1605641404
transform -1 0 22816 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1605641404
transform 1 0 21896 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_224
timestamp 1605641404
transform 1 0 21712 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_231
timestamp 1605641404
transform 1 0 22356 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 1380 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 2392 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1605641404
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_12
timestamp 1605641404
transform 1 0 2208 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 4048 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 5060 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 3404 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1605641404
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1605641404
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1605641404
transform 1 0 3772 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1605641404
transform 1 0 4876 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 6348 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_32_52
timestamp 1605641404
transform 1 0 5888 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_56
timestamp 1605641404
transform 1 0 6256 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1605641404
transform 1 0 8464 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_32_78
timestamp 1605641404
transform 1 0 8280 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1605641404
transform 1 0 10672 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1605641404
transform 1 0 9660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1605641404
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_89
timestamp 1605641404
transform 1 0 9292 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_102
timestamp 1605641404
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1605641404
transform 1 0 12788 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_125
timestamp 1605641404
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_131
timestamp 1605641404
transform 1 0 13156 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1605641404
transform 1 0 13524 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1605641404
transform 1 0 14996 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1605641404
transform 1 0 16284 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1605641404
transform 1 0 16928 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1605641404
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1605641404
transform 1 0 16100 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1605641404
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1605641404
transform 1 0 18584 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1605641404
transform 1 0 19136 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_32_188
timestamp 1605641404
transform 1 0 18400 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1605641404
transform 1 0 18952 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1605641404
transform 1 0 20884 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1605641404
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_212
timestamp 1605641404
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1605641404
transform -1 0 22816 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_231
timestamp 1605641404
transform 1 0 22356 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1605641404
transform 1 0 1564 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 1380 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 2116 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1605641404
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1605641404
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_19
timestamp 1605641404
transform 1 0 2852 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1605641404
transform 1 0 1380 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_9
timestamp 1605641404
transform 1 0 1932 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1605641404
transform 1 0 4048 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 3128 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 4784 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 4968 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1605641404
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_38
timestamp 1605641404
transform 1 0 4600 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1605641404
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_36
timestamp 1605641404
transform 1 0 4416 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 6808 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 6624 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1605641404
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_56
timestamp 1605641404
transform 1 0 6256 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1605641404
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_58
timestamp 1605641404
transform 1 0 6440 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 7912 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 8556 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_33_78
timestamp 1605641404
transform 1 0 8280 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_69
timestamp 1605641404
transform 1 0 7452 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1605641404
transform 1 0 7820 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_93
timestamp 1605641404
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_90
timestamp 1605641404
transform 1 0 9384 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_97
timestamp 1605641404
transform 1 0 10028 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1605641404
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 10028 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_106
timestamp 1605641404
transform 1 0 10856 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_102
timestamp 1605641404
transform 1 0 10488 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _51_
timestamp 1605641404
transform 1 0 10212 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 11040 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 10672 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 12420 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 12880 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1605641404
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1605641404
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_124
timestamp 1605641404
transform 1 0 12512 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1605641404
transform 1 0 14628 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1605641404
transform 1 0 14352 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1605641404
transform 1 0 14904 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_33_139
timestamp 1605641404
transform 1 0 13892 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_143
timestamp 1605641404
transform 1 0 14260 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1605641404
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_144
timestamp 1605641404
transform 1 0 14352 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1605641404
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1605641404
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1605641404
transform 1 0 16560 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1605641404
transform 1 0 15824 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1605641404
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1605641404
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_158
timestamp 1605641404
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _43_
timestamp 1605641404
transform 1 0 18032 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1605641404
transform 1 0 18492 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1605641404
transform 1 0 19136 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1605641404
transform 1 0 17480 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1605641404
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_177
timestamp 1605641404
transform 1 0 17388 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1605641404
transform 1 0 18308 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_176
timestamp 1605641404
transform 1 0 17296 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1605641404
transform 1 0 18952 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1605641404
transform 1 0 21160 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1605641404
transform 1 0 20884 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1605641404
transform 1 0 19504 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1605641404
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_198
timestamp 1605641404
transform 1 0 19320 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_216
timestamp 1605641404
transform 1 0 20976 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_212
timestamp 1605641404
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1605641404
transform 1 0 21896 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1605641404
transform -1 0 22816 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1605641404
transform -1 0 22816 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_227
timestamp 1605641404
transform 1 0 21988 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_224
timestamp 1605641404
transform 1 0 21712 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_230
timestamp 1605641404
transform 1 0 22264 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1605641404
transform 1 0 1380 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1605641404
transform 1 0 2944 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1605641404
transform 1 0 1932 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1605641404
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_7
timestamp 1605641404
transform 1 0 1748 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_18
timestamp 1605641404
transform 1 0 2760 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 4048 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 5060 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1605641404
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_29
timestamp 1605641404
transform 1 0 3772 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1605641404
transform 1 0 4876 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1605641404
transform 1 0 6072 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1605641404
transform 1 0 6900 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1605641404
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_52
timestamp 1605641404
transform 1 0 5888 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_58
timestamp 1605641404
transform 1 0 6440 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 8556 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_35_79
timestamp 1605641404
transform 1 0 8372 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1605641404
transform 1 0 9752 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1605641404
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_90
timestamp 1605641404
transform 1 0 9384 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _79_
timestamp 1605641404
transform 1 0 12604 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1605641404
transform 1 0 11408 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1605641404
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1605641404
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_121
timestamp 1605641404
transform 1 0 12236 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_129
timestamp 1605641404
transform 1 0 12972 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1605641404
transform 1 0 13432 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_35_133
timestamp 1605641404
transform 1 0 13340 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_150
timestamp 1605641404
transform 1 0 14904 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1605641404
transform 1 0 15456 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1605641404
transform 1 0 16468 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1605641404
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_154
timestamp 1605641404
transform 1 0 15272 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_165
timestamp 1605641404
transform 1 0 16284 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1605641404
transform 1 0 17664 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1605641404
transform 1 0 18308 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1605641404
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_176
timestamp 1605641404
transform 1 0 17296 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1605641404
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_196
timestamp 1605641404
transform 1 0 19136 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1605641404
transform 1 0 21160 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1605641404
transform 1 0 19688 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1605641404
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1605641404
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1605641404
transform -1 0 22816 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1605641404
transform 1 0 21988 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_229
timestamp 1605641404
transform 1 0 22172 0 1 21216
box -38 -48 406 592
<< labels >>
rlabel metal2 s 19982 0 20038 480 6 Test_en
port 0 nsew default input
rlabel metal2 s 3974 0 4030 480 6 bottom_width_0_height_0__pin_50_
port 1 nsew default tristate
rlabel metal2 s 11978 0 12034 480 6 bottom_width_0_height_0__pin_51_
port 2 nsew default tristate
rlabel metal3 s 0 11840 480 11960 6 ccff_head
port 3 nsew default input
rlabel metal3 s 23520 5992 24000 6112 6 ccff_tail
port 4 nsew default tristate
rlabel metal3 s 0 19864 480 19984 6 left_width_0_height_0__pin_52_
port 5 nsew default input
rlabel metal3 s 0 3952 480 4072 6 prog_clk
port 6 nsew default input
rlabel metal3 s 23520 6808 24000 6928 6 right_width_0_height_0__pin_16_
port 7 nsew default input
rlabel metal3 s 23520 7488 24000 7608 6 right_width_0_height_0__pin_17_
port 8 nsew default input
rlabel metal3 s 23520 8168 24000 8288 6 right_width_0_height_0__pin_18_
port 9 nsew default input
rlabel metal3 s 23520 8984 24000 9104 6 right_width_0_height_0__pin_19_
port 10 nsew default input
rlabel metal3 s 23520 9664 24000 9784 6 right_width_0_height_0__pin_20_
port 11 nsew default input
rlabel metal3 s 23520 10344 24000 10464 6 right_width_0_height_0__pin_21_
port 12 nsew default input
rlabel metal3 s 23520 11160 24000 11280 6 right_width_0_height_0__pin_22_
port 13 nsew default input
rlabel metal3 s 23520 11840 24000 11960 6 right_width_0_height_0__pin_23_
port 14 nsew default input
rlabel metal3 s 23520 12520 24000 12640 6 right_width_0_height_0__pin_24_
port 15 nsew default input
rlabel metal3 s 23520 13336 24000 13456 6 right_width_0_height_0__pin_25_
port 16 nsew default input
rlabel metal3 s 23520 14016 24000 14136 6 right_width_0_height_0__pin_26_
port 17 nsew default input
rlabel metal3 s 23520 14696 24000 14816 6 right_width_0_height_0__pin_27_
port 18 nsew default input
rlabel metal3 s 23520 15512 24000 15632 6 right_width_0_height_0__pin_28_
port 19 nsew default input
rlabel metal3 s 23520 16192 24000 16312 6 right_width_0_height_0__pin_29_
port 20 nsew default input
rlabel metal3 s 23520 16872 24000 16992 6 right_width_0_height_0__pin_30_
port 21 nsew default input
rlabel metal3 s 23520 17688 24000 17808 6 right_width_0_height_0__pin_31_
port 22 nsew default input
rlabel metal3 s 23520 280 24000 400 6 right_width_0_height_0__pin_42_lower
port 23 nsew default tristate
rlabel metal3 s 23520 18368 24000 18488 6 right_width_0_height_0__pin_42_upper
port 24 nsew default tristate
rlabel metal3 s 23520 960 24000 1080 6 right_width_0_height_0__pin_43_lower
port 25 nsew default tristate
rlabel metal3 s 23520 19048 24000 19168 6 right_width_0_height_0__pin_43_upper
port 26 nsew default tristate
rlabel metal3 s 23520 1640 24000 1760 6 right_width_0_height_0__pin_44_lower
port 27 nsew default tristate
rlabel metal3 s 23520 19864 24000 19984 6 right_width_0_height_0__pin_44_upper
port 28 nsew default tristate
rlabel metal3 s 23520 2456 24000 2576 6 right_width_0_height_0__pin_45_lower
port 29 nsew default tristate
rlabel metal3 s 23520 20544 24000 20664 6 right_width_0_height_0__pin_45_upper
port 30 nsew default tristate
rlabel metal3 s 23520 3136 24000 3256 6 right_width_0_height_0__pin_46_lower
port 31 nsew default tristate
rlabel metal3 s 23520 21224 24000 21344 6 right_width_0_height_0__pin_46_upper
port 32 nsew default tristate
rlabel metal3 s 23520 3816 24000 3936 6 right_width_0_height_0__pin_47_lower
port 33 nsew default tristate
rlabel metal3 s 23520 22040 24000 22160 6 right_width_0_height_0__pin_47_upper
port 34 nsew default tristate
rlabel metal3 s 23520 4632 24000 4752 6 right_width_0_height_0__pin_48_lower
port 35 nsew default tristate
rlabel metal3 s 23520 22720 24000 22840 6 right_width_0_height_0__pin_48_upper
port 36 nsew default tristate
rlabel metal3 s 23520 5312 24000 5432 6 right_width_0_height_0__pin_49_lower
port 37 nsew default tristate
rlabel metal3 s 23520 23400 24000 23520 6 right_width_0_height_0__pin_49_upper
port 38 nsew default tristate
rlabel metal2 s 5906 23520 5962 24000 6 top_width_0_height_0__pin_0_
port 39 nsew default input
rlabel metal2 s 12990 23520 13046 24000 6 top_width_0_height_0__pin_10_
port 40 nsew default input
rlabel metal2 s 13634 23520 13690 24000 6 top_width_0_height_0__pin_11_
port 41 nsew default input
rlabel metal2 s 14370 23520 14426 24000 6 top_width_0_height_0__pin_12_
port 42 nsew default input
rlabel metal2 s 15106 23520 15162 24000 6 top_width_0_height_0__pin_13_
port 43 nsew default input
rlabel metal2 s 15750 23520 15806 24000 6 top_width_0_height_0__pin_14_
port 44 nsew default input
rlabel metal2 s 16486 23520 16542 24000 6 top_width_0_height_0__pin_15_
port 45 nsew default input
rlabel metal2 s 6642 23520 6698 24000 6 top_width_0_height_0__pin_1_
port 46 nsew default input
rlabel metal2 s 7286 23520 7342 24000 6 top_width_0_height_0__pin_2_
port 47 nsew default input
rlabel metal2 s 17222 23520 17278 24000 6 top_width_0_height_0__pin_32_
port 48 nsew default input
rlabel metal2 s 17866 23520 17922 24000 6 top_width_0_height_0__pin_33_
port 49 nsew default input
rlabel metal2 s 18602 23520 18658 24000 6 top_width_0_height_0__pin_34_lower
port 50 nsew default tristate
rlabel metal2 s 294 23520 350 24000 6 top_width_0_height_0__pin_34_upper
port 51 nsew default tristate
rlabel metal2 s 19338 23520 19394 24000 6 top_width_0_height_0__pin_35_lower
port 52 nsew default tristate
rlabel metal2 s 938 23520 994 24000 6 top_width_0_height_0__pin_35_upper
port 53 nsew default tristate
rlabel metal2 s 19982 23520 20038 24000 6 top_width_0_height_0__pin_36_lower
port 54 nsew default tristate
rlabel metal2 s 1674 23520 1730 24000 6 top_width_0_height_0__pin_36_upper
port 55 nsew default tristate
rlabel metal2 s 20718 23520 20774 24000 6 top_width_0_height_0__pin_37_lower
port 56 nsew default tristate
rlabel metal2 s 2410 23520 2466 24000 6 top_width_0_height_0__pin_37_upper
port 57 nsew default tristate
rlabel metal2 s 21454 23520 21510 24000 6 top_width_0_height_0__pin_38_lower
port 58 nsew default tristate
rlabel metal2 s 3054 23520 3110 24000 6 top_width_0_height_0__pin_38_upper
port 59 nsew default tristate
rlabel metal2 s 22098 23520 22154 24000 6 top_width_0_height_0__pin_39_lower
port 60 nsew default tristate
rlabel metal2 s 3790 23520 3846 24000 6 top_width_0_height_0__pin_39_upper
port 61 nsew default tristate
rlabel metal2 s 8022 23520 8078 24000 6 top_width_0_height_0__pin_3_
port 62 nsew default input
rlabel metal2 s 22834 23520 22890 24000 6 top_width_0_height_0__pin_40_lower
port 63 nsew default tristate
rlabel metal2 s 4526 23520 4582 24000 6 top_width_0_height_0__pin_40_upper
port 64 nsew default tristate
rlabel metal2 s 23570 23520 23626 24000 6 top_width_0_height_0__pin_41_lower
port 65 nsew default tristate
rlabel metal2 s 5170 23520 5226 24000 6 top_width_0_height_0__pin_41_upper
port 66 nsew default tristate
rlabel metal2 s 8758 23520 8814 24000 6 top_width_0_height_0__pin_4_
port 67 nsew default input
rlabel metal2 s 9402 23520 9458 24000 6 top_width_0_height_0__pin_5_
port 68 nsew default input
rlabel metal2 s 10138 23520 10194 24000 6 top_width_0_height_0__pin_6_
port 69 nsew default input
rlabel metal2 s 10874 23520 10930 24000 6 top_width_0_height_0__pin_7_
port 70 nsew default input
rlabel metal2 s 11518 23520 11574 24000 6 top_width_0_height_0__pin_8_
port 71 nsew default input
rlabel metal2 s 12254 23520 12310 24000 6 top_width_0_height_0__pin_9_
port 72 nsew default input
rlabel metal4 s 4576 2128 4896 21808 6 VPWR
port 73 nsew default input
rlabel metal4 s 8208 2128 8528 21808 6 VGND
port 74 nsew default input
<< properties >>
string FIXED_BBOX 0 0 24000 24000
<< end >>
