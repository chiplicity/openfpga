VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__0_
  CLASS BLOCK ;
  FOREIGN sb_2__0_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 114.000 BY 114.000 ;
  PIN ccff_head
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 110.000 57.160 114.000 57.760 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.720 4.000 103.320 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 86.400 4.000 87.000 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.120 4.000 89.720 ;
    END
  END chanx_left_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.950 110.000 19.230 114.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.950 110.000 42.230 114.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 110.000 44.530 114.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.550 110.000 46.830 114.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.850 110.000 49.130 114.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 110.000 51.430 114.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 110.000 53.730 114.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.750 110.000 56.030 114.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 110.000 58.330 114.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 110.000 60.170 114.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 110.000 62.470 114.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.250 110.000 21.530 114.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.550 110.000 23.830 114.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.850 110.000 26.130 114.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 110.000 28.430 114.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 110.000 30.730 114.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.750 110.000 33.030 114.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 110.000 35.330 114.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 110.000 37.630 114.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.650 110.000 39.930 114.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 110.000 64.770 114.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 110.000 87.770 114.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 110.000 90.070 114.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 92.090 110.000 92.370 114.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 110.000 94.670 114.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 96.690 110.000 96.970 114.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 110.000 99.270 114.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 110.000 101.570 114.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.590 110.000 103.870 114.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 110.000 106.170 114.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 110.000 108.470 114.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 66.790 110.000 67.070 114.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 110.000 69.370 114.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 71.390 110.000 71.670 114.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 110.000 73.970 114.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 110.000 76.270 114.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 110.000 78.570 114.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 110.000 80.870 114.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 110.000 83.170 114.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 110.000 85.470 114.000 ;
    END
  END chany_top_out[9]
  PIN left_bottom_grid_pin_11_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_11_
  PIN left_bottom_grid_pin_13_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_13_
  PIN left_bottom_grid_pin_15_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END left_bottom_grid_pin_15_
  PIN left_bottom_grid_pin_17_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END left_bottom_grid_pin_17_
  PIN left_bottom_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END left_bottom_grid_pin_1_
  PIN left_bottom_grid_pin_3_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END left_bottom_grid_pin_3_
  PIN left_bottom_grid_pin_5_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END left_bottom_grid_pin_5_
  PIN left_bottom_grid_pin_7_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END left_bottom_grid_pin_7_
  PIN left_bottom_grid_pin_9_
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END left_bottom_grid_pin_9_
  PIN prog_clk_0_N_in
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 110.000 110.770 114.000 ;
    END
  END prog_clk_0_N_in
  PIN top_left_grid_pin_42_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.010 110.000 1.290 114.000 ;
    END
  END top_left_grid_pin_42_
  PIN top_left_grid_pin_43_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 110.000 3.130 114.000 ;
    END
  END top_left_grid_pin_43_
  PIN top_left_grid_pin_44_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 110.000 5.430 114.000 ;
    END
  END top_left_grid_pin_44_
  PIN top_left_grid_pin_45_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 110.000 7.730 114.000 ;
    END
  END top_left_grid_pin_45_
  PIN top_left_grid_pin_46_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.750 110.000 10.030 114.000 ;
    END
  END top_left_grid_pin_46_
  PIN top_left_grid_pin_47_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.050 110.000 12.330 114.000 ;
    END
  END top_left_grid_pin_47_
  PIN top_left_grid_pin_48_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 110.000 14.630 114.000 ;
    END
  END top_left_grid_pin_48_
  PIN top_left_grid_pin_49_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 110.000 16.930 114.000 ;
    END
  END top_left_grid_pin_49_
  PIN top_right_grid_pin_1_
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 110.000 113.070 114.000 ;
    END
  END top_right_grid_pin_1_
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.880 10.640 23.480 100.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.040 10.640 40.640 100.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 108.100 100.725 ;
      LAYER met1 ;
        RECT 0.990 2.760 113.090 103.660 ;
      LAYER met2 ;
        RECT 1.570 109.720 2.570 112.725 ;
        RECT 3.410 109.720 4.870 112.725 ;
        RECT 5.710 109.720 7.170 112.725 ;
        RECT 8.010 109.720 9.470 112.725 ;
        RECT 10.310 109.720 11.770 112.725 ;
        RECT 12.610 109.720 14.070 112.725 ;
        RECT 14.910 109.720 16.370 112.725 ;
        RECT 17.210 109.720 18.670 112.725 ;
        RECT 19.510 109.720 20.970 112.725 ;
        RECT 21.810 109.720 23.270 112.725 ;
        RECT 24.110 109.720 25.570 112.725 ;
        RECT 26.410 109.720 27.870 112.725 ;
        RECT 28.710 109.720 30.170 112.725 ;
        RECT 31.010 109.720 32.470 112.725 ;
        RECT 33.310 109.720 34.770 112.725 ;
        RECT 35.610 109.720 37.070 112.725 ;
        RECT 37.910 109.720 39.370 112.725 ;
        RECT 40.210 109.720 41.670 112.725 ;
        RECT 42.510 109.720 43.970 112.725 ;
        RECT 44.810 109.720 46.270 112.725 ;
        RECT 47.110 109.720 48.570 112.725 ;
        RECT 49.410 109.720 50.870 112.725 ;
        RECT 51.710 109.720 53.170 112.725 ;
        RECT 54.010 109.720 55.470 112.725 ;
        RECT 56.310 109.720 57.770 112.725 ;
        RECT 58.610 109.720 59.610 112.725 ;
        RECT 60.450 109.720 61.910 112.725 ;
        RECT 62.750 109.720 64.210 112.725 ;
        RECT 65.050 109.720 66.510 112.725 ;
        RECT 67.350 109.720 68.810 112.725 ;
        RECT 69.650 109.720 71.110 112.725 ;
        RECT 71.950 109.720 73.410 112.725 ;
        RECT 74.250 109.720 75.710 112.725 ;
        RECT 76.550 109.720 78.010 112.725 ;
        RECT 78.850 109.720 80.310 112.725 ;
        RECT 81.150 109.720 82.610 112.725 ;
        RECT 83.450 109.720 84.910 112.725 ;
        RECT 85.750 109.720 87.210 112.725 ;
        RECT 88.050 109.720 89.510 112.725 ;
        RECT 90.350 109.720 91.810 112.725 ;
        RECT 92.650 109.720 94.110 112.725 ;
        RECT 94.950 109.720 96.410 112.725 ;
        RECT 97.250 109.720 98.710 112.725 ;
        RECT 99.550 109.720 101.010 112.725 ;
        RECT 101.850 109.720 103.310 112.725 ;
        RECT 104.150 109.720 105.610 112.725 ;
        RECT 106.450 109.720 107.910 112.725 ;
        RECT 108.750 109.720 110.210 112.725 ;
        RECT 111.050 109.720 112.510 112.725 ;
        RECT 1.020 4.280 113.060 109.720 ;
        RECT 1.020 0.835 56.850 4.280 ;
        RECT 57.690 0.835 113.060 4.280 ;
      LAYER met3 ;
        RECT 4.400 111.840 110.000 112.705 ;
        RECT 4.000 111.200 110.000 111.840 ;
        RECT 4.400 109.800 110.000 111.200 ;
        RECT 4.000 108.480 110.000 109.800 ;
        RECT 4.400 107.080 110.000 108.480 ;
        RECT 4.000 106.440 110.000 107.080 ;
        RECT 4.400 105.040 110.000 106.440 ;
        RECT 4.000 103.720 110.000 105.040 ;
        RECT 4.400 102.320 110.000 103.720 ;
        RECT 4.000 101.680 110.000 102.320 ;
        RECT 4.400 100.280 110.000 101.680 ;
        RECT 4.000 99.640 110.000 100.280 ;
        RECT 4.400 98.240 110.000 99.640 ;
        RECT 4.000 96.920 110.000 98.240 ;
        RECT 4.400 95.520 110.000 96.920 ;
        RECT 4.000 94.880 110.000 95.520 ;
        RECT 4.400 93.480 110.000 94.880 ;
        RECT 4.000 92.160 110.000 93.480 ;
        RECT 4.400 90.760 110.000 92.160 ;
        RECT 4.000 90.120 110.000 90.760 ;
        RECT 4.400 88.720 110.000 90.120 ;
        RECT 4.000 87.400 110.000 88.720 ;
        RECT 4.400 86.000 110.000 87.400 ;
        RECT 4.000 85.360 110.000 86.000 ;
        RECT 4.400 83.960 110.000 85.360 ;
        RECT 4.000 83.320 110.000 83.960 ;
        RECT 4.400 81.920 110.000 83.320 ;
        RECT 4.000 80.600 110.000 81.920 ;
        RECT 4.400 79.200 110.000 80.600 ;
        RECT 4.000 78.560 110.000 79.200 ;
        RECT 4.400 77.160 110.000 78.560 ;
        RECT 4.000 75.840 110.000 77.160 ;
        RECT 4.400 74.440 110.000 75.840 ;
        RECT 4.000 73.800 110.000 74.440 ;
        RECT 4.400 72.400 110.000 73.800 ;
        RECT 4.000 71.080 110.000 72.400 ;
        RECT 4.400 69.680 110.000 71.080 ;
        RECT 4.000 69.040 110.000 69.680 ;
        RECT 4.400 67.640 110.000 69.040 ;
        RECT 4.000 67.000 110.000 67.640 ;
        RECT 4.400 65.600 110.000 67.000 ;
        RECT 4.000 64.280 110.000 65.600 ;
        RECT 4.400 62.880 110.000 64.280 ;
        RECT 4.000 62.240 110.000 62.880 ;
        RECT 4.400 60.840 110.000 62.240 ;
        RECT 4.000 59.520 110.000 60.840 ;
        RECT 4.400 58.160 110.000 59.520 ;
        RECT 4.400 58.120 109.600 58.160 ;
        RECT 4.000 57.480 109.600 58.120 ;
        RECT 4.400 56.760 109.600 57.480 ;
        RECT 4.400 56.080 110.000 56.760 ;
        RECT 4.000 54.760 110.000 56.080 ;
        RECT 4.400 53.360 110.000 54.760 ;
        RECT 4.000 52.720 110.000 53.360 ;
        RECT 4.400 51.320 110.000 52.720 ;
        RECT 4.000 50.680 110.000 51.320 ;
        RECT 4.400 49.280 110.000 50.680 ;
        RECT 4.000 47.960 110.000 49.280 ;
        RECT 4.400 46.560 110.000 47.960 ;
        RECT 4.000 45.920 110.000 46.560 ;
        RECT 4.400 44.520 110.000 45.920 ;
        RECT 4.000 43.200 110.000 44.520 ;
        RECT 4.400 41.800 110.000 43.200 ;
        RECT 4.000 41.160 110.000 41.800 ;
        RECT 4.400 39.760 110.000 41.160 ;
        RECT 4.000 38.440 110.000 39.760 ;
        RECT 4.400 37.040 110.000 38.440 ;
        RECT 4.000 36.400 110.000 37.040 ;
        RECT 4.400 35.000 110.000 36.400 ;
        RECT 4.000 34.360 110.000 35.000 ;
        RECT 4.400 32.960 110.000 34.360 ;
        RECT 4.000 31.640 110.000 32.960 ;
        RECT 4.400 30.240 110.000 31.640 ;
        RECT 4.000 29.600 110.000 30.240 ;
        RECT 4.400 28.200 110.000 29.600 ;
        RECT 4.000 26.880 110.000 28.200 ;
        RECT 4.400 25.480 110.000 26.880 ;
        RECT 4.000 24.840 110.000 25.480 ;
        RECT 4.400 23.440 110.000 24.840 ;
        RECT 4.000 22.120 110.000 23.440 ;
        RECT 4.400 20.720 110.000 22.120 ;
        RECT 4.000 20.080 110.000 20.720 ;
        RECT 4.400 18.680 110.000 20.080 ;
        RECT 4.000 18.040 110.000 18.680 ;
        RECT 4.400 16.640 110.000 18.040 ;
        RECT 4.000 15.320 110.000 16.640 ;
        RECT 4.400 13.920 110.000 15.320 ;
        RECT 4.000 13.280 110.000 13.920 ;
        RECT 4.400 11.880 110.000 13.280 ;
        RECT 4.000 10.560 110.000 11.880 ;
        RECT 4.400 9.160 110.000 10.560 ;
        RECT 4.000 8.520 110.000 9.160 ;
        RECT 4.400 7.120 110.000 8.520 ;
        RECT 4.000 5.800 110.000 7.120 ;
        RECT 4.400 4.400 110.000 5.800 ;
        RECT 4.000 3.760 110.000 4.400 ;
        RECT 4.400 2.360 110.000 3.760 ;
        RECT 4.000 1.720 110.000 2.360 ;
        RECT 4.400 0.855 110.000 1.720 ;
      LAYER met4 ;
        RECT 56.200 10.640 92.120 100.880 ;
  END
END sb_2__0_
END LIBRARY

