magic
tech EFS8A
magscale 1 2
timestamp 1603796101
<< locali >>
rect 20453 6647 20487 6749
rect 2605 5083 2639 5321
rect 11621 3927 11655 4097
rect 4905 2975 4939 3145
<< viali >>
rect 1593 9129 1627 9163
rect 1409 8993 1443 9027
rect 6469 8993 6503 9027
rect 6653 8789 6687 8823
rect 1547 8585 1581 8619
rect 20499 8585 20533 8619
rect 6975 8517 7009 8551
rect 2329 8449 2363 8483
rect 1476 8381 1510 8415
rect 6904 8381 6938 8415
rect 16313 8381 16347 8415
rect 17049 8381 17083 8415
rect 20428 8381 20462 8415
rect 1961 8313 1995 8347
rect 6561 8313 6595 8347
rect 7297 8313 7331 8347
rect 20913 8313 20947 8347
rect 16681 8245 16715 8279
rect 1593 8041 1627 8075
rect 16313 8041 16347 8075
rect 35633 8041 35667 8075
rect 7021 7973 7055 8007
rect 16681 7973 16715 8007
rect 21234 7973 21268 8007
rect 28365 7973 28399 8007
rect 1409 7905 1443 7939
rect 5892 7905 5926 7939
rect 13185 7905 13219 7939
rect 14197 7905 14231 7939
rect 15669 7905 15703 7939
rect 17141 7905 17175 7939
rect 35449 7905 35483 7939
rect 6929 7837 6963 7871
rect 7205 7837 7239 7871
rect 20729 7837 20763 7871
rect 20913 7837 20947 7871
rect 28273 7837 28307 7871
rect 28917 7837 28951 7871
rect 5963 7769 5997 7803
rect 5273 7701 5307 7735
rect 6653 7701 6687 7735
rect 13369 7701 13403 7735
rect 14381 7701 14415 7735
rect 15853 7701 15887 7735
rect 17325 7701 17359 7735
rect 19533 7701 19567 7735
rect 21833 7701 21867 7735
rect 22109 7701 22143 7735
rect 25329 7701 25363 7735
rect 1869 7497 1903 7531
rect 7757 7497 7791 7531
rect 8033 7497 8067 7531
rect 16129 7497 16163 7531
rect 16359 7497 16393 7531
rect 17233 7497 17267 7531
rect 21281 7497 21315 7531
rect 28457 7497 28491 7531
rect 28825 7497 28859 7531
rect 29423 7497 29457 7531
rect 15761 7429 15795 7463
rect 16497 7429 16531 7463
rect 16589 7361 16623 7395
rect 21925 7361 21959 7395
rect 27997 7361 28031 7395
rect 5273 7293 5307 7327
rect 6837 7293 6871 7327
rect 8585 7293 8619 7327
rect 12265 7293 12299 7327
rect 13093 7293 13127 7327
rect 15301 7293 15335 7327
rect 18061 7293 18095 7327
rect 18521 7293 18555 7327
rect 19809 7293 19843 7327
rect 19993 7293 20027 7327
rect 20361 7293 20395 7327
rect 20729 7293 20763 7327
rect 25145 7293 25179 7327
rect 25237 7293 25271 7327
rect 25697 7293 25731 7327
rect 26065 7293 26099 7327
rect 26433 7293 26467 7327
rect 29320 7293 29354 7327
rect 29745 7293 29779 7327
rect 35449 7293 35483 7327
rect 5917 7225 5951 7259
rect 7199 7225 7233 7259
rect 13185 7225 13219 7259
rect 14289 7225 14323 7259
rect 16221 7225 16255 7259
rect 16957 7225 16991 7259
rect 19441 7225 19475 7259
rect 22017 7225 22051 7259
rect 22569 7225 22603 7259
rect 26709 7225 26743 7259
rect 1409 7157 1443 7191
rect 4537 7157 4571 7191
rect 5089 7157 5123 7191
rect 6193 7157 6227 7191
rect 6561 7157 6595 7191
rect 8401 7157 8435 7191
rect 8769 7157 8803 7191
rect 9137 7157 9171 7191
rect 13553 7157 13587 7191
rect 13829 7157 13863 7191
rect 14933 7157 14967 7191
rect 18245 7157 18279 7191
rect 18981 7157 19015 7191
rect 20729 7157 20763 7191
rect 21649 7157 21683 7191
rect 24685 7157 24719 7191
rect 5457 6953 5491 6987
rect 13645 6953 13679 6987
rect 14749 6953 14783 6987
rect 15577 6953 15611 6987
rect 21005 6953 21039 6987
rect 24685 6953 24719 6987
rect 25329 6953 25363 6987
rect 28181 6953 28215 6987
rect 7665 6885 7699 6919
rect 27582 6885 27616 6919
rect 29285 6885 29319 6919
rect 1476 6817 1510 6851
rect 5181 6817 5215 6851
rect 5641 6817 5675 6851
rect 6193 6817 6227 6851
rect 6377 6817 6411 6851
rect 11621 6817 11655 6851
rect 11805 6817 11839 6851
rect 12909 6817 12943 6851
rect 13001 6817 13035 6851
rect 15669 6817 15703 6851
rect 17233 6817 17267 6851
rect 18245 6817 18279 6851
rect 19809 6817 19843 6851
rect 21189 6817 21223 6851
rect 21373 6817 21407 6851
rect 21925 6817 21959 6851
rect 22109 6817 22143 6851
rect 24317 6817 24351 6851
rect 24501 6817 24535 6851
rect 25605 6817 25639 6851
rect 27261 6817 27295 6851
rect 4169 6749 4203 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 9689 6749 9723 6783
rect 13148 6749 13182 6783
rect 13369 6749 13403 6783
rect 15025 6749 15059 6783
rect 15816 6749 15850 6783
rect 16037 6749 16071 6783
rect 16405 6749 16439 6783
rect 20269 6749 20303 6783
rect 20453 6749 20487 6783
rect 29193 6749 29227 6783
rect 29837 6749 29871 6783
rect 12541 6681 12575 6715
rect 15945 6681 15979 6715
rect 1547 6613 1581 6647
rect 4721 6613 4755 6647
rect 5089 6613 5123 6647
rect 6929 6613 6963 6647
rect 7297 6613 7331 6647
rect 11897 6613 11931 6647
rect 13277 6613 13311 6647
rect 14105 6613 14139 6647
rect 17417 6613 17451 6647
rect 18429 6613 18463 6647
rect 19533 6613 19567 6647
rect 20453 6613 20487 6647
rect 20637 6613 20671 6647
rect 25973 6613 26007 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 6285 6409 6319 6443
rect 8677 6409 8711 6443
rect 13369 6409 13403 6443
rect 15761 6409 15795 6443
rect 16129 6409 16163 6443
rect 17233 6409 17267 6443
rect 18521 6409 18555 6443
rect 18889 6409 18923 6443
rect 22109 6409 22143 6443
rect 24225 6409 24259 6443
rect 26893 6409 26927 6443
rect 33425 6409 33459 6443
rect 8217 6341 8251 6375
rect 13645 6341 13679 6375
rect 28733 6341 28767 6375
rect 30205 6341 30239 6375
rect 1409 6205 1443 6239
rect 3985 6205 4019 6239
rect 4721 6205 4755 6239
rect 5181 6205 5215 6239
rect 5457 6205 5491 6239
rect 5825 6205 5859 6239
rect 6837 6205 6871 6239
rect 7573 6205 7607 6239
rect 7849 6205 7883 6239
rect 8217 6205 8251 6239
rect 9045 6205 9079 6239
rect 9229 6205 9263 6239
rect 11380 6205 11414 6239
rect 11805 6205 11839 6239
rect 12633 6205 12667 6239
rect 14105 6205 14139 6239
rect 14565 6205 14599 6239
rect 14749 6205 14783 6239
rect 15117 6205 15151 6239
rect 16589 6205 16623 6239
rect 18061 6205 18095 6239
rect 20269 6205 20303 6239
rect 20453 6205 20487 6239
rect 20821 6205 20855 6239
rect 21189 6205 21223 6239
rect 23673 6205 23707 6239
rect 25145 6205 25179 6239
rect 25605 6205 25639 6239
rect 26065 6205 26099 6239
rect 26433 6205 26467 6239
rect 27756 6205 27790 6239
rect 28181 6205 28215 6239
rect 29285 6205 29319 6239
rect 30481 6205 30515 6239
rect 33241 6205 33275 6239
rect 33793 6205 33827 6239
rect 3433 6137 3467 6171
rect 6653 6137 6687 6171
rect 9137 6137 9171 6171
rect 11253 6137 11287 6171
rect 12173 6137 12207 6171
rect 12449 6137 12483 6171
rect 19533 6137 19567 6171
rect 22477 6137 22511 6171
rect 24961 6137 24995 6171
rect 29606 6137 29640 6171
rect 2053 6069 2087 6103
rect 4353 6069 4387 6103
rect 4537 6069 4571 6103
rect 10149 6069 10183 6103
rect 10885 6069 10919 6103
rect 11483 6069 11517 6103
rect 12725 6069 12759 6103
rect 14197 6069 14231 6103
rect 16681 6069 16715 6103
rect 18245 6069 18279 6103
rect 19809 6069 19843 6103
rect 21373 6069 21407 6103
rect 21833 6069 21867 6103
rect 23857 6069 23891 6103
rect 24593 6069 24627 6103
rect 26341 6069 26375 6103
rect 27261 6069 27295 6103
rect 27859 6069 27893 6103
rect 29009 6069 29043 6103
rect 30849 6069 30883 6103
rect 7941 5865 7975 5899
rect 10241 5865 10275 5899
rect 11989 5865 12023 5899
rect 12357 5865 12391 5899
rect 13737 5865 13771 5899
rect 15577 5865 15611 5899
rect 16313 5865 16347 5899
rect 20269 5865 20303 5899
rect 28273 5865 28307 5899
rect 2145 5797 2179 5831
rect 8309 5797 8343 5831
rect 10057 5797 10091 5831
rect 15025 5797 15059 5831
rect 21275 5797 21309 5831
rect 28641 5797 28675 5831
rect 29146 5797 29180 5831
rect 5273 5729 5307 5763
rect 6469 5729 6503 5763
rect 6929 5729 6963 5763
rect 7205 5729 7239 5763
rect 7389 5729 7423 5763
rect 8560 5729 8594 5763
rect 10333 5729 10367 5763
rect 10609 5729 10643 5763
rect 10977 5729 11011 5763
rect 11345 5729 11379 5763
rect 12817 5729 12851 5763
rect 13001 5729 13035 5763
rect 13369 5729 13403 5763
rect 13921 5729 13955 5763
rect 14657 5729 14691 5763
rect 15853 5729 15887 5763
rect 17325 5729 17359 5763
rect 17601 5729 17635 5763
rect 17969 5729 18003 5763
rect 18337 5729 18371 5763
rect 19752 5729 19786 5763
rect 20913 5729 20947 5763
rect 24133 5729 24167 5763
rect 24593 5729 24627 5763
rect 24961 5729 24995 5763
rect 25513 5729 25547 5763
rect 26801 5729 26835 5763
rect 26985 5729 27019 5763
rect 27353 5729 27387 5763
rect 27721 5729 27755 5763
rect 28825 5729 28859 5763
rect 2053 5661 2087 5695
rect 4537 5661 4571 5695
rect 25605 5661 25639 5695
rect 27997 5661 28031 5695
rect 2605 5593 2639 5627
rect 7573 5593 7607 5627
rect 18521 5593 18555 5627
rect 1685 5525 1719 5559
rect 5089 5525 5123 5559
rect 5733 5525 5767 5559
rect 6101 5525 6135 5559
rect 8631 5525 8665 5559
rect 9505 5525 9539 5559
rect 14381 5525 14415 5559
rect 17049 5525 17083 5559
rect 19855 5525 19889 5559
rect 20637 5525 20671 5559
rect 21833 5525 21867 5559
rect 25881 5525 25915 5559
rect 29745 5525 29779 5559
rect 30941 5525 30975 5559
rect 2513 5321 2547 5355
rect 2605 5321 2639 5355
rect 3249 5321 3283 5355
rect 4353 5321 4387 5355
rect 6285 5321 6319 5355
rect 7757 5321 7791 5355
rect 9965 5321 9999 5355
rect 12173 5321 12207 5355
rect 15853 5321 15887 5355
rect 16221 5321 16255 5355
rect 17509 5321 17543 5355
rect 19349 5321 19383 5355
rect 19717 5321 19751 5355
rect 20453 5321 20487 5355
rect 22661 5321 22695 5355
rect 24133 5321 24167 5355
rect 25145 5321 25179 5355
rect 30665 5321 30699 5355
rect 1593 5185 1627 5219
rect 8033 5253 8067 5287
rect 24501 5253 24535 5287
rect 27169 5253 27203 5287
rect 3479 5185 3513 5219
rect 3893 5185 3927 5219
rect 6837 5185 6871 5219
rect 13645 5185 13679 5219
rect 17141 5185 17175 5219
rect 22293 5185 22327 5219
rect 27445 5185 27479 5219
rect 27721 5185 27755 5219
rect 28365 5185 28399 5219
rect 30021 5185 30055 5219
rect 31217 5185 31251 5219
rect 3392 5117 3426 5151
rect 4721 5117 4755 5151
rect 5181 5117 5215 5151
rect 5457 5117 5491 5151
rect 5825 5117 5859 5151
rect 8953 5117 8987 5151
rect 9080 5117 9114 5151
rect 9597 5117 9631 5151
rect 10333 5117 10367 5151
rect 10701 5117 10735 5151
rect 10885 5117 10919 5151
rect 11253 5117 11287 5151
rect 14013 5117 14047 5151
rect 14381 5117 14415 5151
rect 14749 5117 14783 5151
rect 14933 5117 14967 5151
rect 15301 5117 15335 5151
rect 16497 5117 16531 5151
rect 18061 5117 18095 5151
rect 20729 5117 20763 5151
rect 21005 5117 21039 5151
rect 21373 5117 21407 5151
rect 21741 5117 21775 5151
rect 25329 5117 25363 5151
rect 25789 5117 25823 5151
rect 26157 5117 26191 5151
rect 26525 5117 26559 5151
rect 1914 5049 1948 5083
rect 2605 5049 2639 5083
rect 2881 5049 2915 5083
rect 7158 5049 7192 5083
rect 11529 5049 11563 5083
rect 12633 5049 12667 5083
rect 12725 5049 12759 5083
rect 13277 5049 13311 5083
rect 18382 5049 18416 5083
rect 26801 5049 26835 5083
rect 27813 5049 27847 5083
rect 29377 5049 29411 5083
rect 29469 5049 29503 5083
rect 30941 5049 30975 5083
rect 31033 5049 31067 5083
rect 5641 4981 5675 5015
rect 6561 4981 6595 5015
rect 8585 4981 8619 5015
rect 9183 4981 9217 5015
rect 11897 4981 11931 5015
rect 15301 4981 15335 5015
rect 17785 4981 17819 5015
rect 18981 4981 19015 5015
rect 20821 4981 20855 5015
rect 23489 4981 23523 5015
rect 28825 4981 28859 5015
rect 30297 4981 30331 5015
rect 2789 4777 2823 4811
rect 5089 4777 5123 4811
rect 5549 4777 5583 4811
rect 6929 4777 6963 4811
rect 7849 4777 7883 4811
rect 9505 4777 9539 4811
rect 15025 4777 15059 4811
rect 15485 4777 15519 4811
rect 20545 4777 20579 4811
rect 25329 4777 25363 4811
rect 26709 4777 26743 4811
rect 29837 4777 29871 4811
rect 1822 4709 1856 4743
rect 3893 4709 3927 4743
rect 7481 4709 7515 4743
rect 8217 4709 8251 4743
rect 10149 4709 10183 4743
rect 12633 4709 12667 4743
rect 13823 4709 13857 4743
rect 14657 4709 14691 4743
rect 16313 4709 16347 4743
rect 18245 4709 18279 4743
rect 18521 4709 18555 4743
rect 19349 4709 19383 4743
rect 19441 4709 19475 4743
rect 21275 4709 21309 4743
rect 22845 4709 22879 4743
rect 24869 4709 24903 4743
rect 25697 4709 25731 4743
rect 26249 4709 26283 4743
rect 27214 4709 27248 4743
rect 28962 4709 28996 4743
rect 30573 4709 30607 4743
rect 4261 4641 4295 4675
rect 5733 4641 5767 4675
rect 6193 4641 6227 4675
rect 6561 4641 6595 4675
rect 7113 4641 7147 4675
rect 10517 4641 10551 4675
rect 10977 4641 11011 4675
rect 11161 4641 11195 4675
rect 11437 4641 11471 4675
rect 13461 4641 13495 4675
rect 15301 4641 15335 4675
rect 16681 4641 16715 4675
rect 17049 4641 17083 4675
rect 17417 4641 17451 4675
rect 17601 4641 17635 4675
rect 17969 4641 18003 4675
rect 20913 4641 20947 4675
rect 24225 4641 24259 4675
rect 27813 4641 27847 4675
rect 1501 4573 1535 4607
rect 8125 4573 8159 4607
rect 8493 4573 8527 4607
rect 12265 4573 12299 4607
rect 19993 4573 20027 4607
rect 22753 4573 22787 4607
rect 23029 4573 23063 4607
rect 26893 4573 26927 4607
rect 28641 4573 28675 4607
rect 30481 4573 30515 4607
rect 30757 4573 30791 4607
rect 11621 4505 11655 4539
rect 13001 4505 13035 4539
rect 13369 4505 13403 4539
rect 14381 4505 14415 4539
rect 15853 4505 15887 4539
rect 24409 4505 24443 4539
rect 2421 4437 2455 4471
rect 4353 4437 4387 4471
rect 21833 4437 21867 4471
rect 23673 4437 23707 4471
rect 28181 4437 28215 4471
rect 28549 4437 28583 4471
rect 29561 4437 29595 4471
rect 1685 4233 1719 4267
rect 4537 4233 4571 4267
rect 6561 4233 6595 4267
rect 8125 4233 8159 4267
rect 10609 4233 10643 4267
rect 10977 4233 11011 4267
rect 15485 4233 15519 4267
rect 15853 4233 15887 4267
rect 16957 4233 16991 4267
rect 19717 4233 19751 4267
rect 21005 4233 21039 4267
rect 22845 4233 22879 4267
rect 25145 4233 25179 4267
rect 28641 4233 28675 4267
rect 30665 4233 30699 4267
rect 26709 4165 26743 4199
rect 1869 4097 1903 4131
rect 3709 4097 3743 4131
rect 5917 4097 5951 4131
rect 6837 4097 6871 4131
rect 8401 4097 8435 4131
rect 8953 4097 8987 4131
rect 9413 4097 9447 4131
rect 11621 4097 11655 4131
rect 12449 4097 12483 4131
rect 14197 4097 14231 4131
rect 16313 4097 16347 4131
rect 17417 4097 17451 4131
rect 18153 4097 18187 4131
rect 21281 4097 21315 4131
rect 22477 4097 22511 4131
rect 24041 4097 24075 4131
rect 29377 4097 29411 4131
rect 30987 4097 31021 4131
rect 6285 4029 6319 4063
rect 11412 4029 11446 4063
rect 1961 3961 1995 3995
rect 2513 3961 2547 3995
rect 3433 3961 3467 3995
rect 3525 3961 3559 3995
rect 5273 3961 5307 3995
rect 5365 3961 5399 3995
rect 7158 3961 7192 3995
rect 9229 3961 9263 3995
rect 9734 3961 9768 3995
rect 15117 4029 15151 4063
rect 19952 4029 19986 4063
rect 25605 4029 25639 4063
rect 25881 4029 25915 4063
rect 26157 4029 26191 4063
rect 26525 4029 26559 4063
rect 28365 4029 28399 4063
rect 30389 4029 30423 4063
rect 30884 4029 30918 4063
rect 31309 4029 31343 4063
rect 12811 3961 12845 3995
rect 13645 3961 13679 3995
rect 14105 3961 14139 3995
rect 14559 3961 14593 3995
rect 16037 3961 16071 3995
rect 16129 3961 16163 3995
rect 17877 3961 17911 3995
rect 18515 3961 18549 3995
rect 20039 3961 20073 3995
rect 21602 3961 21636 3995
rect 23765 3961 23799 3995
rect 23857 3961 23891 3995
rect 27721 3961 27755 3995
rect 27813 3961 27847 3995
rect 29469 3961 29503 3995
rect 30021 3961 30055 3995
rect 2789 3893 2823 3927
rect 3249 3893 3283 3927
rect 5089 3893 5123 3927
rect 7757 3893 7791 3927
rect 10333 3893 10367 3927
rect 11483 3893 11517 3927
rect 11621 3893 11655 3927
rect 11897 3893 11931 3927
rect 12265 3893 12299 3927
rect 13369 3893 13403 3927
rect 19073 3893 19107 3927
rect 19441 3893 19475 3927
rect 20453 3893 20487 3927
rect 22201 3893 22235 3927
rect 23397 3893 23431 3927
rect 24685 3893 24719 3927
rect 27077 3893 27111 3927
rect 27445 3893 27479 3927
rect 29101 3893 29135 3927
rect 2513 3689 2547 3723
rect 2973 3689 3007 3723
rect 3433 3689 3467 3723
rect 4261 3689 4295 3723
rect 5089 3689 5123 3723
rect 5457 3689 5491 3723
rect 6837 3689 6871 3723
rect 9505 3689 9539 3723
rect 10701 3689 10735 3723
rect 12081 3689 12115 3723
rect 13645 3689 13679 3723
rect 14657 3689 14691 3723
rect 16773 3689 16807 3723
rect 18245 3689 18279 3723
rect 20729 3689 20763 3723
rect 21281 3689 21315 3723
rect 22753 3689 22787 3723
rect 25421 3689 25455 3723
rect 27721 3689 27755 3723
rect 29975 3689 30009 3723
rect 30481 3689 30515 3723
rect 30987 3689 31021 3723
rect 1593 3621 1627 3655
rect 1685 3621 1719 3655
rect 3893 3621 3927 3655
rect 5870 3621 5904 3655
rect 7481 3621 7515 3655
rect 10241 3621 10275 3655
rect 11206 3621 11240 3655
rect 12725 3621 12759 3655
rect 12817 3621 12851 3655
rect 15663 3621 15697 3655
rect 17233 3621 17267 3655
rect 19441 3621 19475 3655
rect 19993 3621 20027 3655
rect 21925 3621 21959 3655
rect 25697 3621 25731 3655
rect 26846 3621 26880 3655
rect 28457 3621 28491 3655
rect 4604 3553 4638 3587
rect 5549 3553 5583 3587
rect 9689 3553 9723 3587
rect 10885 3553 10919 3587
rect 12449 3553 12483 3587
rect 14232 3553 14266 3587
rect 15301 3553 15335 3587
rect 23340 3553 23374 3587
rect 26065 3553 26099 3587
rect 27445 3553 27479 3587
rect 29872 3553 29906 3587
rect 30916 3553 30950 3587
rect 2237 3485 2271 3519
rect 7389 3485 7423 3519
rect 8033 3485 8067 3519
rect 8309 3485 8343 3519
rect 13369 3485 13403 3519
rect 17141 3485 17175 3519
rect 17417 3485 17451 3519
rect 19349 3485 19383 3519
rect 21833 3485 21867 3519
rect 23443 3485 23477 3519
rect 26525 3485 26559 3519
rect 28365 3485 28399 3519
rect 9873 3417 9907 3451
rect 14335 3417 14369 3451
rect 22385 3417 22419 3451
rect 28917 3417 28951 3451
rect 4675 3349 4709 3383
rect 6469 3349 6503 3383
rect 11805 3349 11839 3383
rect 14013 3349 14047 3383
rect 15025 3349 15059 3383
rect 16221 3349 16255 3383
rect 20269 3349 20303 3383
rect 28089 3349 28123 3383
rect 29561 3349 29595 3383
rect 2881 3145 2915 3179
rect 4721 3145 4755 3179
rect 4905 3145 4939 3179
rect 6193 3145 6227 3179
rect 8309 3145 8343 3179
rect 10885 3145 10919 3179
rect 12081 3145 12115 3179
rect 13369 3145 13403 3179
rect 14473 3145 14507 3179
rect 16405 3145 16439 3179
rect 17417 3145 17451 3179
rect 17785 3145 17819 3179
rect 18613 3145 18647 3179
rect 19533 3145 19567 3179
rect 22293 3145 22327 3179
rect 26893 3145 26927 3179
rect 27215 3145 27249 3179
rect 27997 3145 28031 3179
rect 29009 3145 29043 3179
rect 30113 3145 30147 3179
rect 30941 3145 30975 3179
rect 2237 3009 2271 3043
rect 2513 3009 2547 3043
rect 5825 3077 5859 3111
rect 7481 3077 7515 3111
rect 14105 3077 14139 3111
rect 16129 3077 16163 3111
rect 18843 3077 18877 3111
rect 21925 3077 21959 3111
rect 26617 3077 26651 3111
rect 29745 3077 29779 3111
rect 6561 3009 6595 3043
rect 6929 3009 6963 3043
rect 9689 3009 9723 3043
rect 10333 3009 10367 3043
rect 11805 3009 11839 3043
rect 13553 3009 13587 3043
rect 15117 3009 15151 3043
rect 15393 3009 15427 3043
rect 19809 3009 19843 3043
rect 20269 3009 20303 3043
rect 21373 3009 21407 3043
rect 22661 3009 22695 3043
rect 2053 2941 2087 2975
rect 3525 2941 3559 2975
rect 3709 2941 3743 2975
rect 4905 2941 4939 2975
rect 8401 2941 8435 2975
rect 8953 2941 8987 2975
rect 9505 2941 9539 2975
rect 11161 2941 11195 2975
rect 12516 2941 12550 2975
rect 16656 2941 16690 2975
rect 17049 2941 17083 2975
rect 18772 2941 18806 2975
rect 23305 2941 23339 2975
rect 27112 2941 27146 2975
rect 27537 2941 27571 2975
rect 28089 2941 28123 2975
rect 28641 2941 28675 2975
rect 29561 2941 29595 2975
rect 4353 2873 4387 2907
rect 4997 2873 5031 2907
rect 5273 2873 5307 2907
rect 5365 2873 5399 2907
rect 7021 2873 7055 2907
rect 9781 2873 9815 2907
rect 13001 2873 13035 2907
rect 13645 2873 13679 2907
rect 15209 2873 15243 2907
rect 19901 2873 19935 2907
rect 20729 2873 20763 2907
rect 21465 2873 21499 2907
rect 7849 2805 7883 2839
rect 8585 2805 8619 2839
rect 11345 2805 11379 2839
rect 12587 2805 12621 2839
rect 14933 2805 14967 2839
rect 16727 2805 16761 2839
rect 19165 2805 19199 2839
rect 21189 2805 21223 2839
rect 28273 2805 28307 2839
rect 1639 2601 1673 2635
rect 3065 2601 3099 2635
rect 3893 2601 3927 2635
rect 4353 2601 4387 2635
rect 6285 2601 6319 2635
rect 9597 2601 9631 2635
rect 13737 2601 13771 2635
rect 14335 2601 14369 2635
rect 15117 2601 15151 2635
rect 19441 2601 19475 2635
rect 21327 2601 21361 2635
rect 22109 2601 22143 2635
rect 22339 2601 22373 2635
rect 27675 2601 27709 2635
rect 28733 2601 28767 2635
rect 31585 2601 31619 2635
rect 32781 2601 32815 2635
rect 2329 2533 2363 2567
rect 7389 2533 7423 2567
rect 7941 2533 7975 2567
rect 10885 2533 10919 2567
rect 11161 2533 11195 2567
rect 11713 2533 11747 2567
rect 12449 2533 12483 2567
rect 12817 2533 12851 2567
rect 13369 2533 13403 2567
rect 14657 2533 14691 2567
rect 19073 2533 19107 2567
rect 19625 2533 19659 2567
rect 19717 2533 19751 2567
rect 20269 2533 20303 2567
rect 1568 2465 1602 2499
rect 2053 2465 2087 2499
rect 2881 2465 2915 2499
rect 4169 2465 4203 2499
rect 5181 2465 5215 2499
rect 5917 2465 5951 2499
rect 9781 2465 9815 2499
rect 10425 2465 10459 2499
rect 14264 2465 14298 2499
rect 15520 2465 15554 2499
rect 15945 2465 15979 2499
rect 21256 2465 21290 2499
rect 22268 2465 22302 2499
rect 22753 2465 22787 2499
rect 27604 2465 27638 2499
rect 27997 2465 28031 2499
rect 28549 2465 28583 2499
rect 29101 2465 29135 2499
rect 30297 2465 30331 2499
rect 30849 2465 30883 2499
rect 31401 2465 31435 2499
rect 31953 2465 31987 2499
rect 32597 2465 32631 2499
rect 33149 2465 33183 2499
rect 3525 2397 3559 2431
rect 6009 2397 6043 2431
rect 6653 2397 6687 2431
rect 7297 2397 7331 2431
rect 11069 2397 11103 2431
rect 12725 2397 12759 2431
rect 14013 2397 14047 2431
rect 4813 2261 4847 2295
rect 8309 2261 8343 2295
rect 9965 2261 9999 2295
rect 12081 2261 12115 2295
rect 15623 2261 15657 2295
rect 21741 2261 21775 2295
rect 30481 2261 30515 2295
<< metal1 >>
rect 3418 13812 3424 13864
rect 3476 13852 3482 13864
rect 19334 13852 19340 13864
rect 3476 13824 19340 13852
rect 3476 13812 3482 13824
rect 19334 13812 19340 13824
rect 19392 13812 19398 13864
rect 1104 13626 38824 13648
rect 1104 13574 14315 13626
rect 14367 13574 14379 13626
rect 14431 13574 14443 13626
rect 14495 13574 14507 13626
rect 14559 13574 27648 13626
rect 27700 13574 27712 13626
rect 27764 13574 27776 13626
rect 27828 13574 27840 13626
rect 27892 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 7648 13082
rect 7700 13030 7712 13082
rect 7764 13030 7776 13082
rect 7828 13030 7840 13082
rect 7892 13030 20982 13082
rect 21034 13030 21046 13082
rect 21098 13030 21110 13082
rect 21162 13030 21174 13082
rect 21226 13030 34315 13082
rect 34367 13030 34379 13082
rect 34431 13030 34443 13082
rect 34495 13030 34507 13082
rect 34559 13030 38824 13082
rect 1104 13008 38824 13030
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 16206 12628 16212 12640
rect 15252 12600 16212 12628
rect 15252 12588 15258 12600
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 1104 12538 38824 12560
rect 1104 12486 14315 12538
rect 14367 12486 14379 12538
rect 14431 12486 14443 12538
rect 14495 12486 14507 12538
rect 14559 12486 27648 12538
rect 27700 12486 27712 12538
rect 27764 12486 27776 12538
rect 27828 12486 27840 12538
rect 27892 12486 38824 12538
rect 1104 12464 38824 12486
rect 1104 11994 38824 12016
rect 1104 11942 7648 11994
rect 7700 11942 7712 11994
rect 7764 11942 7776 11994
rect 7828 11942 7840 11994
rect 7892 11942 20982 11994
rect 21034 11942 21046 11994
rect 21098 11942 21110 11994
rect 21162 11942 21174 11994
rect 21226 11942 34315 11994
rect 34367 11942 34379 11994
rect 34431 11942 34443 11994
rect 34495 11942 34507 11994
rect 34559 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 14315 11450
rect 14367 11398 14379 11450
rect 14431 11398 14443 11450
rect 14495 11398 14507 11450
rect 14559 11398 27648 11450
rect 27700 11398 27712 11450
rect 27764 11398 27776 11450
rect 27828 11398 27840 11450
rect 27892 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 7648 10906
rect 7700 10854 7712 10906
rect 7764 10854 7776 10906
rect 7828 10854 7840 10906
rect 7892 10854 20982 10906
rect 21034 10854 21046 10906
rect 21098 10854 21110 10906
rect 21162 10854 21174 10906
rect 21226 10854 34315 10906
rect 34367 10854 34379 10906
rect 34431 10854 34443 10906
rect 34495 10854 34507 10906
rect 34559 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 14315 10362
rect 14367 10310 14379 10362
rect 14431 10310 14443 10362
rect 14495 10310 14507 10362
rect 14559 10310 27648 10362
rect 27700 10310 27712 10362
rect 27764 10310 27776 10362
rect 27828 10310 27840 10362
rect 27892 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 7648 9818
rect 7700 9766 7712 9818
rect 7764 9766 7776 9818
rect 7828 9766 7840 9818
rect 7892 9766 20982 9818
rect 21034 9766 21046 9818
rect 21098 9766 21110 9818
rect 21162 9766 21174 9818
rect 21226 9766 34315 9818
rect 34367 9766 34379 9818
rect 34431 9766 34443 9818
rect 34495 9766 34507 9818
rect 34559 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 14315 9274
rect 14367 9222 14379 9274
rect 14431 9222 14443 9274
rect 14495 9222 14507 9274
rect 14559 9222 27648 9274
rect 27700 9222 27712 9274
rect 27764 9222 27776 9274
rect 27828 9222 27840 9274
rect 27892 9222 38824 9274
rect 1104 9200 38824 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 1946 9024 1952 9036
rect 1443 8996 1952 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 9024 6515 9027
rect 6546 9024 6552 9036
rect 6503 8996 6552 9024
rect 6503 8993 6515 8996
rect 6457 8987 6515 8993
rect 6546 8984 6552 8996
rect 6604 8984 6610 9036
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6512 8792 6653 8820
rect 6512 8780 6518 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6641 8783 6699 8789
rect 1104 8730 38824 8752
rect 1104 8678 7648 8730
rect 7700 8678 7712 8730
rect 7764 8678 7776 8730
rect 7828 8678 7840 8730
rect 7892 8678 20982 8730
rect 21034 8678 21046 8730
rect 21098 8678 21110 8730
rect 21162 8678 21174 8730
rect 21226 8678 34315 8730
rect 34367 8678 34379 8730
rect 34431 8678 34443 8730
rect 34495 8678 34507 8730
rect 34559 8678 38824 8730
rect 1104 8656 38824 8678
rect 1394 8576 1400 8628
rect 1452 8616 1458 8628
rect 1535 8619 1593 8625
rect 1535 8616 1547 8619
rect 1452 8588 1547 8616
rect 1452 8576 1458 8588
rect 1535 8585 1547 8588
rect 1581 8585 1593 8619
rect 1535 8579 1593 8585
rect 19334 8576 19340 8628
rect 19392 8616 19398 8628
rect 20487 8619 20545 8625
rect 20487 8616 20499 8619
rect 19392 8588 20499 8616
rect 19392 8576 19398 8588
rect 20487 8585 20499 8588
rect 20533 8585 20545 8619
rect 20487 8579 20545 8585
rect 6914 8508 6920 8560
rect 6972 8557 6978 8560
rect 6972 8551 7021 8557
rect 6972 8517 6975 8551
rect 7009 8517 7021 8551
rect 6972 8511 7021 8517
rect 6972 8508 6978 8511
rect 2314 8480 2320 8492
rect 2275 8452 2320 8480
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 1464 8415 1522 8421
rect 1464 8381 1476 8415
rect 1510 8412 1522 8415
rect 2332 8412 2360 8440
rect 1510 8384 2360 8412
rect 6892 8415 6950 8421
rect 1510 8381 1522 8384
rect 1464 8375 1522 8381
rect 6892 8381 6904 8415
rect 6938 8412 6950 8415
rect 16301 8415 16359 8421
rect 6938 8384 7236 8412
rect 6938 8381 6950 8384
rect 6892 8375 6950 8381
rect 7208 8356 7236 8384
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 17034 8412 17040 8424
rect 16347 8384 17040 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 17034 8372 17040 8384
rect 17092 8372 17098 8424
rect 20416 8415 20474 8421
rect 20416 8381 20428 8415
rect 20462 8412 20474 8415
rect 20462 8384 20944 8412
rect 20462 8381 20474 8384
rect 20416 8375 20474 8381
rect 1946 8344 1952 8356
rect 1907 8316 1952 8344
rect 1946 8304 1952 8316
rect 2004 8304 2010 8356
rect 6546 8344 6552 8356
rect 6507 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 7190 8304 7196 8356
rect 7248 8344 7254 8356
rect 20916 8353 20944 8384
rect 7285 8347 7343 8353
rect 7285 8344 7297 8347
rect 7248 8316 7297 8344
rect 7248 8304 7254 8316
rect 7285 8313 7297 8316
rect 7331 8313 7343 8347
rect 7285 8307 7343 8313
rect 20901 8347 20959 8353
rect 20901 8313 20913 8347
rect 20947 8344 20959 8347
rect 20947 8316 22140 8344
rect 20947 8313 20959 8316
rect 20901 8307 20959 8313
rect 16666 8276 16672 8288
rect 16627 8248 16672 8276
rect 16666 8236 16672 8248
rect 16724 8236 16730 8288
rect 22112 8276 22140 8316
rect 22554 8276 22560 8288
rect 22112 8248 22560 8276
rect 22554 8236 22560 8248
rect 22612 8236 22618 8288
rect 1104 8186 38824 8208
rect 1104 8134 14315 8186
rect 14367 8134 14379 8186
rect 14431 8134 14443 8186
rect 14495 8134 14507 8186
rect 14559 8134 27648 8186
rect 27700 8134 27712 8186
rect 27764 8134 27776 8186
rect 27828 8134 27840 8186
rect 27892 8134 38824 8186
rect 1104 8112 38824 8134
rect 1578 8072 1584 8084
rect 1539 8044 1584 8072
rect 1578 8032 1584 8044
rect 1636 8032 1642 8084
rect 16301 8075 16359 8081
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16574 8072 16580 8084
rect 16347 8044 16580 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16574 8032 16580 8044
rect 16632 8072 16638 8084
rect 17862 8072 17868 8084
rect 16632 8044 17868 8072
rect 16632 8032 16638 8044
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 35618 8072 35624 8084
rect 35579 8044 35624 8072
rect 35618 8032 35624 8044
rect 35676 8032 35682 8084
rect 5258 7964 5264 8016
rect 5316 8004 5322 8016
rect 7006 8004 7012 8016
rect 5316 7976 7012 8004
rect 5316 7964 5322 7976
rect 7006 7964 7012 7976
rect 7064 7964 7070 8016
rect 16666 8004 16672 8016
rect 16627 7976 16672 8004
rect 16666 7964 16672 7976
rect 16724 7964 16730 8016
rect 19794 7964 19800 8016
rect 19852 8004 19858 8016
rect 21266 8013 21272 8016
rect 21222 8007 21272 8013
rect 21222 8004 21234 8007
rect 19852 7976 21234 8004
rect 19852 7964 19858 7976
rect 21222 7973 21234 7976
rect 21268 7973 21272 8007
rect 21222 7967 21272 7973
rect 21266 7964 21272 7967
rect 21324 8004 21330 8016
rect 28353 8007 28411 8013
rect 21324 7976 21370 8004
rect 21324 7964 21330 7976
rect 28353 7973 28365 8007
rect 28399 8004 28411 8007
rect 28718 8004 28724 8016
rect 28399 7976 28724 8004
rect 28399 7973 28411 7976
rect 28353 7967 28411 7973
rect 28718 7964 28724 7976
rect 28776 7964 28782 8016
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7936 1455 7939
rect 1854 7936 1860 7948
rect 1443 7908 1860 7936
rect 1443 7905 1455 7908
rect 1397 7899 1455 7905
rect 1854 7896 1860 7908
rect 1912 7896 1918 7948
rect 5880 7939 5938 7945
rect 5880 7905 5892 7939
rect 5926 7936 5938 7939
rect 6086 7936 6092 7948
rect 5926 7908 6092 7936
rect 5926 7905 5938 7908
rect 5880 7899 5938 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 13173 7939 13231 7945
rect 13173 7905 13185 7939
rect 13219 7936 13231 7939
rect 13630 7936 13636 7948
rect 13219 7908 13636 7936
rect 13219 7905 13231 7908
rect 13173 7899 13231 7905
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 14182 7936 14188 7948
rect 14143 7908 14188 7936
rect 14182 7896 14188 7908
rect 14240 7896 14246 7948
rect 15654 7936 15660 7948
rect 15615 7908 15660 7936
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 17126 7936 17132 7948
rect 17087 7908 17132 7936
rect 17126 7896 17132 7908
rect 17184 7896 17190 7948
rect 35434 7936 35440 7948
rect 35395 7908 35440 7936
rect 35434 7896 35440 7908
rect 35492 7896 35498 7948
rect 6917 7871 6975 7877
rect 6917 7837 6929 7871
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 5951 7803 6009 7809
rect 5951 7769 5963 7803
rect 5997 7800 6009 7803
rect 6730 7800 6736 7812
rect 5997 7772 6736 7800
rect 5997 7769 6009 7772
rect 5951 7763 6009 7769
rect 6730 7760 6736 7772
rect 6788 7760 6794 7812
rect 5258 7732 5264 7744
rect 5219 7704 5264 7732
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 6638 7732 6644 7744
rect 6599 7704 6644 7732
rect 6638 7692 6644 7704
rect 6696 7732 6702 7744
rect 6932 7732 6960 7831
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 7156 7840 7205 7868
rect 7156 7828 7162 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7868 20775 7871
rect 20806 7868 20812 7880
rect 20763 7840 20812 7868
rect 20763 7837 20775 7840
rect 20717 7831 20775 7837
rect 20806 7828 20812 7840
rect 20864 7868 20870 7880
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 20864 7840 20913 7868
rect 20864 7828 20870 7840
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7868 28319 7871
rect 28442 7868 28448 7880
rect 28307 7840 28448 7868
rect 28307 7837 28319 7840
rect 28261 7831 28319 7837
rect 28442 7828 28448 7840
rect 28500 7828 28506 7880
rect 28902 7868 28908 7880
rect 28863 7840 28908 7868
rect 28902 7828 28908 7840
rect 28960 7828 28966 7880
rect 6696 7704 6960 7732
rect 13357 7735 13415 7741
rect 6696 7692 6702 7704
rect 13357 7701 13369 7735
rect 13403 7732 13415 7735
rect 13722 7732 13728 7744
rect 13403 7704 13728 7732
rect 13403 7701 13415 7704
rect 13357 7695 13415 7701
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 14369 7735 14427 7741
rect 14369 7732 14381 7735
rect 13872 7704 14381 7732
rect 13872 7692 13878 7704
rect 14369 7701 14381 7704
rect 14415 7701 14427 7735
rect 14369 7695 14427 7701
rect 15841 7735 15899 7741
rect 15841 7701 15853 7735
rect 15887 7732 15899 7735
rect 16390 7732 16396 7744
rect 15887 7704 16396 7732
rect 15887 7701 15899 7704
rect 15841 7695 15899 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17310 7732 17316 7744
rect 17271 7704 17316 7732
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 19518 7732 19524 7744
rect 19479 7704 19524 7732
rect 19518 7692 19524 7704
rect 19576 7692 19582 7744
rect 21821 7735 21879 7741
rect 21821 7701 21833 7735
rect 21867 7732 21879 7735
rect 22002 7732 22008 7744
rect 21867 7704 22008 7732
rect 21867 7701 21879 7704
rect 21821 7695 21879 7701
rect 22002 7692 22008 7704
rect 22060 7732 22066 7744
rect 22097 7735 22155 7741
rect 22097 7732 22109 7735
rect 22060 7704 22109 7732
rect 22060 7692 22066 7704
rect 22097 7701 22109 7704
rect 22143 7701 22155 7735
rect 22097 7695 22155 7701
rect 25317 7735 25375 7741
rect 25317 7701 25329 7735
rect 25363 7732 25375 7735
rect 26050 7732 26056 7744
rect 25363 7704 26056 7732
rect 25363 7701 25375 7704
rect 25317 7695 25375 7701
rect 26050 7692 26056 7704
rect 26108 7692 26114 7744
rect 1104 7642 38824 7664
rect 1104 7590 7648 7642
rect 7700 7590 7712 7642
rect 7764 7590 7776 7642
rect 7828 7590 7840 7642
rect 7892 7590 20982 7642
rect 21034 7590 21046 7642
rect 21098 7590 21110 7642
rect 21162 7590 21174 7642
rect 21226 7590 34315 7642
rect 34367 7590 34379 7642
rect 34431 7590 34443 7642
rect 34495 7590 34507 7642
rect 34559 7590 38824 7642
rect 1104 7568 38824 7590
rect 1854 7528 1860 7540
rect 1815 7500 1860 7528
rect 1854 7488 1860 7500
rect 1912 7528 1918 7540
rect 2222 7528 2228 7540
rect 1912 7500 2228 7528
rect 1912 7488 1918 7500
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7745 7531 7803 7537
rect 7745 7528 7757 7531
rect 7064 7500 7757 7528
rect 7064 7488 7070 7500
rect 7745 7497 7757 7500
rect 7791 7528 7803 7531
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 7791 7500 8033 7528
rect 7791 7497 7803 7500
rect 7745 7491 7803 7497
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7528 16175 7531
rect 16347 7531 16405 7537
rect 16347 7528 16359 7531
rect 16163 7500 16359 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16347 7497 16359 7500
rect 16393 7528 16405 7531
rect 16942 7528 16948 7540
rect 16393 7500 16948 7528
rect 16393 7497 16405 7500
rect 16347 7491 16405 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 17184 7500 17233 7528
rect 17184 7488 17190 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 21266 7528 21272 7540
rect 21227 7500 21272 7528
rect 17221 7491 17279 7497
rect 21266 7488 21272 7500
rect 21324 7488 21330 7540
rect 28442 7528 28448 7540
rect 28403 7500 28448 7528
rect 28442 7488 28448 7500
rect 28500 7488 28506 7540
rect 28718 7488 28724 7540
rect 28776 7528 28782 7540
rect 28813 7531 28871 7537
rect 28813 7528 28825 7531
rect 28776 7500 28825 7528
rect 28776 7488 28782 7500
rect 28813 7497 28825 7500
rect 28859 7497 28871 7531
rect 28813 7491 28871 7497
rect 28994 7488 29000 7540
rect 29052 7528 29058 7540
rect 29411 7531 29469 7537
rect 29411 7528 29423 7531
rect 29052 7500 29423 7528
rect 29052 7488 29058 7500
rect 29411 7497 29423 7500
rect 29457 7497 29469 7531
rect 29411 7491 29469 7497
rect 15746 7460 15752 7472
rect 15659 7432 15752 7460
rect 15746 7420 15752 7432
rect 15804 7460 15810 7472
rect 16482 7460 16488 7472
rect 15804 7432 16488 7460
rect 15804 7420 15810 7432
rect 16482 7420 16488 7432
rect 16540 7420 16546 7472
rect 16574 7392 16580 7404
rect 15304 7364 16580 7392
rect 5258 7324 5264 7336
rect 5219 7296 5264 7324
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 8573 7327 8631 7333
rect 7024 7296 7236 7324
rect 5905 7259 5963 7265
rect 5905 7225 5917 7259
rect 5951 7256 5963 7259
rect 6914 7256 6920 7268
rect 5951 7228 6920 7256
rect 5951 7225 5963 7228
rect 5905 7219 5963 7225
rect 6914 7216 6920 7228
rect 6972 7216 6978 7268
rect 1397 7191 1455 7197
rect 1397 7157 1409 7191
rect 1443 7188 1455 7191
rect 1486 7188 1492 7200
rect 1443 7160 1492 7188
rect 1443 7157 1455 7160
rect 1397 7151 1455 7157
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 4525 7191 4583 7197
rect 4525 7157 4537 7191
rect 4571 7188 4583 7191
rect 5074 7188 5080 7200
rect 4571 7160 5080 7188
rect 4571 7157 4583 7160
rect 4525 7151 4583 7157
rect 5074 7148 5080 7160
rect 5132 7148 5138 7200
rect 6086 7148 6092 7200
rect 6144 7188 6150 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 6144 7160 6193 7188
rect 6144 7148 6150 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 6546 7188 6552 7200
rect 6507 7160 6552 7188
rect 6181 7151 6239 7157
rect 6546 7148 6552 7160
rect 6604 7188 6610 7200
rect 7024 7188 7052 7296
rect 7208 7265 7236 7296
rect 8573 7293 8585 7327
rect 8619 7324 8631 7327
rect 12253 7327 12311 7333
rect 8619 7296 9168 7324
rect 8619 7293 8631 7296
rect 8573 7287 8631 7293
rect 7187 7259 7245 7265
rect 7187 7225 7199 7259
rect 7233 7225 7245 7259
rect 7187 7219 7245 7225
rect 9140 7200 9168 7296
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 13078 7324 13084 7336
rect 12299 7296 13084 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 14734 7284 14740 7336
rect 14792 7324 14798 7336
rect 15304 7333 15332 7364
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 19518 7352 19524 7404
rect 19576 7392 19582 7404
rect 19576 7364 20392 7392
rect 19576 7352 19582 7364
rect 15289 7327 15347 7333
rect 15289 7324 15301 7327
rect 14792 7296 15301 7324
rect 14792 7284 14798 7296
rect 15289 7293 15301 7296
rect 15335 7293 15347 7327
rect 15289 7287 15347 7293
rect 16298 7284 16304 7336
rect 16356 7324 16362 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 16356 7296 18061 7324
rect 16356 7284 16362 7296
rect 18049 7293 18061 7296
rect 18095 7324 18107 7327
rect 18506 7324 18512 7336
rect 18095 7296 18512 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 19797 7327 19855 7333
rect 19797 7293 19809 7327
rect 19843 7293 19855 7327
rect 19978 7324 19984 7336
rect 19939 7296 19984 7324
rect 19797 7287 19855 7293
rect 13170 7256 13176 7268
rect 13131 7228 13176 7256
rect 13170 7216 13176 7228
rect 13228 7216 13234 7268
rect 14182 7216 14188 7268
rect 14240 7256 14246 7268
rect 14277 7259 14335 7265
rect 14277 7256 14289 7259
rect 14240 7228 14289 7256
rect 14240 7216 14246 7228
rect 14277 7225 14289 7228
rect 14323 7256 14335 7259
rect 14826 7256 14832 7268
rect 14323 7228 14832 7256
rect 14323 7225 14335 7228
rect 14277 7219 14335 7225
rect 14826 7216 14832 7228
rect 14884 7216 14890 7268
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16209 7259 16267 7265
rect 16209 7256 16221 7259
rect 15988 7228 16221 7256
rect 15988 7216 15994 7228
rect 16209 7225 16221 7228
rect 16255 7256 16267 7259
rect 16666 7256 16672 7268
rect 16255 7228 16672 7256
rect 16255 7225 16267 7228
rect 16209 7219 16267 7225
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 16942 7256 16948 7268
rect 16903 7228 16948 7256
rect 16942 7216 16948 7228
rect 17000 7216 17006 7268
rect 19429 7259 19487 7265
rect 19429 7256 19441 7259
rect 18248 7228 19441 7256
rect 6604 7160 7052 7188
rect 6604 7148 6610 7160
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8260 7160 8401 7188
rect 8260 7148 8266 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8754 7188 8760 7200
rect 8715 7160 8760 7188
rect 8389 7151 8447 7157
rect 8754 7148 8760 7160
rect 8812 7148 8818 7200
rect 9122 7188 9128 7200
rect 9083 7160 9128 7188
rect 9122 7148 9128 7160
rect 9180 7148 9186 7200
rect 13541 7191 13599 7197
rect 13541 7157 13553 7191
rect 13587 7188 13599 7191
rect 13630 7188 13636 7200
rect 13587 7160 13636 7188
rect 13587 7157 13599 7160
rect 13541 7151 13599 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13814 7188 13820 7200
rect 13775 7160 13820 7188
rect 13814 7148 13820 7160
rect 13872 7148 13878 7200
rect 14918 7188 14924 7200
rect 14879 7160 14924 7188
rect 14918 7148 14924 7160
rect 14976 7148 14982 7200
rect 18248 7197 18276 7228
rect 19429 7225 19441 7228
rect 19475 7256 19487 7259
rect 19812 7256 19840 7287
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 20364 7333 20392 7364
rect 21634 7352 21640 7404
rect 21692 7392 21698 7404
rect 21913 7395 21971 7401
rect 21913 7392 21925 7395
rect 21692 7364 21925 7392
rect 21692 7352 21698 7364
rect 21913 7361 21925 7364
rect 21959 7361 21971 7395
rect 21913 7355 21971 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7392 28043 7395
rect 28460 7392 28488 7488
rect 28031 7364 28488 7392
rect 28031 7361 28043 7364
rect 27985 7355 28043 7361
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20714 7324 20720 7336
rect 20675 7296 20720 7324
rect 20349 7287 20407 7293
rect 20714 7284 20720 7296
rect 20772 7284 20778 7336
rect 25130 7324 25136 7336
rect 25043 7296 25136 7324
rect 25130 7284 25136 7296
rect 25188 7324 25194 7336
rect 25225 7327 25283 7333
rect 25225 7324 25237 7327
rect 25188 7296 25237 7324
rect 25188 7284 25194 7296
rect 25225 7293 25237 7296
rect 25271 7293 25283 7327
rect 25682 7324 25688 7336
rect 25643 7296 25688 7324
rect 25225 7287 25283 7293
rect 25682 7284 25688 7296
rect 25740 7284 25746 7336
rect 26050 7324 26056 7336
rect 26011 7296 26056 7324
rect 26050 7284 26056 7296
rect 26108 7284 26114 7336
rect 26418 7324 26424 7336
rect 26379 7296 26424 7324
rect 26418 7284 26424 7296
rect 26476 7284 26482 7336
rect 28902 7284 28908 7336
rect 28960 7324 28966 7336
rect 29308 7327 29366 7333
rect 29308 7324 29320 7327
rect 28960 7296 29320 7324
rect 28960 7284 28966 7296
rect 29308 7293 29320 7296
rect 29354 7324 29366 7327
rect 29733 7327 29791 7333
rect 29733 7324 29745 7327
rect 29354 7296 29745 7324
rect 29354 7293 29366 7296
rect 29308 7287 29366 7293
rect 29733 7293 29745 7296
rect 29779 7324 29791 7327
rect 29822 7324 29828 7336
rect 29779 7296 29828 7324
rect 29779 7293 29791 7296
rect 29733 7287 29791 7293
rect 29822 7284 29828 7296
rect 29880 7284 29886 7336
rect 35434 7324 35440 7336
rect 35395 7296 35440 7324
rect 35434 7284 35440 7296
rect 35492 7284 35498 7336
rect 20530 7256 20536 7268
rect 19475 7228 20536 7256
rect 19475 7225 19487 7228
rect 19429 7219 19487 7225
rect 20530 7216 20536 7228
rect 20588 7216 20594 7268
rect 22002 7256 22008 7268
rect 21963 7228 22008 7256
rect 22002 7216 22008 7228
rect 22060 7216 22066 7268
rect 22554 7256 22560 7268
rect 22515 7228 22560 7256
rect 22554 7216 22560 7228
rect 22612 7216 22618 7268
rect 26694 7256 26700 7268
rect 26655 7228 26700 7256
rect 26694 7216 26700 7228
rect 26752 7216 26758 7268
rect 18233 7191 18291 7197
rect 18233 7157 18245 7191
rect 18279 7157 18291 7191
rect 18966 7188 18972 7200
rect 18927 7160 18972 7188
rect 18233 7151 18291 7157
rect 18966 7148 18972 7160
rect 19024 7148 19030 7200
rect 20622 7148 20628 7200
rect 20680 7188 20686 7200
rect 20717 7191 20775 7197
rect 20717 7188 20729 7191
rect 20680 7160 20729 7188
rect 20680 7148 20686 7160
rect 20717 7157 20729 7160
rect 20763 7157 20775 7191
rect 21634 7188 21640 7200
rect 21595 7160 21640 7188
rect 20717 7151 20775 7157
rect 21634 7148 21640 7160
rect 21692 7148 21698 7200
rect 24670 7188 24676 7200
rect 24631 7160 24676 7188
rect 24670 7148 24676 7160
rect 24728 7148 24734 7200
rect 1104 7098 38824 7120
rect 1104 7046 14315 7098
rect 14367 7046 14379 7098
rect 14431 7046 14443 7098
rect 14495 7046 14507 7098
rect 14559 7046 27648 7098
rect 27700 7046 27712 7098
rect 27764 7046 27776 7098
rect 27828 7046 27840 7098
rect 27892 7046 38824 7098
rect 1104 7024 38824 7046
rect 5445 6987 5503 6993
rect 5445 6953 5457 6987
rect 5491 6984 5503 6987
rect 5534 6984 5540 6996
rect 5491 6956 5540 6984
rect 5491 6953 5503 6956
rect 5445 6947 5503 6953
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 13630 6984 13636 6996
rect 13591 6956 13636 6984
rect 13630 6944 13636 6956
rect 13688 6944 13694 6996
rect 14734 6984 14740 6996
rect 14695 6956 14740 6984
rect 14734 6944 14740 6956
rect 14792 6944 14798 6996
rect 15565 6987 15623 6993
rect 15565 6953 15577 6987
rect 15611 6984 15623 6987
rect 15654 6984 15660 6996
rect 15611 6956 15660 6984
rect 15611 6953 15623 6956
rect 15565 6947 15623 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 20806 6944 20812 6996
rect 20864 6984 20870 6996
rect 20993 6987 21051 6993
rect 20993 6984 21005 6987
rect 20864 6956 21005 6984
rect 20864 6944 20870 6956
rect 20993 6953 21005 6956
rect 21039 6953 21051 6987
rect 24670 6984 24676 6996
rect 24631 6956 24676 6984
rect 20993 6947 21051 6953
rect 24670 6944 24676 6956
rect 24728 6944 24734 6996
rect 25314 6984 25320 6996
rect 25227 6956 25320 6984
rect 25314 6944 25320 6956
rect 25372 6984 25378 6996
rect 25682 6984 25688 6996
rect 25372 6956 25688 6984
rect 25372 6944 25378 6956
rect 25682 6944 25688 6956
rect 25740 6944 25746 6996
rect 28169 6987 28227 6993
rect 28169 6953 28181 6987
rect 28215 6984 28227 6987
rect 28718 6984 28724 6996
rect 28215 6956 28724 6984
rect 28215 6953 28227 6956
rect 28169 6947 28227 6953
rect 28718 6944 28724 6956
rect 28776 6944 28782 6996
rect 7653 6919 7711 6925
rect 7653 6916 7665 6919
rect 7392 6888 7665 6916
rect 7392 6860 7420 6888
rect 7653 6885 7665 6888
rect 7699 6885 7711 6919
rect 11974 6916 11980 6928
rect 7653 6879 7711 6885
rect 11808 6888 11980 6916
rect 1464 6851 1522 6857
rect 1464 6817 1476 6851
rect 1510 6848 1522 6851
rect 2314 6848 2320 6860
rect 1510 6820 2320 6848
rect 1510 6817 1522 6820
rect 1464 6811 1522 6817
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 5169 6851 5227 6857
rect 5169 6817 5181 6851
rect 5215 6817 5227 6851
rect 5169 6811 5227 6817
rect 4154 6780 4160 6792
rect 4115 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4798 6672 4804 6724
rect 4856 6712 4862 6724
rect 5184 6712 5212 6811
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5629 6851 5687 6857
rect 5629 6848 5641 6851
rect 5316 6820 5641 6848
rect 5316 6808 5322 6820
rect 5629 6817 5641 6820
rect 5675 6817 5687 6851
rect 6178 6848 6184 6860
rect 6139 6820 6184 6848
rect 5629 6811 5687 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6365 6851 6423 6857
rect 6365 6848 6377 6851
rect 6328 6820 6377 6848
rect 6328 6808 6334 6820
rect 6365 6817 6377 6820
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7374 6848 7380 6860
rect 6972 6820 7380 6848
rect 6972 6808 6978 6820
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 11808 6857 11836 6888
rect 11974 6876 11980 6888
rect 12032 6916 12038 6928
rect 13170 6916 13176 6928
rect 12032 6888 13176 6916
rect 12032 6876 12038 6888
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 15746 6916 15752 6928
rect 15672 6888 15752 6916
rect 11609 6851 11667 6857
rect 11609 6817 11621 6851
rect 11655 6817 11667 6851
rect 11609 6811 11667 6817
rect 11793 6851 11851 6857
rect 11793 6817 11805 6851
rect 11839 6817 11851 6851
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 11793 6811 11851 6817
rect 11992 6820 12909 6848
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6749 7895 6783
rect 9674 6780 9680 6792
rect 9635 6752 9680 6780
rect 7837 6743 7895 6749
rect 6454 6712 6460 6724
rect 4856 6684 6460 6712
rect 4856 6672 4862 6684
rect 6454 6672 6460 6684
rect 6512 6712 6518 6724
rect 6512 6684 7052 6712
rect 6512 6672 6518 6684
rect 1394 6604 1400 6656
rect 1452 6644 1458 6656
rect 1535 6647 1593 6653
rect 1535 6644 1547 6647
rect 1452 6616 1547 6644
rect 1452 6604 1458 6616
rect 1535 6613 1547 6616
rect 1581 6613 1593 6647
rect 1535 6607 1593 6613
rect 4709 6647 4767 6653
rect 4709 6613 4721 6647
rect 4755 6644 4767 6647
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4755 6616 5089 6644
rect 4755 6613 4767 6616
rect 4709 6607 4767 6613
rect 5077 6613 5089 6616
rect 5123 6644 5135 6647
rect 5166 6644 5172 6656
rect 5123 6616 5172 6644
rect 5123 6613 5135 6616
rect 5077 6607 5135 6613
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7024 6644 7052 6684
rect 7098 6672 7104 6724
rect 7156 6712 7162 6724
rect 7852 6712 7880 6743
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 11624 6780 11652 6811
rect 11992 6780 12020 6820
rect 12897 6817 12909 6820
rect 12943 6848 12955 6851
rect 12986 6848 12992 6860
rect 12943 6820 12992 6848
rect 12943 6817 12955 6820
rect 12897 6811 12955 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 15672 6857 15700 6888
rect 15746 6876 15752 6888
rect 15804 6876 15810 6928
rect 21634 6916 21640 6928
rect 20640 6888 21640 6916
rect 15657 6851 15715 6857
rect 15657 6817 15669 6851
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17221 6851 17279 6857
rect 17221 6848 17233 6851
rect 17184 6820 17233 6848
rect 17184 6808 17190 6820
rect 17221 6817 17233 6820
rect 17267 6817 17279 6851
rect 17221 6811 17279 6817
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6817 18291 6851
rect 18233 6811 18291 6817
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20640 6848 20668 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 19843 6820 20668 6848
rect 21177 6851 21235 6857
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 21177 6817 21189 6851
rect 21223 6817 21235 6851
rect 21358 6848 21364 6860
rect 21319 6820 21364 6848
rect 21177 6811 21235 6817
rect 13170 6789 13176 6792
rect 11624 6752 12020 6780
rect 13136 6783 13176 6789
rect 13136 6749 13148 6783
rect 13136 6743 13176 6749
rect 13170 6740 13176 6743
rect 13228 6740 13234 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 14918 6780 14924 6792
rect 13403 6752 14924 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 7156 6684 7880 6712
rect 12529 6715 12587 6721
rect 7156 6672 7162 6684
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 13372 6712 13400 6743
rect 14918 6740 14924 6752
rect 14976 6780 14982 6792
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14976 6752 15025 6780
rect 14976 6740 14982 6752
rect 15013 6749 15025 6752
rect 15059 6780 15071 6783
rect 15804 6783 15862 6789
rect 15804 6780 15816 6783
rect 15059 6752 15816 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 15804 6749 15816 6752
rect 15850 6749 15862 6783
rect 16022 6780 16028 6792
rect 15983 6752 16028 6780
rect 15804 6743 15862 6749
rect 16022 6740 16028 6752
rect 16080 6740 16086 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6780 16451 6783
rect 18248 6780 18276 6811
rect 18874 6780 18880 6792
rect 16439 6752 18880 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 20257 6783 20315 6789
rect 20257 6780 20269 6783
rect 19024 6752 20269 6780
rect 19024 6740 19030 6752
rect 20257 6749 20269 6752
rect 20303 6780 20315 6783
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 20303 6752 20453 6780
rect 20303 6749 20315 6752
rect 20257 6743 20315 6749
rect 20441 6749 20453 6752
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20530 6740 20536 6792
rect 20588 6780 20594 6792
rect 21192 6780 21220 6811
rect 21358 6808 21364 6820
rect 21416 6808 21422 6860
rect 21910 6848 21916 6860
rect 21871 6820 21916 6848
rect 21910 6808 21916 6820
rect 21968 6808 21974 6860
rect 22097 6851 22155 6857
rect 22097 6817 22109 6851
rect 22143 6817 22155 6851
rect 24302 6848 24308 6860
rect 24263 6820 24308 6848
rect 22097 6811 22155 6817
rect 21818 6780 21824 6792
rect 20588 6752 21824 6780
rect 20588 6740 20594 6752
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 22112 6780 22140 6811
rect 24302 6808 24308 6820
rect 24360 6848 24366 6860
rect 24489 6851 24547 6857
rect 24489 6848 24501 6851
rect 24360 6820 24501 6848
rect 24360 6808 24366 6820
rect 24489 6817 24501 6820
rect 24535 6817 24547 6851
rect 24688 6848 24716 6944
rect 27570 6919 27628 6925
rect 27570 6885 27582 6919
rect 27616 6885 27628 6919
rect 27570 6879 27628 6885
rect 25593 6851 25651 6857
rect 25593 6848 25605 6851
rect 24688 6820 25605 6848
rect 24489 6811 24547 6817
rect 25593 6817 25605 6820
rect 25639 6848 25651 6851
rect 26418 6848 26424 6860
rect 25639 6820 26424 6848
rect 25639 6817 25651 6820
rect 25593 6811 25651 6817
rect 26418 6808 26424 6820
rect 26476 6808 26482 6860
rect 26694 6808 26700 6860
rect 26752 6848 26758 6860
rect 27249 6851 27307 6857
rect 27249 6848 27261 6851
rect 26752 6820 27261 6848
rect 26752 6808 26758 6820
rect 27249 6817 27261 6820
rect 27295 6817 27307 6851
rect 27249 6811 27307 6817
rect 21928 6752 22140 6780
rect 15930 6712 15936 6724
rect 12575 6684 13400 6712
rect 15891 6684 15936 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 21358 6712 21364 6724
rect 19996 6684 21364 6712
rect 19996 6656 20024 6684
rect 21358 6672 21364 6684
rect 21416 6672 21422 6724
rect 21726 6672 21732 6724
rect 21784 6712 21790 6724
rect 21928 6712 21956 6752
rect 27154 6740 27160 6792
rect 27212 6780 27218 6792
rect 27585 6780 27613 6879
rect 29178 6876 29184 6928
rect 29236 6916 29242 6928
rect 29273 6919 29331 6925
rect 29273 6916 29285 6919
rect 29236 6888 29285 6916
rect 29236 6876 29242 6888
rect 29273 6885 29285 6888
rect 29319 6885 29331 6919
rect 29273 6879 29331 6885
rect 27212 6752 27613 6780
rect 29181 6783 29239 6789
rect 27212 6740 27218 6752
rect 29181 6749 29193 6783
rect 29227 6749 29239 6783
rect 29822 6780 29828 6792
rect 29735 6752 29828 6780
rect 29181 6743 29239 6749
rect 21784 6684 21956 6712
rect 29196 6712 29224 6743
rect 29822 6740 29828 6752
rect 29880 6780 29886 6792
rect 30282 6780 30288 6792
rect 29880 6752 30288 6780
rect 29880 6740 29886 6752
rect 30282 6740 30288 6752
rect 30340 6740 30346 6792
rect 30006 6712 30012 6724
rect 29196 6684 30012 6712
rect 21784 6672 21790 6684
rect 30006 6672 30012 6684
rect 30064 6672 30070 6724
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 7024 6616 7297 6644
rect 7285 6613 7297 6616
rect 7331 6613 7343 6647
rect 11882 6644 11888 6656
rect 11843 6616 11888 6644
rect 7285 6607 7343 6613
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 13265 6647 13323 6653
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13630 6644 13636 6656
rect 13311 6616 13636 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13630 6604 13636 6616
rect 13688 6604 13694 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 17402 6644 17408 6656
rect 17363 6616 17408 6644
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 18046 6604 18052 6656
rect 18104 6644 18110 6656
rect 18417 6647 18475 6653
rect 18417 6644 18429 6647
rect 18104 6616 18429 6644
rect 18104 6604 18110 6616
rect 18417 6613 18429 6616
rect 18463 6644 18475 6647
rect 18966 6644 18972 6656
rect 18463 6616 18972 6644
rect 18463 6613 18475 6616
rect 18417 6607 18475 6613
rect 18966 6604 18972 6616
rect 19024 6604 19030 6656
rect 19426 6604 19432 6656
rect 19484 6644 19490 6656
rect 19521 6647 19579 6653
rect 19521 6644 19533 6647
rect 19484 6616 19533 6644
rect 19484 6604 19490 6616
rect 19521 6613 19533 6616
rect 19567 6644 19579 6647
rect 19978 6644 19984 6656
rect 19567 6616 19984 6644
rect 19567 6613 19579 6616
rect 19521 6607 19579 6613
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20441 6647 20499 6653
rect 20441 6613 20453 6647
rect 20487 6644 20499 6647
rect 20625 6647 20683 6653
rect 20625 6644 20637 6647
rect 20487 6616 20637 6644
rect 20487 6613 20499 6616
rect 20441 6607 20499 6613
rect 20625 6613 20637 6616
rect 20671 6644 20683 6647
rect 20714 6644 20720 6656
rect 20671 6616 20720 6644
rect 20671 6613 20683 6616
rect 20625 6607 20683 6613
rect 20714 6604 20720 6616
rect 20772 6604 20778 6656
rect 21376 6644 21404 6672
rect 22094 6644 22100 6656
rect 21376 6616 22100 6644
rect 22094 6604 22100 6616
rect 22152 6604 22158 6656
rect 25590 6604 25596 6656
rect 25648 6644 25654 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 25648 6616 25973 6644
rect 25648 6604 25654 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 1104 6554 38824 6576
rect 1104 6502 7648 6554
rect 7700 6502 7712 6554
rect 7764 6502 7776 6554
rect 7828 6502 7840 6554
rect 7892 6502 20982 6554
rect 21034 6502 21046 6554
rect 21098 6502 21110 6554
rect 21162 6502 21174 6554
rect 21226 6502 34315 6554
rect 34367 6502 34379 6554
rect 34431 6502 34443 6554
rect 34495 6502 34507 6554
rect 34559 6502 38824 6554
rect 1104 6480 38824 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2314 6440 2320 6452
rect 2275 6412 2320 6440
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 6273 6443 6331 6449
rect 6273 6409 6285 6443
rect 6319 6440 6331 6443
rect 6454 6440 6460 6452
rect 6319 6412 6460 6440
rect 6319 6409 6331 6412
rect 6273 6403 6331 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8665 6443 8723 6449
rect 8665 6440 8677 6443
rect 8076 6412 8677 6440
rect 8076 6400 8082 6412
rect 8665 6409 8677 6412
rect 8711 6440 8723 6443
rect 8754 6440 8760 6452
rect 8711 6412 8760 6440
rect 8711 6409 8723 6412
rect 8665 6403 8723 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13357 6443 13415 6449
rect 13357 6440 13369 6443
rect 13136 6412 13369 6440
rect 13136 6400 13142 6412
rect 13357 6409 13369 6412
rect 13403 6440 13415 6443
rect 15749 6443 15807 6449
rect 15749 6440 15761 6443
rect 13403 6412 15761 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 15749 6409 15761 6412
rect 15795 6440 15807 6443
rect 16022 6440 16028 6452
rect 15795 6412 16028 6440
rect 15795 6409 15807 6412
rect 15749 6403 15807 6409
rect 16022 6400 16028 6412
rect 16080 6400 16086 6452
rect 16117 6443 16175 6449
rect 16117 6409 16129 6443
rect 16163 6440 16175 6443
rect 17126 6440 17132 6452
rect 16163 6412 17132 6440
rect 16163 6409 16175 6412
rect 16117 6403 16175 6409
rect 8202 6372 8208 6384
rect 8163 6344 8208 6372
rect 8202 6332 8208 6344
rect 8260 6332 8266 6384
rect 13630 6372 13636 6384
rect 13591 6344 13636 6372
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 5074 6264 5080 6316
rect 5132 6304 5138 6316
rect 6178 6304 6184 6316
rect 5132 6276 6184 6304
rect 5132 6264 5138 6276
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 3973 6239 4031 6245
rect 1443 6208 2084 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2056 6112 2084 6208
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4709 6239 4767 6245
rect 4709 6236 4721 6239
rect 4019 6208 4721 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4709 6205 4721 6208
rect 4755 6236 4767 6239
rect 4798 6236 4804 6248
rect 4755 6208 4804 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5166 6236 5172 6248
rect 5127 6208 5172 6236
rect 5166 6196 5172 6208
rect 5224 6196 5230 6248
rect 5460 6245 5488 6276
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6914 6304 6920 6316
rect 6288 6276 6920 6304
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5810 6236 5816 6248
rect 5723 6208 5816 6236
rect 5445 6199 5503 6205
rect 5810 6196 5816 6208
rect 5868 6236 5874 6248
rect 6288 6236 6316 6276
rect 6914 6264 6920 6276
rect 6972 6304 6978 6316
rect 6972 6276 8248 6304
rect 6972 6264 6978 6276
rect 5868 6208 6316 6236
rect 5868 6196 5874 6208
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6825 6239 6883 6245
rect 6825 6236 6837 6239
rect 6512 6208 6837 6236
rect 6512 6196 6518 6208
rect 6825 6205 6837 6208
rect 6871 6205 6883 6239
rect 7558 6236 7564 6248
rect 7519 6208 7564 6236
rect 6825 6199 6883 6205
rect 7558 6196 7564 6208
rect 7616 6196 7622 6248
rect 7837 6239 7895 6245
rect 7837 6205 7849 6239
rect 7883 6236 7895 6239
rect 8018 6236 8024 6248
rect 7883 6208 8024 6236
rect 7883 6205 7895 6208
rect 7837 6199 7895 6205
rect 8018 6196 8024 6208
rect 8076 6196 8082 6248
rect 8220 6245 8248 6276
rect 8205 6239 8263 6245
rect 8205 6205 8217 6239
rect 8251 6205 8263 6239
rect 8205 6199 8263 6205
rect 3421 6171 3479 6177
rect 3421 6137 3433 6171
rect 3467 6168 3479 6171
rect 4062 6168 4068 6180
rect 3467 6140 4068 6168
rect 3467 6137 3479 6140
rect 3421 6131 3479 6137
rect 4062 6128 4068 6140
rect 4120 6128 4126 6180
rect 6641 6171 6699 6177
rect 6641 6137 6653 6171
rect 6687 6168 6699 6171
rect 6914 6168 6920 6180
rect 6687 6140 6920 6168
rect 6687 6137 6699 6140
rect 6641 6131 6699 6137
rect 6914 6128 6920 6140
rect 6972 6168 6978 6180
rect 7576 6168 7604 6196
rect 6972 6140 7604 6168
rect 8220 6168 8248 6199
rect 8294 6196 8300 6248
rect 8352 6236 8358 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8352 6208 9045 6236
rect 8352 6196 8358 6208
rect 9033 6205 9045 6208
rect 9079 6236 9091 6239
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 9079 6208 9229 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9217 6205 9229 6208
rect 9263 6205 9275 6239
rect 9217 6199 9275 6205
rect 11330 6196 11336 6248
rect 11388 6245 11394 6248
rect 11388 6239 11426 6245
rect 11414 6236 11426 6239
rect 11793 6239 11851 6245
rect 11793 6236 11805 6239
rect 11414 6208 11805 6236
rect 11414 6205 11426 6208
rect 11388 6199 11426 6205
rect 11793 6205 11805 6208
rect 11839 6236 11851 6239
rect 12066 6236 12072 6248
rect 11839 6208 12072 6236
rect 11839 6205 11851 6208
rect 11793 6199 11851 6205
rect 11388 6196 11394 6199
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 13078 6236 13084 6248
rect 12667 6208 13084 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 14090 6236 14096 6248
rect 14051 6208 14096 6236
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6205 14611 6239
rect 14734 6236 14740 6248
rect 14695 6208 14740 6236
rect 14553 6199 14611 6205
rect 9122 6168 9128 6180
rect 8220 6140 8708 6168
rect 9083 6140 9128 6168
rect 6972 6128 6978 6140
rect 2038 6100 2044 6112
rect 1999 6072 2044 6100
rect 2038 6060 2044 6072
rect 2096 6060 2102 6112
rect 4338 6100 4344 6112
rect 4299 6072 4344 6100
rect 4338 6060 4344 6072
rect 4396 6060 4402 6112
rect 4522 6100 4528 6112
rect 4483 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 8680 6100 8708 6140
rect 9122 6128 9128 6140
rect 9180 6128 9186 6180
rect 11241 6171 11299 6177
rect 11241 6137 11253 6171
rect 11287 6168 11299 6171
rect 12161 6171 12219 6177
rect 12161 6168 12173 6171
rect 11287 6140 12173 6168
rect 11287 6137 11299 6140
rect 11241 6131 11299 6137
rect 12161 6137 12173 6140
rect 12207 6168 12219 6171
rect 12437 6171 12495 6177
rect 12437 6168 12449 6171
rect 12207 6140 12449 6168
rect 12207 6137 12219 6140
rect 12161 6131 12219 6137
rect 12437 6137 12449 6140
rect 12483 6168 12495 6171
rect 12986 6168 12992 6180
rect 12483 6140 12992 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 12986 6128 12992 6140
rect 13044 6128 13050 6180
rect 14568 6168 14596 6199
rect 14734 6196 14740 6208
rect 14792 6196 14798 6248
rect 15102 6236 15108 6248
rect 15063 6208 15108 6236
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 16592 6245 16620 6412
rect 17126 6400 17132 6412
rect 17184 6440 17190 6452
rect 17221 6443 17279 6449
rect 17221 6440 17233 6443
rect 17184 6412 17233 6440
rect 17184 6400 17190 6412
rect 17221 6409 17233 6412
rect 17267 6409 17279 6443
rect 18506 6440 18512 6452
rect 18467 6412 18512 6440
rect 17221 6403 17279 6409
rect 18506 6400 18512 6412
rect 18564 6400 18570 6452
rect 18874 6440 18880 6452
rect 18835 6412 18880 6440
rect 18874 6400 18880 6412
rect 18932 6400 18938 6452
rect 22094 6440 22100 6452
rect 22055 6412 22100 6440
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 24210 6440 24216 6452
rect 24171 6412 24216 6440
rect 24210 6400 24216 6412
rect 24268 6400 24274 6452
rect 26694 6400 26700 6452
rect 26752 6440 26758 6452
rect 26881 6443 26939 6449
rect 26881 6440 26893 6443
rect 26752 6412 26893 6440
rect 26752 6400 26758 6412
rect 26881 6409 26893 6412
rect 26927 6409 26939 6443
rect 33410 6440 33416 6452
rect 33371 6412 33416 6440
rect 26881 6403 26939 6409
rect 33410 6400 33416 6412
rect 33468 6400 33474 6452
rect 28721 6375 28779 6381
rect 28721 6341 28733 6375
rect 28767 6372 28779 6375
rect 29178 6372 29184 6384
rect 28767 6344 29184 6372
rect 28767 6341 28779 6344
rect 28721 6335 28779 6341
rect 29178 6332 29184 6344
rect 29236 6372 29242 6384
rect 30193 6375 30251 6381
rect 30193 6372 30205 6375
rect 29236 6344 30205 6372
rect 29236 6332 29242 6344
rect 30193 6341 30205 6344
rect 30239 6341 30251 6375
rect 30193 6335 30251 6341
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 20772 6276 21220 6304
rect 20772 6264 20778 6276
rect 16577 6239 16635 6245
rect 16577 6205 16589 6239
rect 16623 6205 16635 6239
rect 16577 6199 16635 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6236 18107 6239
rect 18506 6236 18512 6248
rect 18095 6208 18512 6236
rect 18095 6205 18107 6208
rect 18049 6199 18107 6205
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 20257 6239 20315 6245
rect 20257 6205 20269 6239
rect 20303 6205 20315 6239
rect 20438 6236 20444 6248
rect 20399 6208 20444 6236
rect 20257 6199 20315 6205
rect 14642 6168 14648 6180
rect 14568 6140 14648 6168
rect 14642 6128 14648 6140
rect 14700 6128 14706 6180
rect 19521 6171 19579 6177
rect 19521 6137 19533 6171
rect 19567 6168 19579 6171
rect 20272 6168 20300 6199
rect 20438 6196 20444 6208
rect 20496 6196 20502 6248
rect 21192 6245 21220 6276
rect 20809 6239 20867 6245
rect 20809 6205 20821 6239
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 21177 6239 21235 6245
rect 21177 6205 21189 6239
rect 21223 6236 21235 6239
rect 21726 6236 21732 6248
rect 21223 6208 21732 6236
rect 21223 6205 21235 6208
rect 21177 6199 21235 6205
rect 20530 6168 20536 6180
rect 19567 6140 20536 6168
rect 19567 6137 19579 6140
rect 19521 6131 19579 6137
rect 20530 6128 20536 6140
rect 20588 6128 20594 6180
rect 20824 6168 20852 6199
rect 21726 6196 21732 6208
rect 21784 6196 21790 6248
rect 23661 6239 23719 6245
rect 23661 6205 23673 6239
rect 23707 6236 23719 6239
rect 24210 6236 24216 6248
rect 23707 6208 24216 6236
rect 23707 6205 23719 6208
rect 23661 6199 23719 6205
rect 24210 6196 24216 6208
rect 24268 6196 24274 6248
rect 25130 6236 25136 6248
rect 25043 6208 25136 6236
rect 25130 6196 25136 6208
rect 25188 6196 25194 6248
rect 25590 6236 25596 6248
rect 25551 6208 25596 6236
rect 25590 6196 25596 6208
rect 25648 6196 25654 6248
rect 26050 6196 26056 6248
rect 26108 6236 26114 6248
rect 26418 6236 26424 6248
rect 26108 6208 26201 6236
rect 26379 6208 26424 6236
rect 26108 6196 26114 6208
rect 26418 6196 26424 6208
rect 26476 6236 26482 6248
rect 27522 6236 27528 6248
rect 26476 6208 27528 6236
rect 26476 6196 26482 6208
rect 27522 6196 27528 6208
rect 27580 6196 27586 6248
rect 27706 6196 27712 6248
rect 27764 6245 27770 6248
rect 27764 6239 27802 6245
rect 27790 6236 27802 6239
rect 27982 6236 27988 6248
rect 27790 6208 27988 6236
rect 27790 6205 27802 6208
rect 27764 6199 27802 6205
rect 27764 6196 27770 6199
rect 27982 6196 27988 6208
rect 28040 6236 28046 6248
rect 28169 6239 28227 6245
rect 28169 6236 28181 6239
rect 28040 6208 28181 6236
rect 28040 6196 28046 6208
rect 28169 6205 28181 6208
rect 28215 6205 28227 6239
rect 29270 6236 29276 6248
rect 29231 6208 29276 6236
rect 28169 6199 28227 6205
rect 29270 6196 29276 6208
rect 29328 6236 29334 6248
rect 30469 6239 30527 6245
rect 30469 6236 30481 6239
rect 29328 6208 30481 6236
rect 29328 6196 29334 6208
rect 30469 6205 30481 6208
rect 30515 6205 30527 6239
rect 33226 6236 33232 6248
rect 33187 6208 33232 6236
rect 30469 6199 30527 6205
rect 33226 6196 33232 6208
rect 33284 6236 33290 6248
rect 33781 6239 33839 6245
rect 33781 6236 33793 6239
rect 33284 6208 33793 6236
rect 33284 6196 33290 6208
rect 33781 6205 33793 6208
rect 33827 6205 33839 6239
rect 33781 6199 33839 6205
rect 21910 6168 21916 6180
rect 20824 6140 21916 6168
rect 10134 6100 10140 6112
rect 8680 6072 10140 6100
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10873 6103 10931 6109
rect 10873 6069 10885 6103
rect 10919 6100 10931 6103
rect 10962 6100 10968 6112
rect 10919 6072 10968 6100
rect 10919 6069 10931 6072
rect 10873 6063 10931 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 11471 6103 11529 6109
rect 11471 6069 11483 6103
rect 11517 6100 11529 6103
rect 11698 6100 11704 6112
rect 11517 6072 11704 6100
rect 11517 6069 11529 6072
rect 11471 6063 11529 6069
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 12710 6100 12716 6112
rect 12671 6072 12716 6100
rect 12710 6060 12716 6072
rect 12768 6060 12774 6112
rect 14182 6100 14188 6112
rect 14143 6072 14188 6100
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 16666 6100 16672 6112
rect 16627 6072 16672 6100
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 17310 6060 17316 6112
rect 17368 6100 17374 6112
rect 18233 6103 18291 6109
rect 18233 6100 18245 6103
rect 17368 6072 18245 6100
rect 17368 6060 17374 6072
rect 18233 6069 18245 6072
rect 18279 6069 18291 6103
rect 19794 6100 19800 6112
rect 19755 6072 19800 6100
rect 18233 6063 18291 6069
rect 19794 6060 19800 6072
rect 19852 6100 19858 6112
rect 20824 6100 20852 6140
rect 21910 6128 21916 6140
rect 21968 6168 21974 6180
rect 22465 6171 22523 6177
rect 22465 6168 22477 6171
rect 21968 6140 22477 6168
rect 21968 6128 21974 6140
rect 22465 6137 22477 6140
rect 22511 6168 22523 6171
rect 22511 6140 23980 6168
rect 22511 6137 22523 6140
rect 22465 6131 22523 6137
rect 21358 6100 21364 6112
rect 19852 6072 20852 6100
rect 21319 6072 21364 6100
rect 19852 6060 19858 6072
rect 21358 6060 21364 6072
rect 21416 6060 21422 6112
rect 21818 6100 21824 6112
rect 21779 6072 21824 6100
rect 21818 6060 21824 6072
rect 21876 6060 21882 6112
rect 23842 6100 23848 6112
rect 23803 6072 23848 6100
rect 23842 6060 23848 6072
rect 23900 6060 23906 6112
rect 23952 6100 23980 6140
rect 24118 6128 24124 6180
rect 24176 6168 24182 6180
rect 24949 6171 25007 6177
rect 24949 6168 24961 6171
rect 24176 6140 24961 6168
rect 24176 6128 24182 6140
rect 24949 6137 24961 6140
rect 24995 6168 25007 6171
rect 25148 6168 25176 6196
rect 24995 6140 25176 6168
rect 26068 6168 26096 6196
rect 27338 6168 27344 6180
rect 26068 6140 27344 6168
rect 24995 6137 25007 6140
rect 24949 6131 25007 6137
rect 24581 6103 24639 6109
rect 24581 6100 24593 6103
rect 23952 6072 24593 6100
rect 24581 6069 24593 6072
rect 24627 6100 24639 6103
rect 26068 6100 26096 6140
rect 27338 6128 27344 6140
rect 27396 6128 27402 6180
rect 29594 6171 29652 6177
rect 29594 6168 29606 6171
rect 29012 6140 29606 6168
rect 24627 6072 26096 6100
rect 24627 6069 24639 6072
rect 24581 6063 24639 6069
rect 26142 6060 26148 6112
rect 26200 6100 26206 6112
rect 26329 6103 26387 6109
rect 26329 6100 26341 6103
rect 26200 6072 26341 6100
rect 26200 6060 26206 6072
rect 26329 6069 26341 6072
rect 26375 6069 26387 6103
rect 26329 6063 26387 6069
rect 27154 6060 27160 6112
rect 27212 6100 27218 6112
rect 27249 6103 27307 6109
rect 27249 6100 27261 6103
rect 27212 6072 27261 6100
rect 27212 6060 27218 6072
rect 27249 6069 27261 6072
rect 27295 6069 27307 6103
rect 27249 6063 27307 6069
rect 27847 6103 27905 6109
rect 27847 6069 27859 6103
rect 27893 6100 27905 6103
rect 28074 6100 28080 6112
rect 27893 6072 28080 6100
rect 27893 6069 27905 6072
rect 27847 6063 27905 6069
rect 28074 6060 28080 6072
rect 28132 6060 28138 6112
rect 28810 6060 28816 6112
rect 28868 6100 28874 6112
rect 29012 6109 29040 6140
rect 29594 6137 29606 6140
rect 29640 6137 29652 6171
rect 29594 6131 29652 6137
rect 28997 6103 29055 6109
rect 28997 6100 29009 6103
rect 28868 6072 29009 6100
rect 28868 6060 28874 6072
rect 28997 6069 29009 6072
rect 29043 6069 29055 6103
rect 28997 6063 29055 6069
rect 30006 6060 30012 6112
rect 30064 6100 30070 6112
rect 30837 6103 30895 6109
rect 30837 6100 30849 6103
rect 30064 6072 30849 6100
rect 30064 6060 30070 6072
rect 30837 6069 30849 6072
rect 30883 6069 30895 6103
rect 30837 6063 30895 6069
rect 1104 6010 38824 6032
rect 1104 5958 14315 6010
rect 14367 5958 14379 6010
rect 14431 5958 14443 6010
rect 14495 5958 14507 6010
rect 14559 5958 27648 6010
rect 27700 5958 27712 6010
rect 27764 5958 27776 6010
rect 27828 5958 27840 6010
rect 27892 5958 38824 6010
rect 1104 5936 38824 5958
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7432 5868 7941 5896
rect 7432 5856 7438 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 9582 5856 9588 5908
rect 9640 5896 9646 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 9640 5868 10241 5896
rect 9640 5856 9646 5868
rect 10229 5865 10241 5868
rect 10275 5865 10287 5899
rect 11974 5896 11980 5908
rect 11935 5868 11980 5896
rect 10229 5859 10287 5865
rect 11974 5856 11980 5868
rect 12032 5896 12038 5908
rect 12345 5899 12403 5905
rect 12345 5896 12357 5899
rect 12032 5868 12357 5896
rect 12032 5856 12038 5868
rect 12345 5865 12357 5868
rect 12391 5865 12403 5899
rect 12345 5859 12403 5865
rect 12986 5856 12992 5908
rect 13044 5896 13050 5908
rect 13044 5868 13124 5896
rect 13044 5856 13050 5868
rect 2130 5828 2136 5840
rect 2091 5800 2136 5828
rect 2130 5788 2136 5800
rect 2188 5788 2194 5840
rect 5276 5800 6960 5828
rect 5276 5769 5304 5800
rect 6932 5772 6960 5800
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 7524 5800 8309 5828
rect 7524 5788 7530 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 8297 5791 8355 5797
rect 10045 5831 10103 5837
rect 10045 5797 10057 5831
rect 10091 5828 10103 5831
rect 10134 5828 10140 5840
rect 10091 5800 10140 5828
rect 10091 5797 10103 5800
rect 10045 5791 10103 5797
rect 10134 5788 10140 5800
rect 10192 5828 10198 5840
rect 13096 5828 13124 5868
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 13725 5899 13783 5905
rect 13725 5896 13737 5899
rect 13504 5868 13737 5896
rect 13504 5856 13510 5868
rect 13725 5865 13737 5868
rect 13771 5865 13783 5899
rect 13725 5859 13783 5865
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15654 5896 15660 5908
rect 15611 5868 15660 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 16301 5899 16359 5905
rect 16301 5896 16313 5899
rect 15804 5868 16313 5896
rect 15804 5856 15810 5868
rect 16301 5865 16313 5868
rect 16347 5865 16359 5899
rect 16301 5859 16359 5865
rect 20257 5899 20315 5905
rect 20257 5865 20269 5899
rect 20303 5896 20315 5899
rect 20438 5896 20444 5908
rect 20303 5868 20444 5896
rect 20303 5865 20315 5868
rect 20257 5859 20315 5865
rect 20438 5856 20444 5868
rect 20496 5896 20502 5908
rect 20806 5896 20812 5908
rect 20496 5868 20812 5896
rect 20496 5856 20502 5868
rect 20806 5856 20812 5868
rect 20864 5856 20870 5908
rect 28074 5856 28080 5908
rect 28132 5896 28138 5908
rect 28261 5899 28319 5905
rect 28261 5896 28273 5899
rect 28132 5868 28273 5896
rect 28132 5856 28138 5868
rect 28261 5865 28273 5868
rect 28307 5865 28319 5899
rect 28261 5859 28319 5865
rect 28810 5856 28816 5908
rect 28868 5856 28874 5908
rect 15013 5831 15071 5837
rect 15013 5828 15025 5831
rect 10192 5800 10916 5828
rect 13096 5800 15025 5828
rect 10192 5788 10198 5800
rect 10888 5772 10916 5800
rect 15013 5797 15025 5800
rect 15059 5828 15071 5831
rect 15930 5828 15936 5840
rect 15059 5800 15936 5828
rect 15059 5797 15071 5800
rect 15013 5791 15071 5797
rect 15930 5788 15936 5800
rect 15988 5788 15994 5840
rect 21266 5837 21272 5840
rect 21263 5828 21272 5837
rect 21227 5800 21272 5828
rect 21263 5791 21272 5800
rect 21266 5788 21272 5791
rect 21324 5788 21330 5840
rect 23842 5788 23848 5840
rect 23900 5828 23906 5840
rect 24854 5828 24860 5840
rect 23900 5800 24860 5828
rect 23900 5788 23906 5800
rect 24854 5788 24860 5800
rect 24912 5828 24918 5840
rect 28629 5831 28687 5837
rect 28629 5828 28641 5831
rect 24912 5800 24992 5828
rect 24912 5788 24918 5800
rect 5261 5763 5319 5769
rect 5261 5729 5273 5763
rect 5307 5729 5319 5763
rect 6454 5760 6460 5772
rect 6415 5732 6460 5760
rect 5261 5723 5319 5729
rect 6454 5720 6460 5732
rect 6512 5720 6518 5772
rect 6914 5760 6920 5772
rect 6875 5732 6920 5760
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5729 7251 5763
rect 7374 5760 7380 5772
rect 7335 5732 7380 5760
rect 7193 5723 7251 5729
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 2774 5692 2780 5704
rect 2087 5664 2780 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4396 5664 4537 5692
rect 4396 5652 4402 5664
rect 4525 5661 4537 5664
rect 4571 5692 4583 5695
rect 5810 5692 5816 5704
rect 4571 5664 5816 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 5810 5652 5816 5664
rect 5868 5652 5874 5704
rect 7208 5692 7236 5723
rect 7374 5720 7380 5732
rect 7432 5720 7438 5772
rect 8570 5769 8576 5772
rect 8548 5763 8576 5769
rect 8548 5729 8560 5763
rect 8548 5723 8576 5729
rect 8570 5720 8576 5723
rect 8628 5720 8634 5772
rect 10318 5760 10324 5772
rect 10279 5732 10324 5760
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 10594 5760 10600 5772
rect 10555 5732 10600 5760
rect 10594 5720 10600 5732
rect 10652 5720 10658 5772
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10928 5732 10977 5760
rect 10928 5720 10934 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 11238 5720 11244 5772
rect 11296 5760 11302 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11296 5732 11345 5760
rect 11296 5720 11302 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 11333 5723 11391 5729
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 12986 5760 12992 5772
rect 12899 5732 12992 5760
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5729 13415 5763
rect 13357 5723 13415 5729
rect 8018 5692 8024 5704
rect 7208 5664 8024 5692
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 12342 5652 12348 5704
rect 12400 5692 12406 5704
rect 13004 5692 13032 5720
rect 12400 5664 13032 5692
rect 13372 5692 13400 5723
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 13909 5763 13967 5769
rect 13909 5760 13921 5763
rect 13780 5732 13921 5760
rect 13780 5720 13786 5732
rect 13909 5729 13921 5732
rect 13955 5760 13967 5763
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 13955 5732 14657 5760
rect 13955 5729 13967 5732
rect 13909 5723 13967 5729
rect 14645 5729 14657 5732
rect 14691 5760 14703 5763
rect 15102 5760 15108 5772
rect 14691 5732 15108 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 15838 5760 15844 5772
rect 15799 5732 15844 5760
rect 15838 5720 15844 5732
rect 15896 5720 15902 5772
rect 17310 5760 17316 5772
rect 17271 5732 17316 5760
rect 17310 5720 17316 5732
rect 17368 5720 17374 5772
rect 17402 5720 17408 5772
rect 17460 5760 17466 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17460 5732 17601 5760
rect 17460 5720 17466 5732
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 17954 5760 17960 5772
rect 17915 5732 17960 5760
rect 17589 5723 17647 5729
rect 17954 5720 17960 5732
rect 18012 5720 18018 5772
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18325 5763 18383 5769
rect 18325 5760 18337 5763
rect 18104 5732 18337 5760
rect 18104 5720 18110 5732
rect 18325 5729 18337 5732
rect 18371 5729 18383 5763
rect 18325 5723 18383 5729
rect 19702 5720 19708 5772
rect 19760 5769 19766 5772
rect 19760 5763 19798 5769
rect 19786 5729 19798 5763
rect 19760 5723 19798 5729
rect 19760 5720 19766 5723
rect 20714 5720 20720 5772
rect 20772 5760 20778 5772
rect 20901 5763 20959 5769
rect 20901 5760 20913 5763
rect 20772 5732 20913 5760
rect 20772 5720 20778 5732
rect 20901 5729 20913 5732
rect 20947 5760 20959 5763
rect 22002 5760 22008 5772
rect 20947 5732 22008 5760
rect 20947 5729 20959 5732
rect 20901 5723 20959 5729
rect 22002 5720 22008 5732
rect 22060 5720 22066 5772
rect 22094 5720 22100 5772
rect 22152 5720 22158 5772
rect 24118 5760 24124 5772
rect 24079 5732 24124 5760
rect 24118 5720 24124 5732
rect 24176 5720 24182 5772
rect 24964 5769 24992 5800
rect 26436 5800 28641 5828
rect 24581 5763 24639 5769
rect 24581 5729 24593 5763
rect 24627 5729 24639 5763
rect 24581 5723 24639 5729
rect 24949 5763 25007 5769
rect 24949 5729 24961 5763
rect 24995 5729 25007 5763
rect 24949 5723 25007 5729
rect 25501 5763 25559 5769
rect 25501 5729 25513 5763
rect 25547 5760 25559 5763
rect 26326 5760 26332 5772
rect 25547 5732 26332 5760
rect 25547 5729 25559 5732
rect 25501 5723 25559 5729
rect 13814 5692 13820 5704
rect 13372 5664 13820 5692
rect 12400 5652 12406 5664
rect 2590 5624 2596 5636
rect 2551 5596 2596 5624
rect 2590 5584 2596 5596
rect 2648 5584 2654 5636
rect 6914 5584 6920 5636
rect 6972 5624 6978 5636
rect 7561 5627 7619 5633
rect 7561 5624 7573 5627
rect 6972 5596 7573 5624
rect 6972 5584 6978 5596
rect 7561 5593 7573 5596
rect 7607 5593 7619 5627
rect 7561 5587 7619 5593
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 13372 5624 13400 5664
rect 13814 5652 13820 5664
rect 13872 5692 13878 5704
rect 14734 5692 14740 5704
rect 13872 5664 14740 5692
rect 13872 5652 13878 5664
rect 14734 5652 14740 5664
rect 14792 5652 14798 5704
rect 17972 5692 18000 5720
rect 19518 5692 19524 5704
rect 17972 5664 19524 5692
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 22112 5692 22140 5720
rect 24486 5692 24492 5704
rect 22112 5664 24492 5692
rect 24486 5652 24492 5664
rect 24544 5692 24550 5704
rect 24596 5692 24624 5723
rect 26326 5720 26332 5732
rect 26384 5720 26390 5772
rect 25314 5692 25320 5704
rect 24544 5664 25320 5692
rect 24544 5652 24550 5664
rect 25314 5652 25320 5664
rect 25372 5652 25378 5704
rect 25593 5695 25651 5701
rect 25593 5661 25605 5695
rect 25639 5692 25651 5695
rect 26436 5692 26464 5800
rect 28629 5797 28641 5800
rect 28675 5797 28687 5831
rect 28828 5828 28856 5856
rect 29134 5831 29192 5837
rect 29134 5828 29146 5831
rect 28828 5800 29146 5828
rect 28629 5791 28687 5797
rect 29134 5797 29146 5800
rect 29180 5797 29192 5831
rect 29134 5791 29192 5797
rect 26786 5760 26792 5772
rect 26747 5732 26792 5760
rect 26786 5720 26792 5732
rect 26844 5720 26850 5772
rect 26973 5763 27031 5769
rect 26973 5729 26985 5763
rect 27019 5729 27031 5763
rect 27338 5760 27344 5772
rect 27299 5732 27344 5760
rect 26973 5723 27031 5729
rect 25639 5664 26464 5692
rect 25639 5661 25651 5664
rect 25593 5655 25651 5661
rect 18506 5624 18512 5636
rect 12492 5596 13400 5624
rect 18467 5596 18512 5624
rect 12492 5584 12498 5596
rect 18506 5584 18512 5596
rect 18564 5584 18570 5636
rect 1670 5556 1676 5568
rect 1631 5528 1676 5556
rect 1670 5516 1676 5528
rect 1728 5516 1734 5568
rect 5077 5559 5135 5565
rect 5077 5525 5089 5559
rect 5123 5556 5135 5559
rect 5166 5556 5172 5568
rect 5123 5528 5172 5556
rect 5123 5525 5135 5528
rect 5077 5519 5135 5525
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6089 5559 6147 5565
rect 6089 5556 6101 5559
rect 5767 5528 6101 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6089 5525 6101 5528
rect 6135 5556 6147 5559
rect 6270 5556 6276 5568
rect 6135 5528 6276 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 8386 5516 8392 5568
rect 8444 5556 8450 5568
rect 8619 5559 8677 5565
rect 8619 5556 8631 5559
rect 8444 5528 8631 5556
rect 8444 5516 8450 5528
rect 8619 5525 8631 5528
rect 8665 5525 8677 5559
rect 9490 5556 9496 5568
rect 9451 5528 9496 5556
rect 8619 5519 8677 5525
rect 9490 5516 9496 5528
rect 9548 5516 9554 5568
rect 14369 5559 14427 5565
rect 14369 5525 14381 5559
rect 14415 5556 14427 5559
rect 14642 5556 14648 5568
rect 14415 5528 14648 5556
rect 14415 5525 14427 5528
rect 14369 5519 14427 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 17037 5559 17095 5565
rect 17037 5525 17049 5559
rect 17083 5556 17095 5559
rect 17954 5556 17960 5568
rect 17083 5528 17960 5556
rect 17083 5525 17095 5528
rect 17037 5519 17095 5525
rect 17954 5516 17960 5528
rect 18012 5516 18018 5568
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19843 5559 19901 5565
rect 19843 5556 19855 5559
rect 19392 5528 19855 5556
rect 19392 5516 19398 5528
rect 19843 5525 19855 5528
rect 19889 5525 19901 5559
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 19843 5519 19901 5525
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 21821 5559 21879 5565
rect 21821 5525 21833 5559
rect 21867 5556 21879 5559
rect 22094 5556 22100 5568
rect 21867 5528 22100 5556
rect 21867 5525 21879 5528
rect 21821 5519 21879 5525
rect 22094 5516 22100 5528
rect 22152 5516 22158 5568
rect 25590 5516 25596 5568
rect 25648 5556 25654 5568
rect 25869 5559 25927 5565
rect 25869 5556 25881 5559
rect 25648 5528 25881 5556
rect 25648 5516 25654 5528
rect 25869 5525 25881 5528
rect 25915 5556 25927 5559
rect 26988 5556 27016 5723
rect 27338 5720 27344 5732
rect 27396 5720 27402 5772
rect 27522 5720 27528 5772
rect 27580 5760 27586 5772
rect 27709 5763 27767 5769
rect 27709 5760 27721 5763
rect 27580 5732 27721 5760
rect 27580 5720 27586 5732
rect 27709 5729 27721 5732
rect 27755 5729 27767 5763
rect 28644 5760 28672 5791
rect 28813 5763 28871 5769
rect 28813 5760 28825 5763
rect 28644 5732 28825 5760
rect 27709 5723 27767 5729
rect 28813 5729 28825 5732
rect 28859 5729 28871 5763
rect 28813 5723 28871 5729
rect 27985 5695 28043 5701
rect 27985 5661 27997 5695
rect 28031 5692 28043 5695
rect 29270 5692 29276 5704
rect 28031 5664 29276 5692
rect 28031 5661 28043 5664
rect 27985 5655 28043 5661
rect 29270 5652 29276 5664
rect 29328 5652 29334 5704
rect 25915 5528 27016 5556
rect 29733 5559 29791 5565
rect 25915 5525 25927 5528
rect 25869 5519 25927 5525
rect 29733 5525 29745 5559
rect 29779 5556 29791 5559
rect 30374 5556 30380 5568
rect 29779 5528 30380 5556
rect 29779 5525 29791 5528
rect 29733 5519 29791 5525
rect 30374 5516 30380 5528
rect 30432 5516 30438 5568
rect 30926 5556 30932 5568
rect 30887 5528 30932 5556
rect 30926 5516 30932 5528
rect 30984 5516 30990 5568
rect 1104 5466 38824 5488
rect 1104 5414 7648 5466
rect 7700 5414 7712 5466
rect 7764 5414 7776 5466
rect 7828 5414 7840 5466
rect 7892 5414 20982 5466
rect 21034 5414 21046 5466
rect 21098 5414 21110 5466
rect 21162 5414 21174 5466
rect 21226 5414 34315 5466
rect 34367 5414 34379 5466
rect 34431 5414 34443 5466
rect 34495 5414 34507 5466
rect 34559 5414 38824 5466
rect 1104 5392 38824 5414
rect 2130 5312 2136 5364
rect 2188 5352 2194 5364
rect 2501 5355 2559 5361
rect 2501 5352 2513 5355
rect 2188 5324 2513 5352
rect 2188 5312 2194 5324
rect 2501 5321 2513 5324
rect 2547 5352 2559 5355
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2547 5324 2605 5352
rect 2547 5321 2559 5324
rect 2501 5315 2559 5321
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 3326 5352 3332 5364
rect 3283 5324 3332 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 3252 5284 3280 5315
rect 3326 5312 3332 5324
rect 3384 5312 3390 5364
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 6273 5355 6331 5361
rect 6273 5352 6285 5355
rect 4387 5324 6285 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 6273 5321 6285 5324
rect 6319 5352 6331 5355
rect 6822 5352 6828 5364
rect 6319 5324 6828 5352
rect 6319 5321 6331 5324
rect 6273 5315 6331 5321
rect 6822 5312 6828 5324
rect 6880 5312 6886 5364
rect 7745 5355 7803 5361
rect 7745 5321 7757 5355
rect 7791 5352 7803 5355
rect 8202 5352 8208 5364
rect 7791 5324 8208 5352
rect 7791 5321 7803 5324
rect 7745 5315 7803 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9953 5355 10011 5361
rect 9953 5321 9965 5355
rect 9999 5352 10011 5355
rect 10594 5352 10600 5364
rect 9999 5324 10600 5352
rect 9999 5321 10011 5324
rect 9953 5315 10011 5321
rect 10594 5312 10600 5324
rect 10652 5352 10658 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 10652 5324 12173 5352
rect 10652 5312 10658 5324
rect 12161 5321 12173 5324
rect 12207 5352 12219 5355
rect 12342 5352 12348 5364
rect 12207 5324 12348 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 15838 5352 15844 5364
rect 15799 5324 15844 5352
rect 15838 5312 15844 5324
rect 15896 5312 15902 5364
rect 16206 5352 16212 5364
rect 16167 5324 16212 5352
rect 16206 5312 16212 5324
rect 16264 5312 16270 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17862 5352 17868 5364
rect 17543 5324 17868 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 17954 5312 17960 5364
rect 18012 5352 18018 5364
rect 19337 5355 19395 5361
rect 19337 5352 19349 5355
rect 18012 5324 19349 5352
rect 18012 5312 18018 5324
rect 19337 5321 19349 5324
rect 19383 5321 19395 5355
rect 19702 5352 19708 5364
rect 19663 5324 19708 5352
rect 19337 5315 19395 5321
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5352 20499 5355
rect 21266 5352 21272 5364
rect 20487 5324 21272 5352
rect 20487 5321 20499 5324
rect 20441 5315 20499 5321
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22649 5355 22707 5361
rect 22649 5352 22661 5355
rect 22244 5324 22661 5352
rect 22244 5312 22250 5324
rect 22649 5321 22661 5324
rect 22695 5321 22707 5355
rect 24118 5352 24124 5364
rect 24079 5324 24124 5352
rect 22649 5315 22707 5321
rect 24118 5312 24124 5324
rect 24176 5352 24182 5364
rect 25133 5355 25191 5361
rect 25133 5352 25145 5355
rect 24176 5324 25145 5352
rect 24176 5312 24182 5324
rect 25133 5321 25145 5324
rect 25179 5321 25191 5355
rect 25133 5315 25191 5321
rect 1596 5256 3280 5284
rect 1596 5225 1624 5256
rect 6546 5244 6552 5296
rect 6604 5284 6610 5296
rect 8018 5284 8024 5296
rect 6604 5256 8024 5284
rect 6604 5244 6610 5256
rect 8018 5244 8024 5256
rect 8076 5244 8082 5296
rect 24486 5284 24492 5296
rect 24447 5256 24492 5284
rect 24486 5244 24492 5256
rect 24544 5244 24550 5296
rect 1581 5219 1639 5225
rect 1581 5185 1593 5219
rect 1627 5185 1639 5219
rect 1581 5179 1639 5185
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3467 5219 3525 5225
rect 3467 5216 3479 5219
rect 2832 5188 3479 5216
rect 2832 5176 2838 5188
rect 3467 5185 3479 5188
rect 3513 5185 3525 5219
rect 3878 5216 3884 5228
rect 3839 5188 3884 5216
rect 3467 5179 3525 5185
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 6564 5216 6592 5244
rect 5460 5188 6592 5216
rect 6825 5219 6883 5225
rect 3380 5151 3438 5157
rect 3380 5117 3392 5151
rect 3426 5148 3438 5151
rect 3694 5148 3700 5160
rect 3426 5120 3700 5148
rect 3426 5117 3438 5120
rect 3380 5111 3438 5117
rect 3694 5108 3700 5120
rect 3752 5148 3758 5160
rect 3896 5148 3924 5176
rect 5460 5160 5488 5188
rect 6825 5185 6837 5219
rect 6871 5216 6883 5219
rect 6914 5216 6920 5228
rect 6871 5188 6920 5216
rect 6871 5185 6883 5188
rect 6825 5179 6883 5185
rect 6914 5176 6920 5188
rect 6972 5176 6978 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14642 5216 14648 5228
rect 13679 5188 14648 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 3752 5120 3924 5148
rect 4709 5151 4767 5157
rect 3752 5108 3758 5120
rect 4709 5117 4721 5151
rect 4755 5148 4767 5151
rect 4798 5148 4804 5160
rect 4755 5120 4804 5148
rect 4755 5117 4767 5120
rect 4709 5111 4767 5117
rect 4798 5108 4804 5120
rect 4856 5108 4862 5160
rect 5166 5148 5172 5160
rect 5127 5120 5172 5148
rect 5166 5108 5172 5120
rect 5224 5108 5230 5160
rect 5442 5148 5448 5160
rect 5355 5120 5448 5148
rect 5442 5108 5448 5120
rect 5500 5108 5506 5160
rect 5810 5148 5816 5160
rect 5771 5120 5816 5148
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9068 5151 9126 5157
rect 9068 5148 9080 5151
rect 8987 5120 9080 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9068 5117 9080 5120
rect 9114 5117 9126 5151
rect 9068 5111 9126 5117
rect 9585 5151 9643 5157
rect 9585 5117 9597 5151
rect 9631 5148 9643 5151
rect 10318 5148 10324 5160
rect 9631 5120 10324 5148
rect 9631 5117 9643 5120
rect 9585 5111 9643 5117
rect 1670 5040 1676 5092
rect 1728 5080 1734 5092
rect 1902 5083 1960 5089
rect 1902 5080 1914 5083
rect 1728 5052 1914 5080
rect 1728 5040 1734 5052
rect 1902 5049 1914 5052
rect 1948 5049 1960 5083
rect 1902 5043 1960 5049
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 2869 5083 2927 5089
rect 2869 5080 2881 5083
rect 2639 5052 2881 5080
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 2869 5049 2881 5052
rect 2915 5080 2927 5083
rect 4154 5080 4160 5092
rect 2915 5052 4160 5080
rect 2915 5049 2927 5052
rect 2869 5043 2927 5049
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 7146 5083 7204 5089
rect 7146 5080 7158 5083
rect 6564 5052 7158 5080
rect 5626 5012 5632 5024
rect 5587 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 6454 4972 6460 5024
rect 6512 5012 6518 5024
rect 6564 5021 6592 5052
rect 7146 5049 7158 5052
rect 7192 5049 7204 5083
rect 8956 5080 8984 5111
rect 10318 5108 10324 5120
rect 10376 5108 10382 5160
rect 10689 5151 10747 5157
rect 10689 5117 10701 5151
rect 10735 5117 10747 5151
rect 10870 5148 10876 5160
rect 10831 5120 10876 5148
rect 10689 5111 10747 5117
rect 9858 5080 9864 5092
rect 8956 5052 9864 5080
rect 7146 5043 7204 5049
rect 9858 5040 9864 5052
rect 9916 5040 9922 5092
rect 6549 5015 6607 5021
rect 6549 5012 6561 5015
rect 6512 4984 6561 5012
rect 6512 4972 6518 4984
rect 6549 4981 6561 4984
rect 6595 4981 6607 5015
rect 8570 5012 8576 5024
rect 8531 4984 8576 5012
rect 6549 4975 6607 4981
rect 8570 4972 8576 4984
rect 8628 4972 8634 5024
rect 8938 4972 8944 5024
rect 8996 5012 9002 5024
rect 9171 5015 9229 5021
rect 9171 5012 9183 5015
rect 8996 4984 9183 5012
rect 8996 4972 9002 4984
rect 9171 4981 9183 4984
rect 9217 4981 9229 5015
rect 10704 5012 10732 5111
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 11238 5148 11244 5160
rect 11199 5120 11244 5148
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 11517 5083 11575 5089
rect 11517 5049 11529 5083
rect 11563 5080 11575 5083
rect 12434 5080 12440 5092
rect 11563 5052 12440 5080
rect 11563 5049 11575 5052
rect 11517 5043 11575 5049
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 12618 5080 12624 5092
rect 12579 5052 12624 5080
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 13265 5083 13323 5089
rect 12768 5052 12813 5080
rect 12768 5040 12774 5052
rect 13265 5049 13277 5083
rect 13311 5080 13323 5083
rect 13630 5080 13636 5092
rect 13311 5052 13636 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 13630 5040 13636 5052
rect 13688 5040 13694 5092
rect 10962 5012 10968 5024
rect 10704 4984 10968 5012
rect 9171 4975 9229 4981
rect 10962 4972 10968 4984
rect 11020 5012 11026 5024
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11020 4984 11897 5012
rect 11020 4972 11026 4984
rect 11885 4981 11897 4984
rect 11931 5012 11943 5015
rect 13740 5012 13768 5188
rect 14642 5176 14648 5188
rect 14700 5216 14706 5228
rect 15838 5216 15844 5228
rect 14700 5188 15844 5216
rect 14700 5176 14706 5188
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14090 5148 14096 5160
rect 14047 5120 14096 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 14090 5108 14096 5120
rect 14148 5148 14154 5160
rect 14366 5148 14372 5160
rect 14148 5120 14372 5148
rect 14148 5108 14154 5120
rect 14366 5108 14372 5120
rect 14424 5108 14430 5160
rect 14752 5157 14780 5188
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 17126 5216 17132 5228
rect 17087 5188 17132 5216
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 22278 5216 22284 5228
rect 21008 5188 22284 5216
rect 14737 5151 14795 5157
rect 14737 5117 14749 5151
rect 14783 5117 14795 5151
rect 14918 5148 14924 5160
rect 14879 5120 14924 5148
rect 14737 5111 14795 5117
rect 14918 5108 14924 5120
rect 14976 5108 14982 5160
rect 15194 5108 15200 5160
rect 15252 5148 15258 5160
rect 15289 5151 15347 5157
rect 15289 5148 15301 5151
rect 15252 5120 15301 5148
rect 15252 5108 15258 5120
rect 15289 5117 15301 5120
rect 15335 5117 15347 5151
rect 15289 5111 15347 5117
rect 16206 5108 16212 5160
rect 16264 5148 16270 5160
rect 16485 5151 16543 5157
rect 16485 5148 16497 5151
rect 16264 5120 16497 5148
rect 16264 5108 16270 5120
rect 16485 5117 16497 5120
rect 16531 5117 16543 5151
rect 18046 5148 18052 5160
rect 18007 5120 18052 5148
rect 16485 5111 16543 5117
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 20714 5148 20720 5160
rect 20675 5120 20720 5148
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 20806 5108 20812 5160
rect 20864 5148 20870 5160
rect 21008 5157 21036 5188
rect 22278 5176 22284 5188
rect 22336 5176 22342 5228
rect 20993 5151 21051 5157
rect 20993 5148 21005 5151
rect 20864 5120 21005 5148
rect 20864 5108 20870 5120
rect 20993 5117 21005 5120
rect 21039 5117 21051 5151
rect 20993 5111 21051 5117
rect 21082 5108 21088 5160
rect 21140 5148 21146 5160
rect 21361 5151 21419 5157
rect 21361 5148 21373 5151
rect 21140 5120 21373 5148
rect 21140 5108 21146 5120
rect 21361 5117 21373 5120
rect 21407 5148 21419 5151
rect 21450 5148 21456 5160
rect 21407 5120 21456 5148
rect 21407 5117 21419 5120
rect 21361 5111 21419 5117
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 21726 5148 21732 5160
rect 21687 5120 21732 5148
rect 21726 5108 21732 5120
rect 21784 5108 21790 5160
rect 25148 5148 25176 5315
rect 30374 5312 30380 5364
rect 30432 5352 30438 5364
rect 30653 5355 30711 5361
rect 30653 5352 30665 5355
rect 30432 5324 30665 5352
rect 30432 5312 30438 5324
rect 30653 5321 30665 5324
rect 30699 5352 30711 5355
rect 31018 5352 31024 5364
rect 30699 5324 31024 5352
rect 30699 5321 30711 5324
rect 30653 5315 30711 5321
rect 31018 5312 31024 5324
rect 31076 5312 31082 5364
rect 25682 5244 25688 5296
rect 25740 5284 25746 5296
rect 27157 5287 27215 5293
rect 25740 5256 26832 5284
rect 25740 5244 25746 5256
rect 26804 5228 26832 5256
rect 27157 5253 27169 5287
rect 27203 5284 27215 5287
rect 27338 5284 27344 5296
rect 27203 5256 27344 5284
rect 27203 5253 27215 5256
rect 27157 5247 27215 5253
rect 27338 5244 27344 5256
rect 27396 5244 27402 5296
rect 28902 5244 28908 5296
rect 28960 5284 28966 5296
rect 28960 5256 30052 5284
rect 28960 5244 28966 5256
rect 30024 5228 30052 5256
rect 26786 5176 26792 5228
rect 26844 5216 26850 5228
rect 27433 5219 27491 5225
rect 27433 5216 27445 5219
rect 26844 5188 27445 5216
rect 26844 5176 26850 5188
rect 27433 5185 27445 5188
rect 27479 5185 27491 5219
rect 27433 5179 27491 5185
rect 27709 5219 27767 5225
rect 27709 5185 27721 5219
rect 27755 5216 27767 5219
rect 28074 5216 28080 5228
rect 27755 5188 28080 5216
rect 27755 5185 27767 5188
rect 27709 5179 27767 5185
rect 28074 5176 28080 5188
rect 28132 5176 28138 5228
rect 28353 5219 28411 5225
rect 28353 5185 28365 5219
rect 28399 5216 28411 5219
rect 29638 5216 29644 5228
rect 28399 5188 29644 5216
rect 28399 5185 28411 5188
rect 28353 5179 28411 5185
rect 29638 5176 29644 5188
rect 29696 5176 29702 5228
rect 30006 5216 30012 5228
rect 29967 5188 30012 5216
rect 30006 5176 30012 5188
rect 30064 5176 30070 5228
rect 30282 5176 30288 5228
rect 30340 5216 30346 5228
rect 31205 5219 31263 5225
rect 31205 5216 31217 5219
rect 30340 5188 31217 5216
rect 30340 5176 30346 5188
rect 31205 5185 31217 5188
rect 31251 5185 31263 5219
rect 31205 5179 31263 5185
rect 25317 5151 25375 5157
rect 25317 5148 25329 5151
rect 25148 5120 25329 5148
rect 25317 5117 25329 5120
rect 25363 5117 25375 5151
rect 25317 5111 25375 5117
rect 25590 5108 25596 5160
rect 25648 5148 25654 5160
rect 25777 5151 25835 5157
rect 25777 5148 25789 5151
rect 25648 5120 25789 5148
rect 25648 5108 25654 5120
rect 25777 5117 25789 5120
rect 25823 5117 25835 5151
rect 25777 5111 25835 5117
rect 26050 5108 26056 5160
rect 26108 5148 26114 5160
rect 26145 5151 26203 5157
rect 26145 5148 26157 5151
rect 26108 5120 26157 5148
rect 26108 5108 26114 5120
rect 26145 5117 26157 5120
rect 26191 5117 26203 5151
rect 26145 5111 26203 5117
rect 26326 5108 26332 5160
rect 26384 5148 26390 5160
rect 26513 5151 26571 5157
rect 26513 5148 26525 5151
rect 26384 5120 26525 5148
rect 26384 5108 26390 5120
rect 26513 5117 26525 5120
rect 26559 5117 26571 5151
rect 26513 5111 26571 5117
rect 18370 5083 18428 5089
rect 18370 5080 18382 5083
rect 17788 5052 18382 5080
rect 17788 5024 17816 5052
rect 18370 5049 18382 5052
rect 18416 5049 18428 5083
rect 18370 5043 18428 5049
rect 26789 5083 26847 5089
rect 26789 5049 26801 5083
rect 26835 5080 26847 5083
rect 27522 5080 27528 5092
rect 26835 5052 27528 5080
rect 26835 5049 26847 5052
rect 26789 5043 26847 5049
rect 27522 5040 27528 5052
rect 27580 5040 27586 5092
rect 27801 5083 27859 5089
rect 27801 5049 27813 5083
rect 27847 5080 27859 5083
rect 28166 5080 28172 5092
rect 27847 5052 28172 5080
rect 27847 5049 27859 5052
rect 27801 5043 27859 5049
rect 28166 5040 28172 5052
rect 28224 5040 28230 5092
rect 29362 5080 29368 5092
rect 29323 5052 29368 5080
rect 29362 5040 29368 5052
rect 29420 5040 29426 5092
rect 29454 5040 29460 5092
rect 29512 5080 29518 5092
rect 30926 5080 30932 5092
rect 29512 5052 29557 5080
rect 30887 5052 30932 5080
rect 29512 5040 29518 5052
rect 30926 5040 30932 5052
rect 30984 5040 30990 5092
rect 31018 5040 31024 5092
rect 31076 5080 31082 5092
rect 31076 5052 31121 5080
rect 31076 5040 31082 5052
rect 15286 5012 15292 5024
rect 11931 4984 13768 5012
rect 15247 4984 15292 5012
rect 11931 4981 11943 4984
rect 11885 4975 11943 4981
rect 15286 4972 15292 4984
rect 15344 4972 15350 5024
rect 17770 5012 17776 5024
rect 17731 4984 17776 5012
rect 17770 4972 17776 4984
rect 17828 4972 17834 5024
rect 18969 5015 19027 5021
rect 18969 4981 18981 5015
rect 19015 5012 19027 5015
rect 19242 5012 19248 5024
rect 19015 4984 19248 5012
rect 19015 4981 19027 4984
rect 18969 4975 19027 4981
rect 19242 4972 19248 4984
rect 19300 4972 19306 5024
rect 20806 5012 20812 5024
rect 20767 4984 20812 5012
rect 20806 4972 20812 4984
rect 20864 4972 20870 5024
rect 23474 5012 23480 5024
rect 23435 4984 23480 5012
rect 23474 4972 23480 4984
rect 23532 4972 23538 5024
rect 28810 5012 28816 5024
rect 28771 4984 28816 5012
rect 28810 4972 28816 4984
rect 28868 4972 28874 5024
rect 29472 5012 29500 5040
rect 30285 5015 30343 5021
rect 30285 5012 30297 5015
rect 29472 4984 30297 5012
rect 30285 4981 30297 4984
rect 30331 5012 30343 5015
rect 30558 5012 30564 5024
rect 30331 4984 30564 5012
rect 30331 4981 30343 4984
rect 30285 4975 30343 4981
rect 30558 4972 30564 4984
rect 30616 4972 30622 5024
rect 1104 4922 38824 4944
rect 1104 4870 14315 4922
rect 14367 4870 14379 4922
rect 14431 4870 14443 4922
rect 14495 4870 14507 4922
rect 14559 4870 27648 4922
rect 27700 4870 27712 4922
rect 27764 4870 27776 4922
rect 27828 4870 27840 4922
rect 27892 4870 38824 4922
rect 1104 4848 38824 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 2832 4780 2877 4808
rect 2832 4768 2838 4780
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4856 4780 5089 4808
rect 4856 4768 4862 4780
rect 5077 4777 5089 4780
rect 5123 4808 5135 4811
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 5123 4780 5549 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5537 4777 5549 4780
rect 5583 4808 5595 4811
rect 5718 4808 5724 4820
rect 5583 4780 5724 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5718 4768 5724 4780
rect 5776 4808 5782 4820
rect 5776 4780 6316 4808
rect 5776 4768 5782 4780
rect 1670 4700 1676 4752
rect 1728 4740 1734 4752
rect 1810 4743 1868 4749
rect 1810 4740 1822 4743
rect 1728 4712 1822 4740
rect 1728 4700 1734 4712
rect 1810 4709 1822 4712
rect 1856 4709 1868 4743
rect 1810 4703 1868 4709
rect 3881 4743 3939 4749
rect 3881 4709 3893 4743
rect 3927 4740 3939 4743
rect 5166 4740 5172 4752
rect 3927 4712 5172 4740
rect 3927 4709 3939 4712
rect 3881 4703 3939 4709
rect 5166 4700 5172 4712
rect 5224 4740 5230 4752
rect 6288 4740 6316 4780
rect 6822 4768 6828 4820
rect 6880 4808 6886 4820
rect 6917 4811 6975 4817
rect 6917 4808 6929 4811
rect 6880 4780 6929 4808
rect 6880 4768 6886 4780
rect 6917 4777 6929 4780
rect 6963 4777 6975 4811
rect 6917 4771 6975 4777
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7837 4811 7895 4817
rect 7837 4808 7849 4811
rect 7064 4780 7849 4808
rect 7064 4768 7070 4780
rect 7837 4777 7849 4780
rect 7883 4777 7895 4811
rect 9490 4808 9496 4820
rect 9451 4780 9496 4808
rect 7837 4771 7895 4777
rect 9490 4768 9496 4780
rect 9548 4768 9554 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12710 4808 12716 4820
rect 12308 4780 12716 4808
rect 12308 4768 12314 4780
rect 12710 4768 12716 4780
rect 12768 4808 12774 4820
rect 15013 4811 15071 4817
rect 15013 4808 15025 4811
rect 12768 4780 15025 4808
rect 12768 4768 12774 4780
rect 15013 4777 15025 4780
rect 15059 4777 15071 4811
rect 15013 4771 15071 4777
rect 15473 4811 15531 4817
rect 15473 4777 15485 4811
rect 15519 4777 15531 4811
rect 15473 4771 15531 4777
rect 7469 4743 7527 4749
rect 7469 4740 7481 4743
rect 5224 4712 6224 4740
rect 6288 4712 7481 4740
rect 5224 4700 5230 4712
rect 4246 4672 4252 4684
rect 4207 4644 4252 4672
rect 4246 4632 4252 4644
rect 4304 4632 4310 4684
rect 5718 4672 5724 4684
rect 5679 4644 5724 4672
rect 5718 4632 5724 4644
rect 5776 4632 5782 4684
rect 6196 4681 6224 4712
rect 7469 4709 7481 4712
rect 7515 4709 7527 4743
rect 8202 4740 8208 4752
rect 8163 4712 8208 4740
rect 7469 4703 7527 4709
rect 8202 4700 8208 4712
rect 8260 4700 8266 4752
rect 10137 4743 10195 4749
rect 10137 4709 10149 4743
rect 10183 4740 10195 4743
rect 10318 4740 10324 4752
rect 10183 4712 10324 4740
rect 10183 4709 10195 4712
rect 10137 4703 10195 4709
rect 10318 4700 10324 4712
rect 10376 4740 10382 4752
rect 12621 4743 12679 4749
rect 12621 4740 12633 4743
rect 10376 4712 12633 4740
rect 10376 4700 10382 4712
rect 6181 4675 6239 4681
rect 6181 4641 6193 4675
rect 6227 4641 6239 4675
rect 6546 4672 6552 4684
rect 6507 4644 6552 4672
rect 6181 4635 6239 4641
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 7101 4675 7159 4681
rect 7101 4641 7113 4675
rect 7147 4672 7159 4675
rect 7282 4672 7288 4684
rect 7147 4644 7288 4672
rect 7147 4641 7159 4644
rect 7101 4635 7159 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 10520 4681 10548 4712
rect 12621 4709 12633 4712
rect 12667 4740 12679 4743
rect 12802 4740 12808 4752
rect 12667 4712 12808 4740
rect 12667 4709 12679 4712
rect 12621 4703 12679 4709
rect 12802 4700 12808 4712
rect 12860 4700 12866 4752
rect 13814 4749 13820 4752
rect 13811 4740 13820 4749
rect 13775 4712 13820 4740
rect 13811 4703 13820 4712
rect 13814 4700 13820 4703
rect 13872 4700 13878 4752
rect 14090 4700 14096 4752
rect 14148 4740 14154 4752
rect 14645 4743 14703 4749
rect 14645 4740 14657 4743
rect 14148 4712 14657 4740
rect 14148 4700 14154 4712
rect 14645 4709 14657 4712
rect 14691 4740 14703 4743
rect 14918 4740 14924 4752
rect 14691 4712 14924 4740
rect 14691 4709 14703 4712
rect 14645 4703 14703 4709
rect 14918 4700 14924 4712
rect 14976 4740 14982 4752
rect 15488 4740 15516 4771
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 20533 4811 20591 4817
rect 20533 4808 20545 4811
rect 19576 4780 20545 4808
rect 19576 4768 19582 4780
rect 20533 4777 20545 4780
rect 20579 4808 20591 4811
rect 21082 4808 21088 4820
rect 20579 4780 21088 4808
rect 20579 4777 20591 4780
rect 20533 4771 20591 4777
rect 21082 4768 21088 4780
rect 21140 4768 21146 4820
rect 23474 4768 23480 4820
rect 23532 4808 23538 4820
rect 25130 4808 25136 4820
rect 23532 4780 25136 4808
rect 23532 4768 23538 4780
rect 25130 4768 25136 4780
rect 25188 4808 25194 4820
rect 25317 4811 25375 4817
rect 25317 4808 25329 4811
rect 25188 4780 25329 4808
rect 25188 4768 25194 4780
rect 25317 4777 25329 4780
rect 25363 4808 25375 4811
rect 26326 4808 26332 4820
rect 25363 4780 26332 4808
rect 25363 4777 25375 4780
rect 25317 4771 25375 4777
rect 26326 4768 26332 4780
rect 26384 4808 26390 4820
rect 26697 4811 26755 4817
rect 26697 4808 26709 4811
rect 26384 4780 26709 4808
rect 26384 4768 26390 4780
rect 26697 4777 26709 4780
rect 26743 4777 26755 4811
rect 26697 4771 26755 4777
rect 29362 4768 29368 4820
rect 29420 4808 29426 4820
rect 29822 4808 29828 4820
rect 29420 4780 29828 4808
rect 29420 4768 29426 4780
rect 29822 4768 29828 4780
rect 29880 4768 29886 4820
rect 14976 4712 15516 4740
rect 14976 4700 14982 4712
rect 15838 4700 15844 4752
rect 15896 4740 15902 4752
rect 16301 4743 16359 4749
rect 16301 4740 16313 4743
rect 15896 4712 16313 4740
rect 15896 4700 15902 4712
rect 16301 4709 16313 4712
rect 16347 4740 16359 4743
rect 16347 4712 17448 4740
rect 16347 4709 16359 4712
rect 16301 4703 16359 4709
rect 17420 4684 17448 4712
rect 18046 4700 18052 4752
rect 18104 4740 18110 4752
rect 18233 4743 18291 4749
rect 18233 4740 18245 4743
rect 18104 4712 18245 4740
rect 18104 4700 18110 4712
rect 18233 4709 18245 4712
rect 18279 4740 18291 4743
rect 18509 4743 18567 4749
rect 18509 4740 18521 4743
rect 18279 4712 18521 4740
rect 18279 4709 18291 4712
rect 18233 4703 18291 4709
rect 18509 4709 18521 4712
rect 18555 4709 18567 4743
rect 19334 4740 19340 4752
rect 19295 4712 19340 4740
rect 18509 4703 18567 4709
rect 19334 4700 19340 4712
rect 19392 4700 19398 4752
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 21266 4749 21272 4752
rect 21263 4740 21272 4749
rect 19484 4712 19529 4740
rect 21227 4712 21272 4740
rect 19484 4700 19490 4712
rect 21263 4703 21272 4712
rect 21266 4700 21272 4703
rect 21324 4700 21330 4752
rect 22094 4700 22100 4752
rect 22152 4740 22158 4752
rect 22830 4740 22836 4752
rect 22152 4712 22836 4740
rect 22152 4700 22158 4712
rect 22830 4700 22836 4712
rect 22888 4700 22894 4752
rect 24854 4740 24860 4752
rect 24815 4712 24860 4740
rect 24854 4700 24860 4712
rect 24912 4740 24918 4752
rect 25685 4743 25743 4749
rect 25685 4740 25697 4743
rect 24912 4712 25697 4740
rect 24912 4700 24918 4712
rect 25685 4709 25697 4712
rect 25731 4740 25743 4743
rect 26050 4740 26056 4752
rect 25731 4712 26056 4740
rect 25731 4709 25743 4712
rect 25685 4703 25743 4709
rect 26050 4700 26056 4712
rect 26108 4700 26114 4752
rect 26237 4743 26295 4749
rect 26237 4740 26249 4743
rect 26160 4712 26249 4740
rect 10505 4675 10563 4681
rect 10505 4641 10517 4675
rect 10551 4641 10563 4675
rect 10962 4672 10968 4684
rect 10923 4644 10968 4672
rect 10505 4635 10563 4641
rect 10962 4632 10968 4644
rect 11020 4632 11026 4684
rect 11149 4675 11207 4681
rect 11149 4641 11161 4675
rect 11195 4641 11207 4675
rect 11149 4635 11207 4641
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 2498 4604 2504 4616
rect 1535 4576 2504 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 6788 4576 8125 4604
rect 6788 4564 6794 4576
rect 8113 4573 8125 4576
rect 8159 4604 8171 4607
rect 8294 4604 8300 4616
rect 8159 4576 8300 4604
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 8478 4604 8484 4616
rect 8439 4576 8484 4604
rect 8478 4564 8484 4576
rect 8536 4564 8542 4616
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 11164 4604 11192 4635
rect 11238 4632 11244 4684
rect 11296 4672 11302 4684
rect 11425 4675 11483 4681
rect 11425 4672 11437 4675
rect 11296 4644 11437 4672
rect 11296 4632 11302 4644
rect 11425 4641 11437 4644
rect 11471 4672 11483 4675
rect 13446 4672 13452 4684
rect 11471 4644 12940 4672
rect 13407 4644 13452 4672
rect 11471 4641 11483 4644
rect 11425 4635 11483 4641
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 10928 4576 12265 4604
rect 10928 4564 10934 4576
rect 12253 4573 12265 4576
rect 12299 4604 12311 4607
rect 12342 4604 12348 4616
rect 12299 4576 12348 4604
rect 12299 4573 12311 4576
rect 12253 4567 12311 4573
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 11606 4536 11612 4548
rect 11567 4508 11612 4536
rect 11606 4496 11612 4508
rect 11664 4496 11670 4548
rect 12912 4536 12940 4644
rect 13446 4632 13452 4644
rect 13504 4632 13510 4684
rect 15289 4675 15347 4681
rect 15289 4641 15301 4675
rect 15335 4672 15347 4675
rect 15654 4672 15660 4684
rect 15335 4644 15660 4672
rect 15335 4641 15347 4644
rect 15289 4635 15347 4641
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 16669 4675 16727 4681
rect 16669 4641 16681 4675
rect 16715 4672 16727 4675
rect 16758 4672 16764 4684
rect 16715 4644 16764 4672
rect 16715 4641 16727 4644
rect 16669 4635 16727 4641
rect 16758 4632 16764 4644
rect 16816 4672 16822 4684
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16816 4644 17049 4672
rect 16816 4632 16822 4644
rect 17037 4641 17049 4644
rect 17083 4672 17095 4675
rect 17218 4672 17224 4684
rect 17083 4644 17224 4672
rect 17083 4641 17095 4644
rect 17037 4635 17095 4641
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 17402 4672 17408 4684
rect 17363 4644 17408 4672
rect 17402 4632 17408 4644
rect 17460 4632 17466 4684
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4641 17647 4675
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 17589 4635 17647 4641
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 17604 4604 17632 4635
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 20714 4632 20720 4684
rect 20772 4672 20778 4684
rect 20901 4675 20959 4681
rect 20901 4672 20913 4675
rect 20772 4644 20913 4672
rect 20772 4632 20778 4644
rect 20901 4641 20913 4644
rect 20947 4672 20959 4675
rect 21358 4672 21364 4684
rect 20947 4644 21364 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 24213 4675 24271 4681
rect 24213 4641 24225 4675
rect 24259 4672 24271 4675
rect 24670 4672 24676 4684
rect 24259 4644 24676 4672
rect 24259 4641 24271 4644
rect 24213 4635 24271 4641
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 19978 4604 19984 4616
rect 16632 4576 17632 4604
rect 19891 4576 19984 4604
rect 16632 4564 16638 4576
rect 19978 4564 19984 4576
rect 20036 4604 20042 4616
rect 22738 4604 22744 4616
rect 20036 4576 22744 4604
rect 20036 4564 20042 4576
rect 22738 4564 22744 4576
rect 22796 4564 22802 4616
rect 23017 4607 23075 4613
rect 23017 4573 23029 4607
rect 23063 4573 23075 4607
rect 23017 4567 23075 4573
rect 12989 4539 13047 4545
rect 12989 4536 13001 4539
rect 12912 4508 13001 4536
rect 12989 4505 13001 4508
rect 13035 4536 13047 4539
rect 13357 4539 13415 4545
rect 13357 4536 13369 4539
rect 13035 4508 13369 4536
rect 13035 4505 13047 4508
rect 12989 4499 13047 4505
rect 13357 4505 13369 4508
rect 13403 4536 13415 4539
rect 13722 4536 13728 4548
rect 13403 4508 13728 4536
rect 13403 4505 13415 4508
rect 13357 4499 13415 4505
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 14369 4539 14427 4545
rect 14369 4505 14381 4539
rect 14415 4536 14427 4539
rect 15841 4539 15899 4545
rect 15841 4536 15853 4539
rect 14415 4508 15853 4536
rect 14415 4505 14427 4508
rect 14369 4499 14427 4505
rect 15841 4505 15853 4508
rect 15887 4536 15899 4539
rect 16114 4536 16120 4548
rect 15887 4508 16120 4536
rect 15887 4505 15899 4508
rect 15841 4499 15899 4505
rect 16114 4496 16120 4508
rect 16172 4496 16178 4548
rect 22094 4496 22100 4548
rect 22152 4536 22158 4548
rect 22554 4536 22560 4548
rect 22152 4508 22560 4536
rect 22152 4496 22158 4508
rect 22554 4496 22560 4508
rect 22612 4536 22618 4548
rect 23032 4536 23060 4567
rect 25590 4564 25596 4616
rect 25648 4604 25654 4616
rect 25866 4604 25872 4616
rect 25648 4576 25872 4604
rect 25648 4564 25654 4576
rect 25866 4564 25872 4576
rect 25924 4604 25930 4616
rect 26160 4604 26188 4712
rect 26237 4709 26249 4712
rect 26283 4709 26295 4743
rect 26237 4703 26295 4709
rect 27154 4700 27160 4752
rect 27212 4749 27218 4752
rect 27212 4743 27260 4749
rect 27212 4709 27214 4743
rect 27248 4709 27260 4743
rect 27212 4703 27260 4709
rect 27212 4700 27218 4703
rect 28810 4700 28816 4752
rect 28868 4740 28874 4752
rect 28950 4743 29008 4749
rect 28950 4740 28962 4743
rect 28868 4712 28962 4740
rect 28868 4700 28874 4712
rect 28950 4709 28962 4712
rect 28996 4709 29008 4743
rect 30558 4740 30564 4752
rect 30519 4712 30564 4740
rect 28950 4703 29008 4709
rect 30558 4700 30564 4712
rect 30616 4700 30622 4752
rect 27801 4675 27859 4681
rect 27801 4641 27813 4675
rect 27847 4672 27859 4675
rect 29454 4672 29460 4684
rect 27847 4644 29460 4672
rect 27847 4641 27859 4644
rect 27801 4635 27859 4641
rect 29454 4632 29460 4644
rect 29512 4632 29518 4684
rect 26878 4604 26884 4616
rect 25924 4576 26188 4604
rect 26839 4576 26884 4604
rect 25924 4564 25930 4576
rect 26878 4564 26884 4576
rect 26936 4564 26942 4616
rect 27522 4564 27528 4616
rect 27580 4604 27586 4616
rect 28626 4604 28632 4616
rect 27580 4576 28632 4604
rect 27580 4564 27586 4576
rect 28626 4564 28632 4576
rect 28684 4564 28690 4616
rect 30466 4604 30472 4616
rect 30427 4576 30472 4604
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 30745 4607 30803 4613
rect 30745 4573 30757 4607
rect 30791 4604 30803 4607
rect 30926 4604 30932 4616
rect 30791 4576 30932 4604
rect 30791 4573 30803 4576
rect 30745 4567 30803 4573
rect 24394 4536 24400 4548
rect 22612 4508 23060 4536
rect 24355 4508 24400 4536
rect 22612 4496 22618 4508
rect 24394 4496 24400 4508
rect 24452 4496 24458 4548
rect 30374 4496 30380 4548
rect 30432 4536 30438 4548
rect 30760 4536 30788 4567
rect 30926 4564 30932 4576
rect 30984 4564 30990 4616
rect 30432 4508 30788 4536
rect 30432 4496 30438 4508
rect 1946 4428 1952 4480
rect 2004 4468 2010 4480
rect 2409 4471 2467 4477
rect 2409 4468 2421 4471
rect 2004 4440 2421 4468
rect 2004 4428 2010 4440
rect 2409 4437 2421 4440
rect 2455 4437 2467 4471
rect 2409 4431 2467 4437
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 4341 4471 4399 4477
rect 4341 4468 4353 4471
rect 3936 4440 4353 4468
rect 3936 4428 3942 4440
rect 4341 4437 4353 4440
rect 4387 4437 4399 4471
rect 21818 4468 21824 4480
rect 21779 4440 21824 4468
rect 4341 4431 4399 4437
rect 21818 4428 21824 4440
rect 21876 4428 21882 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 23661 4471 23719 4477
rect 23661 4468 23673 4471
rect 23532 4440 23673 4468
rect 23532 4428 23538 4440
rect 23661 4437 23673 4440
rect 23707 4437 23719 4471
rect 28166 4468 28172 4480
rect 28127 4440 28172 4468
rect 23661 4431 23719 4437
rect 28166 4428 28172 4440
rect 28224 4428 28230 4480
rect 28534 4468 28540 4480
rect 28495 4440 28540 4468
rect 28534 4428 28540 4440
rect 28592 4428 28598 4480
rect 29546 4468 29552 4480
rect 29507 4440 29552 4468
rect 29546 4428 29552 4440
rect 29604 4428 29610 4480
rect 1104 4378 38824 4400
rect 1104 4326 7648 4378
rect 7700 4326 7712 4378
rect 7764 4326 7776 4378
rect 7828 4326 7840 4378
rect 7892 4326 20982 4378
rect 21034 4326 21046 4378
rect 21098 4326 21110 4378
rect 21162 4326 21174 4378
rect 21226 4326 34315 4378
rect 34367 4326 34379 4378
rect 34431 4326 34443 4378
rect 34495 4326 34507 4378
rect 34559 4326 38824 4378
rect 1104 4304 38824 4326
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 5442 4264 5448 4276
rect 4571 4236 5448 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 5442 4224 5448 4236
rect 5500 4224 5506 4276
rect 6454 4264 6460 4276
rect 5828 4236 6460 4264
rect 1688 4196 1716 4224
rect 5828 4208 5856 4236
rect 6454 4224 6460 4236
rect 6512 4264 6518 4276
rect 6549 4267 6607 4273
rect 6549 4264 6561 4267
rect 6512 4236 6561 4264
rect 6512 4224 6518 4236
rect 6549 4233 6561 4236
rect 6595 4233 6607 4267
rect 6549 4227 6607 4233
rect 8113 4267 8171 4273
rect 8113 4233 8125 4267
rect 8159 4264 8171 4267
rect 8202 4264 8208 4276
rect 8159 4236 8208 4264
rect 8159 4233 8171 4236
rect 8113 4227 8171 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 10318 4224 10324 4276
rect 10376 4264 10382 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10376 4236 10609 4264
rect 10376 4224 10382 4236
rect 10597 4233 10609 4236
rect 10643 4233 10655 4267
rect 10962 4264 10968 4276
rect 10923 4236 10968 4264
rect 10597 4227 10655 4233
rect 10962 4224 10968 4236
rect 11020 4224 11026 4276
rect 15473 4267 15531 4273
rect 15473 4233 15485 4267
rect 15519 4264 15531 4267
rect 15654 4264 15660 4276
rect 15519 4236 15660 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 15654 4224 15660 4236
rect 15712 4224 15718 4276
rect 15838 4264 15844 4276
rect 15799 4236 15844 4264
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 16574 4224 16580 4276
rect 16632 4264 16638 4276
rect 16945 4267 17003 4273
rect 16945 4264 16957 4267
rect 16632 4236 16957 4264
rect 16632 4224 16638 4236
rect 16945 4233 16957 4236
rect 16991 4233 17003 4267
rect 16945 4227 17003 4233
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19392 4236 19717 4264
rect 19392 4224 19398 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 20993 4267 21051 4273
rect 20993 4233 21005 4267
rect 21039 4264 21051 4267
rect 21266 4264 21272 4276
rect 21039 4236 21272 4264
rect 21039 4233 21051 4236
rect 20993 4227 21051 4233
rect 5810 4196 5816 4208
rect 1688 4168 5816 4196
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6638 4196 6644 4208
rect 6551 4168 6644 4196
rect 6638 4156 6644 4168
rect 6696 4196 6702 4208
rect 8478 4196 8484 4208
rect 6696 4168 8484 4196
rect 6696 4156 6702 4168
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 12618 4196 12624 4208
rect 12360 4168 12624 4196
rect 1857 4131 1915 4137
rect 1857 4097 1869 4131
rect 1903 4128 1915 4131
rect 2590 4128 2596 4140
rect 1903 4100 2596 4128
rect 1903 4097 1915 4100
rect 1857 4091 1915 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3016 4100 3709 4128
rect 3016 4088 3022 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 5905 4131 5963 4137
rect 5905 4097 5917 4131
rect 5951 4128 5963 4131
rect 6656 4128 6684 4156
rect 6822 4128 6828 4140
rect 5951 4100 6684 4128
rect 6783 4100 6828 4128
rect 5951 4097 5963 4100
rect 5905 4091 5963 4097
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 8294 4088 8300 4140
rect 8352 4128 8358 4140
rect 8389 4131 8447 4137
rect 8389 4128 8401 4131
rect 8352 4100 8401 4128
rect 8352 4088 8358 4100
rect 8389 4097 8401 4100
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8941 4131 8999 4137
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9401 4131 9459 4137
rect 9401 4128 9413 4131
rect 8987 4100 9413 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9401 4097 9413 4100
rect 9447 4128 9459 4131
rect 9582 4128 9588 4140
rect 9447 4100 9588 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4128 11667 4131
rect 12360 4128 12388 4168
rect 12618 4156 12624 4168
rect 12676 4156 12682 4208
rect 21008 4196 21036 4227
rect 21266 4224 21272 4236
rect 21324 4224 21330 4276
rect 22830 4264 22836 4276
rect 22791 4236 22836 4264
rect 22830 4224 22836 4236
rect 22888 4224 22894 4276
rect 25130 4264 25136 4276
rect 25091 4236 25136 4264
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 27154 4224 27160 4276
rect 27212 4264 27218 4276
rect 28629 4267 28687 4273
rect 28629 4264 28641 4267
rect 27212 4236 28641 4264
rect 27212 4224 27218 4236
rect 28629 4233 28641 4236
rect 28675 4264 28687 4267
rect 28810 4264 28816 4276
rect 28675 4236 28816 4264
rect 28675 4233 28687 4236
rect 28629 4227 28687 4233
rect 28810 4224 28816 4236
rect 28868 4224 28874 4276
rect 30558 4224 30564 4276
rect 30616 4264 30622 4276
rect 30653 4267 30711 4273
rect 30653 4264 30665 4267
rect 30616 4236 30665 4264
rect 30616 4224 30622 4236
rect 30653 4233 30665 4236
rect 30699 4233 30711 4267
rect 30653 4227 30711 4233
rect 18616 4168 21036 4196
rect 26697 4199 26755 4205
rect 11655 4100 12388 4128
rect 11655 4097 11667 4100
rect 11609 4091 11667 4097
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 14182 4128 14188 4140
rect 12492 4100 12537 4128
rect 14143 4100 14188 4128
rect 12492 4088 12498 4100
rect 14182 4088 14188 4100
rect 14240 4088 14246 4140
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 15436 4100 16313 4128
rect 15436 4088 15442 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4128 17463 4131
rect 17862 4128 17868 4140
rect 17451 4100 17868 4128
rect 17451 4097 17463 4100
rect 17405 4091 17463 4097
rect 17862 4088 17868 4100
rect 17920 4088 17926 4140
rect 18141 4131 18199 4137
rect 18141 4097 18153 4131
rect 18187 4128 18199 4131
rect 18506 4128 18512 4140
rect 18187 4100 18512 4128
rect 18187 4097 18199 4100
rect 18141 4091 18199 4097
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 6270 4060 6276 4072
rect 6231 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 11400 4063 11458 4069
rect 11400 4029 11412 4063
rect 11446 4060 11458 4063
rect 11446 4032 11928 4060
rect 11446 4029 11458 4032
rect 11400 4023 11458 4029
rect 1946 3992 1952 4004
rect 1907 3964 1952 3992
rect 1946 3952 1952 3964
rect 2004 3952 2010 4004
rect 2314 3952 2320 4004
rect 2372 3992 2378 4004
rect 2501 3995 2559 4001
rect 2501 3992 2513 3995
rect 2372 3964 2513 3992
rect 2372 3952 2378 3964
rect 2501 3961 2513 3964
rect 2547 3961 2559 3995
rect 3418 3992 3424 4004
rect 3379 3964 3424 3992
rect 2501 3955 2559 3961
rect 3418 3952 3424 3964
rect 3476 3952 3482 4004
rect 3513 3995 3571 4001
rect 3513 3961 3525 3995
rect 3559 3992 3571 3995
rect 3878 3992 3884 4004
rect 3559 3964 3884 3992
rect 3559 3961 3571 3964
rect 3513 3955 3571 3961
rect 1964 3924 1992 3952
rect 2777 3927 2835 3933
rect 2777 3924 2789 3927
rect 1964 3896 2789 3924
rect 2777 3893 2789 3896
rect 2823 3924 2835 3927
rect 2866 3924 2872 3936
rect 2823 3896 2872 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3528 3924 3556 3955
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 5258 3992 5264 4004
rect 5219 3964 5264 3992
rect 5258 3952 5264 3964
rect 5316 3952 5322 4004
rect 5350 3952 5356 4004
rect 5408 3992 5414 4004
rect 5408 3964 5453 3992
rect 5408 3952 5414 3964
rect 6454 3952 6460 4004
rect 6512 3992 6518 4004
rect 7146 3995 7204 4001
rect 7146 3992 7158 3995
rect 6512 3964 7158 3992
rect 6512 3952 6518 3964
rect 7146 3961 7158 3964
rect 7192 3992 7204 3995
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 7192 3964 9229 3992
rect 7192 3961 7204 3964
rect 7146 3955 7204 3961
rect 9217 3961 9229 3964
rect 9263 3992 9275 3995
rect 9722 3995 9780 4001
rect 9722 3992 9734 3995
rect 9263 3964 9734 3992
rect 9263 3961 9275 3964
rect 9217 3955 9275 3961
rect 9722 3961 9734 3964
rect 9768 3992 9780 3995
rect 10778 3992 10784 4004
rect 9768 3964 10784 3992
rect 9768 3961 9780 3964
rect 9722 3955 9780 3961
rect 10778 3952 10784 3964
rect 10836 3952 10842 4004
rect 3283 3896 3556 3924
rect 5077 3927 5135 3933
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5368 3924 5396 3952
rect 11900 3936 11928 4032
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 15102 4060 15108 4072
rect 13780 4032 15108 4060
rect 13780 4020 13786 4032
rect 15102 4020 15108 4032
rect 15160 4020 15166 4072
rect 12799 3995 12857 4001
rect 12799 3992 12811 3995
rect 12268 3964 12811 3992
rect 5123 3896 5396 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7524 3896 7757 3924
rect 7524 3884 7530 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 10318 3924 10324 3936
rect 10279 3896 10324 3924
rect 7745 3887 7803 3893
rect 10318 3884 10324 3896
rect 10376 3884 10382 3936
rect 11054 3884 11060 3936
rect 11112 3924 11118 3936
rect 11471 3927 11529 3933
rect 11471 3924 11483 3927
rect 11112 3896 11483 3924
rect 11112 3884 11118 3896
rect 11471 3893 11483 3896
rect 11517 3924 11529 3927
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 11517 3896 11621 3924
rect 11517 3893 11529 3896
rect 11471 3887 11529 3893
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11882 3924 11888 3936
rect 11843 3896 11888 3924
rect 11609 3887 11667 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12268 3933 12296 3964
rect 12799 3961 12811 3964
rect 12845 3992 12857 3995
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 12845 3964 13645 3992
rect 12845 3961 12857 3964
rect 12799 3955 12857 3961
rect 13633 3961 13645 3964
rect 13679 3992 13691 3995
rect 13814 3992 13820 4004
rect 13679 3964 13820 3992
rect 13679 3961 13691 3964
rect 13633 3955 13691 3961
rect 13814 3952 13820 3964
rect 13872 3992 13878 4004
rect 14093 3995 14151 4001
rect 14093 3992 14105 3995
rect 13872 3964 14105 3992
rect 13872 3952 13878 3964
rect 14093 3961 14105 3964
rect 14139 3992 14151 3995
rect 14547 3995 14605 4001
rect 14547 3992 14559 3995
rect 14139 3964 14559 3992
rect 14139 3961 14151 3964
rect 14093 3955 14151 3961
rect 14547 3961 14559 3964
rect 14593 3992 14605 3995
rect 14734 3992 14740 4004
rect 14593 3964 14740 3992
rect 14593 3961 14605 3964
rect 14547 3955 14605 3961
rect 14734 3952 14740 3964
rect 14792 3952 14798 4004
rect 15010 3952 15016 4004
rect 15068 3992 15074 4004
rect 16025 3995 16083 4001
rect 16025 3992 16037 3995
rect 15068 3964 16037 3992
rect 15068 3952 15074 3964
rect 16025 3961 16037 3964
rect 16071 3961 16083 3995
rect 16025 3955 16083 3961
rect 16114 3952 16120 4004
rect 16172 3992 16178 4004
rect 16172 3964 16217 3992
rect 16172 3952 16178 3964
rect 17770 3952 17776 4004
rect 17828 3992 17834 4004
rect 17865 3995 17923 4001
rect 17865 3992 17877 3995
rect 17828 3964 17877 3992
rect 17828 3952 17834 3964
rect 17865 3961 17877 3964
rect 17911 3992 17923 3995
rect 18503 3995 18561 4001
rect 18503 3992 18515 3995
rect 17911 3964 18515 3992
rect 17911 3961 17923 3964
rect 17865 3955 17923 3961
rect 18503 3961 18515 3964
rect 18549 3992 18561 3995
rect 18616 3992 18644 4168
rect 26697 4165 26709 4199
rect 26743 4196 26755 4199
rect 26878 4196 26884 4208
rect 26743 4168 26884 4196
rect 26743 4165 26755 4168
rect 26697 4159 26755 4165
rect 26878 4156 26884 4168
rect 26936 4196 26942 4208
rect 27430 4196 27436 4208
rect 26936 4168 27436 4196
rect 26936 4156 26942 4168
rect 27430 4156 27436 4168
rect 27488 4156 27494 4208
rect 28534 4156 28540 4208
rect 28592 4196 28598 4208
rect 28592 4168 28948 4196
rect 28592 4156 28598 4168
rect 20806 4088 20812 4140
rect 20864 4128 20870 4140
rect 21269 4131 21327 4137
rect 21269 4128 21281 4131
rect 20864 4100 21281 4128
rect 20864 4088 20870 4100
rect 21269 4097 21281 4100
rect 21315 4128 21327 4131
rect 22465 4131 22523 4137
rect 22465 4128 22477 4131
rect 21315 4100 22477 4128
rect 21315 4097 21327 4100
rect 21269 4091 21327 4097
rect 22465 4097 22477 4100
rect 22511 4097 22523 4131
rect 22465 4091 22523 4097
rect 22738 4088 22744 4140
rect 22796 4128 22802 4140
rect 24029 4131 24087 4137
rect 24029 4128 24041 4131
rect 22796 4100 24041 4128
rect 22796 4088 22802 4100
rect 24029 4097 24041 4100
rect 24075 4097 24087 4131
rect 28920 4128 28948 4168
rect 29365 4131 29423 4137
rect 29365 4128 29377 4131
rect 28920 4100 29377 4128
rect 24029 4091 24087 4097
rect 29365 4097 29377 4100
rect 29411 4128 29423 4131
rect 30975 4131 31033 4137
rect 30975 4128 30987 4131
rect 29411 4100 30987 4128
rect 29411 4097 29423 4100
rect 29365 4091 29423 4097
rect 30975 4097 30987 4100
rect 31021 4097 31033 4131
rect 30975 4091 31033 4097
rect 19940 4063 19998 4069
rect 19940 4029 19952 4063
rect 19986 4060 19998 4063
rect 25590 4060 25596 4072
rect 19986 4032 20484 4060
rect 25551 4032 25596 4060
rect 19986 4029 19998 4032
rect 19940 4023 19998 4029
rect 18549 3964 18644 3992
rect 18549 3961 18561 3964
rect 18503 3955 18561 3961
rect 19610 3952 19616 4004
rect 19668 3992 19674 4004
rect 20027 3995 20085 4001
rect 20027 3992 20039 3995
rect 19668 3964 20039 3992
rect 19668 3952 19674 3964
rect 20027 3961 20039 3964
rect 20073 3961 20085 3995
rect 20027 3955 20085 3961
rect 20456 3936 20484 4032
rect 25590 4020 25596 4032
rect 25648 4020 25654 4072
rect 25866 4060 25872 4072
rect 25827 4032 25872 4060
rect 25866 4020 25872 4032
rect 25924 4020 25930 4072
rect 26050 4020 26056 4072
rect 26108 4060 26114 4072
rect 26145 4063 26203 4069
rect 26145 4060 26157 4063
rect 26108 4032 26157 4060
rect 26108 4020 26114 4032
rect 26145 4029 26157 4032
rect 26191 4029 26203 4063
rect 26145 4023 26203 4029
rect 26326 4020 26332 4072
rect 26384 4060 26390 4072
rect 26513 4063 26571 4069
rect 26513 4060 26525 4063
rect 26384 4032 26525 4060
rect 26384 4020 26390 4032
rect 26513 4029 26525 4032
rect 26559 4029 26571 4063
rect 26513 4023 26571 4029
rect 28353 4063 28411 4069
rect 28353 4029 28365 4063
rect 28399 4060 28411 4063
rect 28902 4060 28908 4072
rect 28399 4032 28908 4060
rect 28399 4029 28411 4032
rect 28353 4023 28411 4029
rect 28902 4020 28908 4032
rect 28960 4020 28966 4072
rect 30282 4060 30288 4072
rect 30024 4032 30288 4060
rect 21266 3952 21272 4004
rect 21324 3992 21330 4004
rect 21590 3995 21648 4001
rect 21590 3992 21602 3995
rect 21324 3964 21602 3992
rect 21324 3952 21330 3964
rect 21590 3961 21602 3964
rect 21636 3961 21648 3995
rect 21590 3955 21648 3961
rect 23474 3952 23480 4004
rect 23532 3992 23538 4004
rect 23753 3995 23811 4001
rect 23753 3992 23765 3995
rect 23532 3964 23765 3992
rect 23532 3952 23538 3964
rect 23753 3961 23765 3964
rect 23799 3961 23811 3995
rect 23753 3955 23811 3961
rect 23845 3995 23903 4001
rect 23845 3961 23857 3995
rect 23891 3961 23903 3995
rect 23845 3955 23903 3961
rect 12253 3927 12311 3933
rect 12253 3924 12265 3927
rect 12032 3896 12265 3924
rect 12032 3884 12038 3896
rect 12253 3893 12265 3896
rect 12299 3893 12311 3927
rect 13354 3924 13360 3936
rect 13315 3896 13360 3924
rect 12253 3887 12311 3893
rect 13354 3884 13360 3896
rect 13412 3884 13418 3936
rect 19061 3927 19119 3933
rect 19061 3893 19073 3927
rect 19107 3924 19119 3927
rect 19426 3924 19432 3936
rect 19107 3896 19432 3924
rect 19107 3893 19119 3896
rect 19061 3887 19119 3893
rect 19426 3884 19432 3896
rect 19484 3884 19490 3936
rect 20438 3924 20444 3936
rect 20399 3896 20444 3924
rect 20438 3884 20444 3896
rect 20496 3884 20502 3936
rect 22002 3884 22008 3936
rect 22060 3924 22066 3936
rect 22189 3927 22247 3933
rect 22189 3924 22201 3927
rect 22060 3896 22201 3924
rect 22060 3884 22066 3896
rect 22189 3893 22201 3896
rect 22235 3924 22247 3927
rect 23385 3927 23443 3933
rect 23385 3924 23397 3927
rect 22235 3896 23397 3924
rect 22235 3893 22247 3896
rect 22189 3887 22247 3893
rect 23385 3893 23397 3896
rect 23431 3924 23443 3927
rect 23860 3924 23888 3955
rect 27522 3952 27528 4004
rect 27580 3992 27586 4004
rect 27709 3995 27767 4001
rect 27709 3992 27721 3995
rect 27580 3964 27721 3992
rect 27580 3952 27586 3964
rect 27709 3961 27721 3964
rect 27755 3961 27767 3995
rect 27709 3955 27767 3961
rect 27801 3995 27859 4001
rect 27801 3961 27813 3995
rect 27847 3961 27859 3995
rect 29457 3995 29515 4001
rect 27801 3955 27859 3961
rect 28460 3964 29132 3992
rect 24670 3924 24676 3936
rect 23431 3896 23888 3924
rect 24631 3896 24676 3924
rect 23431 3893 23443 3896
rect 23385 3887 23443 3893
rect 24670 3884 24676 3896
rect 24728 3884 24734 3936
rect 26602 3884 26608 3936
rect 26660 3924 26666 3936
rect 27065 3927 27123 3933
rect 27065 3924 27077 3927
rect 26660 3896 27077 3924
rect 26660 3884 26666 3896
rect 27065 3893 27077 3896
rect 27111 3924 27123 3927
rect 27154 3924 27160 3936
rect 27111 3896 27160 3924
rect 27111 3893 27123 3896
rect 27065 3887 27123 3893
rect 27154 3884 27160 3896
rect 27212 3884 27218 3936
rect 27433 3927 27491 3933
rect 27433 3893 27445 3927
rect 27479 3924 27491 3927
rect 27816 3924 27844 3955
rect 28460 3924 28488 3964
rect 29104 3933 29132 3964
rect 29457 3961 29469 3995
rect 29503 3992 29515 3995
rect 29546 3992 29552 4004
rect 29503 3964 29552 3992
rect 29503 3961 29515 3964
rect 29457 3955 29515 3961
rect 27479 3896 28488 3924
rect 29089 3927 29147 3933
rect 27479 3893 27491 3896
rect 27433 3887 27491 3893
rect 29089 3893 29101 3927
rect 29135 3924 29147 3927
rect 29472 3924 29500 3955
rect 29546 3952 29552 3964
rect 29604 3952 29610 4004
rect 29638 3952 29644 4004
rect 29696 3992 29702 4004
rect 30024 4001 30052 4032
rect 30282 4020 30288 4032
rect 30340 4020 30346 4072
rect 30374 4020 30380 4072
rect 30432 4060 30438 4072
rect 30432 4032 30477 4060
rect 30432 4020 30438 4032
rect 30834 4020 30840 4072
rect 30892 4069 30898 4072
rect 30892 4063 30930 4069
rect 30918 4060 30930 4063
rect 31297 4063 31355 4069
rect 31297 4060 31309 4063
rect 30918 4032 31309 4060
rect 30918 4029 30930 4032
rect 30892 4023 30930 4029
rect 31297 4029 31309 4032
rect 31343 4029 31355 4063
rect 31297 4023 31355 4029
rect 30892 4020 30898 4023
rect 30009 3995 30067 4001
rect 30009 3992 30021 3995
rect 29696 3964 30021 3992
rect 29696 3952 29702 3964
rect 30009 3961 30021 3964
rect 30055 3961 30067 3995
rect 30009 3955 30067 3961
rect 29135 3896 29500 3924
rect 29135 3893 29147 3896
rect 29089 3887 29147 3893
rect 1104 3834 38824 3856
rect 1104 3782 14315 3834
rect 14367 3782 14379 3834
rect 14431 3782 14443 3834
rect 14495 3782 14507 3834
rect 14559 3782 27648 3834
rect 27700 3782 27712 3834
rect 27764 3782 27776 3834
rect 27828 3782 27840 3834
rect 27892 3782 38824 3834
rect 1104 3760 38824 3782
rect 1486 3680 1492 3732
rect 1544 3680 1550 3732
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 2590 3680 2596 3732
rect 2648 3720 2654 3732
rect 2958 3720 2964 3732
rect 2648 3692 2964 3720
rect 2648 3680 2654 3692
rect 2958 3680 2964 3692
rect 3016 3680 3022 3732
rect 3418 3720 3424 3732
rect 3379 3692 3424 3720
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 4246 3720 4252 3732
rect 4207 3692 4252 3720
rect 4246 3680 4252 3692
rect 4304 3680 4310 3732
rect 5077 3723 5135 3729
rect 5077 3689 5089 3723
rect 5123 3720 5135 3723
rect 5166 3720 5172 3732
rect 5123 3692 5172 3720
rect 5123 3689 5135 3692
rect 5077 3683 5135 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5442 3720 5448 3732
rect 5403 3692 5448 3720
rect 5442 3680 5448 3692
rect 5500 3680 5506 3732
rect 6822 3720 6828 3732
rect 6783 3692 6828 3720
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 9493 3723 9551 3729
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9766 3720 9772 3732
rect 9539 3692 9772 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 9766 3680 9772 3692
rect 9824 3720 9830 3732
rect 10318 3720 10324 3732
rect 9824 3692 10324 3720
rect 9824 3680 9830 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 10689 3723 10747 3729
rect 10689 3689 10701 3723
rect 10735 3720 10747 3723
rect 10870 3720 10876 3732
rect 10735 3692 10876 3720
rect 10735 3689 10747 3692
rect 10689 3683 10747 3689
rect 10870 3680 10876 3692
rect 10928 3680 10934 3732
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 12069 3723 12127 3729
rect 12069 3720 12081 3723
rect 11756 3692 12081 3720
rect 11756 3680 11762 3692
rect 12069 3689 12081 3692
rect 12115 3720 12127 3723
rect 12115 3692 12756 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 1504 3652 1532 3680
rect 1581 3655 1639 3661
rect 1581 3652 1593 3655
rect 1504 3624 1593 3652
rect 1581 3621 1593 3624
rect 1627 3621 1639 3655
rect 1581 3615 1639 3621
rect 1670 3612 1676 3664
rect 1728 3652 1734 3664
rect 3881 3655 3939 3661
rect 1728 3624 1773 3652
rect 1728 3612 1734 3624
rect 3881 3621 3893 3655
rect 3927 3652 3939 3655
rect 5258 3652 5264 3664
rect 3927 3624 5264 3652
rect 3927 3621 3939 3624
rect 3881 3615 3939 3621
rect 5258 3612 5264 3624
rect 5316 3612 5322 3664
rect 5810 3612 5816 3664
rect 5868 3661 5874 3664
rect 5868 3655 5916 3661
rect 5868 3621 5870 3655
rect 5904 3621 5916 3655
rect 7466 3652 7472 3664
rect 7427 3624 7472 3652
rect 5868 3615 5916 3621
rect 5868 3612 5874 3615
rect 7466 3612 7472 3624
rect 7524 3612 7530 3664
rect 10226 3652 10232 3664
rect 10187 3624 10232 3652
rect 10226 3612 10232 3624
rect 10284 3612 10290 3664
rect 10778 3612 10784 3664
rect 10836 3652 10842 3664
rect 11194 3655 11252 3661
rect 11194 3652 11206 3655
rect 10836 3624 11206 3652
rect 10836 3612 10842 3624
rect 11194 3621 11206 3624
rect 11240 3652 11252 3655
rect 11974 3652 11980 3664
rect 11240 3624 11980 3652
rect 11240 3621 11252 3624
rect 11194 3615 11252 3621
rect 11974 3612 11980 3624
rect 12032 3612 12038 3664
rect 12728 3661 12756 3692
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 13633 3723 13691 3729
rect 13633 3720 13645 3723
rect 13504 3692 13645 3720
rect 13504 3680 13510 3692
rect 13633 3689 13645 3692
rect 13679 3689 13691 3723
rect 13633 3683 13691 3689
rect 14182 3680 14188 3732
rect 14240 3720 14246 3732
rect 14645 3723 14703 3729
rect 14645 3720 14657 3723
rect 14240 3692 14657 3720
rect 14240 3680 14246 3692
rect 14645 3689 14657 3692
rect 14691 3689 14703 3723
rect 16758 3720 16764 3732
rect 16719 3692 16764 3720
rect 14645 3683 14703 3689
rect 16758 3680 16764 3692
rect 16816 3680 16822 3732
rect 17770 3720 17776 3732
rect 17052 3692 17776 3720
rect 12713 3655 12771 3661
rect 12713 3621 12725 3655
rect 12759 3621 12771 3655
rect 12713 3615 12771 3621
rect 12805 3655 12863 3661
rect 12805 3621 12817 3655
rect 12851 3652 12863 3655
rect 13354 3652 13360 3664
rect 12851 3624 13360 3652
rect 12851 3621 12863 3624
rect 12805 3615 12863 3621
rect 13354 3612 13360 3624
rect 13412 3612 13418 3664
rect 14734 3612 14740 3664
rect 14792 3652 14798 3664
rect 15651 3655 15709 3661
rect 15651 3652 15663 3655
rect 14792 3624 15663 3652
rect 14792 3612 14798 3624
rect 15651 3621 15663 3624
rect 15697 3652 15709 3655
rect 16114 3652 16120 3664
rect 15697 3624 16120 3652
rect 15697 3621 15709 3624
rect 15651 3615 15709 3621
rect 16114 3612 16120 3624
rect 16172 3652 16178 3664
rect 17052 3652 17080 3692
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 18233 3723 18291 3729
rect 18233 3689 18245 3723
rect 18279 3720 18291 3723
rect 18506 3720 18512 3732
rect 18279 3692 18512 3720
rect 18279 3689 18291 3692
rect 18233 3683 18291 3689
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 20714 3720 20720 3732
rect 20675 3692 20720 3720
rect 20714 3680 20720 3692
rect 20772 3680 20778 3732
rect 21266 3720 21272 3732
rect 21227 3692 21272 3720
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 22738 3720 22744 3732
rect 22699 3692 22744 3720
rect 22738 3680 22744 3692
rect 22796 3680 22802 3732
rect 25409 3723 25467 3729
rect 25409 3689 25421 3723
rect 25455 3720 25467 3723
rect 26050 3720 26056 3732
rect 25455 3692 26056 3720
rect 25455 3689 25467 3692
rect 25409 3683 25467 3689
rect 26050 3680 26056 3692
rect 26108 3680 26114 3732
rect 27430 3680 27436 3732
rect 27488 3720 27494 3732
rect 27709 3723 27767 3729
rect 27709 3720 27721 3723
rect 27488 3692 27721 3720
rect 27488 3680 27494 3692
rect 27709 3689 27721 3692
rect 27755 3689 27767 3723
rect 27709 3683 27767 3689
rect 29822 3680 29828 3732
rect 29880 3720 29886 3732
rect 29963 3723 30021 3729
rect 29963 3720 29975 3723
rect 29880 3692 29975 3720
rect 29880 3680 29886 3692
rect 29963 3689 29975 3692
rect 30009 3689 30021 3723
rect 30466 3720 30472 3732
rect 30427 3692 30472 3720
rect 29963 3683 30021 3689
rect 30466 3680 30472 3692
rect 30524 3720 30530 3732
rect 30975 3723 31033 3729
rect 30975 3720 30987 3723
rect 30524 3692 30987 3720
rect 30524 3680 30530 3692
rect 30975 3689 30987 3692
rect 31021 3689 31033 3723
rect 30975 3683 31033 3689
rect 17218 3652 17224 3664
rect 16172 3624 17080 3652
rect 17179 3624 17224 3652
rect 16172 3612 16178 3624
rect 17218 3612 17224 3624
rect 17276 3612 17282 3664
rect 19334 3612 19340 3664
rect 19392 3652 19398 3664
rect 19429 3655 19487 3661
rect 19429 3652 19441 3655
rect 19392 3624 19441 3652
rect 19392 3612 19398 3624
rect 19429 3621 19441 3624
rect 19475 3621 19487 3655
rect 19978 3652 19984 3664
rect 19939 3624 19984 3652
rect 19429 3615 19487 3621
rect 19978 3612 19984 3624
rect 20036 3612 20042 3664
rect 21913 3655 21971 3661
rect 21913 3621 21925 3655
rect 21959 3652 21971 3655
rect 22002 3652 22008 3664
rect 21959 3624 22008 3652
rect 21959 3621 21971 3624
rect 21913 3615 21971 3621
rect 22002 3612 22008 3624
rect 22060 3612 22066 3664
rect 25590 3612 25596 3664
rect 25648 3652 25654 3664
rect 25685 3655 25743 3661
rect 25685 3652 25697 3655
rect 25648 3624 25697 3652
rect 25648 3612 25654 3624
rect 25685 3621 25697 3624
rect 25731 3621 25743 3655
rect 25685 3615 25743 3621
rect 26602 3612 26608 3664
rect 26660 3652 26666 3664
rect 26834 3655 26892 3661
rect 26834 3652 26846 3655
rect 26660 3624 26846 3652
rect 26660 3612 26666 3624
rect 26834 3621 26846 3624
rect 26880 3621 26892 3655
rect 28166 3652 28172 3664
rect 26834 3615 26892 3621
rect 27448 3624 28172 3652
rect 4614 3593 4620 3596
rect 4592 3587 4620 3593
rect 4592 3553 4604 3587
rect 4592 3547 4620 3553
rect 4614 3544 4620 3547
rect 4672 3544 4678 3596
rect 5537 3587 5595 3593
rect 5537 3553 5549 3587
rect 5583 3584 5595 3587
rect 5626 3584 5632 3596
rect 5583 3556 5632 3584
rect 5583 3553 5595 3556
rect 5537 3547 5595 3553
rect 5626 3544 5632 3556
rect 5684 3544 5690 3596
rect 9490 3544 9496 3596
rect 9548 3584 9554 3596
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9548 3556 9689 3584
rect 9548 3544 9554 3556
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 9677 3547 9735 3553
rect 10873 3587 10931 3593
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11606 3584 11612 3596
rect 10919 3556 11612 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12492 3556 12537 3584
rect 12492 3544 12498 3556
rect 14182 3544 14188 3596
rect 14240 3593 14246 3596
rect 14240 3587 14278 3593
rect 14266 3553 14278 3587
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 14240 3547 14278 3553
rect 14240 3544 14246 3547
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 23290 3544 23296 3596
rect 23348 3593 23354 3596
rect 23348 3587 23386 3593
rect 23374 3584 23386 3587
rect 24670 3584 24676 3596
rect 23374 3556 24676 3584
rect 23374 3553 23386 3556
rect 23348 3547 23386 3553
rect 23348 3544 23354 3547
rect 24670 3544 24676 3556
rect 24728 3544 24734 3596
rect 25866 3544 25872 3596
rect 25924 3584 25930 3596
rect 27448 3593 27476 3624
rect 28166 3612 28172 3624
rect 28224 3652 28230 3664
rect 28445 3655 28503 3661
rect 28445 3652 28457 3655
rect 28224 3624 28457 3652
rect 28224 3612 28230 3624
rect 28445 3621 28457 3624
rect 28491 3652 28503 3655
rect 28994 3652 29000 3664
rect 28491 3624 29000 3652
rect 28491 3621 28503 3624
rect 28445 3615 28503 3621
rect 28994 3612 29000 3624
rect 29052 3612 29058 3664
rect 26053 3587 26111 3593
rect 26053 3584 26065 3587
rect 25924 3556 26065 3584
rect 25924 3544 25930 3556
rect 26053 3553 26065 3556
rect 26099 3553 26111 3587
rect 26053 3547 26111 3553
rect 27433 3587 27491 3593
rect 27433 3553 27445 3587
rect 27479 3553 27491 3587
rect 27433 3547 27491 3553
rect 29730 3544 29736 3596
rect 29788 3584 29794 3596
rect 29860 3587 29918 3593
rect 29860 3584 29872 3587
rect 29788 3556 29872 3584
rect 29788 3544 29794 3556
rect 29860 3553 29872 3556
rect 29906 3553 29918 3587
rect 29860 3547 29918 3553
rect 30904 3587 30962 3593
rect 30904 3553 30916 3587
rect 30950 3584 30962 3587
rect 31110 3584 31116 3596
rect 30950 3556 31116 3584
rect 30950 3553 30962 3556
rect 30904 3547 30962 3553
rect 31110 3544 31116 3556
rect 31168 3544 31174 3596
rect 2225 3519 2283 3525
rect 2225 3485 2237 3519
rect 2271 3516 2283 3519
rect 2314 3516 2320 3528
rect 2271 3488 2320 3516
rect 2271 3485 2283 3488
rect 2225 3479 2283 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 8018 3516 8024 3528
rect 7931 3488 8024 3516
rect 7377 3479 7435 3485
rect 2682 3408 2688 3460
rect 2740 3448 2746 3460
rect 3418 3448 3424 3460
rect 2740 3420 3424 3448
rect 2740 3408 2746 3420
rect 3418 3408 3424 3420
rect 3476 3408 3482 3460
rect 7392 3448 7420 3479
rect 8018 3476 8024 3488
rect 8076 3516 8082 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8076 3488 8309 3516
rect 8076 3476 8082 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 13357 3519 13415 3525
rect 13357 3485 13369 3519
rect 13403 3516 13415 3519
rect 14090 3516 14096 3528
rect 13403 3488 14096 3516
rect 13403 3485 13415 3488
rect 13357 3479 13415 3485
rect 8386 3448 8392 3460
rect 7392 3420 8392 3448
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 9214 3408 9220 3460
rect 9272 3448 9278 3460
rect 9861 3451 9919 3457
rect 9861 3448 9873 3451
rect 9272 3420 9873 3448
rect 9272 3408 9278 3420
rect 9861 3417 9873 3420
rect 9907 3417 9919 3451
rect 12250 3448 12256 3460
rect 9861 3411 9919 3417
rect 11808 3420 12256 3448
rect 4154 3340 4160 3392
rect 4212 3380 4218 3392
rect 4663 3383 4721 3389
rect 4663 3380 4675 3383
rect 4212 3352 4675 3380
rect 4212 3340 4218 3352
rect 4663 3349 4675 3352
rect 4709 3349 4721 3383
rect 6454 3380 6460 3392
rect 6415 3352 6460 3380
rect 4663 3343 4721 3349
rect 6454 3340 6460 3352
rect 6512 3340 6518 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11808 3389 11836 3420
rect 12250 3408 12256 3420
rect 12308 3408 12314 3460
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13372 3448 13400 3479
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17402 3516 17408 3528
rect 17363 3488 17408 3516
rect 17129 3479 17187 3485
rect 12492 3420 13400 3448
rect 14323 3451 14381 3457
rect 12492 3408 12498 3420
rect 14323 3417 14335 3451
rect 14369 3448 14381 3451
rect 17144 3448 17172 3479
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 18656 3488 19349 3516
rect 18656 3476 18662 3488
rect 19337 3485 19349 3488
rect 19383 3516 19395 3519
rect 20622 3516 20628 3528
rect 19383 3488 20628 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 21821 3519 21879 3525
rect 21821 3485 21833 3519
rect 21867 3516 21879 3519
rect 22094 3516 22100 3528
rect 21867 3488 22100 3516
rect 21867 3485 21879 3488
rect 21821 3479 21879 3485
rect 22094 3476 22100 3488
rect 22152 3516 22158 3528
rect 23431 3519 23489 3525
rect 23431 3516 23443 3519
rect 22152 3488 23443 3516
rect 22152 3476 22158 3488
rect 23431 3485 23443 3488
rect 23477 3485 23489 3519
rect 23431 3479 23489 3485
rect 26234 3476 26240 3528
rect 26292 3516 26298 3528
rect 26510 3516 26516 3528
rect 26292 3488 26516 3516
rect 26292 3476 26298 3488
rect 26510 3476 26516 3488
rect 26568 3476 26574 3528
rect 27982 3476 27988 3528
rect 28040 3516 28046 3528
rect 28353 3519 28411 3525
rect 28353 3516 28365 3519
rect 28040 3488 28365 3516
rect 28040 3476 28046 3488
rect 28353 3485 28365 3488
rect 28399 3485 28411 3519
rect 28353 3479 28411 3485
rect 17770 3448 17776 3460
rect 14369 3420 17776 3448
rect 14369 3417 14381 3420
rect 14323 3411 14381 3417
rect 17770 3408 17776 3420
rect 17828 3408 17834 3460
rect 22370 3448 22376 3460
rect 22331 3420 22376 3448
rect 22370 3408 22376 3420
rect 22428 3408 22434 3460
rect 28902 3448 28908 3460
rect 28863 3420 28908 3448
rect 28902 3408 28908 3420
rect 28960 3408 28966 3460
rect 11793 3383 11851 3389
rect 11793 3380 11805 3383
rect 11204 3352 11805 3380
rect 11204 3340 11210 3352
rect 11793 3349 11805 3352
rect 11839 3349 11851 3383
rect 13998 3380 14004 3392
rect 13959 3352 14004 3380
rect 11793 3343 11851 3349
rect 13998 3340 14004 3352
rect 14056 3340 14062 3392
rect 15010 3380 15016 3392
rect 14971 3352 15016 3380
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 15194 3340 15200 3392
rect 15252 3380 15258 3392
rect 16209 3383 16267 3389
rect 16209 3380 16221 3383
rect 15252 3352 16221 3380
rect 15252 3340 15258 3352
rect 16209 3349 16221 3352
rect 16255 3349 16267 3383
rect 16209 3343 16267 3349
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 20257 3383 20315 3389
rect 20257 3380 20269 3383
rect 19852 3352 20269 3380
rect 19852 3340 19858 3352
rect 20257 3349 20269 3352
rect 20303 3349 20315 3383
rect 20257 3343 20315 3349
rect 27798 3340 27804 3392
rect 27856 3380 27862 3392
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 27856 3352 28089 3380
rect 27856 3340 27862 3352
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 29546 3380 29552 3392
rect 29507 3352 29552 3380
rect 28077 3343 28135 3349
rect 29546 3340 29552 3352
rect 29604 3340 29610 3392
rect 1104 3290 38824 3312
rect 1104 3238 7648 3290
rect 7700 3238 7712 3290
rect 7764 3238 7776 3290
rect 7828 3238 7840 3290
rect 7892 3238 20982 3290
rect 21034 3238 21046 3290
rect 21098 3238 21110 3290
rect 21162 3238 21174 3290
rect 21226 3238 34315 3290
rect 34367 3238 34379 3290
rect 34431 3238 34443 3290
rect 34495 3238 34507 3290
rect 34559 3238 38824 3290
rect 1104 3216 38824 3238
rect 2866 3176 2872 3188
rect 2827 3148 2872 3176
rect 2866 3136 2872 3148
rect 2924 3136 2930 3188
rect 4246 3136 4252 3188
rect 4304 3176 4310 3188
rect 4709 3179 4767 3185
rect 4709 3176 4721 3179
rect 4304 3148 4721 3176
rect 4304 3136 4310 3148
rect 4709 3145 4721 3148
rect 4755 3176 4767 3179
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4755 3148 4905 3176
rect 4755 3145 4767 3148
rect 4709 3139 4767 3145
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5960 3148 6193 3176
rect 5960 3136 5966 3148
rect 6181 3145 6193 3148
rect 6227 3145 6239 3179
rect 6181 3139 6239 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8386 3176 8392 3188
rect 8343 3148 8392 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8386 3136 8392 3148
rect 8444 3136 8450 3188
rect 10778 3136 10784 3188
rect 10836 3176 10842 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10836 3148 10885 3176
rect 10836 3136 10842 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 11606 3136 11612 3188
rect 11664 3176 11670 3188
rect 12069 3179 12127 3185
rect 12069 3176 12081 3179
rect 11664 3148 12081 3176
rect 11664 3136 11670 3148
rect 12069 3145 12081 3148
rect 12115 3145 12127 3179
rect 13354 3176 13360 3188
rect 13315 3148 13360 3176
rect 12069 3139 12127 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14461 3179 14519 3185
rect 14461 3176 14473 3179
rect 14240 3148 14473 3176
rect 14240 3136 14246 3148
rect 14461 3145 14473 3148
rect 14507 3176 14519 3179
rect 14918 3176 14924 3188
rect 14507 3148 14924 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15286 3136 15292 3188
rect 15344 3176 15350 3188
rect 16393 3179 16451 3185
rect 16393 3176 16405 3179
rect 15344 3148 16405 3176
rect 15344 3136 15350 3148
rect 16393 3145 16405 3148
rect 16439 3145 16451 3179
rect 16393 3139 16451 3145
rect 17218 3136 17224 3188
rect 17276 3176 17282 3188
rect 17405 3179 17463 3185
rect 17405 3176 17417 3179
rect 17276 3148 17417 3176
rect 17276 3136 17282 3148
rect 17405 3145 17417 3148
rect 17451 3145 17463 3179
rect 17770 3176 17776 3188
rect 17731 3148 17776 3176
rect 17405 3139 17463 3145
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18598 3176 18604 3188
rect 18559 3148 18604 3176
rect 18598 3136 18604 3148
rect 18656 3136 18662 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19521 3179 19579 3185
rect 19521 3176 19533 3179
rect 19392 3148 19533 3176
rect 19392 3136 19398 3148
rect 19521 3145 19533 3148
rect 19567 3145 19579 3179
rect 19521 3139 19579 3145
rect 22002 3136 22008 3188
rect 22060 3176 22066 3188
rect 22281 3179 22339 3185
rect 22281 3176 22293 3179
rect 22060 3148 22293 3176
rect 22060 3136 22066 3148
rect 22281 3145 22293 3148
rect 22327 3145 22339 3179
rect 22281 3139 22339 3145
rect 26510 3136 26516 3188
rect 26568 3176 26574 3188
rect 26881 3179 26939 3185
rect 26881 3176 26893 3179
rect 26568 3148 26893 3176
rect 26568 3136 26574 3148
rect 26881 3145 26893 3148
rect 26927 3145 26939 3179
rect 26881 3139 26939 3145
rect 27203 3179 27261 3185
rect 27203 3145 27215 3179
rect 27249 3176 27261 3179
rect 27522 3176 27528 3188
rect 27249 3148 27528 3176
rect 27249 3145 27261 3148
rect 27203 3139 27261 3145
rect 27522 3136 27528 3148
rect 27580 3176 27586 3188
rect 27798 3176 27804 3188
rect 27580 3148 27804 3176
rect 27580 3136 27586 3148
rect 27798 3136 27804 3148
rect 27856 3136 27862 3188
rect 27982 3176 27988 3188
rect 27943 3148 27988 3176
rect 27982 3136 27988 3148
rect 28040 3136 28046 3188
rect 28994 3176 29000 3188
rect 28955 3148 29000 3176
rect 28994 3136 29000 3148
rect 29052 3136 29058 3188
rect 29822 3136 29828 3188
rect 29880 3176 29886 3188
rect 30101 3179 30159 3185
rect 30101 3176 30113 3179
rect 29880 3148 30113 3176
rect 29880 3136 29886 3148
rect 30101 3145 30113 3148
rect 30147 3145 30159 3179
rect 30101 3139 30159 3145
rect 30929 3179 30987 3185
rect 30929 3145 30941 3179
rect 30975 3176 30987 3179
rect 31110 3176 31116 3188
rect 30975 3148 31116 3176
rect 30975 3145 30987 3148
rect 30929 3139 30987 3145
rect 31110 3136 31116 3148
rect 31168 3136 31174 3188
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 4614 3108 4620 3120
rect 4120 3080 4620 3108
rect 4120 3068 4126 3080
rect 4614 3068 4620 3080
rect 4672 3108 4678 3120
rect 5813 3111 5871 3117
rect 5813 3108 5825 3111
rect 4672 3080 5825 3108
rect 4672 3068 4678 3080
rect 5813 3077 5825 3080
rect 5859 3108 5871 3111
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 5859 3080 7481 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 13630 3068 13636 3120
rect 13688 3108 13694 3120
rect 14093 3111 14151 3117
rect 14093 3108 14105 3111
rect 13688 3080 14105 3108
rect 13688 3068 13694 3080
rect 14093 3077 14105 3080
rect 14139 3108 14151 3111
rect 15010 3108 15016 3120
rect 14139 3080 15016 3108
rect 14139 3077 14151 3080
rect 14093 3071 14151 3077
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 16114 3108 16120 3120
rect 16075 3080 16120 3108
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 18831 3111 18889 3117
rect 18831 3077 18843 3111
rect 18877 3108 18889 3111
rect 21910 3108 21916 3120
rect 18877 3080 19840 3108
rect 21871 3080 21916 3108
rect 18877 3077 18889 3080
rect 18831 3071 18889 3077
rect 19812 3052 19840 3080
rect 21910 3068 21916 3080
rect 21968 3068 21974 3120
rect 26602 3108 26608 3120
rect 26563 3080 26608 3108
rect 26602 3068 26608 3080
rect 26660 3068 26666 3120
rect 29730 3108 29736 3120
rect 29691 3080 29736 3108
rect 29730 3068 29736 3080
rect 29788 3068 29794 3120
rect 1670 3000 1676 3052
rect 1728 3040 1734 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 1728 3012 2237 3040
rect 1728 3000 1734 3012
rect 2225 3009 2237 3012
rect 2271 3040 2283 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 2271 3012 2513 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 6454 3040 6460 3052
rect 2501 3003 2559 3009
rect 3712 3012 6460 3040
rect 3712 2981 3740 3012
rect 6454 3000 6460 3012
rect 6512 3040 6518 3052
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 6512 3012 6561 3040
rect 6512 3000 6518 3012
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 8018 3040 8024 3052
rect 6963 3012 8024 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2941 2099 2975
rect 2041 2935 2099 2941
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3559 2944 3709 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 4939 2944 5120 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 2056 2904 2084 2935
rect 2866 2904 2872 2916
rect 2056 2876 2872 2904
rect 2866 2864 2872 2876
rect 2924 2864 2930 2916
rect 4341 2907 4399 2913
rect 4341 2873 4353 2907
rect 4387 2904 4399 2907
rect 4985 2907 5043 2913
rect 4985 2904 4997 2907
rect 4387 2876 4997 2904
rect 4387 2873 4399 2876
rect 4341 2867 4399 2873
rect 4985 2873 4997 2876
rect 5031 2873 5043 2907
rect 5092 2904 5120 2944
rect 5261 2907 5319 2913
rect 5261 2904 5273 2907
rect 5092 2876 5273 2904
rect 4985 2867 5043 2873
rect 5261 2873 5273 2876
rect 5307 2873 5319 2907
rect 5261 2867 5319 2873
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2873 5411 2907
rect 6564 2904 6592 3003
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 9674 3040 9680 3052
rect 9635 3012 9680 3040
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 11790 3040 11796 3052
rect 11164 3012 11796 3040
rect 8389 2975 8447 2981
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 8938 2972 8944 2984
rect 8435 2944 8944 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9490 2972 9496 2984
rect 9451 2944 9496 2972
rect 9490 2932 9496 2944
rect 9548 2932 9554 2984
rect 11164 2981 11192 3012
rect 11790 3000 11796 3012
rect 11848 3000 11854 3052
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3040 13599 3043
rect 13998 3040 14004 3052
rect 13587 3012 14004 3040
rect 13587 3009 13599 3012
rect 13541 3003 13599 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 19794 3040 19800 3052
rect 19755 3012 19800 3040
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 20254 3040 20260 3052
rect 20215 3012 20260 3040
rect 20254 3000 20260 3012
rect 20312 3040 20318 3052
rect 21361 3043 21419 3049
rect 21361 3040 21373 3043
rect 20312 3012 21373 3040
rect 20312 3000 20318 3012
rect 21361 3009 21373 3012
rect 21407 3040 21419 3043
rect 22370 3040 22376 3052
rect 21407 3012 22376 3040
rect 21407 3009 21419 3012
rect 21361 3003 21419 3009
rect 22370 3000 22376 3012
rect 22428 3040 22434 3052
rect 22649 3043 22707 3049
rect 22649 3040 22661 3043
rect 22428 3012 22661 3040
rect 22428 3000 22434 3012
rect 22649 3009 22661 3012
rect 22695 3009 22707 3043
rect 22649 3003 22707 3009
rect 16666 2981 16672 2984
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 12504 2975 12562 2981
rect 12504 2941 12516 2975
rect 12550 2972 12562 2975
rect 16644 2975 16672 2981
rect 16644 2972 16656 2975
rect 12550 2944 13032 2972
rect 16579 2944 16656 2972
rect 12550 2941 12562 2944
rect 12504 2935 12562 2941
rect 7009 2907 7067 2913
rect 7009 2904 7021 2907
rect 6564 2876 7021 2904
rect 5353 2867 5411 2873
rect 7009 2873 7021 2876
rect 7055 2873 7067 2907
rect 9766 2904 9772 2916
rect 9727 2876 9772 2904
rect 7009 2867 7067 2873
rect 5000 2836 5028 2867
rect 5368 2836 5396 2867
rect 9766 2864 9772 2876
rect 9824 2864 9830 2916
rect 13004 2913 13032 2944
rect 16644 2941 16656 2944
rect 16724 2972 16730 2984
rect 17037 2975 17095 2981
rect 17037 2972 17049 2975
rect 16724 2944 17049 2972
rect 16644 2935 16672 2941
rect 16666 2932 16672 2935
rect 16724 2932 16730 2944
rect 17037 2941 17049 2944
rect 17083 2941 17095 2975
rect 17037 2935 17095 2941
rect 18760 2975 18818 2981
rect 18760 2941 18772 2975
rect 18806 2972 18818 2975
rect 23290 2972 23296 2984
rect 18806 2944 19196 2972
rect 23251 2944 23296 2972
rect 18806 2941 18818 2944
rect 18760 2935 18818 2941
rect 12989 2907 13047 2913
rect 12989 2873 13001 2907
rect 13035 2904 13047 2907
rect 13538 2904 13544 2916
rect 13035 2876 13544 2904
rect 13035 2873 13047 2876
rect 12989 2867 13047 2873
rect 13538 2864 13544 2876
rect 13596 2864 13602 2916
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13722 2904 13728 2916
rect 13679 2876 13728 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13722 2864 13728 2876
rect 13780 2864 13786 2916
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 15252 2876 15297 2904
rect 15252 2864 15258 2876
rect 5000 2808 5396 2836
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7466 2836 7472 2848
rect 7156 2808 7472 2836
rect 7156 2796 7162 2808
rect 7466 2796 7472 2808
rect 7524 2836 7530 2848
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 7524 2808 7849 2836
rect 7524 2796 7530 2808
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 7837 2799 7895 2805
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8573 2839 8631 2845
rect 8573 2836 8585 2839
rect 8352 2808 8585 2836
rect 8352 2796 8358 2808
rect 8573 2805 8585 2808
rect 8619 2805 8631 2839
rect 8573 2799 8631 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11333 2839 11391 2845
rect 11333 2836 11345 2839
rect 11112 2808 11345 2836
rect 11112 2796 11118 2808
rect 11333 2805 11345 2808
rect 11379 2805 11391 2839
rect 11333 2799 11391 2805
rect 12575 2839 12633 2845
rect 12575 2805 12587 2839
rect 12621 2836 12633 2839
rect 12710 2836 12716 2848
rect 12621 2808 12716 2836
rect 12621 2805 12633 2808
rect 12575 2799 12633 2805
rect 12710 2796 12716 2808
rect 12768 2796 12774 2848
rect 14921 2839 14979 2845
rect 14921 2805 14933 2839
rect 14967 2836 14979 2839
rect 15212 2836 15240 2864
rect 19168 2848 19196 2944
rect 23290 2932 23296 2944
rect 23348 2932 23354 2984
rect 27062 2932 27068 2984
rect 27120 2981 27126 2984
rect 27120 2975 27158 2981
rect 27146 2972 27158 2975
rect 27525 2975 27583 2981
rect 27525 2972 27537 2975
rect 27146 2944 27537 2972
rect 27146 2941 27158 2944
rect 27120 2935 27158 2941
rect 27525 2941 27537 2944
rect 27571 2941 27583 2975
rect 28074 2972 28080 2984
rect 28035 2944 28080 2972
rect 27525 2935 27583 2941
rect 27120 2932 27126 2935
rect 28074 2932 28080 2944
rect 28132 2972 28138 2984
rect 28629 2975 28687 2981
rect 28629 2972 28641 2975
rect 28132 2944 28641 2972
rect 28132 2932 28138 2944
rect 28629 2941 28641 2944
rect 28675 2941 28687 2975
rect 29546 2972 29552 2984
rect 29507 2944 29552 2972
rect 28629 2935 28687 2941
rect 29546 2932 29552 2944
rect 29604 2932 29610 2984
rect 19334 2864 19340 2916
rect 19392 2904 19398 2916
rect 19889 2907 19947 2913
rect 19889 2904 19901 2907
rect 19392 2876 19901 2904
rect 19392 2864 19398 2876
rect 19889 2873 19901 2876
rect 19935 2904 19947 2907
rect 20717 2907 20775 2913
rect 20717 2904 20729 2907
rect 19935 2876 20729 2904
rect 19935 2873 19947 2876
rect 19889 2867 19947 2873
rect 20717 2873 20729 2876
rect 20763 2873 20775 2907
rect 20717 2867 20775 2873
rect 21453 2907 21511 2913
rect 21453 2873 21465 2907
rect 21499 2904 21511 2907
rect 21818 2904 21824 2916
rect 21499 2876 21824 2904
rect 21499 2873 21511 2876
rect 21453 2867 21511 2873
rect 14967 2808 15240 2836
rect 14967 2805 14979 2808
rect 14921 2799 14979 2805
rect 16574 2796 16580 2848
rect 16632 2836 16638 2848
rect 16715 2839 16773 2845
rect 16715 2836 16727 2839
rect 16632 2808 16727 2836
rect 16632 2796 16638 2808
rect 16715 2805 16727 2808
rect 16761 2805 16773 2839
rect 19150 2836 19156 2848
rect 19111 2808 19156 2836
rect 16715 2799 16773 2805
rect 19150 2796 19156 2808
rect 19208 2796 19214 2848
rect 21177 2839 21235 2845
rect 21177 2805 21189 2839
rect 21223 2836 21235 2839
rect 21468 2836 21496 2867
rect 21818 2864 21824 2876
rect 21876 2864 21882 2916
rect 28258 2836 28264 2848
rect 21223 2808 21496 2836
rect 28219 2808 28264 2836
rect 21223 2805 21235 2808
rect 21177 2799 21235 2805
rect 28258 2796 28264 2808
rect 28316 2796 28322 2848
rect 1104 2746 38824 2768
rect 1104 2694 14315 2746
rect 14367 2694 14379 2746
rect 14431 2694 14443 2746
rect 14495 2694 14507 2746
rect 14559 2694 27648 2746
rect 27700 2694 27712 2746
rect 27764 2694 27776 2746
rect 27828 2694 27840 2746
rect 27892 2694 38824 2746
rect 1104 2672 38824 2694
rect 1486 2592 1492 2644
rect 1544 2592 1550 2644
rect 1627 2635 1685 2641
rect 1627 2601 1639 2635
rect 1673 2632 1685 2635
rect 2682 2632 2688 2644
rect 1673 2604 2688 2632
rect 1673 2601 1685 2604
rect 1627 2595 1685 2601
rect 2682 2592 2688 2604
rect 2740 2592 2746 2644
rect 3050 2632 3056 2644
rect 3011 2604 3056 2632
rect 3050 2592 3056 2604
rect 3108 2592 3114 2644
rect 3881 2635 3939 2641
rect 3881 2601 3893 2635
rect 3927 2632 3939 2635
rect 4062 2632 4068 2644
rect 3927 2604 4068 2632
rect 3927 2601 3939 2604
rect 3881 2595 3939 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4338 2632 4344 2644
rect 4299 2604 4344 2632
rect 4338 2592 4344 2604
rect 4396 2592 4402 2644
rect 5626 2592 5632 2644
rect 5684 2632 5690 2644
rect 6273 2635 6331 2641
rect 6273 2632 6285 2635
rect 5684 2604 6285 2632
rect 5684 2592 5690 2604
rect 6273 2601 6285 2604
rect 6319 2601 6331 2635
rect 7098 2632 7104 2644
rect 6273 2595 6331 2601
rect 6380 2604 7104 2632
rect 1504 2564 1532 2592
rect 2317 2567 2375 2573
rect 2317 2564 2329 2567
rect 1504 2536 2329 2564
rect 2317 2533 2329 2536
rect 2363 2533 2375 2567
rect 2317 2527 2375 2533
rect 1556 2499 1614 2505
rect 1556 2465 1568 2499
rect 1602 2496 1614 2499
rect 2038 2496 2044 2508
rect 1602 2468 2044 2496
rect 1602 2465 1614 2468
rect 1556 2459 1614 2465
rect 2038 2456 2044 2468
rect 2096 2456 2102 2508
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2465 2927 2499
rect 2869 2459 2927 2465
rect 4157 2499 4215 2505
rect 4157 2465 4169 2499
rect 4203 2496 4215 2499
rect 4798 2496 4804 2508
rect 4203 2468 4804 2496
rect 4203 2465 4215 2468
rect 4157 2459 4215 2465
rect 2884 2428 2912 2459
rect 4798 2456 4804 2468
rect 4856 2456 4862 2508
rect 5169 2499 5227 2505
rect 5169 2465 5181 2499
rect 5215 2496 5227 2499
rect 5905 2499 5963 2505
rect 5905 2496 5917 2499
rect 5215 2468 5917 2496
rect 5215 2465 5227 2468
rect 5169 2459 5227 2465
rect 5905 2465 5917 2468
rect 5951 2496 5963 2499
rect 6380 2496 6408 2604
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 9582 2632 9588 2644
rect 9543 2604 9588 2632
rect 9582 2592 9588 2604
rect 9640 2592 9646 2644
rect 13722 2632 13728 2644
rect 13683 2604 13728 2632
rect 13722 2592 13728 2604
rect 13780 2592 13786 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14323 2635 14381 2641
rect 14323 2632 14335 2635
rect 14056 2604 14335 2632
rect 14056 2592 14062 2604
rect 14323 2601 14335 2604
rect 14369 2601 14381 2635
rect 15102 2632 15108 2644
rect 15063 2604 15108 2632
rect 14323 2595 14381 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 19426 2632 19432 2644
rect 19387 2604 19432 2632
rect 19426 2592 19432 2604
rect 19484 2632 19490 2644
rect 19484 2604 19748 2632
rect 19484 2592 19490 2604
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 5951 2468 6408 2496
rect 6656 2536 7389 2564
rect 5951 2465 5963 2468
rect 5905 2459 5963 2465
rect 3510 2428 3516 2440
rect 2884 2400 3516 2428
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 6656 2437 6684 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 7929 2567 7987 2573
rect 7929 2533 7941 2567
rect 7975 2564 7987 2567
rect 8018 2564 8024 2576
rect 7975 2536 8024 2564
rect 7975 2533 7987 2536
rect 7929 2527 7987 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 10873 2567 10931 2573
rect 10873 2533 10885 2567
rect 10919 2564 10931 2567
rect 11146 2564 11152 2576
rect 10919 2536 11152 2564
rect 10919 2533 10931 2536
rect 10873 2527 10931 2533
rect 11146 2524 11152 2536
rect 11204 2524 11210 2576
rect 11701 2567 11759 2573
rect 11701 2533 11713 2567
rect 11747 2564 11759 2567
rect 12342 2564 12348 2576
rect 11747 2536 12348 2564
rect 11747 2533 11759 2536
rect 11701 2527 11759 2533
rect 12342 2524 12348 2536
rect 12400 2524 12406 2576
rect 12437 2567 12495 2573
rect 12437 2533 12449 2567
rect 12483 2564 12495 2567
rect 12805 2567 12863 2573
rect 12805 2564 12817 2567
rect 12483 2536 12817 2564
rect 12483 2533 12495 2536
rect 12437 2527 12495 2533
rect 12805 2533 12817 2536
rect 12851 2564 12863 2567
rect 13170 2564 13176 2576
rect 12851 2536 13176 2564
rect 12851 2533 12863 2536
rect 12805 2527 12863 2533
rect 13170 2524 13176 2536
rect 13228 2524 13234 2576
rect 13357 2567 13415 2573
rect 13357 2533 13369 2567
rect 13403 2564 13415 2567
rect 13630 2564 13636 2576
rect 13403 2536 13636 2564
rect 13403 2533 13415 2536
rect 13357 2527 13415 2533
rect 13630 2524 13636 2536
rect 13688 2524 13694 2576
rect 13906 2524 13912 2576
rect 13964 2564 13970 2576
rect 14645 2567 14703 2573
rect 14645 2564 14657 2567
rect 13964 2536 14657 2564
rect 13964 2524 13970 2536
rect 9769 2499 9827 2505
rect 9769 2465 9781 2499
rect 9815 2496 9827 2499
rect 10410 2496 10416 2508
rect 9815 2468 10416 2496
rect 9815 2465 9827 2468
rect 9769 2459 9827 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 14292 2505 14320 2536
rect 14645 2533 14657 2536
rect 14691 2564 14703 2567
rect 14734 2564 14740 2576
rect 14691 2536 14740 2564
rect 14691 2533 14703 2536
rect 14645 2527 14703 2533
rect 14734 2524 14740 2536
rect 14792 2524 14798 2576
rect 19061 2567 19119 2573
rect 19061 2533 19073 2567
rect 19107 2564 19119 2567
rect 19610 2564 19616 2576
rect 19107 2536 19616 2564
rect 19107 2533 19119 2536
rect 19061 2527 19119 2533
rect 19610 2524 19616 2536
rect 19668 2524 19674 2576
rect 19720 2573 19748 2604
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 21315 2635 21373 2641
rect 21315 2632 21327 2635
rect 20772 2604 21327 2632
rect 20772 2592 20778 2604
rect 21315 2601 21327 2604
rect 21361 2601 21373 2635
rect 21315 2595 21373 2601
rect 22094 2592 22100 2644
rect 22152 2632 22158 2644
rect 22327 2635 22385 2641
rect 22152 2604 22197 2632
rect 22152 2592 22158 2604
rect 22327 2601 22339 2635
rect 22373 2632 22385 2635
rect 23382 2632 23388 2644
rect 22373 2604 23388 2632
rect 22373 2601 22385 2604
rect 22327 2595 22385 2601
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 27663 2635 27721 2641
rect 27663 2601 27675 2635
rect 27709 2632 27721 2635
rect 27982 2632 27988 2644
rect 27709 2604 27988 2632
rect 27709 2601 27721 2604
rect 27663 2595 27721 2601
rect 27982 2592 27988 2604
rect 28040 2592 28046 2644
rect 28718 2632 28724 2644
rect 28679 2604 28724 2632
rect 28718 2592 28724 2604
rect 28776 2592 28782 2644
rect 31570 2632 31576 2644
rect 31531 2604 31576 2632
rect 31570 2592 31576 2604
rect 31628 2592 31634 2644
rect 32766 2632 32772 2644
rect 32727 2604 32772 2632
rect 32766 2592 32772 2604
rect 32824 2592 32830 2644
rect 19705 2567 19763 2573
rect 19705 2533 19717 2567
rect 19751 2533 19763 2567
rect 20254 2564 20260 2576
rect 20215 2536 20260 2564
rect 19705 2527 19763 2533
rect 20254 2524 20260 2536
rect 20312 2524 20318 2576
rect 14252 2499 14320 2505
rect 14252 2465 14264 2499
rect 14298 2468 14320 2499
rect 14298 2465 14310 2468
rect 14252 2459 14310 2465
rect 15470 2456 15476 2508
rect 15528 2505 15534 2508
rect 15528 2499 15566 2505
rect 15554 2496 15566 2499
rect 15933 2499 15991 2505
rect 15933 2496 15945 2499
rect 15554 2468 15945 2496
rect 15554 2465 15566 2468
rect 15528 2459 15566 2465
rect 15933 2465 15945 2468
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 15528 2456 15534 2459
rect 20806 2456 20812 2508
rect 20864 2496 20870 2508
rect 21244 2499 21302 2505
rect 21244 2496 21256 2499
rect 20864 2468 21256 2496
rect 20864 2456 20870 2468
rect 21244 2465 21256 2468
rect 21290 2496 21302 2499
rect 21726 2496 21732 2508
rect 21290 2468 21732 2496
rect 21290 2465 21302 2468
rect 21244 2459 21302 2465
rect 21726 2456 21732 2468
rect 21784 2456 21790 2508
rect 22256 2499 22314 2505
rect 22256 2465 22268 2499
rect 22302 2496 22314 2499
rect 22741 2499 22799 2505
rect 22741 2496 22753 2499
rect 22302 2468 22753 2496
rect 22302 2465 22314 2468
rect 22256 2459 22314 2465
rect 22741 2465 22753 2468
rect 22787 2496 22799 2499
rect 23290 2496 23296 2508
rect 22787 2468 23296 2496
rect 22787 2465 22799 2468
rect 22741 2459 22799 2465
rect 23290 2456 23296 2468
rect 23348 2456 23354 2508
rect 27614 2505 27620 2508
rect 27592 2499 27620 2505
rect 27592 2465 27604 2499
rect 27672 2496 27678 2508
rect 27985 2499 28043 2505
rect 27985 2496 27997 2499
rect 27672 2468 27997 2496
rect 27592 2459 27620 2465
rect 27614 2456 27620 2459
rect 27672 2456 27678 2468
rect 27985 2465 27997 2468
rect 28031 2465 28043 2499
rect 28534 2496 28540 2508
rect 28495 2468 28540 2496
rect 27985 2459 28043 2465
rect 28534 2456 28540 2468
rect 28592 2496 28598 2508
rect 29089 2499 29147 2505
rect 29089 2496 29101 2499
rect 28592 2468 29101 2496
rect 28592 2456 28598 2468
rect 29089 2465 29101 2468
rect 29135 2465 29147 2499
rect 30282 2496 30288 2508
rect 30243 2468 30288 2496
rect 29089 2459 29147 2465
rect 30282 2456 30288 2468
rect 30340 2496 30346 2508
rect 30837 2499 30895 2505
rect 30837 2496 30849 2499
rect 30340 2468 30849 2496
rect 30340 2456 30346 2468
rect 30837 2465 30849 2468
rect 30883 2465 30895 2499
rect 31386 2496 31392 2508
rect 31347 2468 31392 2496
rect 30837 2459 30895 2465
rect 31386 2456 31392 2468
rect 31444 2496 31450 2508
rect 31941 2499 31999 2505
rect 31941 2496 31953 2499
rect 31444 2468 31953 2496
rect 31444 2456 31450 2468
rect 31941 2465 31953 2468
rect 31987 2465 31999 2499
rect 32582 2496 32588 2508
rect 32495 2468 32588 2496
rect 31941 2459 31999 2465
rect 32582 2456 32588 2468
rect 32640 2496 32646 2508
rect 33137 2499 33195 2505
rect 33137 2496 33149 2499
rect 32640 2468 33149 2496
rect 32640 2456 32646 2468
rect 33137 2465 33149 2468
rect 33183 2465 33195 2499
rect 33137 2459 33195 2465
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2428 6055 2431
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 6043 2400 6653 2428
rect 6043 2397 6055 2400
rect 5997 2391 6055 2397
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 6641 2391 6699 2397
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 11057 2431 11115 2437
rect 7331 2400 8340 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 8312 2301 8340 2400
rect 11057 2397 11069 2431
rect 11103 2428 11115 2431
rect 12710 2428 12716 2440
rect 11103 2400 12112 2428
rect 12623 2400 12716 2428
rect 11103 2397 11115 2400
rect 11057 2391 11115 2397
rect 12084 2304 12112 2400
rect 12710 2388 12716 2400
rect 12768 2428 12774 2440
rect 14001 2431 14059 2437
rect 14001 2428 14013 2431
rect 12768 2400 14013 2428
rect 12768 2388 12774 2400
rect 14001 2397 14013 2400
rect 14047 2397 14059 2431
rect 14001 2391 14059 2397
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 15102 2428 15108 2440
rect 14148 2400 15108 2428
rect 14148 2388 14154 2400
rect 15102 2388 15108 2400
rect 15160 2388 15166 2440
rect 33042 2428 33048 2440
rect 30392 2400 33048 2428
rect 8297 2295 8355 2301
rect 8297 2261 8309 2295
rect 8343 2292 8355 2295
rect 8386 2292 8392 2304
rect 8343 2264 8392 2292
rect 8343 2261 8355 2264
rect 8297 2255 8355 2261
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 10134 2292 10140 2304
rect 9999 2264 10140 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 10134 2252 10140 2264
rect 10192 2252 10198 2304
rect 12066 2292 12072 2304
rect 12027 2264 12072 2292
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15611 2295 15669 2301
rect 15611 2292 15623 2295
rect 15252 2264 15623 2292
rect 15252 2252 15258 2264
rect 15611 2261 15623 2264
rect 15657 2261 15669 2295
rect 21726 2292 21732 2304
rect 21687 2264 21732 2292
rect 15611 2255 15669 2261
rect 21726 2252 21732 2264
rect 21784 2252 21790 2304
rect 30392 2292 30420 2400
rect 33042 2388 33048 2400
rect 33100 2388 33106 2440
rect 30469 2295 30527 2301
rect 30469 2292 30481 2295
rect 30392 2264 30481 2292
rect 30469 2261 30481 2264
rect 30515 2261 30527 2295
rect 30469 2255 30527 2261
rect 1104 2202 38824 2224
rect 1104 2150 7648 2202
rect 7700 2150 7712 2202
rect 7764 2150 7776 2202
rect 7828 2150 7840 2202
rect 7892 2150 20982 2202
rect 21034 2150 21046 2202
rect 21098 2150 21110 2202
rect 21162 2150 21174 2202
rect 21226 2150 34315 2202
rect 34367 2150 34379 2202
rect 34431 2150 34443 2202
rect 34495 2150 34507 2202
rect 34559 2150 38824 2202
rect 1104 2128 38824 2150
rect 12434 1844 12440 1896
rect 12492 1884 12498 1896
rect 15378 1884 15384 1896
rect 12492 1856 15384 1884
rect 12492 1844 12498 1856
rect 15378 1844 15384 1856
rect 15436 1844 15442 1896
<< via1 >>
rect 3424 13812 3476 13864
rect 19340 13812 19392 13864
rect 14315 13574 14367 13626
rect 14379 13574 14431 13626
rect 14443 13574 14495 13626
rect 14507 13574 14559 13626
rect 27648 13574 27700 13626
rect 27712 13574 27764 13626
rect 27776 13574 27828 13626
rect 27840 13574 27892 13626
rect 7648 13030 7700 13082
rect 7712 13030 7764 13082
rect 7776 13030 7828 13082
rect 7840 13030 7892 13082
rect 20982 13030 21034 13082
rect 21046 13030 21098 13082
rect 21110 13030 21162 13082
rect 21174 13030 21226 13082
rect 34315 13030 34367 13082
rect 34379 13030 34431 13082
rect 34443 13030 34495 13082
rect 34507 13030 34559 13082
rect 15200 12588 15252 12640
rect 16212 12588 16264 12640
rect 14315 12486 14367 12538
rect 14379 12486 14431 12538
rect 14443 12486 14495 12538
rect 14507 12486 14559 12538
rect 27648 12486 27700 12538
rect 27712 12486 27764 12538
rect 27776 12486 27828 12538
rect 27840 12486 27892 12538
rect 7648 11942 7700 11994
rect 7712 11942 7764 11994
rect 7776 11942 7828 11994
rect 7840 11942 7892 11994
rect 20982 11942 21034 11994
rect 21046 11942 21098 11994
rect 21110 11942 21162 11994
rect 21174 11942 21226 11994
rect 34315 11942 34367 11994
rect 34379 11942 34431 11994
rect 34443 11942 34495 11994
rect 34507 11942 34559 11994
rect 14315 11398 14367 11450
rect 14379 11398 14431 11450
rect 14443 11398 14495 11450
rect 14507 11398 14559 11450
rect 27648 11398 27700 11450
rect 27712 11398 27764 11450
rect 27776 11398 27828 11450
rect 27840 11398 27892 11450
rect 7648 10854 7700 10906
rect 7712 10854 7764 10906
rect 7776 10854 7828 10906
rect 7840 10854 7892 10906
rect 20982 10854 21034 10906
rect 21046 10854 21098 10906
rect 21110 10854 21162 10906
rect 21174 10854 21226 10906
rect 34315 10854 34367 10906
rect 34379 10854 34431 10906
rect 34443 10854 34495 10906
rect 34507 10854 34559 10906
rect 14315 10310 14367 10362
rect 14379 10310 14431 10362
rect 14443 10310 14495 10362
rect 14507 10310 14559 10362
rect 27648 10310 27700 10362
rect 27712 10310 27764 10362
rect 27776 10310 27828 10362
rect 27840 10310 27892 10362
rect 7648 9766 7700 9818
rect 7712 9766 7764 9818
rect 7776 9766 7828 9818
rect 7840 9766 7892 9818
rect 20982 9766 21034 9818
rect 21046 9766 21098 9818
rect 21110 9766 21162 9818
rect 21174 9766 21226 9818
rect 34315 9766 34367 9818
rect 34379 9766 34431 9818
rect 34443 9766 34495 9818
rect 34507 9766 34559 9818
rect 14315 9222 14367 9274
rect 14379 9222 14431 9274
rect 14443 9222 14495 9274
rect 14507 9222 14559 9274
rect 27648 9222 27700 9274
rect 27712 9222 27764 9274
rect 27776 9222 27828 9274
rect 27840 9222 27892 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 1952 8984 2004 9036
rect 6552 8984 6604 9036
rect 6460 8780 6512 8832
rect 7648 8678 7700 8730
rect 7712 8678 7764 8730
rect 7776 8678 7828 8730
rect 7840 8678 7892 8730
rect 20982 8678 21034 8730
rect 21046 8678 21098 8730
rect 21110 8678 21162 8730
rect 21174 8678 21226 8730
rect 34315 8678 34367 8730
rect 34379 8678 34431 8730
rect 34443 8678 34495 8730
rect 34507 8678 34559 8730
rect 1400 8576 1452 8628
rect 19340 8576 19392 8628
rect 6920 8508 6972 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 17040 8415 17092 8424
rect 17040 8381 17049 8415
rect 17049 8381 17083 8415
rect 17083 8381 17092 8415
rect 17040 8372 17092 8381
rect 1952 8347 2004 8356
rect 1952 8313 1961 8347
rect 1961 8313 1995 8347
rect 1995 8313 2004 8347
rect 1952 8304 2004 8313
rect 6552 8347 6604 8356
rect 6552 8313 6561 8347
rect 6561 8313 6595 8347
rect 6595 8313 6604 8347
rect 6552 8304 6604 8313
rect 7196 8304 7248 8356
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 22560 8236 22612 8288
rect 14315 8134 14367 8186
rect 14379 8134 14431 8186
rect 14443 8134 14495 8186
rect 14507 8134 14559 8186
rect 27648 8134 27700 8186
rect 27712 8134 27764 8186
rect 27776 8134 27828 8186
rect 27840 8134 27892 8186
rect 1584 8075 1636 8084
rect 1584 8041 1593 8075
rect 1593 8041 1627 8075
rect 1627 8041 1636 8075
rect 1584 8032 1636 8041
rect 16580 8032 16632 8084
rect 17868 8032 17920 8084
rect 35624 8075 35676 8084
rect 35624 8041 35633 8075
rect 35633 8041 35667 8075
rect 35667 8041 35676 8075
rect 35624 8032 35676 8041
rect 5264 7964 5316 8016
rect 7012 8007 7064 8016
rect 7012 7973 7021 8007
rect 7021 7973 7055 8007
rect 7055 7973 7064 8007
rect 7012 7964 7064 7973
rect 16672 8007 16724 8016
rect 16672 7973 16681 8007
rect 16681 7973 16715 8007
rect 16715 7973 16724 8007
rect 16672 7964 16724 7973
rect 19800 7964 19852 8016
rect 21272 7964 21324 8016
rect 28724 7964 28776 8016
rect 1860 7896 1912 7948
rect 6092 7896 6144 7948
rect 13636 7896 13688 7948
rect 14188 7939 14240 7948
rect 14188 7905 14197 7939
rect 14197 7905 14231 7939
rect 14231 7905 14240 7939
rect 14188 7896 14240 7905
rect 15660 7939 15712 7948
rect 15660 7905 15669 7939
rect 15669 7905 15703 7939
rect 15703 7905 15712 7939
rect 15660 7896 15712 7905
rect 17132 7939 17184 7948
rect 17132 7905 17141 7939
rect 17141 7905 17175 7939
rect 17175 7905 17184 7939
rect 17132 7896 17184 7905
rect 35440 7939 35492 7948
rect 35440 7905 35449 7939
rect 35449 7905 35483 7939
rect 35483 7905 35492 7939
rect 35440 7896 35492 7905
rect 6736 7760 6788 7812
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 7104 7828 7156 7880
rect 20812 7828 20864 7880
rect 28448 7828 28500 7880
rect 28908 7871 28960 7880
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 6644 7692 6696 7701
rect 13728 7692 13780 7744
rect 13820 7692 13872 7744
rect 16396 7692 16448 7744
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 19524 7735 19576 7744
rect 19524 7701 19533 7735
rect 19533 7701 19567 7735
rect 19567 7701 19576 7735
rect 19524 7692 19576 7701
rect 22008 7692 22060 7744
rect 26056 7692 26108 7744
rect 7648 7590 7700 7642
rect 7712 7590 7764 7642
rect 7776 7590 7828 7642
rect 7840 7590 7892 7642
rect 20982 7590 21034 7642
rect 21046 7590 21098 7642
rect 21110 7590 21162 7642
rect 21174 7590 21226 7642
rect 34315 7590 34367 7642
rect 34379 7590 34431 7642
rect 34443 7590 34495 7642
rect 34507 7590 34559 7642
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 2228 7488 2280 7540
rect 7012 7488 7064 7540
rect 16028 7488 16080 7540
rect 16948 7488 17000 7540
rect 17132 7488 17184 7540
rect 21272 7531 21324 7540
rect 21272 7497 21281 7531
rect 21281 7497 21315 7531
rect 21315 7497 21324 7531
rect 21272 7488 21324 7497
rect 28448 7531 28500 7540
rect 28448 7497 28457 7531
rect 28457 7497 28491 7531
rect 28491 7497 28500 7531
rect 28448 7488 28500 7497
rect 28724 7488 28776 7540
rect 29000 7488 29052 7540
rect 15752 7463 15804 7472
rect 15752 7429 15761 7463
rect 15761 7429 15795 7463
rect 15795 7429 15804 7463
rect 16488 7463 16540 7472
rect 15752 7420 15804 7429
rect 16488 7429 16497 7463
rect 16497 7429 16531 7463
rect 16531 7429 16540 7463
rect 16488 7420 16540 7429
rect 16580 7395 16632 7404
rect 5264 7327 5316 7336
rect 5264 7293 5273 7327
rect 5273 7293 5307 7327
rect 5307 7293 5316 7327
rect 5264 7284 5316 7293
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 6920 7216 6972 7268
rect 1492 7148 1544 7200
rect 5080 7191 5132 7200
rect 5080 7157 5089 7191
rect 5089 7157 5123 7191
rect 5123 7157 5132 7191
rect 5080 7148 5132 7157
rect 6092 7148 6144 7200
rect 6552 7191 6604 7200
rect 6552 7157 6561 7191
rect 6561 7157 6595 7191
rect 6595 7157 6604 7191
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 14740 7284 14792 7336
rect 16580 7361 16589 7395
rect 16589 7361 16623 7395
rect 16623 7361 16632 7395
rect 16580 7352 16632 7361
rect 19524 7352 19576 7404
rect 16304 7284 16356 7336
rect 18512 7327 18564 7336
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 19984 7327 20036 7336
rect 13176 7259 13228 7268
rect 13176 7225 13185 7259
rect 13185 7225 13219 7259
rect 13219 7225 13228 7259
rect 13176 7216 13228 7225
rect 14188 7216 14240 7268
rect 14832 7216 14884 7268
rect 15936 7216 15988 7268
rect 16672 7216 16724 7268
rect 16948 7259 17000 7268
rect 16948 7225 16957 7259
rect 16957 7225 16991 7259
rect 16991 7225 17000 7259
rect 16948 7216 17000 7225
rect 6552 7148 6604 7157
rect 8208 7148 8260 7200
rect 8760 7191 8812 7200
rect 8760 7157 8769 7191
rect 8769 7157 8803 7191
rect 8803 7157 8812 7191
rect 8760 7148 8812 7157
rect 9128 7191 9180 7200
rect 9128 7157 9137 7191
rect 9137 7157 9171 7191
rect 9171 7157 9180 7191
rect 9128 7148 9180 7157
rect 13636 7148 13688 7200
rect 13820 7191 13872 7200
rect 13820 7157 13829 7191
rect 13829 7157 13863 7191
rect 13863 7157 13872 7191
rect 13820 7148 13872 7157
rect 14924 7191 14976 7200
rect 14924 7157 14933 7191
rect 14933 7157 14967 7191
rect 14967 7157 14976 7191
rect 14924 7148 14976 7157
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 21640 7352 21692 7404
rect 20720 7327 20772 7336
rect 20720 7293 20729 7327
rect 20729 7293 20763 7327
rect 20763 7293 20772 7327
rect 20720 7284 20772 7293
rect 25136 7327 25188 7336
rect 25136 7293 25145 7327
rect 25145 7293 25179 7327
rect 25179 7293 25188 7327
rect 25136 7284 25188 7293
rect 25688 7327 25740 7336
rect 25688 7293 25697 7327
rect 25697 7293 25731 7327
rect 25731 7293 25740 7327
rect 25688 7284 25740 7293
rect 26056 7327 26108 7336
rect 26056 7293 26065 7327
rect 26065 7293 26099 7327
rect 26099 7293 26108 7327
rect 26056 7284 26108 7293
rect 26424 7327 26476 7336
rect 26424 7293 26433 7327
rect 26433 7293 26467 7327
rect 26467 7293 26476 7327
rect 26424 7284 26476 7293
rect 28908 7284 28960 7336
rect 29828 7284 29880 7336
rect 35440 7327 35492 7336
rect 35440 7293 35449 7327
rect 35449 7293 35483 7327
rect 35483 7293 35492 7327
rect 35440 7284 35492 7293
rect 20536 7216 20588 7268
rect 22008 7259 22060 7268
rect 22008 7225 22017 7259
rect 22017 7225 22051 7259
rect 22051 7225 22060 7259
rect 22008 7216 22060 7225
rect 22560 7259 22612 7268
rect 22560 7225 22569 7259
rect 22569 7225 22603 7259
rect 22603 7225 22612 7259
rect 22560 7216 22612 7225
rect 26700 7259 26752 7268
rect 26700 7225 26709 7259
rect 26709 7225 26743 7259
rect 26743 7225 26752 7259
rect 26700 7216 26752 7225
rect 18972 7191 19024 7200
rect 18972 7157 18981 7191
rect 18981 7157 19015 7191
rect 19015 7157 19024 7191
rect 18972 7148 19024 7157
rect 20628 7148 20680 7200
rect 21640 7191 21692 7200
rect 21640 7157 21649 7191
rect 21649 7157 21683 7191
rect 21683 7157 21692 7191
rect 21640 7148 21692 7157
rect 24676 7191 24728 7200
rect 24676 7157 24685 7191
rect 24685 7157 24719 7191
rect 24719 7157 24728 7191
rect 24676 7148 24728 7157
rect 14315 7046 14367 7098
rect 14379 7046 14431 7098
rect 14443 7046 14495 7098
rect 14507 7046 14559 7098
rect 27648 7046 27700 7098
rect 27712 7046 27764 7098
rect 27776 7046 27828 7098
rect 27840 7046 27892 7098
rect 5540 6944 5592 6996
rect 13636 6987 13688 6996
rect 13636 6953 13645 6987
rect 13645 6953 13679 6987
rect 13679 6953 13688 6987
rect 13636 6944 13688 6953
rect 14740 6987 14792 6996
rect 14740 6953 14749 6987
rect 14749 6953 14783 6987
rect 14783 6953 14792 6987
rect 14740 6944 14792 6953
rect 15660 6944 15712 6996
rect 20812 6944 20864 6996
rect 24676 6987 24728 6996
rect 24676 6953 24685 6987
rect 24685 6953 24719 6987
rect 24719 6953 24728 6987
rect 24676 6944 24728 6953
rect 25320 6987 25372 6996
rect 25320 6953 25329 6987
rect 25329 6953 25363 6987
rect 25363 6953 25372 6987
rect 25320 6944 25372 6953
rect 25688 6944 25740 6996
rect 28724 6944 28776 6996
rect 2320 6808 2372 6860
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4804 6672 4856 6724
rect 5264 6808 5316 6860
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 6276 6808 6328 6860
rect 6920 6808 6972 6860
rect 7380 6808 7432 6860
rect 11980 6876 12032 6928
rect 13176 6876 13228 6928
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 9680 6783 9732 6792
rect 6460 6672 6512 6724
rect 1400 6604 1452 6656
rect 5172 6604 5224 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7104 6672 7156 6724
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 12992 6851 13044 6860
rect 12992 6817 13001 6851
rect 13001 6817 13035 6851
rect 13035 6817 13044 6851
rect 12992 6808 13044 6817
rect 15752 6876 15804 6928
rect 17132 6808 17184 6860
rect 21640 6876 21692 6928
rect 21364 6851 21416 6860
rect 13176 6783 13228 6792
rect 13176 6749 13182 6783
rect 13182 6749 13228 6783
rect 13176 6740 13228 6749
rect 14924 6740 14976 6792
rect 16028 6783 16080 6792
rect 16028 6749 16037 6783
rect 16037 6749 16071 6783
rect 16071 6749 16080 6783
rect 16028 6740 16080 6749
rect 18880 6740 18932 6792
rect 18972 6740 19024 6792
rect 20536 6740 20588 6792
rect 21364 6817 21373 6851
rect 21373 6817 21407 6851
rect 21407 6817 21416 6851
rect 21364 6808 21416 6817
rect 21916 6851 21968 6860
rect 21916 6817 21925 6851
rect 21925 6817 21959 6851
rect 21959 6817 21968 6851
rect 21916 6808 21968 6817
rect 24308 6851 24360 6860
rect 21824 6740 21876 6792
rect 24308 6817 24317 6851
rect 24317 6817 24351 6851
rect 24351 6817 24360 6851
rect 24308 6808 24360 6817
rect 26424 6808 26476 6860
rect 26700 6808 26752 6860
rect 15936 6715 15988 6724
rect 15936 6681 15945 6715
rect 15945 6681 15979 6715
rect 15979 6681 15988 6715
rect 15936 6672 15988 6681
rect 21364 6672 21416 6724
rect 21732 6672 21784 6724
rect 27160 6740 27212 6792
rect 29184 6876 29236 6928
rect 29828 6783 29880 6792
rect 29828 6749 29837 6783
rect 29837 6749 29871 6783
rect 29871 6749 29880 6783
rect 29828 6740 29880 6749
rect 30288 6740 30340 6792
rect 30012 6672 30064 6724
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 13636 6604 13688 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 17408 6647 17460 6656
rect 17408 6613 17417 6647
rect 17417 6613 17451 6647
rect 17451 6613 17460 6647
rect 17408 6604 17460 6613
rect 18052 6604 18104 6656
rect 18972 6604 19024 6656
rect 19432 6604 19484 6656
rect 19984 6604 20036 6656
rect 20720 6604 20772 6656
rect 22100 6604 22152 6656
rect 25596 6604 25648 6656
rect 7648 6502 7700 6554
rect 7712 6502 7764 6554
rect 7776 6502 7828 6554
rect 7840 6502 7892 6554
rect 20982 6502 21034 6554
rect 21046 6502 21098 6554
rect 21110 6502 21162 6554
rect 21174 6502 21226 6554
rect 34315 6502 34367 6554
rect 34379 6502 34431 6554
rect 34443 6502 34495 6554
rect 34507 6502 34559 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 6460 6400 6512 6452
rect 8024 6400 8076 6452
rect 8760 6400 8812 6452
rect 13084 6400 13136 6452
rect 16028 6400 16080 6452
rect 8208 6375 8260 6384
rect 8208 6341 8217 6375
rect 8217 6341 8251 6375
rect 8251 6341 8260 6375
rect 8208 6332 8260 6341
rect 13636 6375 13688 6384
rect 13636 6341 13645 6375
rect 13645 6341 13679 6375
rect 13679 6341 13688 6375
rect 13636 6332 13688 6341
rect 5080 6264 5132 6316
rect 4804 6196 4856 6248
rect 5172 6239 5224 6248
rect 5172 6205 5181 6239
rect 5181 6205 5215 6239
rect 5215 6205 5224 6239
rect 5172 6196 5224 6205
rect 6184 6264 6236 6316
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 6920 6264 6972 6316
rect 5816 6196 5868 6205
rect 6460 6196 6512 6248
rect 7564 6239 7616 6248
rect 7564 6205 7573 6239
rect 7573 6205 7607 6239
rect 7607 6205 7616 6239
rect 7564 6196 7616 6205
rect 8024 6196 8076 6248
rect 4068 6128 4120 6180
rect 6920 6128 6972 6180
rect 8300 6196 8352 6248
rect 11336 6239 11388 6248
rect 11336 6205 11380 6239
rect 11380 6205 11388 6239
rect 11336 6196 11388 6205
rect 12072 6196 12124 6248
rect 13084 6196 13136 6248
rect 14096 6239 14148 6248
rect 14096 6205 14105 6239
rect 14105 6205 14139 6239
rect 14139 6205 14148 6239
rect 14096 6196 14148 6205
rect 14740 6239 14792 6248
rect 9128 6171 9180 6180
rect 2044 6103 2096 6112
rect 2044 6069 2053 6103
rect 2053 6069 2087 6103
rect 2087 6069 2096 6103
rect 2044 6060 2096 6069
rect 4344 6103 4396 6112
rect 4344 6069 4353 6103
rect 4353 6069 4387 6103
rect 4387 6069 4396 6103
rect 4344 6060 4396 6069
rect 4528 6103 4580 6112
rect 4528 6069 4537 6103
rect 4537 6069 4571 6103
rect 4571 6069 4580 6103
rect 4528 6060 4580 6069
rect 9128 6137 9137 6171
rect 9137 6137 9171 6171
rect 9171 6137 9180 6171
rect 9128 6128 9180 6137
rect 12992 6128 13044 6180
rect 14740 6205 14749 6239
rect 14749 6205 14783 6239
rect 14783 6205 14792 6239
rect 14740 6196 14792 6205
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 17132 6400 17184 6452
rect 18512 6443 18564 6452
rect 18512 6409 18521 6443
rect 18521 6409 18555 6443
rect 18555 6409 18564 6443
rect 18512 6400 18564 6409
rect 18880 6443 18932 6452
rect 18880 6409 18889 6443
rect 18889 6409 18923 6443
rect 18923 6409 18932 6443
rect 18880 6400 18932 6409
rect 22100 6443 22152 6452
rect 22100 6409 22109 6443
rect 22109 6409 22143 6443
rect 22143 6409 22152 6443
rect 22100 6400 22152 6409
rect 24216 6443 24268 6452
rect 24216 6409 24225 6443
rect 24225 6409 24259 6443
rect 24259 6409 24268 6443
rect 24216 6400 24268 6409
rect 26700 6400 26752 6452
rect 33416 6443 33468 6452
rect 33416 6409 33425 6443
rect 33425 6409 33459 6443
rect 33459 6409 33468 6443
rect 33416 6400 33468 6409
rect 29184 6332 29236 6384
rect 20720 6264 20772 6316
rect 18512 6196 18564 6248
rect 20444 6239 20496 6248
rect 14648 6128 14700 6180
rect 20444 6205 20453 6239
rect 20453 6205 20487 6239
rect 20487 6205 20496 6239
rect 20444 6196 20496 6205
rect 20536 6128 20588 6180
rect 21732 6196 21784 6248
rect 24216 6196 24268 6248
rect 25136 6239 25188 6248
rect 25136 6205 25145 6239
rect 25145 6205 25179 6239
rect 25179 6205 25188 6239
rect 25136 6196 25188 6205
rect 25596 6239 25648 6248
rect 25596 6205 25605 6239
rect 25605 6205 25639 6239
rect 25639 6205 25648 6239
rect 25596 6196 25648 6205
rect 26056 6239 26108 6248
rect 26056 6205 26065 6239
rect 26065 6205 26099 6239
rect 26099 6205 26108 6239
rect 26424 6239 26476 6248
rect 26056 6196 26108 6205
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 27528 6196 27580 6248
rect 27712 6239 27764 6248
rect 27712 6205 27756 6239
rect 27756 6205 27764 6239
rect 27712 6196 27764 6205
rect 27988 6196 28040 6248
rect 29276 6239 29328 6248
rect 29276 6205 29285 6239
rect 29285 6205 29319 6239
rect 29319 6205 29328 6239
rect 29276 6196 29328 6205
rect 33232 6239 33284 6248
rect 33232 6205 33241 6239
rect 33241 6205 33275 6239
rect 33275 6205 33284 6239
rect 33232 6196 33284 6205
rect 10140 6103 10192 6112
rect 10140 6069 10149 6103
rect 10149 6069 10183 6103
rect 10183 6069 10192 6103
rect 10140 6060 10192 6069
rect 10968 6060 11020 6112
rect 11704 6060 11756 6112
rect 12716 6103 12768 6112
rect 12716 6069 12725 6103
rect 12725 6069 12759 6103
rect 12759 6069 12768 6103
rect 12716 6060 12768 6069
rect 14188 6103 14240 6112
rect 14188 6069 14197 6103
rect 14197 6069 14231 6103
rect 14231 6069 14240 6103
rect 14188 6060 14240 6069
rect 16672 6103 16724 6112
rect 16672 6069 16681 6103
rect 16681 6069 16715 6103
rect 16715 6069 16724 6103
rect 16672 6060 16724 6069
rect 17316 6060 17368 6112
rect 19800 6103 19852 6112
rect 19800 6069 19809 6103
rect 19809 6069 19843 6103
rect 19843 6069 19852 6103
rect 21916 6128 21968 6180
rect 21364 6103 21416 6112
rect 19800 6060 19852 6069
rect 21364 6069 21373 6103
rect 21373 6069 21407 6103
rect 21407 6069 21416 6103
rect 21364 6060 21416 6069
rect 21824 6103 21876 6112
rect 21824 6069 21833 6103
rect 21833 6069 21867 6103
rect 21867 6069 21876 6103
rect 21824 6060 21876 6069
rect 23848 6103 23900 6112
rect 23848 6069 23857 6103
rect 23857 6069 23891 6103
rect 23891 6069 23900 6103
rect 23848 6060 23900 6069
rect 24124 6128 24176 6180
rect 27344 6128 27396 6180
rect 26148 6060 26200 6112
rect 27160 6060 27212 6112
rect 28080 6060 28132 6112
rect 28816 6060 28868 6112
rect 30012 6060 30064 6112
rect 14315 5958 14367 6010
rect 14379 5958 14431 6010
rect 14443 5958 14495 6010
rect 14507 5958 14559 6010
rect 27648 5958 27700 6010
rect 27712 5958 27764 6010
rect 27776 5958 27828 6010
rect 27840 5958 27892 6010
rect 7380 5856 7432 5908
rect 9588 5856 9640 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 12992 5856 13044 5908
rect 2136 5831 2188 5840
rect 2136 5797 2145 5831
rect 2145 5797 2179 5831
rect 2179 5797 2188 5831
rect 2136 5788 2188 5797
rect 7472 5788 7524 5840
rect 10140 5788 10192 5840
rect 13452 5856 13504 5908
rect 15660 5856 15712 5908
rect 15752 5856 15804 5908
rect 20444 5856 20496 5908
rect 20812 5856 20864 5908
rect 28080 5856 28132 5908
rect 28816 5856 28868 5908
rect 15936 5788 15988 5840
rect 21272 5831 21324 5840
rect 21272 5797 21275 5831
rect 21275 5797 21309 5831
rect 21309 5797 21324 5831
rect 21272 5788 21324 5797
rect 23848 5788 23900 5840
rect 24860 5788 24912 5840
rect 6460 5763 6512 5772
rect 6460 5729 6469 5763
rect 6469 5729 6503 5763
rect 6503 5729 6512 5763
rect 6460 5720 6512 5729
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 7380 5763 7432 5772
rect 2780 5652 2832 5704
rect 4344 5652 4396 5704
rect 5816 5652 5868 5704
rect 7380 5729 7389 5763
rect 7389 5729 7423 5763
rect 7423 5729 7432 5763
rect 7380 5720 7432 5729
rect 8576 5763 8628 5772
rect 8576 5729 8594 5763
rect 8594 5729 8628 5763
rect 8576 5720 8628 5729
rect 10324 5763 10376 5772
rect 10324 5729 10333 5763
rect 10333 5729 10367 5763
rect 10367 5729 10376 5763
rect 10324 5720 10376 5729
rect 10600 5763 10652 5772
rect 10600 5729 10609 5763
rect 10609 5729 10643 5763
rect 10643 5729 10652 5763
rect 10600 5720 10652 5729
rect 10876 5720 10928 5772
rect 11244 5720 11296 5772
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 12992 5763 13044 5772
rect 12992 5729 13001 5763
rect 13001 5729 13035 5763
rect 13035 5729 13044 5763
rect 12992 5720 13044 5729
rect 8024 5652 8076 5704
rect 12348 5652 12400 5704
rect 13728 5720 13780 5772
rect 15108 5720 15160 5772
rect 15844 5763 15896 5772
rect 15844 5729 15853 5763
rect 15853 5729 15887 5763
rect 15887 5729 15896 5763
rect 15844 5720 15896 5729
rect 17316 5763 17368 5772
rect 17316 5729 17325 5763
rect 17325 5729 17359 5763
rect 17359 5729 17368 5763
rect 17316 5720 17368 5729
rect 17408 5720 17460 5772
rect 17960 5763 18012 5772
rect 17960 5729 17969 5763
rect 17969 5729 18003 5763
rect 18003 5729 18012 5763
rect 17960 5720 18012 5729
rect 18052 5720 18104 5772
rect 19708 5763 19760 5772
rect 19708 5729 19752 5763
rect 19752 5729 19760 5763
rect 19708 5720 19760 5729
rect 20720 5720 20772 5772
rect 22008 5720 22060 5772
rect 22100 5720 22152 5772
rect 24124 5763 24176 5772
rect 24124 5729 24133 5763
rect 24133 5729 24167 5763
rect 24167 5729 24176 5763
rect 24124 5720 24176 5729
rect 2596 5627 2648 5636
rect 2596 5593 2605 5627
rect 2605 5593 2639 5627
rect 2639 5593 2648 5627
rect 2596 5584 2648 5593
rect 6920 5584 6972 5636
rect 12440 5584 12492 5636
rect 13820 5652 13872 5704
rect 14740 5652 14792 5704
rect 19524 5652 19576 5704
rect 24492 5652 24544 5704
rect 26332 5720 26384 5772
rect 25320 5652 25372 5704
rect 26792 5763 26844 5772
rect 26792 5729 26801 5763
rect 26801 5729 26835 5763
rect 26835 5729 26844 5763
rect 26792 5720 26844 5729
rect 27344 5763 27396 5772
rect 18512 5627 18564 5636
rect 18512 5593 18521 5627
rect 18521 5593 18555 5627
rect 18555 5593 18564 5627
rect 18512 5584 18564 5593
rect 1676 5559 1728 5568
rect 1676 5525 1685 5559
rect 1685 5525 1719 5559
rect 1719 5525 1728 5559
rect 1676 5516 1728 5525
rect 5172 5516 5224 5568
rect 6276 5516 6328 5568
rect 8392 5516 8444 5568
rect 9496 5559 9548 5568
rect 9496 5525 9505 5559
rect 9505 5525 9539 5559
rect 9539 5525 9548 5559
rect 9496 5516 9548 5525
rect 14648 5516 14700 5568
rect 17960 5516 18012 5568
rect 19340 5516 19392 5568
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 22100 5516 22152 5568
rect 25596 5516 25648 5568
rect 27344 5729 27353 5763
rect 27353 5729 27387 5763
rect 27387 5729 27396 5763
rect 27344 5720 27396 5729
rect 27528 5720 27580 5772
rect 29276 5652 29328 5704
rect 30380 5516 30432 5568
rect 30932 5559 30984 5568
rect 30932 5525 30941 5559
rect 30941 5525 30975 5559
rect 30975 5525 30984 5559
rect 30932 5516 30984 5525
rect 7648 5414 7700 5466
rect 7712 5414 7764 5466
rect 7776 5414 7828 5466
rect 7840 5414 7892 5466
rect 20982 5414 21034 5466
rect 21046 5414 21098 5466
rect 21110 5414 21162 5466
rect 21174 5414 21226 5466
rect 34315 5414 34367 5466
rect 34379 5414 34431 5466
rect 34443 5414 34495 5466
rect 34507 5414 34559 5466
rect 2136 5312 2188 5364
rect 3332 5312 3384 5364
rect 6828 5312 6880 5364
rect 8208 5312 8260 5364
rect 10600 5312 10652 5364
rect 12348 5312 12400 5364
rect 15844 5355 15896 5364
rect 15844 5321 15853 5355
rect 15853 5321 15887 5355
rect 15887 5321 15896 5355
rect 15844 5312 15896 5321
rect 16212 5355 16264 5364
rect 16212 5321 16221 5355
rect 16221 5321 16255 5355
rect 16255 5321 16264 5355
rect 16212 5312 16264 5321
rect 17868 5312 17920 5364
rect 17960 5312 18012 5364
rect 19708 5355 19760 5364
rect 19708 5321 19717 5355
rect 19717 5321 19751 5355
rect 19751 5321 19760 5355
rect 19708 5312 19760 5321
rect 21272 5312 21324 5364
rect 22192 5312 22244 5364
rect 24124 5355 24176 5364
rect 24124 5321 24133 5355
rect 24133 5321 24167 5355
rect 24167 5321 24176 5355
rect 24124 5312 24176 5321
rect 6552 5244 6604 5296
rect 8024 5287 8076 5296
rect 8024 5253 8033 5287
rect 8033 5253 8067 5287
rect 8067 5253 8076 5287
rect 8024 5244 8076 5253
rect 24492 5287 24544 5296
rect 24492 5253 24501 5287
rect 24501 5253 24535 5287
rect 24535 5253 24544 5287
rect 24492 5244 24544 5253
rect 2780 5176 2832 5228
rect 3884 5219 3936 5228
rect 3884 5185 3893 5219
rect 3893 5185 3927 5219
rect 3927 5185 3936 5219
rect 3884 5176 3936 5185
rect 3700 5108 3752 5160
rect 6920 5176 6972 5228
rect 4804 5108 4856 5160
rect 5172 5151 5224 5160
rect 5172 5117 5181 5151
rect 5181 5117 5215 5151
rect 5215 5117 5224 5151
rect 5172 5108 5224 5117
rect 5448 5151 5500 5160
rect 5448 5117 5457 5151
rect 5457 5117 5491 5151
rect 5491 5117 5500 5151
rect 5448 5108 5500 5117
rect 5816 5151 5868 5160
rect 5816 5117 5825 5151
rect 5825 5117 5859 5151
rect 5859 5117 5868 5151
rect 5816 5108 5868 5117
rect 10324 5151 10376 5160
rect 1676 5040 1728 5092
rect 4160 5040 4212 5092
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6460 4972 6512 5024
rect 10324 5117 10333 5151
rect 10333 5117 10367 5151
rect 10367 5117 10376 5151
rect 10324 5108 10376 5117
rect 10876 5151 10928 5160
rect 9864 5040 9916 5092
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 8944 4972 8996 5024
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 10876 5108 10928 5117
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 12440 5040 12492 5092
rect 12624 5083 12676 5092
rect 12624 5049 12633 5083
rect 12633 5049 12667 5083
rect 12667 5049 12676 5083
rect 12624 5040 12676 5049
rect 12716 5083 12768 5092
rect 12716 5049 12725 5083
rect 12725 5049 12759 5083
rect 12759 5049 12768 5083
rect 12716 5040 12768 5049
rect 13636 5040 13688 5092
rect 10968 4972 11020 5024
rect 14648 5176 14700 5228
rect 14096 5108 14148 5160
rect 14372 5151 14424 5160
rect 14372 5117 14381 5151
rect 14381 5117 14415 5151
rect 14415 5117 14424 5151
rect 14372 5108 14424 5117
rect 15844 5176 15896 5228
rect 17132 5219 17184 5228
rect 17132 5185 17141 5219
rect 17141 5185 17175 5219
rect 17175 5185 17184 5219
rect 17132 5176 17184 5185
rect 22284 5219 22336 5228
rect 14924 5151 14976 5160
rect 14924 5117 14933 5151
rect 14933 5117 14967 5151
rect 14967 5117 14976 5151
rect 14924 5108 14976 5117
rect 15200 5108 15252 5160
rect 16212 5108 16264 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 20720 5108 20772 5117
rect 20812 5108 20864 5160
rect 22284 5185 22293 5219
rect 22293 5185 22327 5219
rect 22327 5185 22336 5219
rect 22284 5176 22336 5185
rect 21088 5108 21140 5160
rect 21456 5108 21508 5160
rect 21732 5151 21784 5160
rect 21732 5117 21741 5151
rect 21741 5117 21775 5151
rect 21775 5117 21784 5151
rect 21732 5108 21784 5117
rect 30380 5312 30432 5364
rect 31024 5312 31076 5364
rect 25688 5244 25740 5296
rect 27344 5244 27396 5296
rect 28908 5244 28960 5296
rect 26792 5176 26844 5228
rect 28080 5176 28132 5228
rect 29644 5176 29696 5228
rect 30012 5219 30064 5228
rect 30012 5185 30021 5219
rect 30021 5185 30055 5219
rect 30055 5185 30064 5219
rect 30012 5176 30064 5185
rect 30288 5176 30340 5228
rect 25596 5108 25648 5160
rect 26056 5108 26108 5160
rect 26332 5108 26384 5160
rect 27528 5040 27580 5092
rect 28172 5040 28224 5092
rect 29368 5083 29420 5092
rect 29368 5049 29377 5083
rect 29377 5049 29411 5083
rect 29411 5049 29420 5083
rect 29368 5040 29420 5049
rect 29460 5083 29512 5092
rect 29460 5049 29469 5083
rect 29469 5049 29503 5083
rect 29503 5049 29512 5083
rect 30932 5083 30984 5092
rect 29460 5040 29512 5049
rect 30932 5049 30941 5083
rect 30941 5049 30975 5083
rect 30975 5049 30984 5083
rect 30932 5040 30984 5049
rect 31024 5083 31076 5092
rect 31024 5049 31033 5083
rect 31033 5049 31067 5083
rect 31067 5049 31076 5083
rect 31024 5040 31076 5049
rect 15292 5015 15344 5024
rect 15292 4981 15301 5015
rect 15301 4981 15335 5015
rect 15335 4981 15344 5015
rect 15292 4972 15344 4981
rect 17776 5015 17828 5024
rect 17776 4981 17785 5015
rect 17785 4981 17819 5015
rect 17819 4981 17828 5015
rect 17776 4972 17828 4981
rect 19248 4972 19300 5024
rect 20812 5015 20864 5024
rect 20812 4981 20821 5015
rect 20821 4981 20855 5015
rect 20855 4981 20864 5015
rect 20812 4972 20864 4981
rect 23480 5015 23532 5024
rect 23480 4981 23489 5015
rect 23489 4981 23523 5015
rect 23523 4981 23532 5015
rect 23480 4972 23532 4981
rect 28816 5015 28868 5024
rect 28816 4981 28825 5015
rect 28825 4981 28859 5015
rect 28859 4981 28868 5015
rect 28816 4972 28868 4981
rect 30564 4972 30616 5024
rect 14315 4870 14367 4922
rect 14379 4870 14431 4922
rect 14443 4870 14495 4922
rect 14507 4870 14559 4922
rect 27648 4870 27700 4922
rect 27712 4870 27764 4922
rect 27776 4870 27828 4922
rect 27840 4870 27892 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 4804 4768 4856 4820
rect 5724 4768 5776 4820
rect 1676 4700 1728 4752
rect 5172 4700 5224 4752
rect 6828 4768 6880 4820
rect 7012 4768 7064 4820
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 12256 4768 12308 4820
rect 12716 4768 12768 4820
rect 4252 4675 4304 4684
rect 4252 4641 4261 4675
rect 4261 4641 4295 4675
rect 4295 4641 4304 4675
rect 4252 4632 4304 4641
rect 5724 4675 5776 4684
rect 5724 4641 5733 4675
rect 5733 4641 5767 4675
rect 5767 4641 5776 4675
rect 5724 4632 5776 4641
rect 8208 4743 8260 4752
rect 8208 4709 8217 4743
rect 8217 4709 8251 4743
rect 8251 4709 8260 4743
rect 8208 4700 8260 4709
rect 10324 4700 10376 4752
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 7288 4632 7340 4684
rect 12808 4700 12860 4752
rect 13820 4743 13872 4752
rect 13820 4709 13823 4743
rect 13823 4709 13857 4743
rect 13857 4709 13872 4743
rect 13820 4700 13872 4709
rect 14096 4700 14148 4752
rect 14924 4700 14976 4752
rect 19524 4768 19576 4820
rect 21088 4768 21140 4820
rect 23480 4768 23532 4820
rect 25136 4768 25188 4820
rect 26332 4768 26384 4820
rect 29368 4768 29420 4820
rect 29828 4811 29880 4820
rect 29828 4777 29837 4811
rect 29837 4777 29871 4811
rect 29871 4777 29880 4811
rect 29828 4768 29880 4777
rect 15844 4700 15896 4752
rect 18052 4700 18104 4752
rect 19340 4743 19392 4752
rect 19340 4709 19349 4743
rect 19349 4709 19383 4743
rect 19383 4709 19392 4743
rect 19340 4700 19392 4709
rect 19432 4743 19484 4752
rect 19432 4709 19441 4743
rect 19441 4709 19475 4743
rect 19475 4709 19484 4743
rect 21272 4743 21324 4752
rect 19432 4700 19484 4709
rect 21272 4709 21275 4743
rect 21275 4709 21309 4743
rect 21309 4709 21324 4743
rect 21272 4700 21324 4709
rect 22100 4700 22152 4752
rect 22836 4743 22888 4752
rect 22836 4709 22845 4743
rect 22845 4709 22879 4743
rect 22879 4709 22888 4743
rect 22836 4700 22888 4709
rect 24860 4743 24912 4752
rect 24860 4709 24869 4743
rect 24869 4709 24903 4743
rect 24903 4709 24912 4743
rect 24860 4700 24912 4709
rect 26056 4700 26108 4752
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 2504 4564 2556 4616
rect 6736 4564 6788 4616
rect 8300 4564 8352 4616
rect 8484 4607 8536 4616
rect 8484 4573 8493 4607
rect 8493 4573 8527 4607
rect 8527 4573 8536 4607
rect 8484 4564 8536 4573
rect 10876 4564 10928 4616
rect 11244 4632 11296 4684
rect 13452 4675 13504 4684
rect 12348 4564 12400 4616
rect 11612 4539 11664 4548
rect 11612 4505 11621 4539
rect 11621 4505 11655 4539
rect 11655 4505 11664 4539
rect 11612 4496 11664 4505
rect 13452 4641 13461 4675
rect 13461 4641 13495 4675
rect 13495 4641 13504 4675
rect 13452 4632 13504 4641
rect 15660 4632 15712 4684
rect 16764 4632 16816 4684
rect 17224 4632 17276 4684
rect 17408 4675 17460 4684
rect 17408 4641 17417 4675
rect 17417 4641 17451 4675
rect 17451 4641 17460 4675
rect 17408 4632 17460 4641
rect 17960 4675 18012 4684
rect 16580 4564 16632 4616
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 20720 4632 20772 4684
rect 21364 4632 21416 4684
rect 24676 4632 24728 4684
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 22744 4607 22796 4616
rect 19984 4564 20036 4573
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 13728 4496 13780 4548
rect 16120 4496 16172 4548
rect 22100 4496 22152 4548
rect 22560 4496 22612 4548
rect 25596 4564 25648 4616
rect 25872 4564 25924 4616
rect 27160 4700 27212 4752
rect 28816 4700 28868 4752
rect 30564 4743 30616 4752
rect 30564 4709 30573 4743
rect 30573 4709 30607 4743
rect 30607 4709 30616 4743
rect 30564 4700 30616 4709
rect 29460 4632 29512 4684
rect 26884 4607 26936 4616
rect 26884 4573 26893 4607
rect 26893 4573 26927 4607
rect 26927 4573 26936 4607
rect 26884 4564 26936 4573
rect 27528 4564 27580 4616
rect 28632 4607 28684 4616
rect 28632 4573 28641 4607
rect 28641 4573 28675 4607
rect 28675 4573 28684 4607
rect 28632 4564 28684 4573
rect 30472 4607 30524 4616
rect 30472 4573 30481 4607
rect 30481 4573 30515 4607
rect 30515 4573 30524 4607
rect 30472 4564 30524 4573
rect 24400 4539 24452 4548
rect 24400 4505 24409 4539
rect 24409 4505 24443 4539
rect 24443 4505 24452 4539
rect 24400 4496 24452 4505
rect 30380 4496 30432 4548
rect 30932 4564 30984 4616
rect 1952 4428 2004 4480
rect 3884 4428 3936 4480
rect 21824 4471 21876 4480
rect 21824 4437 21833 4471
rect 21833 4437 21867 4471
rect 21867 4437 21876 4471
rect 21824 4428 21876 4437
rect 23480 4428 23532 4480
rect 28172 4471 28224 4480
rect 28172 4437 28181 4471
rect 28181 4437 28215 4471
rect 28215 4437 28224 4471
rect 28172 4428 28224 4437
rect 28540 4471 28592 4480
rect 28540 4437 28549 4471
rect 28549 4437 28583 4471
rect 28583 4437 28592 4471
rect 28540 4428 28592 4437
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 7648 4326 7700 4378
rect 7712 4326 7764 4378
rect 7776 4326 7828 4378
rect 7840 4326 7892 4378
rect 20982 4326 21034 4378
rect 21046 4326 21098 4378
rect 21110 4326 21162 4378
rect 21174 4326 21226 4378
rect 34315 4326 34367 4378
rect 34379 4326 34431 4378
rect 34443 4326 34495 4378
rect 34507 4326 34559 4378
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 5448 4224 5500 4276
rect 6460 4224 6512 4276
rect 8208 4224 8260 4276
rect 10324 4224 10376 4276
rect 10968 4267 11020 4276
rect 10968 4233 10977 4267
rect 10977 4233 11011 4267
rect 11011 4233 11020 4267
rect 10968 4224 11020 4233
rect 15660 4224 15712 4276
rect 15844 4267 15896 4276
rect 15844 4233 15853 4267
rect 15853 4233 15887 4267
rect 15887 4233 15896 4267
rect 15844 4224 15896 4233
rect 16580 4224 16632 4276
rect 19340 4224 19392 4276
rect 5816 4156 5868 4208
rect 6644 4156 6696 4208
rect 8484 4156 8536 4208
rect 2596 4088 2648 4140
rect 2964 4088 3016 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 8300 4088 8352 4140
rect 9588 4088 9640 4140
rect 12624 4156 12676 4208
rect 21272 4224 21324 4276
rect 22836 4267 22888 4276
rect 22836 4233 22845 4267
rect 22845 4233 22879 4267
rect 22879 4233 22888 4267
rect 22836 4224 22888 4233
rect 25136 4267 25188 4276
rect 25136 4233 25145 4267
rect 25145 4233 25179 4267
rect 25179 4233 25188 4267
rect 25136 4224 25188 4233
rect 27160 4224 27212 4276
rect 28816 4224 28868 4276
rect 30564 4224 30616 4276
rect 12440 4131 12492 4140
rect 12440 4097 12449 4131
rect 12449 4097 12483 4131
rect 12483 4097 12492 4131
rect 14188 4131 14240 4140
rect 12440 4088 12492 4097
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 15384 4088 15436 4140
rect 17868 4088 17920 4140
rect 18512 4088 18564 4140
rect 6276 4063 6328 4072
rect 6276 4029 6285 4063
rect 6285 4029 6319 4063
rect 6319 4029 6328 4063
rect 6276 4020 6328 4029
rect 1952 3995 2004 4004
rect 1952 3961 1961 3995
rect 1961 3961 1995 3995
rect 1995 3961 2004 3995
rect 1952 3952 2004 3961
rect 2320 3952 2372 4004
rect 3424 3995 3476 4004
rect 3424 3961 3433 3995
rect 3433 3961 3467 3995
rect 3467 3961 3476 3995
rect 3424 3952 3476 3961
rect 2872 3884 2924 3936
rect 3884 3952 3936 4004
rect 5264 3995 5316 4004
rect 5264 3961 5273 3995
rect 5273 3961 5307 3995
rect 5307 3961 5316 3995
rect 5264 3952 5316 3961
rect 5356 3995 5408 4004
rect 5356 3961 5365 3995
rect 5365 3961 5399 3995
rect 5399 3961 5408 3995
rect 5356 3952 5408 3961
rect 6460 3952 6512 4004
rect 10784 3952 10836 4004
rect 13728 4020 13780 4072
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 7472 3884 7524 3936
rect 10324 3927 10376 3936
rect 10324 3893 10333 3927
rect 10333 3893 10367 3927
rect 10367 3893 10376 3927
rect 10324 3884 10376 3893
rect 11060 3884 11112 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 11980 3884 12032 3936
rect 13820 3952 13872 4004
rect 14740 3952 14792 4004
rect 15016 3952 15068 4004
rect 16120 3995 16172 4004
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 17776 3952 17828 4004
rect 26884 4156 26936 4208
rect 27436 4156 27488 4208
rect 28540 4156 28592 4208
rect 20812 4088 20864 4140
rect 22744 4088 22796 4140
rect 25596 4063 25648 4072
rect 19616 3952 19668 4004
rect 25596 4029 25605 4063
rect 25605 4029 25639 4063
rect 25639 4029 25648 4063
rect 25596 4020 25648 4029
rect 25872 4063 25924 4072
rect 25872 4029 25881 4063
rect 25881 4029 25915 4063
rect 25915 4029 25924 4063
rect 25872 4020 25924 4029
rect 26056 4020 26108 4072
rect 26332 4020 26384 4072
rect 28908 4020 28960 4072
rect 21272 3952 21324 4004
rect 23480 3952 23532 4004
rect 13360 3927 13412 3936
rect 13360 3893 13369 3927
rect 13369 3893 13403 3927
rect 13403 3893 13412 3927
rect 13360 3884 13412 3893
rect 19432 3927 19484 3936
rect 19432 3893 19441 3927
rect 19441 3893 19475 3927
rect 19475 3893 19484 3927
rect 19432 3884 19484 3893
rect 20444 3927 20496 3936
rect 20444 3893 20453 3927
rect 20453 3893 20487 3927
rect 20487 3893 20496 3927
rect 20444 3884 20496 3893
rect 22008 3884 22060 3936
rect 27528 3952 27580 4004
rect 24676 3927 24728 3936
rect 24676 3893 24685 3927
rect 24685 3893 24719 3927
rect 24719 3893 24728 3927
rect 24676 3884 24728 3893
rect 26608 3884 26660 3936
rect 27160 3884 27212 3936
rect 29552 3952 29604 4004
rect 29644 3952 29696 4004
rect 30288 4020 30340 4072
rect 30380 4063 30432 4072
rect 30380 4029 30389 4063
rect 30389 4029 30423 4063
rect 30423 4029 30432 4063
rect 30380 4020 30432 4029
rect 30840 4063 30892 4072
rect 30840 4029 30884 4063
rect 30884 4029 30892 4063
rect 30840 4020 30892 4029
rect 14315 3782 14367 3834
rect 14379 3782 14431 3834
rect 14443 3782 14495 3834
rect 14507 3782 14559 3834
rect 27648 3782 27700 3834
rect 27712 3782 27764 3834
rect 27776 3782 27828 3834
rect 27840 3782 27892 3834
rect 1492 3680 1544 3732
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2596 3680 2648 3732
rect 2964 3723 3016 3732
rect 2964 3689 2973 3723
rect 2973 3689 3007 3723
rect 3007 3689 3016 3723
rect 2964 3680 3016 3689
rect 3424 3723 3476 3732
rect 3424 3689 3433 3723
rect 3433 3689 3467 3723
rect 3467 3689 3476 3723
rect 3424 3680 3476 3689
rect 4252 3723 4304 3732
rect 4252 3689 4261 3723
rect 4261 3689 4295 3723
rect 4295 3689 4304 3723
rect 4252 3680 4304 3689
rect 5172 3680 5224 3732
rect 5448 3723 5500 3732
rect 5448 3689 5457 3723
rect 5457 3689 5491 3723
rect 5491 3689 5500 3723
rect 5448 3680 5500 3689
rect 6828 3723 6880 3732
rect 6828 3689 6837 3723
rect 6837 3689 6871 3723
rect 6871 3689 6880 3723
rect 6828 3680 6880 3689
rect 9772 3680 9824 3732
rect 10324 3680 10376 3732
rect 10876 3680 10928 3732
rect 11704 3680 11756 3732
rect 1676 3655 1728 3664
rect 1676 3621 1685 3655
rect 1685 3621 1719 3655
rect 1719 3621 1728 3655
rect 1676 3612 1728 3621
rect 5264 3612 5316 3664
rect 5816 3612 5868 3664
rect 7472 3655 7524 3664
rect 7472 3621 7481 3655
rect 7481 3621 7515 3655
rect 7515 3621 7524 3655
rect 7472 3612 7524 3621
rect 10232 3655 10284 3664
rect 10232 3621 10241 3655
rect 10241 3621 10275 3655
rect 10275 3621 10284 3655
rect 10232 3612 10284 3621
rect 10784 3612 10836 3664
rect 11980 3612 12032 3664
rect 13452 3680 13504 3732
rect 14188 3680 14240 3732
rect 16764 3723 16816 3732
rect 16764 3689 16773 3723
rect 16773 3689 16807 3723
rect 16807 3689 16816 3723
rect 16764 3680 16816 3689
rect 13360 3612 13412 3664
rect 14740 3612 14792 3664
rect 16120 3612 16172 3664
rect 17776 3680 17828 3732
rect 18512 3680 18564 3732
rect 20720 3723 20772 3732
rect 20720 3689 20729 3723
rect 20729 3689 20763 3723
rect 20763 3689 20772 3723
rect 20720 3680 20772 3689
rect 21272 3723 21324 3732
rect 21272 3689 21281 3723
rect 21281 3689 21315 3723
rect 21315 3689 21324 3723
rect 21272 3680 21324 3689
rect 22744 3723 22796 3732
rect 22744 3689 22753 3723
rect 22753 3689 22787 3723
rect 22787 3689 22796 3723
rect 22744 3680 22796 3689
rect 26056 3680 26108 3732
rect 27436 3680 27488 3732
rect 29828 3680 29880 3732
rect 30472 3723 30524 3732
rect 30472 3689 30481 3723
rect 30481 3689 30515 3723
rect 30515 3689 30524 3723
rect 30472 3680 30524 3689
rect 17224 3655 17276 3664
rect 17224 3621 17233 3655
rect 17233 3621 17267 3655
rect 17267 3621 17276 3655
rect 17224 3612 17276 3621
rect 19340 3612 19392 3664
rect 19984 3655 20036 3664
rect 19984 3621 19993 3655
rect 19993 3621 20027 3655
rect 20027 3621 20036 3655
rect 19984 3612 20036 3621
rect 22008 3612 22060 3664
rect 25596 3612 25648 3664
rect 26608 3612 26660 3664
rect 4620 3587 4672 3596
rect 4620 3553 4638 3587
rect 4638 3553 4672 3587
rect 4620 3544 4672 3553
rect 5632 3544 5684 3596
rect 9496 3544 9548 3596
rect 11612 3544 11664 3596
rect 12440 3587 12492 3596
rect 12440 3553 12449 3587
rect 12449 3553 12483 3587
rect 12483 3553 12492 3587
rect 12440 3544 12492 3553
rect 14188 3587 14240 3596
rect 14188 3553 14232 3587
rect 14232 3553 14240 3587
rect 15292 3587 15344 3596
rect 14188 3544 14240 3553
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 23296 3587 23348 3596
rect 23296 3553 23340 3587
rect 23340 3553 23348 3587
rect 23296 3544 23348 3553
rect 24676 3544 24728 3596
rect 25872 3544 25924 3596
rect 28172 3612 28224 3664
rect 29000 3612 29052 3664
rect 29736 3544 29788 3596
rect 31116 3544 31168 3596
rect 2320 3476 2372 3528
rect 8024 3519 8076 3528
rect 2688 3408 2740 3460
rect 3424 3408 3476 3460
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 8392 3408 8444 3460
rect 9220 3408 9272 3460
rect 4160 3340 4212 3392
rect 6460 3383 6512 3392
rect 6460 3349 6469 3383
rect 6469 3349 6503 3383
rect 6503 3349 6512 3383
rect 6460 3340 6512 3349
rect 11152 3340 11204 3392
rect 12256 3408 12308 3460
rect 12440 3408 12492 3460
rect 14096 3476 14148 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 18604 3476 18656 3528
rect 20628 3476 20680 3528
rect 22100 3476 22152 3528
rect 26240 3476 26292 3528
rect 26516 3519 26568 3528
rect 26516 3485 26525 3519
rect 26525 3485 26559 3519
rect 26559 3485 26568 3519
rect 26516 3476 26568 3485
rect 27988 3476 28040 3528
rect 17776 3408 17828 3460
rect 22376 3451 22428 3460
rect 22376 3417 22385 3451
rect 22385 3417 22419 3451
rect 22419 3417 22428 3451
rect 22376 3408 22428 3417
rect 28908 3451 28960 3460
rect 28908 3417 28917 3451
rect 28917 3417 28951 3451
rect 28951 3417 28960 3451
rect 28908 3408 28960 3417
rect 14004 3383 14056 3392
rect 14004 3349 14013 3383
rect 14013 3349 14047 3383
rect 14047 3349 14056 3383
rect 14004 3340 14056 3349
rect 15016 3383 15068 3392
rect 15016 3349 15025 3383
rect 15025 3349 15059 3383
rect 15059 3349 15068 3383
rect 15016 3340 15068 3349
rect 15200 3340 15252 3392
rect 19800 3340 19852 3392
rect 27804 3340 27856 3392
rect 29552 3383 29604 3392
rect 29552 3349 29561 3383
rect 29561 3349 29595 3383
rect 29595 3349 29604 3383
rect 29552 3340 29604 3349
rect 7648 3238 7700 3290
rect 7712 3238 7764 3290
rect 7776 3238 7828 3290
rect 7840 3238 7892 3290
rect 20982 3238 21034 3290
rect 21046 3238 21098 3290
rect 21110 3238 21162 3290
rect 21174 3238 21226 3290
rect 34315 3238 34367 3290
rect 34379 3238 34431 3290
rect 34443 3238 34495 3290
rect 34507 3238 34559 3290
rect 2872 3179 2924 3188
rect 2872 3145 2881 3179
rect 2881 3145 2915 3179
rect 2915 3145 2924 3179
rect 2872 3136 2924 3145
rect 4252 3136 4304 3188
rect 5908 3136 5960 3188
rect 8392 3136 8444 3188
rect 10784 3136 10836 3188
rect 11612 3136 11664 3188
rect 13360 3179 13412 3188
rect 13360 3145 13369 3179
rect 13369 3145 13403 3179
rect 13403 3145 13412 3179
rect 13360 3136 13412 3145
rect 14188 3136 14240 3188
rect 14924 3136 14976 3188
rect 15292 3136 15344 3188
rect 17224 3136 17276 3188
rect 17776 3179 17828 3188
rect 17776 3145 17785 3179
rect 17785 3145 17819 3179
rect 17819 3145 17828 3179
rect 17776 3136 17828 3145
rect 18604 3179 18656 3188
rect 18604 3145 18613 3179
rect 18613 3145 18647 3179
rect 18647 3145 18656 3179
rect 18604 3136 18656 3145
rect 19340 3136 19392 3188
rect 22008 3136 22060 3188
rect 26516 3136 26568 3188
rect 27528 3136 27580 3188
rect 27804 3136 27856 3188
rect 27988 3179 28040 3188
rect 27988 3145 27997 3179
rect 27997 3145 28031 3179
rect 28031 3145 28040 3179
rect 27988 3136 28040 3145
rect 29000 3179 29052 3188
rect 29000 3145 29009 3179
rect 29009 3145 29043 3179
rect 29043 3145 29052 3179
rect 29000 3136 29052 3145
rect 29828 3136 29880 3188
rect 31116 3136 31168 3188
rect 4068 3068 4120 3120
rect 4620 3068 4672 3120
rect 13636 3068 13688 3120
rect 15016 3068 15068 3120
rect 16120 3111 16172 3120
rect 16120 3077 16129 3111
rect 16129 3077 16163 3111
rect 16163 3077 16172 3111
rect 16120 3068 16172 3077
rect 21916 3111 21968 3120
rect 21916 3077 21925 3111
rect 21925 3077 21959 3111
rect 21959 3077 21968 3111
rect 21916 3068 21968 3077
rect 26608 3111 26660 3120
rect 26608 3077 26617 3111
rect 26617 3077 26651 3111
rect 26651 3077 26660 3111
rect 26608 3068 26660 3077
rect 29736 3111 29788 3120
rect 29736 3077 29745 3111
rect 29745 3077 29779 3111
rect 29779 3077 29788 3111
rect 29736 3068 29788 3077
rect 1676 3000 1728 3052
rect 6460 3000 6512 3052
rect 2872 2864 2924 2916
rect 8024 3000 8076 3052
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 11796 3043 11848 3052
rect 8944 2975 8996 2984
rect 8944 2941 8953 2975
rect 8953 2941 8987 2975
rect 8987 2941 8996 2975
rect 8944 2932 8996 2941
rect 9496 2975 9548 2984
rect 9496 2941 9505 2975
rect 9505 2941 9539 2975
rect 9539 2941 9548 2975
rect 9496 2932 9548 2941
rect 11796 3009 11805 3043
rect 11805 3009 11839 3043
rect 11839 3009 11848 3043
rect 11796 3000 11848 3009
rect 14004 3000 14056 3052
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 20260 3043 20312 3052
rect 20260 3009 20269 3043
rect 20269 3009 20303 3043
rect 20303 3009 20312 3043
rect 20260 3000 20312 3009
rect 22376 3000 22428 3052
rect 16672 2975 16724 2984
rect 9772 2907 9824 2916
rect 9772 2873 9781 2907
rect 9781 2873 9815 2907
rect 9815 2873 9824 2907
rect 9772 2864 9824 2873
rect 16672 2941 16690 2975
rect 16690 2941 16724 2975
rect 16672 2932 16724 2941
rect 23296 2975 23348 2984
rect 13544 2864 13596 2916
rect 13728 2864 13780 2916
rect 15200 2907 15252 2916
rect 15200 2873 15209 2907
rect 15209 2873 15243 2907
rect 15243 2873 15252 2907
rect 15200 2864 15252 2873
rect 7104 2796 7156 2848
rect 7472 2796 7524 2848
rect 8300 2796 8352 2848
rect 11060 2796 11112 2848
rect 12716 2796 12768 2848
rect 23296 2941 23305 2975
rect 23305 2941 23339 2975
rect 23339 2941 23348 2975
rect 23296 2932 23348 2941
rect 27068 2975 27120 2984
rect 27068 2941 27112 2975
rect 27112 2941 27120 2975
rect 27068 2932 27120 2941
rect 28080 2975 28132 2984
rect 28080 2941 28089 2975
rect 28089 2941 28123 2975
rect 28123 2941 28132 2975
rect 28080 2932 28132 2941
rect 29552 2975 29604 2984
rect 29552 2941 29561 2975
rect 29561 2941 29595 2975
rect 29595 2941 29604 2975
rect 29552 2932 29604 2941
rect 19340 2864 19392 2916
rect 16580 2796 16632 2848
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 19156 2796 19208 2805
rect 21824 2864 21876 2916
rect 28264 2839 28316 2848
rect 28264 2805 28273 2839
rect 28273 2805 28307 2839
rect 28307 2805 28316 2839
rect 28264 2796 28316 2805
rect 14315 2694 14367 2746
rect 14379 2694 14431 2746
rect 14443 2694 14495 2746
rect 14507 2694 14559 2746
rect 27648 2694 27700 2746
rect 27712 2694 27764 2746
rect 27776 2694 27828 2746
rect 27840 2694 27892 2746
rect 1492 2592 1544 2644
rect 2688 2592 2740 2644
rect 3056 2635 3108 2644
rect 3056 2601 3065 2635
rect 3065 2601 3099 2635
rect 3099 2601 3108 2635
rect 3056 2592 3108 2601
rect 4068 2592 4120 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 5632 2592 5684 2644
rect 2044 2499 2096 2508
rect 2044 2465 2053 2499
rect 2053 2465 2087 2499
rect 2087 2465 2096 2499
rect 2044 2456 2096 2465
rect 4804 2456 4856 2508
rect 7104 2592 7156 2644
rect 9588 2635 9640 2644
rect 9588 2601 9597 2635
rect 9597 2601 9631 2635
rect 9631 2601 9640 2635
rect 9588 2592 9640 2601
rect 13728 2635 13780 2644
rect 13728 2601 13737 2635
rect 13737 2601 13771 2635
rect 13771 2601 13780 2635
rect 13728 2592 13780 2601
rect 14004 2592 14056 2644
rect 15108 2635 15160 2644
rect 15108 2601 15117 2635
rect 15117 2601 15151 2635
rect 15151 2601 15160 2635
rect 15108 2592 15160 2601
rect 19432 2635 19484 2644
rect 19432 2601 19441 2635
rect 19441 2601 19475 2635
rect 19475 2601 19484 2635
rect 19432 2592 19484 2601
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 8024 2524 8076 2576
rect 11152 2567 11204 2576
rect 11152 2533 11161 2567
rect 11161 2533 11195 2567
rect 11195 2533 11204 2567
rect 11152 2524 11204 2533
rect 12348 2524 12400 2576
rect 13176 2524 13228 2576
rect 13636 2524 13688 2576
rect 13912 2524 13964 2576
rect 10416 2499 10468 2508
rect 10416 2465 10425 2499
rect 10425 2465 10459 2499
rect 10459 2465 10468 2499
rect 10416 2456 10468 2465
rect 14740 2524 14792 2576
rect 19616 2567 19668 2576
rect 19616 2533 19625 2567
rect 19625 2533 19659 2567
rect 19659 2533 19668 2567
rect 19616 2524 19668 2533
rect 20720 2592 20772 2644
rect 22100 2635 22152 2644
rect 22100 2601 22109 2635
rect 22109 2601 22143 2635
rect 22143 2601 22152 2635
rect 22100 2592 22152 2601
rect 23388 2592 23440 2644
rect 27988 2592 28040 2644
rect 28724 2635 28776 2644
rect 28724 2601 28733 2635
rect 28733 2601 28767 2635
rect 28767 2601 28776 2635
rect 28724 2592 28776 2601
rect 31576 2635 31628 2644
rect 31576 2601 31585 2635
rect 31585 2601 31619 2635
rect 31619 2601 31628 2635
rect 31576 2592 31628 2601
rect 32772 2635 32824 2644
rect 32772 2601 32781 2635
rect 32781 2601 32815 2635
rect 32815 2601 32824 2635
rect 32772 2592 32824 2601
rect 20260 2567 20312 2576
rect 20260 2533 20269 2567
rect 20269 2533 20303 2567
rect 20303 2533 20312 2567
rect 20260 2524 20312 2533
rect 15476 2499 15528 2508
rect 15476 2465 15520 2499
rect 15520 2465 15528 2499
rect 15476 2456 15528 2465
rect 20812 2456 20864 2508
rect 21732 2456 21784 2508
rect 23296 2456 23348 2508
rect 27620 2499 27672 2508
rect 27620 2465 27638 2499
rect 27638 2465 27672 2499
rect 27620 2456 27672 2465
rect 28540 2499 28592 2508
rect 28540 2465 28549 2499
rect 28549 2465 28583 2499
rect 28583 2465 28592 2499
rect 28540 2456 28592 2465
rect 30288 2499 30340 2508
rect 30288 2465 30297 2499
rect 30297 2465 30331 2499
rect 30331 2465 30340 2499
rect 30288 2456 30340 2465
rect 31392 2499 31444 2508
rect 31392 2465 31401 2499
rect 31401 2465 31435 2499
rect 31435 2465 31444 2499
rect 31392 2456 31444 2465
rect 32588 2499 32640 2508
rect 32588 2465 32597 2499
rect 32597 2465 32631 2499
rect 32631 2465 32640 2499
rect 32588 2456 32640 2465
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 12716 2431 12768 2440
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 14096 2388 14148 2440
rect 15108 2388 15160 2440
rect 8392 2252 8444 2304
rect 10140 2252 10192 2304
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 15200 2252 15252 2304
rect 21732 2295 21784 2304
rect 21732 2261 21741 2295
rect 21741 2261 21775 2295
rect 21775 2261 21784 2295
rect 21732 2252 21784 2261
rect 33048 2388 33100 2440
rect 7648 2150 7700 2202
rect 7712 2150 7764 2202
rect 7776 2150 7828 2202
rect 7840 2150 7892 2202
rect 20982 2150 21034 2202
rect 21046 2150 21098 2202
rect 21110 2150 21162 2202
rect 21174 2150 21226 2202
rect 34315 2150 34367 2202
rect 34379 2150 34431 2202
rect 34443 2150 34495 2202
rect 34507 2150 34559 2202
rect 12440 1844 12492 1896
rect 15384 1844 15436 1896
<< metal2 >>
rect 478 15200 534 16000
rect 1398 15200 1454 16000
rect 3422 15736 3478 15745
rect 3422 15671 3478 15680
rect 492 11665 520 15200
rect 478 11656 534 11665
rect 478 11591 534 11600
rect 1412 8634 1440 15200
rect 3436 13870 3464 15671
rect 15198 15200 15254 16000
rect 16118 15200 16174 16000
rect 17038 15200 17094 16000
rect 17958 15200 18014 16000
rect 18878 15200 18934 16000
rect 19798 15200 19854 16000
rect 27158 15200 27214 16000
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 14289 13628 14585 13648
rect 14345 13626 14369 13628
rect 14425 13626 14449 13628
rect 14505 13626 14529 13628
rect 14367 13574 14369 13626
rect 14431 13574 14443 13626
rect 14505 13574 14507 13626
rect 14345 13572 14369 13574
rect 14425 13572 14449 13574
rect 14505 13572 14529 13574
rect 14289 13552 14585 13572
rect 7622 13084 7918 13104
rect 7678 13082 7702 13084
rect 7758 13082 7782 13084
rect 7838 13082 7862 13084
rect 7700 13030 7702 13082
rect 7764 13030 7776 13082
rect 7838 13030 7840 13082
rect 7678 13028 7702 13030
rect 7758 13028 7782 13030
rect 7838 13028 7862 13030
rect 7622 13008 7918 13028
rect 15212 12646 15240 15200
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 14289 12540 14585 12560
rect 14345 12538 14369 12540
rect 14425 12538 14449 12540
rect 14505 12538 14529 12540
rect 14367 12486 14369 12538
rect 14431 12486 14443 12538
rect 14505 12486 14507 12538
rect 14345 12484 14369 12486
rect 14425 12484 14449 12486
rect 14505 12484 14529 12486
rect 14289 12464 14585 12484
rect 16132 12458 16160 15200
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 15212 12430 16160 12458
rect 7622 11996 7918 12016
rect 7678 11994 7702 11996
rect 7758 11994 7782 11996
rect 7838 11994 7862 11996
rect 7700 11942 7702 11994
rect 7764 11942 7776 11994
rect 7838 11942 7840 11994
rect 7678 11940 7702 11942
rect 7758 11940 7782 11942
rect 7838 11940 7862 11942
rect 7622 11920 7918 11940
rect 15106 11656 15162 11665
rect 15106 11591 15162 11600
rect 14289 11452 14585 11472
rect 14345 11450 14369 11452
rect 14425 11450 14449 11452
rect 14505 11450 14529 11452
rect 14367 11398 14369 11450
rect 14431 11398 14443 11450
rect 14505 11398 14507 11450
rect 14345 11396 14369 11398
rect 14425 11396 14449 11398
rect 14505 11396 14529 11398
rect 14289 11376 14585 11396
rect 7622 10908 7918 10928
rect 7678 10906 7702 10908
rect 7758 10906 7782 10908
rect 7838 10906 7862 10908
rect 7700 10854 7702 10906
rect 7764 10854 7776 10906
rect 7838 10854 7840 10906
rect 7678 10852 7702 10854
rect 7758 10852 7782 10854
rect 7838 10852 7862 10854
rect 7622 10832 7918 10852
rect 14289 10364 14585 10384
rect 14345 10362 14369 10364
rect 14425 10362 14449 10364
rect 14505 10362 14529 10364
rect 14367 10310 14369 10362
rect 14431 10310 14443 10362
rect 14505 10310 14507 10362
rect 14345 10308 14369 10310
rect 14425 10308 14449 10310
rect 14505 10308 14529 10310
rect 1582 10296 1638 10305
rect 14289 10288 14585 10308
rect 1582 10231 1638 10240
rect 1596 9178 1624 10231
rect 7622 9820 7918 9840
rect 7678 9818 7702 9820
rect 7758 9818 7782 9820
rect 7838 9818 7862 9820
rect 7700 9766 7702 9818
rect 7764 9766 7776 9818
rect 7838 9766 7840 9818
rect 7678 9764 7702 9766
rect 7758 9764 7782 9766
rect 7838 9764 7862 9766
rect 7622 9744 7918 9764
rect 14289 9276 14585 9296
rect 14345 9274 14369 9276
rect 14425 9274 14449 9276
rect 14505 9274 14529 9276
rect 14367 9222 14369 9274
rect 14431 9222 14443 9274
rect 14505 9222 14507 9274
rect 14345 9220 14369 9222
rect 14425 9220 14449 9222
rect 14505 9220 14529 9222
rect 14289 9200 14585 9220
rect 1584 9172 1636 9178
rect 1584 9114 1636 9120
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1400 8628 1452 8634
rect 1400 8570 1452 8576
rect 1596 8090 1624 8871
rect 1964 8401 1992 8978
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 2318 8528 2374 8537
rect 2318 8463 2320 8472
rect 2372 8463 2374 8472
rect 2320 8434 2372 8440
rect 1950 8392 2006 8401
rect 1950 8327 1952 8336
rect 2004 8327 2006 8336
rect 1952 8298 2004 8304
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 1860 7948 1912 7954
rect 1860 7890 1912 7896
rect 1582 7576 1638 7585
rect 1872 7546 1900 7890
rect 5276 7750 5304 7958
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 1582 7511 1638 7520
rect 1860 7540 1912 7546
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 18 3768 74 3777
rect 18 3703 74 3712
rect 32 800 60 3703
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 952 800 980 2751
rect 18 0 74 800
rect 938 0 994 800
rect 1412 785 1440 6598
rect 1504 3738 1532 7142
rect 1596 6458 1624 7511
rect 1860 7482 1912 7488
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 2044 6112 2096 6118
rect 2042 6080 2044 6089
rect 2096 6080 2098 6089
rect 2042 6015 2098 6024
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 1676 5568 1728 5574
rect 1676 5510 1728 5516
rect 1688 5098 1716 5510
rect 2148 5370 2176 5782
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 1676 5092 1728 5098
rect 1676 5034 1728 5040
rect 1688 4758 1716 5034
rect 2042 4992 2098 5001
rect 2042 4927 2098 4936
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1688 4282 1716 4694
rect 1952 4480 2004 4486
rect 1952 4422 2004 4428
rect 1676 4276 1728 4282
rect 1676 4218 1728 4224
rect 1964 4010 1992 4422
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 2056 3890 2084 4927
rect 1964 3862 2084 3890
rect 1492 3732 1544 3738
rect 1492 3674 1544 3680
rect 1504 2650 1532 3674
rect 1676 3664 1728 3670
rect 1676 3606 1728 3612
rect 1688 3058 1716 3606
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1964 2530 1992 3862
rect 2240 3754 2268 7482
rect 5276 7342 5304 7686
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 6104 7206 6132 7890
rect 5080 7200 5132 7206
rect 5080 7142 5132 7148
rect 6092 7200 6144 7206
rect 6092 7142 6144 7148
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2332 6458 2360 6802
rect 4160 6792 4212 6798
rect 4158 6760 4160 6769
rect 4212 6760 4214 6769
rect 4158 6695 4214 6704
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2332 4010 2360 6394
rect 4816 6254 4844 6666
rect 5092 6322 5120 7142
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5264 6860 5316 6866
rect 5184 6820 5264 6848
rect 5184 6662 5212 6820
rect 5264 6802 5316 6808
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5184 6254 5212 6598
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 5172 6248 5224 6254
rect 5172 6190 5224 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2780 5704 2832 5710
rect 2502 5672 2558 5681
rect 2780 5646 2832 5652
rect 2502 5607 2558 5616
rect 2596 5636 2648 5642
rect 2516 4622 2544 5607
rect 2596 5578 2648 5584
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 2056 3726 2268 3754
rect 2056 3369 2084 3726
rect 2332 3534 2360 3946
rect 2516 3738 2544 4558
rect 2608 4146 2636 5578
rect 2792 5234 2820 5646
rect 3330 5400 3386 5409
rect 3330 5335 3332 5344
rect 3384 5335 3386 5344
rect 3332 5306 3384 5312
rect 3882 5264 3938 5273
rect 2780 5228 2832 5234
rect 3882 5199 3884 5208
rect 2780 5170 2832 5176
rect 3936 5199 3938 5208
rect 3884 5170 3936 5176
rect 2792 4826 2820 5170
rect 3700 5160 3752 5166
rect 3700 5102 3752 5108
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2608 3738 2636 4082
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2688 3460 2740 3466
rect 2688 3402 2740 3408
rect 2042 3360 2098 3369
rect 2042 3295 2098 3304
rect 1872 2502 1992 2530
rect 2056 2514 2084 3295
rect 2700 2650 2728 3402
rect 2884 3194 2912 3878
rect 2976 3738 3004 4082
rect 3424 4004 3476 4010
rect 3424 3946 3476 3952
rect 3436 3738 3464 3946
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3436 3466 3464 3674
rect 3424 3460 3476 3466
rect 3424 3402 3476 3408
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 2884 2922 2912 3130
rect 2872 2916 2924 2922
rect 2872 2858 2924 2864
rect 3054 2816 3110 2825
rect 3054 2751 3110 2760
rect 3068 2650 3096 2751
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 3056 2644 3108 2650
rect 3056 2586 3108 2592
rect 2044 2508 2096 2514
rect 1872 800 1900 2502
rect 2044 2450 2096 2456
rect 3516 2440 3568 2446
rect 3514 2408 3516 2417
rect 3568 2408 3570 2417
rect 3514 2343 3570 2352
rect 2778 2000 2834 2009
rect 2778 1935 2834 1944
rect 2792 800 2820 1935
rect 3712 800 3740 5102
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3896 4010 3924 4422
rect 3884 4004 3936 4010
rect 3884 3946 3936 3952
rect 4080 3584 4108 6122
rect 4344 6112 4396 6118
rect 4344 6054 4396 6060
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4356 5710 4384 6054
rect 4344 5704 4396 5710
rect 4540 5681 4568 6054
rect 4344 5646 4396 5652
rect 4526 5672 4582 5681
rect 4526 5607 4582 5616
rect 4816 5166 4844 6190
rect 5184 5574 5212 6190
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5184 5166 5212 5510
rect 5552 5409 5580 6938
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5828 5710 5856 6190
rect 5816 5704 5868 5710
rect 5816 5646 5868 5652
rect 5538 5400 5594 5409
rect 5538 5335 5594 5344
rect 5828 5166 5856 5646
rect 4804 5160 4856 5166
rect 4804 5102 4856 5108
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5448 5160 5500 5166
rect 5448 5102 5500 5108
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 4160 5092 4212 5098
rect 4212 5052 4292 5080
rect 4160 5034 4212 5040
rect 4264 4690 4292 5052
rect 4816 4826 4844 5102
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5184 4758 5212 5102
rect 5172 4752 5224 4758
rect 5172 4694 5224 4700
rect 4252 4684 4304 4690
rect 4252 4626 4304 4632
rect 4264 3738 4292 4626
rect 4710 3904 4766 3913
rect 4710 3839 4766 3848
rect 4252 3732 4304 3738
rect 4252 3674 4304 3680
rect 4620 3596 4672 3602
rect 4080 3556 4292 3584
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4080 2650 4108 3062
rect 4172 2961 4200 3334
rect 4264 3194 4292 3556
rect 4620 3538 4672 3544
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4632 3126 4660 3538
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4158 2952 4214 2961
rect 4158 2887 4214 2896
rect 4342 2952 4398 2961
rect 4724 2938 4752 3839
rect 5184 3738 5212 4694
rect 5354 4584 5410 4593
rect 5354 4519 5410 4528
rect 5262 4040 5318 4049
rect 5368 4010 5396 4519
rect 5460 4282 5488 5102
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5262 3975 5264 3984
rect 5316 3975 5318 3984
rect 5356 4004 5408 4010
rect 5264 3946 5316 3952
rect 5356 3946 5408 3952
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5276 3670 5304 3946
rect 5460 3738 5488 4218
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5644 3602 5672 4966
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5736 4690 5764 4762
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5828 3670 5856 4150
rect 5816 3664 5868 3670
rect 5816 3606 5868 3612
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5538 3088 5594 3097
rect 5538 3023 5594 3032
rect 4342 2887 4398 2896
rect 4632 2910 4752 2938
rect 4356 2650 4384 2887
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4344 2644 4396 2650
rect 4344 2586 4396 2592
rect 4632 800 4660 2910
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 4816 2310 4844 2450
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4816 1737 4844 2246
rect 4802 1728 4858 1737
rect 4802 1663 4858 1672
rect 5552 800 5580 3023
rect 5644 2650 5672 3538
rect 5828 3176 5856 3606
rect 5908 3188 5960 3194
rect 5828 3148 5908 3176
rect 5908 3130 5960 3136
rect 5632 2644 5684 2650
rect 5632 2586 5684 2592
rect 6104 2145 6132 7142
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6196 6322 6224 6802
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6196 5953 6224 6258
rect 6182 5944 6238 5953
rect 6182 5879 6238 5888
rect 6288 5574 6316 6802
rect 6472 6730 6500 8774
rect 6564 8362 6592 8978
rect 15120 8945 15148 11591
rect 15106 8936 15162 8945
rect 15106 8871 15162 8880
rect 7622 8732 7918 8752
rect 7678 8730 7702 8732
rect 7758 8730 7782 8732
rect 7838 8730 7862 8732
rect 7700 8678 7702 8730
rect 7764 8678 7776 8730
rect 7838 8678 7840 8730
rect 7678 8676 7702 8678
rect 7758 8676 7782 8678
rect 7838 8676 7862 8678
rect 7622 8656 7918 8676
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7102 8528 7158 8537
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 7449 6592 8298
rect 6736 7812 6788 7818
rect 6736 7754 6788 7760
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6550 7440 6606 7449
rect 6550 7375 6606 7384
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 6458 6500 6666
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6472 6254 6500 6394
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 5778 6500 6190
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 4729 6316 5510
rect 6564 5386 6592 7142
rect 6472 5358 6592 5386
rect 6472 5030 6500 5358
rect 6552 5296 6604 5302
rect 6552 5238 6604 5244
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 6274 4720 6330 4729
rect 6274 4655 6330 4664
rect 6288 4078 6316 4655
rect 6472 4282 6500 4966
rect 6564 4690 6592 5238
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6472 4010 6500 4218
rect 6656 4214 6684 7686
rect 6748 4622 6776 7754
rect 6932 7426 6960 8502
rect 7102 8463 7158 8472
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 7024 7546 7052 7958
rect 7116 7886 7144 8463
rect 13910 8392 13966 8401
rect 7196 8356 7248 8362
rect 13910 8327 13966 8336
rect 7196 8298 7248 8304
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 6932 7398 7052 7426
rect 6828 7336 6880 7342
rect 6826 7304 6828 7313
rect 6880 7304 6882 7313
rect 6826 7239 6882 7248
rect 6920 7268 6972 7274
rect 6920 7210 6972 7216
rect 6932 6866 6960 7210
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6322 6960 6598
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6932 5794 6960 6122
rect 6840 5778 6960 5794
rect 6840 5772 6972 5778
rect 6840 5766 6920 5772
rect 6840 5370 6868 5766
rect 6920 5714 6972 5720
rect 6920 5636 6972 5642
rect 6920 5578 6972 5584
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6932 5234 6960 5578
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6828 4820 6880 4826
rect 6932 4808 6960 5170
rect 7024 4978 7052 7398
rect 7116 6730 7144 7822
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 7024 4950 7144 4978
rect 7012 4820 7064 4826
rect 6932 4780 7012 4808
rect 6828 4762 6880 4768
rect 7012 4762 7064 4768
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6840 4146 6868 4762
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6460 4004 6512 4010
rect 6460 3946 6512 3952
rect 6840 3738 6868 4082
rect 7116 4049 7144 4950
rect 7102 4040 7158 4049
rect 7102 3975 7158 3984
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6472 3058 6500 3334
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7104 2848 7156 2854
rect 6458 2816 6514 2825
rect 7104 2790 7156 2796
rect 6458 2751 6514 2760
rect 6090 2136 6146 2145
rect 6090 2071 6146 2080
rect 6104 1601 6132 2071
rect 6090 1592 6146 1601
rect 6090 1527 6146 1536
rect 6472 800 6500 2751
rect 7116 2650 7144 2790
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7208 1737 7236 8298
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 7622 7644 7918 7664
rect 7678 7642 7702 7644
rect 7758 7642 7782 7644
rect 7838 7642 7862 7644
rect 7700 7590 7702 7642
rect 7764 7590 7776 7642
rect 7838 7590 7840 7642
rect 7678 7588 7702 7590
rect 7758 7588 7782 7590
rect 7838 7588 7862 7590
rect 7622 7568 7918 7588
rect 13084 7336 13136 7342
rect 8206 7304 8262 7313
rect 13084 7278 13136 7284
rect 13542 7304 13598 7313
rect 8206 7239 8262 7248
rect 8220 7206 8248 7239
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 9128 7200 9180 7206
rect 9128 7142 9180 7148
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 5914 7420 6802
rect 7564 6792 7616 6798
rect 7562 6760 7564 6769
rect 7616 6760 7618 6769
rect 7484 6718 7562 6746
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5846 7512 6718
rect 7562 6695 7618 6704
rect 7622 6556 7918 6576
rect 7678 6554 7702 6556
rect 7758 6554 7782 6556
rect 7838 6554 7862 6556
rect 7700 6502 7702 6554
rect 7764 6502 7776 6554
rect 7838 6502 7840 6554
rect 7678 6500 7702 6502
rect 7758 6500 7782 6502
rect 7838 6500 7862 6502
rect 7622 6480 7918 6500
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7562 6352 7618 6361
rect 7562 6287 7618 6296
rect 7576 6254 7604 6287
rect 8036 6254 8064 6394
rect 8220 6390 8248 7142
rect 8772 6458 8800 7142
rect 9140 6905 9168 7142
rect 11980 6928 12032 6934
rect 9126 6896 9182 6905
rect 9126 6831 9182 6840
rect 11886 6896 11942 6905
rect 11980 6870 12032 6876
rect 12070 6896 12126 6905
rect 11886 6831 11942 6840
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 7564 6248 7616 6254
rect 7564 6190 7616 6196
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8300 6248 8352 6254
rect 8300 6190 8352 6196
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7380 5772 7432 5778
rect 7380 5714 7432 5720
rect 7286 4720 7342 4729
rect 7392 4706 7420 5714
rect 8036 5710 8064 6190
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 7622 5468 7918 5488
rect 7678 5466 7702 5468
rect 7758 5466 7782 5468
rect 7838 5466 7862 5468
rect 7700 5414 7702 5466
rect 7764 5414 7776 5466
rect 7838 5414 7840 5466
rect 7678 5412 7702 5414
rect 7758 5412 7782 5414
rect 7838 5412 7862 5414
rect 7622 5392 7918 5412
rect 8036 5302 8064 5646
rect 8312 5386 8340 6190
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 8576 5772 8628 5778
rect 8576 5714 8628 5720
rect 8392 5568 8444 5574
rect 8392 5510 8444 5516
rect 8220 5370 8340 5386
rect 8208 5364 8340 5370
rect 8260 5358 8340 5364
rect 8208 5306 8260 5312
rect 8024 5296 8076 5302
rect 8024 5238 8076 5244
rect 8220 4758 8248 5306
rect 7342 4678 7420 4706
rect 8208 4752 8260 4758
rect 8208 4694 8260 4700
rect 7286 4655 7288 4664
rect 7340 4655 7342 4664
rect 7288 4626 7340 4632
rect 7622 4380 7918 4400
rect 7678 4378 7702 4380
rect 7758 4378 7782 4380
rect 7838 4378 7862 4380
rect 7700 4326 7702 4378
rect 7764 4326 7776 4378
rect 7838 4326 7840 4378
rect 7678 4324 7702 4326
rect 7758 4324 7782 4326
rect 7838 4324 7862 4326
rect 7622 4304 7918 4324
rect 8220 4282 8248 4694
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8312 4146 8340 4558
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7484 3670 7512 3878
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7378 2952 7434 2961
rect 7378 2887 7434 2896
rect 7194 1728 7250 1737
rect 7194 1663 7250 1672
rect 7392 800 7420 2887
rect 7484 2854 7512 3606
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7622 3292 7918 3312
rect 7678 3290 7702 3292
rect 7758 3290 7782 3292
rect 7838 3290 7862 3292
rect 7700 3238 7702 3290
rect 7764 3238 7776 3290
rect 7838 3238 7840 3290
rect 7678 3236 7702 3238
rect 7758 3236 7782 3238
rect 7838 3236 7862 3238
rect 7622 3216 7918 3236
rect 8036 3058 8064 3470
rect 8404 3466 8432 5510
rect 8588 5030 8616 5714
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8484 4616 8536 4622
rect 8484 4558 8536 4564
rect 8496 4214 8524 4558
rect 8484 4208 8536 4214
rect 8484 4150 8536 4156
rect 8588 3913 8616 4966
rect 8574 3904 8630 3913
rect 8574 3839 8630 3848
rect 8956 3777 8984 4966
rect 9140 4593 9168 6122
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9496 5568 9548 5574
rect 9496 5510 9548 5516
rect 9508 5137 9536 5510
rect 9494 5128 9550 5137
rect 9494 5063 9550 5072
rect 9508 4826 9536 5063
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9126 4584 9182 4593
rect 9126 4519 9182 4528
rect 9600 4146 9628 5850
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 8942 3768 8998 3777
rect 8942 3703 8998 3712
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 8404 3194 8432 3402
rect 8942 3224 8998 3233
rect 8392 3188 8444 3194
rect 8942 3159 8998 3168
rect 8392 3130 8444 3136
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 8036 2582 8064 2994
rect 8956 2990 8984 3159
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 7622 2204 7918 2224
rect 7678 2202 7702 2204
rect 7758 2202 7782 2204
rect 7838 2202 7862 2204
rect 7700 2150 7702 2202
rect 7764 2150 7776 2202
rect 7838 2150 7840 2202
rect 7678 2148 7702 2150
rect 7758 2148 7782 2150
rect 7838 2148 7862 2150
rect 7622 2128 7918 2148
rect 8312 800 8340 2790
rect 8392 2304 8444 2310
rect 8390 2272 8392 2281
rect 8444 2272 8446 2281
rect 8390 2207 8446 2216
rect 9232 800 9260 3402
rect 9508 2990 9536 3538
rect 9692 3058 9720 6734
rect 11900 6662 11928 6831
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10968 6112 11020 6118
rect 11348 6089 11376 6190
rect 11704 6112 11756 6118
rect 10968 6054 11020 6060
rect 11334 6080 11390 6089
rect 10152 5846 10180 6054
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10600 5772 10652 5778
rect 10600 5714 10652 5720
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10336 5166 10364 5714
rect 10612 5370 10640 5714
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10888 5166 10916 5714
rect 10324 5160 10376 5166
rect 10230 5128 10286 5137
rect 9864 5092 9916 5098
rect 10324 5102 10376 5108
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10980 5114 11008 6054
rect 11704 6054 11756 6060
rect 11334 6015 11390 6024
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11256 5166 11284 5714
rect 11244 5160 11296 5166
rect 11242 5128 11244 5137
rect 11296 5128 11298 5137
rect 10230 5063 10286 5072
rect 9864 5034 9916 5040
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9496 2984 9548 2990
rect 9494 2952 9496 2961
rect 9548 2952 9550 2961
rect 9692 2938 9720 2994
rect 9494 2887 9550 2896
rect 9600 2910 9720 2938
rect 9784 2922 9812 3674
rect 9876 3369 9904 5034
rect 10244 3670 10272 5063
rect 10336 4758 10364 5102
rect 10888 5001 10916 5102
rect 10980 5086 11100 5114
rect 10968 5024 11020 5030
rect 10874 4992 10930 5001
rect 10968 4966 11020 4972
rect 10874 4927 10930 4936
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10874 4720 10930 4729
rect 10336 4282 10364 4694
rect 10980 4690 11008 4966
rect 10874 4655 10930 4664
rect 10968 4684 11020 4690
rect 10888 4622 10916 4655
rect 10968 4626 11020 4632
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10784 4004 10836 4010
rect 10784 3946 10836 3952
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3738 10364 3878
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10796 3670 10824 3946
rect 10888 3738 10916 4558
rect 10980 4282 11008 4626
rect 10968 4276 11020 4282
rect 10968 4218 11020 4224
rect 11072 3942 11100 5086
rect 11242 5063 11298 5072
rect 11256 4690 11284 5063
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 11060 3936 11112 3942
rect 11060 3878 11112 3884
rect 10876 3732 10928 3738
rect 10876 3674 10928 3680
rect 10232 3664 10284 3670
rect 10232 3606 10284 3612
rect 10784 3664 10836 3670
rect 10784 3606 10836 3612
rect 9862 3360 9918 3369
rect 9862 3295 9918 3304
rect 10322 3360 10378 3369
rect 10322 3295 10378 3304
rect 10336 3058 10364 3295
rect 10796 3194 10824 3606
rect 11624 3602 11652 4490
rect 11716 3738 11744 6054
rect 11992 5914 12020 6870
rect 12070 6831 12126 6840
rect 12992 6860 13044 6866
rect 12084 6254 12112 6831
rect 12992 6802 13044 6808
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 13004 6186 13032 6802
rect 13096 6458 13124 7278
rect 13176 7268 13228 7274
rect 13542 7239 13598 7248
rect 13176 7210 13228 7216
rect 13188 6934 13216 7210
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13188 6798 13216 6870
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13096 6254 13124 6394
rect 13084 6248 13136 6254
rect 13084 6190 13136 6196
rect 12992 6180 13044 6186
rect 12992 6122 13044 6128
rect 12716 6112 12768 6118
rect 12716 6054 12768 6060
rect 12728 5953 12756 6054
rect 12714 5944 12770 5953
rect 11980 5908 12032 5914
rect 13004 5914 13032 6122
rect 12714 5879 12770 5888
rect 12992 5908 13044 5914
rect 11980 5850 12032 5856
rect 12992 5850 13044 5856
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 12990 5808 13046 5817
rect 12808 5772 12860 5778
rect 12990 5743 12992 5752
rect 12808 5714 12860 5720
rect 13044 5743 13046 5752
rect 12992 5714 13044 5720
rect 12348 5704 12400 5710
rect 12348 5646 12400 5652
rect 12360 5370 12388 5646
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12452 5250 12480 5578
rect 12820 5545 12848 5714
rect 12806 5536 12862 5545
rect 12806 5471 12862 5480
rect 12360 5222 12480 5250
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9772 2916 9824 2922
rect 9600 2650 9628 2910
rect 9772 2858 9824 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 9588 2644 9640 2650
rect 9588 2586 9640 2592
rect 10414 2544 10470 2553
rect 10414 2479 10416 2488
rect 10468 2479 10470 2488
rect 10416 2450 10468 2456
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 800 10180 2246
rect 11072 800 11100 2790
rect 11164 2582 11192 3334
rect 11624 3194 11652 3538
rect 11900 3233 11928 3878
rect 11992 3670 12020 3878
rect 11980 3664 12032 3670
rect 11980 3606 12032 3612
rect 12268 3466 12296 4762
rect 12360 4622 12388 5222
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 12452 4146 12480 5034
rect 12636 4214 12664 5034
rect 12728 4826 12756 5034
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12820 4758 12848 5471
rect 12808 4752 12860 4758
rect 12808 4694 12860 4700
rect 13464 4690 13492 5850
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 12624 4208 12676 4214
rect 12624 4150 12676 4156
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12452 3602 12480 4082
rect 13360 3936 13412 3942
rect 12530 3904 12586 3913
rect 13360 3878 13412 3884
rect 12530 3839 12586 3848
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12360 3466 12480 3482
rect 12256 3460 12308 3466
rect 12256 3402 12308 3408
rect 12360 3460 12492 3466
rect 12360 3454 12440 3460
rect 11886 3224 11942 3233
rect 11612 3188 11664 3194
rect 11886 3159 11942 3168
rect 11612 3130 11664 3136
rect 11794 3088 11850 3097
rect 11794 3023 11796 3032
rect 11848 3023 11850 3032
rect 11796 2994 11848 3000
rect 11152 2576 11204 2582
rect 11152 2518 11204 2524
rect 11900 1329 11928 3159
rect 12360 2582 12388 3454
rect 12440 3402 12492 3408
rect 12348 2576 12400 2582
rect 12348 2518 12400 2524
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12084 2145 12112 2246
rect 12070 2136 12126 2145
rect 12070 2071 12126 2080
rect 12440 1896 12492 1902
rect 12544 1873 12572 3839
rect 13372 3670 13400 3878
rect 13464 3738 13492 4626
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13360 3664 13412 3670
rect 13360 3606 13412 3612
rect 13372 3194 13400 3606
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12716 2848 12768 2854
rect 12716 2790 12768 2796
rect 12728 2446 12756 2790
rect 13176 2576 13228 2582
rect 13372 2564 13400 3130
rect 13556 2922 13584 7239
rect 13648 7206 13676 7890
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13648 7002 13676 7142
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13636 6656 13688 6662
rect 13636 6598 13688 6604
rect 13648 6390 13676 6598
rect 13636 6384 13688 6390
rect 13634 6352 13636 6361
rect 13688 6352 13690 6361
rect 13634 6287 13690 6296
rect 13740 5778 13768 7686
rect 13832 7206 13860 7686
rect 13820 7200 13872 7206
rect 13820 7142 13872 7148
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13636 5092 13688 5098
rect 13636 5034 13688 5040
rect 13648 3126 13676 5034
rect 13740 4554 13768 5714
rect 13832 5710 13860 7142
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13820 4752 13872 4758
rect 13820 4694 13872 4700
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13556 2825 13584 2858
rect 13542 2816 13598 2825
rect 13542 2751 13598 2760
rect 13648 2582 13676 3062
rect 13740 2922 13768 4014
rect 13832 4010 13860 4694
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 13728 2916 13780 2922
rect 13728 2858 13780 2864
rect 13740 2650 13768 2858
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13924 2582 13952 8327
rect 14289 8188 14585 8208
rect 14345 8186 14369 8188
rect 14425 8186 14449 8188
rect 14505 8186 14529 8188
rect 14367 8134 14369 8186
rect 14431 8134 14443 8186
rect 14505 8134 14507 8186
rect 14345 8132 14369 8134
rect 14425 8132 14449 8134
rect 14505 8132 14529 8134
rect 14289 8112 14585 8132
rect 15212 7993 15240 12430
rect 15198 7984 15254 7993
rect 14188 7948 14240 7954
rect 15198 7919 15254 7928
rect 15660 7948 15712 7954
rect 14188 7890 14240 7896
rect 15660 7890 15712 7896
rect 14200 7274 14228 7890
rect 14738 7440 14794 7449
rect 14738 7375 14794 7384
rect 14752 7342 14780 7375
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14188 7268 14240 7274
rect 14188 7210 14240 7216
rect 14289 7100 14585 7120
rect 14345 7098 14369 7100
rect 14425 7098 14449 7100
rect 14505 7098 14529 7100
rect 14367 7046 14369 7098
rect 14431 7046 14443 7098
rect 14505 7046 14507 7098
rect 14345 7044 14369 7046
rect 14425 7044 14449 7046
rect 14505 7044 14529 7046
rect 14289 7024 14585 7044
rect 14752 7002 14780 7278
rect 14832 7268 14884 7274
rect 14832 7210 14884 7216
rect 14844 7177 14872 7210
rect 14924 7200 14976 7206
rect 14830 7168 14886 7177
rect 14924 7142 14976 7148
rect 14830 7103 14886 7112
rect 14740 6996 14792 7002
rect 14740 6938 14792 6944
rect 14936 6798 14964 7142
rect 15672 7002 15700 7890
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 14924 6792 14976 6798
rect 14924 6734 14976 6740
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14108 6254 14136 6598
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14740 6248 14792 6254
rect 14740 6190 14792 6196
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 14108 5166 14136 6190
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14094 4992 14150 5001
rect 14094 4927 14150 4936
rect 14108 4758 14136 4927
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14200 4146 14228 6054
rect 14289 6012 14585 6032
rect 14345 6010 14369 6012
rect 14425 6010 14449 6012
rect 14505 6010 14529 6012
rect 14367 5958 14369 6010
rect 14431 5958 14443 6010
rect 14505 5958 14507 6010
rect 14345 5956 14369 5958
rect 14425 5956 14449 5958
rect 14505 5956 14529 5958
rect 14289 5936 14585 5956
rect 14660 5574 14688 6122
rect 14752 5710 14780 6190
rect 15120 5778 15148 6190
rect 15672 5914 15700 6938
rect 15764 6934 15792 7414
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15842 7168 15898 7177
rect 15842 7103 15898 7112
rect 15752 6928 15804 6934
rect 15752 6870 15804 6876
rect 15764 6361 15792 6870
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 15764 5914 15792 6287
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15108 5772 15160 5778
rect 15160 5732 15240 5760
rect 15108 5714 15160 5720
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14370 5264 14426 5273
rect 14660 5234 14688 5510
rect 14370 5199 14426 5208
rect 14648 5228 14700 5234
rect 14384 5166 14412 5199
rect 14648 5170 14700 5176
rect 15212 5166 15240 5732
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15200 5160 15252 5166
rect 15200 5102 15252 5108
rect 14289 4924 14585 4944
rect 14345 4922 14369 4924
rect 14425 4922 14449 4924
rect 14505 4922 14529 4924
rect 14367 4870 14369 4922
rect 14431 4870 14443 4922
rect 14505 4870 14507 4922
rect 14345 4868 14369 4870
rect 14425 4868 14449 4870
rect 14505 4868 14529 4870
rect 14289 4848 14585 4868
rect 14936 4758 14964 5102
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14200 3738 14228 4082
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 15016 4004 15068 4010
rect 15016 3946 15068 3952
rect 14289 3836 14585 3856
rect 14345 3834 14369 3836
rect 14425 3834 14449 3836
rect 14505 3834 14529 3836
rect 14367 3782 14369 3834
rect 14431 3782 14443 3834
rect 14505 3782 14507 3834
rect 14345 3780 14369 3782
rect 14425 3780 14449 3782
rect 14505 3780 14529 3782
rect 14289 3760 14585 3780
rect 14188 3732 14240 3738
rect 14188 3674 14240 3680
rect 14752 3670 14780 3946
rect 14740 3664 14792 3670
rect 14186 3632 14242 3641
rect 14740 3606 14792 3612
rect 14186 3567 14188 3576
rect 14240 3567 14242 3576
rect 14188 3538 14240 3544
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 14016 3058 14044 3334
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14016 2650 14044 2994
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 13228 2536 13400 2564
rect 13636 2576 13688 2582
rect 13176 2518 13228 2524
rect 13636 2518 13688 2524
rect 13912 2576 13964 2582
rect 13912 2518 13964 2524
rect 14108 2446 14136 3470
rect 14200 3194 14228 3538
rect 15028 3398 15056 3946
rect 15120 3777 15148 4014
rect 15106 3768 15162 3777
rect 15106 3703 15162 3712
rect 15304 3602 15332 4966
rect 15672 4690 15700 5850
rect 15856 5778 15884 7103
rect 15948 6730 15976 7210
rect 16040 6798 16068 7482
rect 16224 7290 16252 12582
rect 16486 11112 16542 11121
rect 16486 11047 16542 11056
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16304 7336 16356 7342
rect 16224 7284 16304 7290
rect 16224 7278 16356 7284
rect 16224 7262 16344 7278
rect 16028 6792 16080 6798
rect 16028 6734 16080 6740
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 5846 15976 6666
rect 16040 6458 16068 6734
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15844 5772 15896 5778
rect 15844 5714 15896 5720
rect 15856 5370 15884 5714
rect 16224 5370 16252 7262
rect 16408 6089 16436 7686
rect 16500 7478 16528 11047
rect 17052 10282 17080 15200
rect 16960 10254 17080 10282
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16488 7472 16540 7478
rect 16488 7414 16540 7420
rect 16592 7410 16620 8026
rect 16684 8022 16712 8230
rect 16672 8016 16724 8022
rect 16672 7958 16724 7964
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16684 7274 16712 7958
rect 16960 7546 16988 10254
rect 17038 10160 17094 10169
rect 17038 10095 17094 10104
rect 17052 8430 17080 10095
rect 17040 8424 17092 8430
rect 17040 8366 17092 8372
rect 17972 8106 18000 15200
rect 18892 11121 18920 15200
rect 19340 13864 19392 13870
rect 19340 13806 19392 13812
rect 18878 11112 18934 11121
rect 18878 11047 18934 11056
rect 19352 8634 19380 13806
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 17880 8090 18000 8106
rect 17868 8084 18000 8090
rect 17920 8078 18000 8084
rect 17868 8026 17920 8032
rect 19812 8022 19840 15200
rect 20956 13084 21252 13104
rect 21012 13082 21036 13084
rect 21092 13082 21116 13084
rect 21172 13082 21196 13084
rect 21034 13030 21036 13082
rect 21098 13030 21110 13082
rect 21172 13030 21174 13082
rect 21012 13028 21036 13030
rect 21092 13028 21116 13030
rect 21172 13028 21196 13030
rect 20956 13008 21252 13028
rect 20956 11996 21252 12016
rect 21012 11994 21036 11996
rect 21092 11994 21116 11996
rect 21172 11994 21196 11996
rect 21034 11942 21036 11994
rect 21098 11942 21110 11994
rect 21172 11942 21174 11994
rect 21012 11940 21036 11942
rect 21092 11940 21116 11942
rect 21172 11940 21196 11942
rect 20956 11920 21252 11940
rect 20956 10908 21252 10928
rect 21012 10906 21036 10908
rect 21092 10906 21116 10908
rect 21172 10906 21196 10908
rect 21034 10854 21036 10906
rect 21098 10854 21110 10906
rect 21172 10854 21174 10906
rect 21012 10852 21036 10854
rect 21092 10852 21116 10854
rect 21172 10852 21196 10854
rect 20956 10832 21252 10852
rect 20956 9820 21252 9840
rect 21012 9818 21036 9820
rect 21092 9818 21116 9820
rect 21172 9818 21196 9820
rect 21034 9766 21036 9818
rect 21098 9766 21110 9818
rect 21172 9766 21174 9818
rect 21012 9764 21036 9766
rect 21092 9764 21116 9766
rect 21172 9764 21196 9766
rect 20956 9744 21252 9764
rect 20956 8732 21252 8752
rect 21012 8730 21036 8732
rect 21092 8730 21116 8732
rect 21172 8730 21196 8732
rect 21034 8678 21036 8730
rect 21098 8678 21110 8730
rect 21172 8678 21174 8730
rect 21012 8676 21036 8678
rect 21092 8676 21116 8678
rect 21172 8676 21196 8678
rect 20956 8656 21252 8676
rect 22560 8288 22612 8294
rect 22560 8230 22612 8236
rect 19800 8016 19852 8022
rect 17130 7984 17186 7993
rect 19800 7958 19852 7964
rect 21272 8016 21324 8022
rect 21272 7958 21324 7964
rect 17130 7919 17132 7928
rect 17184 7919 17186 7928
rect 17132 7890 17184 7896
rect 17144 7546 17172 7890
rect 20812 7880 20864 7886
rect 20812 7822 20864 7828
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 19524 7744 19576 7750
rect 19524 7686 19576 7692
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16948 7268 17000 7274
rect 16948 7210 17000 7216
rect 16960 7041 16988 7210
rect 16946 7032 17002 7041
rect 16946 6967 17002 6976
rect 17144 6866 17172 7482
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17144 6458 17172 6802
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 17328 6361 17356 7686
rect 19536 7410 19564 7686
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 17314 6352 17370 6361
rect 17314 6287 17370 6296
rect 16672 6112 16724 6118
rect 16394 6080 16450 6089
rect 16672 6054 16724 6060
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 16394 6015 16450 6024
rect 16408 5794 16436 6015
rect 16684 5817 16712 6054
rect 16670 5808 16726 5817
rect 16408 5766 16620 5794
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16212 5364 16264 5370
rect 16212 5306 16264 5312
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15856 4758 15884 5170
rect 16224 5166 16252 5306
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 15844 4752 15896 4758
rect 15844 4694 15896 4700
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15672 4282 15700 4626
rect 15856 4282 15884 4694
rect 16592 4622 16620 5766
rect 17328 5778 17356 6054
rect 17420 5778 17448 6598
rect 18064 5778 18092 6598
rect 18524 6458 18552 7278
rect 18972 7200 19024 7206
rect 18972 7142 19024 7148
rect 18984 6798 19012 7142
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18892 6458 18920 6734
rect 18984 6662 19012 6734
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 19432 6656 19484 6662
rect 19432 6598 19484 6604
rect 18512 6452 18564 6458
rect 18512 6394 18564 6400
rect 18880 6452 18932 6458
rect 18880 6394 18932 6400
rect 18524 6254 18552 6394
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 19444 5817 19472 6598
rect 19430 5808 19486 5817
rect 17316 5772 17368 5778
rect 16670 5743 16726 5752
rect 17236 5732 17316 5760
rect 17236 5545 17264 5732
rect 17316 5714 17368 5720
rect 17408 5772 17460 5778
rect 17960 5772 18012 5778
rect 17408 5714 17460 5720
rect 17880 5732 17960 5760
rect 17222 5536 17278 5545
rect 17222 5471 17278 5480
rect 17130 5264 17186 5273
rect 17130 5199 17132 5208
rect 17184 5199 17186 5208
rect 17132 5170 17184 5176
rect 17236 4690 17264 5471
rect 17420 4690 17448 5714
rect 17880 5370 17908 5732
rect 17960 5714 18012 5720
rect 18052 5772 18104 5778
rect 19430 5743 19486 5752
rect 18052 5714 18104 5720
rect 17960 5568 18012 5574
rect 18064 5556 18092 5714
rect 19536 5710 19564 7346
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20720 7336 20772 7342
rect 20720 7278 20772 7284
rect 19706 6896 19762 6905
rect 19706 6831 19762 6840
rect 19720 5778 19748 6831
rect 19996 6662 20024 7278
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20548 6798 20576 7210
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 20442 6352 20498 6361
rect 20442 6287 20498 6296
rect 20456 6254 20484 6287
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 19800 6112 19852 6118
rect 19798 6080 19800 6089
rect 19852 6080 19854 6089
rect 19798 6015 19854 6024
rect 20456 5914 20484 6190
rect 20536 6180 20588 6186
rect 20536 6122 20588 6128
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 18512 5636 18564 5642
rect 18512 5578 18564 5584
rect 18012 5528 18092 5556
rect 17960 5510 18012 5516
rect 17972 5370 18000 5510
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 17776 5024 17828 5030
rect 17776 4966 17828 4972
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17408 4684 17460 4690
rect 17408 4626 17460 4632
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14738 2816 14794 2825
rect 14289 2748 14585 2768
rect 14738 2751 14794 2760
rect 14345 2746 14369 2748
rect 14425 2746 14449 2748
rect 14505 2746 14529 2748
rect 14367 2694 14369 2746
rect 14431 2694 14443 2746
rect 14505 2694 14507 2746
rect 14345 2692 14369 2694
rect 14425 2692 14449 2694
rect 14505 2692 14529 2694
rect 14289 2672 14585 2692
rect 14752 2582 14780 2751
rect 14936 2689 14964 3130
rect 15028 3126 15056 3334
rect 15106 3224 15162 3233
rect 15106 3159 15162 3168
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15120 3058 15148 3159
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 14922 2680 14978 2689
rect 15120 2650 15148 2994
rect 15212 2922 15240 3334
rect 15304 3194 15332 3538
rect 15396 3369 15424 4082
rect 16132 4010 16160 4490
rect 16592 4282 16620 4558
rect 16580 4276 16632 4282
rect 16580 4218 16632 4224
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 16776 3738 16804 4626
rect 17788 4010 17816 4966
rect 17972 4706 18000 5306
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18064 4758 18092 5102
rect 17880 4690 18000 4706
rect 18052 4752 18104 4758
rect 18052 4694 18104 4700
rect 17880 4684 18012 4690
rect 17880 4678 17960 4684
rect 17880 4146 17908 4678
rect 17960 4626 18012 4632
rect 18524 4146 18552 5578
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19248 5024 19300 5030
rect 19248 4966 19300 4972
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 17776 4004 17828 4010
rect 17776 3946 17828 3952
rect 17222 3768 17278 3777
rect 16764 3732 16816 3738
rect 17788 3738 17816 3946
rect 18524 3738 18552 4082
rect 19260 3754 19288 4966
rect 19352 4758 19380 5510
rect 19536 4826 19564 5646
rect 19720 5370 19748 5714
rect 20548 5556 20576 6122
rect 20640 5760 20668 7142
rect 20732 6662 20760 7278
rect 20824 7002 20852 7822
rect 20956 7644 21252 7664
rect 21012 7642 21036 7644
rect 21092 7642 21116 7644
rect 21172 7642 21196 7644
rect 21034 7590 21036 7642
rect 21098 7590 21110 7642
rect 21172 7590 21174 7642
rect 21012 7588 21036 7590
rect 21092 7588 21116 7590
rect 21172 7588 21196 7590
rect 20956 7568 21252 7588
rect 21284 7546 21312 7958
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21272 7540 21324 7546
rect 21272 7482 21324 7488
rect 20812 6996 20864 7002
rect 20812 6938 20864 6944
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 6322 20760 6598
rect 20956 6556 21252 6576
rect 21012 6554 21036 6556
rect 21092 6554 21116 6556
rect 21172 6554 21196 6556
rect 21034 6502 21036 6554
rect 21098 6502 21110 6554
rect 21172 6502 21174 6554
rect 21012 6500 21036 6502
rect 21092 6500 21116 6502
rect 21172 6500 21196 6502
rect 20956 6480 21252 6500
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20812 5908 20864 5914
rect 20812 5850 20864 5856
rect 20720 5772 20772 5778
rect 20640 5732 20720 5760
rect 20720 5714 20772 5720
rect 20628 5568 20680 5574
rect 20548 5528 20628 5556
rect 20628 5510 20680 5516
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19340 4752 19392 4758
rect 19340 4694 19392 4700
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 19352 4282 19380 4694
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19444 3942 19472 4694
rect 19616 4004 19668 4010
rect 19616 3946 19668 3952
rect 19432 3936 19484 3942
rect 19432 3878 19484 3884
rect 17222 3703 17278 3712
rect 17776 3732 17828 3738
rect 16764 3674 16816 3680
rect 17236 3670 17264 3703
rect 17776 3674 17828 3680
rect 18512 3732 18564 3738
rect 19260 3726 19380 3754
rect 18512 3674 18564 3680
rect 19352 3670 19380 3726
rect 16120 3664 16172 3670
rect 16120 3606 16172 3612
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 19340 3664 19392 3670
rect 19340 3606 19392 3612
rect 15474 3496 15530 3505
rect 15474 3431 15530 3440
rect 15382 3360 15438 3369
rect 15382 3295 15438 3304
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15396 3058 15424 3295
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15488 2961 15516 3431
rect 16132 3126 16160 3606
rect 17236 3194 17264 3606
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 17420 3233 17448 3470
rect 17776 3460 17828 3466
rect 17776 3402 17828 3408
rect 17406 3224 17462 3233
rect 17224 3188 17276 3194
rect 17788 3194 17816 3402
rect 18616 3194 18644 3470
rect 19352 3194 19380 3606
rect 17406 3159 17462 3168
rect 17776 3188 17828 3194
rect 17224 3130 17276 3136
rect 17776 3130 17828 3136
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16684 2990 16712 3021
rect 16672 2984 16724 2990
rect 15474 2952 15530 2961
rect 15200 2916 15252 2922
rect 15474 2887 15530 2896
rect 16670 2952 16672 2961
rect 16724 2952 16726 2961
rect 19352 2922 19380 3130
rect 16670 2887 16726 2896
rect 19340 2916 19392 2922
rect 15200 2858 15252 2864
rect 14922 2615 14978 2624
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 15120 2446 15148 2586
rect 15488 2514 15516 2887
rect 16580 2848 16632 2854
rect 16580 2790 16632 2796
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15200 2304 15252 2310
rect 15198 2272 15200 2281
rect 15252 2272 15254 2281
rect 15198 2207 15254 2216
rect 15382 2272 15438 2281
rect 15382 2207 15438 2216
rect 15396 1902 15424 2207
rect 16592 2145 16620 2790
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 16684 2009 16712 2887
rect 19340 2858 19392 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 17038 2680 17094 2689
rect 17038 2615 17094 2624
rect 17052 2530 17080 2615
rect 17314 2544 17370 2553
rect 17052 2502 17314 2530
rect 17314 2479 17370 2488
rect 16670 2000 16726 2009
rect 16670 1935 16726 1944
rect 15384 1896 15436 1902
rect 12440 1838 12492 1844
rect 12530 1864 12586 1873
rect 12452 1601 12480 1838
rect 15384 1838 15436 1844
rect 12530 1799 12586 1808
rect 19168 1737 19196 2790
rect 19444 2650 19472 3878
rect 19432 2644 19484 2650
rect 19432 2586 19484 2592
rect 19628 2582 19656 3946
rect 19720 3641 19748 5306
rect 20640 5250 20668 5510
rect 20718 5264 20774 5273
rect 20640 5222 20718 5250
rect 20718 5199 20774 5208
rect 20732 5166 20760 5199
rect 20824 5166 20852 5850
rect 21284 5846 21312 7482
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 21652 7206 21680 7346
rect 22020 7274 22048 7686
rect 22572 7274 22600 8230
rect 26056 7744 26108 7750
rect 26056 7686 26108 7692
rect 24214 7440 24270 7449
rect 24214 7375 24270 7384
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 22560 7268 22612 7274
rect 22560 7210 22612 7216
rect 21640 7200 21692 7206
rect 21640 7142 21692 7148
rect 21652 6934 21680 7142
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 21364 6860 21416 6866
rect 21364 6802 21416 6808
rect 21916 6860 21968 6866
rect 21916 6802 21968 6808
rect 21376 6730 21404 6802
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21744 6254 21772 6666
rect 21732 6248 21784 6254
rect 21732 6190 21784 6196
rect 21364 6112 21416 6118
rect 21364 6054 21416 6060
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 20956 5468 21252 5488
rect 21012 5466 21036 5468
rect 21092 5466 21116 5468
rect 21172 5466 21196 5468
rect 21034 5414 21036 5466
rect 21098 5414 21110 5466
rect 21172 5414 21174 5466
rect 21012 5412 21036 5414
rect 21092 5412 21116 5414
rect 21172 5412 21196 5414
rect 20956 5392 21252 5412
rect 21284 5370 21312 5782
rect 21272 5364 21324 5370
rect 21272 5306 21324 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 20812 5160 20864 5166
rect 20812 5102 20864 5108
rect 21088 5160 21140 5166
rect 21088 5102 21140 5108
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 3670 20024 4558
rect 20444 3936 20496 3942
rect 20444 3878 20496 3884
rect 19984 3664 20036 3670
rect 19706 3632 19762 3641
rect 19984 3606 20036 3612
rect 19706 3567 19762 3576
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 3058 19840 3334
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20272 2582 20300 2994
rect 19616 2576 19668 2582
rect 19616 2518 19668 2524
rect 20260 2576 20312 2582
rect 20260 2518 20312 2524
rect 20456 2281 20484 3878
rect 20732 3738 20760 4626
rect 20824 4146 20852 4966
rect 21100 4826 21128 5102
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21284 4758 21312 5306
rect 21272 4752 21324 4758
rect 21272 4694 21324 4700
rect 20956 4380 21252 4400
rect 21012 4378 21036 4380
rect 21092 4378 21116 4380
rect 21172 4378 21196 4380
rect 21034 4326 21036 4378
rect 21098 4326 21110 4378
rect 21172 4326 21174 4378
rect 21012 4324 21036 4326
rect 21092 4324 21116 4326
rect 21172 4324 21196 4326
rect 20956 4304 21252 4324
rect 21284 4282 21312 4694
rect 21376 4690 21404 6054
rect 21454 5672 21510 5681
rect 21454 5607 21510 5616
rect 21468 5166 21496 5607
rect 21744 5166 21772 6190
rect 21836 6118 21864 6734
rect 21928 6186 21956 6802
rect 22100 6656 22152 6662
rect 22100 6598 22152 6604
rect 22112 6458 22140 6598
rect 22100 6452 22152 6458
rect 22100 6394 22152 6400
rect 21916 6180 21968 6186
rect 21916 6122 21968 6128
rect 21824 6112 21876 6118
rect 21824 6054 21876 6060
rect 21836 5817 21864 6054
rect 21822 5808 21878 5817
rect 22112 5778 22140 6394
rect 22282 6216 22338 6225
rect 22282 6151 22338 6160
rect 21822 5743 21878 5752
rect 22008 5772 22060 5778
rect 22008 5714 22060 5720
rect 22100 5772 22152 5778
rect 22100 5714 22152 5720
rect 22020 5658 22048 5714
rect 22020 5630 22232 5658
rect 22100 5568 22152 5574
rect 22100 5510 22152 5516
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21732 5160 21784 5166
rect 21732 5102 21784 5108
rect 22112 4758 22140 5510
rect 22204 5370 22232 5630
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 5234 22324 6151
rect 22284 5228 22336 5234
rect 22284 5170 22336 5176
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 22572 4554 22600 7210
rect 24228 7177 24256 7375
rect 26068 7342 26096 7686
rect 27172 7449 27200 15200
rect 27622 13628 27918 13648
rect 27678 13626 27702 13628
rect 27758 13626 27782 13628
rect 27838 13626 27862 13628
rect 27700 13574 27702 13626
rect 27764 13574 27776 13626
rect 27838 13574 27840 13626
rect 27678 13572 27702 13574
rect 27758 13572 27782 13574
rect 27838 13572 27862 13574
rect 27622 13552 27918 13572
rect 34289 13084 34585 13104
rect 34345 13082 34369 13084
rect 34425 13082 34449 13084
rect 34505 13082 34529 13084
rect 34367 13030 34369 13082
rect 34431 13030 34443 13082
rect 34505 13030 34507 13082
rect 34345 13028 34369 13030
rect 34425 13028 34449 13030
rect 34505 13028 34529 13030
rect 34289 13008 34585 13028
rect 27622 12540 27918 12560
rect 27678 12538 27702 12540
rect 27758 12538 27782 12540
rect 27838 12538 27862 12540
rect 27700 12486 27702 12538
rect 27764 12486 27776 12538
rect 27838 12486 27840 12538
rect 27678 12484 27702 12486
rect 27758 12484 27782 12486
rect 27838 12484 27862 12486
rect 27622 12464 27918 12484
rect 34289 11996 34585 12016
rect 34345 11994 34369 11996
rect 34425 11994 34449 11996
rect 34505 11994 34529 11996
rect 34367 11942 34369 11994
rect 34431 11942 34443 11994
rect 34505 11942 34507 11994
rect 34345 11940 34369 11942
rect 34425 11940 34449 11942
rect 34505 11940 34529 11942
rect 34289 11920 34585 11940
rect 27622 11452 27918 11472
rect 27678 11450 27702 11452
rect 27758 11450 27782 11452
rect 27838 11450 27862 11452
rect 27700 11398 27702 11450
rect 27764 11398 27776 11450
rect 27838 11398 27840 11450
rect 27678 11396 27702 11398
rect 27758 11396 27782 11398
rect 27838 11396 27862 11398
rect 27622 11376 27918 11396
rect 34289 10908 34585 10928
rect 34345 10906 34369 10908
rect 34425 10906 34449 10908
rect 34505 10906 34529 10908
rect 34367 10854 34369 10906
rect 34431 10854 34443 10906
rect 34505 10854 34507 10906
rect 34345 10852 34369 10854
rect 34425 10852 34449 10854
rect 34505 10852 34529 10854
rect 34289 10832 34585 10852
rect 27622 10364 27918 10384
rect 27678 10362 27702 10364
rect 27758 10362 27782 10364
rect 27838 10362 27862 10364
rect 27700 10310 27702 10362
rect 27764 10310 27776 10362
rect 27838 10310 27840 10362
rect 27678 10308 27702 10310
rect 27758 10308 27782 10310
rect 27838 10308 27862 10310
rect 27622 10288 27918 10308
rect 34289 9820 34585 9840
rect 34345 9818 34369 9820
rect 34425 9818 34449 9820
rect 34505 9818 34529 9820
rect 34367 9766 34369 9818
rect 34431 9766 34443 9818
rect 34505 9766 34507 9818
rect 34345 9764 34369 9766
rect 34425 9764 34449 9766
rect 34505 9764 34529 9766
rect 34289 9744 34585 9764
rect 27622 9276 27918 9296
rect 27678 9274 27702 9276
rect 27758 9274 27782 9276
rect 27838 9274 27862 9276
rect 27700 9222 27702 9274
rect 27764 9222 27776 9274
rect 27838 9222 27840 9274
rect 27678 9220 27702 9222
rect 27758 9220 27782 9222
rect 27838 9220 27862 9222
rect 27622 9200 27918 9220
rect 28998 8936 29054 8945
rect 28998 8871 29054 8880
rect 35622 8936 35678 8945
rect 35622 8871 35678 8880
rect 27622 8188 27918 8208
rect 27678 8186 27702 8188
rect 27758 8186 27782 8188
rect 27838 8186 27862 8188
rect 27700 8134 27702 8186
rect 27764 8134 27776 8186
rect 27838 8134 27840 8186
rect 27678 8132 27702 8134
rect 27758 8132 27782 8134
rect 27838 8132 27862 8134
rect 27622 8112 27918 8132
rect 28724 8016 28776 8022
rect 28724 7958 28776 7964
rect 28448 7880 28500 7886
rect 28448 7822 28500 7828
rect 28460 7546 28488 7822
rect 28736 7546 28764 7958
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28448 7540 28500 7546
rect 28448 7482 28500 7488
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 27158 7440 27214 7449
rect 27158 7375 27214 7384
rect 25136 7336 25188 7342
rect 25136 7278 25188 7284
rect 25688 7336 25740 7342
rect 25688 7278 25740 7284
rect 26056 7336 26108 7342
rect 26056 7278 26108 7284
rect 26424 7336 26476 7342
rect 26424 7278 26476 7284
rect 24676 7200 24728 7206
rect 24214 7168 24270 7177
rect 24676 7142 24728 7148
rect 24214 7103 24270 7112
rect 24228 6458 24256 7103
rect 24306 7032 24362 7041
rect 24688 7002 24716 7142
rect 24306 6967 24362 6976
rect 24676 6996 24728 7002
rect 24320 6866 24348 6967
rect 24676 6938 24728 6944
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 24216 6452 24268 6458
rect 24216 6394 24268 6400
rect 24228 6254 24256 6394
rect 25148 6254 25176 7278
rect 25700 7002 25728 7278
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25688 6996 25740 7002
rect 25688 6938 25740 6944
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 25136 6248 25188 6254
rect 25136 6190 25188 6196
rect 24124 6180 24176 6186
rect 24124 6122 24176 6128
rect 23848 6112 23900 6118
rect 23848 6054 23900 6060
rect 23860 5846 23888 6054
rect 23848 5840 23900 5846
rect 24136 5817 24164 6122
rect 24860 5840 24912 5846
rect 23848 5782 23900 5788
rect 24122 5808 24178 5817
rect 23860 5681 23888 5782
rect 24860 5782 24912 5788
rect 24122 5743 24124 5752
rect 24176 5743 24178 5752
rect 24124 5714 24176 5720
rect 23846 5672 23902 5681
rect 23846 5607 23902 5616
rect 24136 5370 24164 5714
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24124 5364 24176 5370
rect 24124 5306 24176 5312
rect 24504 5302 24532 5646
rect 24492 5296 24544 5302
rect 24492 5238 24544 5244
rect 23480 5024 23532 5030
rect 23480 4966 23532 4972
rect 23492 4826 23520 4966
rect 23480 4820 23532 4826
rect 23480 4762 23532 4768
rect 24872 4758 24900 5782
rect 25332 5710 25360 6938
rect 25596 6656 25648 6662
rect 25596 6598 25648 6604
rect 25608 6254 25636 6598
rect 26068 6254 26096 7278
rect 26436 6866 26464 7278
rect 26700 7268 26752 7274
rect 26700 7210 26752 7216
rect 26712 6866 26740 7210
rect 27622 7100 27918 7120
rect 27678 7098 27702 7100
rect 27758 7098 27782 7100
rect 27838 7098 27862 7100
rect 27700 7046 27702 7098
rect 27764 7046 27776 7098
rect 27838 7046 27840 7098
rect 27678 7044 27702 7046
rect 27758 7044 27782 7046
rect 27838 7044 27862 7046
rect 27622 7024 27918 7044
rect 28736 7002 28764 7482
rect 28920 7342 28948 7822
rect 29012 7546 29040 8871
rect 34289 8732 34585 8752
rect 34345 8730 34369 8732
rect 34425 8730 34449 8732
rect 34505 8730 34529 8732
rect 34367 8678 34369 8730
rect 34431 8678 34443 8730
rect 34505 8678 34507 8730
rect 34345 8676 34369 8678
rect 34425 8676 34449 8678
rect 34505 8676 34529 8678
rect 34289 8656 34585 8676
rect 35636 8090 35664 8871
rect 35624 8084 35676 8090
rect 35624 8026 35676 8032
rect 35440 7948 35492 7954
rect 35440 7890 35492 7896
rect 34289 7644 34585 7664
rect 34345 7642 34369 7644
rect 34425 7642 34449 7644
rect 34505 7642 34529 7644
rect 34367 7590 34369 7642
rect 34431 7590 34443 7642
rect 34505 7590 34507 7642
rect 34345 7588 34369 7590
rect 34425 7588 34449 7590
rect 34505 7588 34529 7590
rect 34289 7568 34585 7588
rect 29000 7540 29052 7546
rect 29000 7482 29052 7488
rect 33414 7440 33470 7449
rect 33414 7375 33470 7384
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 28724 6996 28776 7002
rect 28724 6938 28776 6944
rect 29184 6928 29236 6934
rect 29184 6870 29236 6876
rect 26424 6860 26476 6866
rect 26424 6802 26476 6808
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26436 6254 26464 6802
rect 26712 6458 26740 6802
rect 27160 6792 27212 6798
rect 27160 6734 27212 6740
rect 26700 6452 26752 6458
rect 26700 6394 26752 6400
rect 25596 6248 25648 6254
rect 25594 6216 25596 6225
rect 26056 6248 26108 6254
rect 25648 6216 25650 6225
rect 26424 6248 26476 6254
rect 26056 6190 26108 6196
rect 26344 6208 26424 6236
rect 25594 6151 25650 6160
rect 25320 5704 25372 5710
rect 25320 5646 25372 5652
rect 25608 5574 25636 6151
rect 26148 6112 26200 6118
rect 26148 6054 26200 6060
rect 25596 5568 25648 5574
rect 25596 5510 25648 5516
rect 25608 5166 25636 5510
rect 25688 5296 25740 5302
rect 25686 5264 25688 5273
rect 25740 5264 25742 5273
rect 25686 5199 25742 5208
rect 25596 5160 25648 5166
rect 25596 5102 25648 5108
rect 25136 4820 25188 4826
rect 25136 4762 25188 4768
rect 22836 4752 22888 4758
rect 22836 4694 22888 4700
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22100 4548 22152 4554
rect 21928 4508 22100 4536
rect 21824 4480 21876 4486
rect 21824 4422 21876 4428
rect 21272 4276 21324 4282
rect 21272 4218 21324 4224
rect 21284 4185 21312 4218
rect 20902 4176 20958 4185
rect 20812 4140 20864 4146
rect 20902 4111 20958 4120
rect 21270 4176 21326 4185
rect 21270 4111 21326 4120
rect 20812 4082 20864 4088
rect 20916 4026 20944 4111
rect 20824 3998 20944 4026
rect 21284 4010 21312 4111
rect 21272 4004 21324 4010
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 20628 3528 20680 3534
rect 20680 3488 20760 3516
rect 20628 3470 20680 3476
rect 20732 2650 20760 3488
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20824 2514 20852 3998
rect 21272 3946 21324 3952
rect 21284 3738 21312 3946
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 20956 3292 21252 3312
rect 21012 3290 21036 3292
rect 21092 3290 21116 3292
rect 21172 3290 21196 3292
rect 21034 3238 21036 3290
rect 21098 3238 21110 3290
rect 21172 3238 21174 3290
rect 21012 3236 21036 3238
rect 21092 3236 21116 3238
rect 21172 3236 21196 3238
rect 20956 3216 21252 3236
rect 21836 2922 21864 4422
rect 21928 3126 21956 4508
rect 22100 4490 22152 4496
rect 22560 4548 22612 4554
rect 22560 4490 22612 4496
rect 22756 4146 22784 4558
rect 22848 4282 22876 4694
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24398 4584 24454 4593
rect 24398 4519 24400 4528
rect 24452 4519 24454 4528
rect 24400 4490 24452 4496
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 22836 4276 22888 4282
rect 22836 4218 22888 4224
rect 22744 4140 22796 4146
rect 22744 4082 22796 4088
rect 22008 3936 22060 3942
rect 22008 3878 22060 3884
rect 22020 3670 22048 3878
rect 22756 3738 22784 4082
rect 23492 4010 23520 4422
rect 23480 4004 23532 4010
rect 23400 3964 23480 3992
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 22008 3664 22060 3670
rect 22008 3606 22060 3612
rect 22020 3194 22048 3606
rect 23296 3596 23348 3602
rect 23296 3538 23348 3544
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21824 2916 21876 2922
rect 21824 2858 21876 2864
rect 22112 2650 22140 3470
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22388 3058 22416 3402
rect 22376 3052 22428 3058
rect 22376 2994 22428 3000
rect 23308 2990 23336 3538
rect 23296 2984 23348 2990
rect 23294 2952 23296 2961
rect 23348 2952 23350 2961
rect 23294 2887 23350 2896
rect 23294 2680 23350 2689
rect 22100 2644 22152 2650
rect 23400 2650 23428 3964
rect 23480 3946 23532 3952
rect 24688 3942 24716 4626
rect 25148 4282 25176 4762
rect 25608 4622 25636 5102
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 25596 4072 25648 4078
rect 25700 4060 25728 5199
rect 26056 5160 26108 5166
rect 26056 5102 26108 5108
rect 26068 4758 26096 5102
rect 26056 4752 26108 4758
rect 26056 4694 26108 4700
rect 25872 4616 25924 4622
rect 25872 4558 25924 4564
rect 25884 4078 25912 4558
rect 26068 4078 26096 4694
rect 25648 4032 25728 4060
rect 25872 4072 25924 4078
rect 25596 4014 25648 4020
rect 25872 4014 25924 4020
rect 26056 4072 26108 4078
rect 26056 4014 26108 4020
rect 24676 3936 24728 3942
rect 24676 3878 24728 3884
rect 24688 3602 24716 3878
rect 25608 3670 25636 4014
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 25884 3602 25912 4014
rect 26068 3738 26096 4014
rect 26056 3732 26108 3738
rect 26056 3674 26108 3680
rect 26160 3618 26188 6054
rect 26344 5778 26372 6208
rect 26424 6190 26476 6196
rect 27172 6118 27200 6734
rect 29196 6390 29224 6870
rect 29840 6798 29868 7278
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 30288 6792 30340 6798
rect 30288 6734 30340 6740
rect 30012 6724 30064 6730
rect 30012 6666 30064 6672
rect 29184 6384 29236 6390
rect 27710 6352 27766 6361
rect 29184 6326 29236 6332
rect 27710 6287 27766 6296
rect 27724 6254 27752 6287
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27988 6248 28040 6254
rect 27988 6190 28040 6196
rect 29276 6248 29328 6254
rect 29276 6190 29328 6196
rect 27344 6180 27396 6186
rect 27344 6122 27396 6128
rect 27160 6112 27212 6118
rect 27160 6054 27212 6060
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26792 5772 26844 5778
rect 26792 5714 26844 5720
rect 26344 5166 26372 5714
rect 26804 5234 26832 5714
rect 26792 5228 26844 5234
rect 26792 5170 26844 5176
rect 26332 5160 26384 5166
rect 26332 5102 26384 5108
rect 26344 4826 26372 5102
rect 26332 4820 26384 4826
rect 26332 4762 26384 4768
rect 26344 4078 26372 4762
rect 27172 4758 27200 6054
rect 27356 5778 27384 6122
rect 27540 5778 27568 6190
rect 27622 6012 27918 6032
rect 27678 6010 27702 6012
rect 27758 6010 27782 6012
rect 27838 6010 27862 6012
rect 27700 5958 27702 6010
rect 27764 5958 27776 6010
rect 27838 5958 27840 6010
rect 27678 5956 27702 5958
rect 27758 5956 27782 5958
rect 27838 5956 27862 5958
rect 27622 5936 27918 5956
rect 27344 5772 27396 5778
rect 27344 5714 27396 5720
rect 27528 5772 27580 5778
rect 27528 5714 27580 5720
rect 27356 5302 27384 5714
rect 27344 5296 27396 5302
rect 27344 5238 27396 5244
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 27160 4752 27212 4758
rect 27160 4694 27212 4700
rect 26884 4616 26936 4622
rect 26884 4558 26936 4564
rect 26896 4214 26924 4558
rect 27066 4448 27122 4457
rect 27066 4383 27122 4392
rect 26884 4208 26936 4214
rect 26606 4176 26662 4185
rect 26884 4150 26936 4156
rect 26606 4111 26662 4120
rect 26332 4072 26384 4078
rect 26332 4014 26384 4020
rect 26620 3942 26648 4111
rect 26608 3936 26660 3942
rect 26608 3878 26660 3884
rect 26620 3670 26648 3878
rect 26608 3664 26660 3670
rect 24676 3596 24728 3602
rect 24676 3538 24728 3544
rect 25872 3596 25924 3602
rect 26160 3590 26280 3618
rect 26608 3606 26660 3612
rect 25872 3538 25924 3544
rect 26252 3534 26280 3590
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 26528 3194 26556 3470
rect 26516 3188 26568 3194
rect 26516 3130 26568 3136
rect 26620 3126 26648 3606
rect 27080 3233 27108 4383
rect 27172 4282 27200 4694
rect 27540 4622 27568 5034
rect 27622 4924 27918 4944
rect 27678 4922 27702 4924
rect 27758 4922 27782 4924
rect 27838 4922 27862 4924
rect 27700 4870 27702 4922
rect 27764 4870 27776 4922
rect 27838 4870 27840 4922
rect 27678 4868 27702 4870
rect 27758 4868 27782 4870
rect 27838 4868 27862 4870
rect 27622 4848 27918 4868
rect 28000 4842 28028 6190
rect 28080 6112 28132 6118
rect 28080 6054 28132 6060
rect 28816 6112 28868 6118
rect 28816 6054 28868 6060
rect 28092 5914 28120 6054
rect 28828 5914 28856 6054
rect 28080 5908 28132 5914
rect 28080 5850 28132 5856
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 28092 5234 28120 5850
rect 28080 5228 28132 5234
rect 28080 5170 28132 5176
rect 28172 5092 28224 5098
rect 28172 5034 28224 5040
rect 28000 4814 28120 4842
rect 27528 4616 27580 4622
rect 27528 4558 27580 4564
rect 27160 4276 27212 4282
rect 27160 4218 27212 4224
rect 27172 3942 27200 4218
rect 27436 4208 27488 4214
rect 27436 4150 27488 4156
rect 27160 3936 27212 3942
rect 27160 3878 27212 3884
rect 27448 3738 27476 4150
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27436 3732 27488 3738
rect 27436 3674 27488 3680
rect 27066 3224 27122 3233
rect 27540 3194 27568 3946
rect 27622 3836 27918 3856
rect 27678 3834 27702 3836
rect 27758 3834 27782 3836
rect 27838 3834 27862 3836
rect 27700 3782 27702 3834
rect 27764 3782 27776 3834
rect 27838 3782 27840 3834
rect 27678 3780 27702 3782
rect 27758 3780 27782 3782
rect 27838 3780 27862 3782
rect 27622 3760 27918 3780
rect 27988 3528 28040 3534
rect 27988 3470 28040 3476
rect 27804 3392 27856 3398
rect 27804 3334 27856 3340
rect 27816 3194 27844 3334
rect 28000 3194 28028 3470
rect 27066 3159 27122 3168
rect 27528 3188 27580 3194
rect 26608 3120 26660 3126
rect 26608 3062 26660 3068
rect 27080 2990 27108 3159
rect 27528 3130 27580 3136
rect 27804 3188 27856 3194
rect 27804 3130 27856 3136
rect 27988 3188 28040 3194
rect 27988 3130 28040 3136
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 27622 2748 27918 2768
rect 27678 2746 27702 2748
rect 27758 2746 27782 2748
rect 27838 2746 27862 2748
rect 27700 2694 27702 2746
rect 27764 2694 27776 2746
rect 27838 2694 27840 2746
rect 27678 2692 27702 2694
rect 27758 2692 27782 2694
rect 27838 2692 27862 2694
rect 27622 2672 27918 2692
rect 28000 2650 28028 3130
rect 28092 2990 28120 4814
rect 28184 4486 28212 5034
rect 28828 5030 28856 5850
rect 29288 5710 29316 6190
rect 30024 6118 30052 6666
rect 30012 6112 30064 6118
rect 30012 6054 30064 6060
rect 29276 5704 29328 5710
rect 29276 5646 29328 5652
rect 28908 5296 28960 5302
rect 28908 5238 28960 5244
rect 28816 5024 28868 5030
rect 28816 4966 28868 4972
rect 28828 4758 28856 4966
rect 28816 4752 28868 4758
rect 28816 4694 28868 4700
rect 28632 4616 28684 4622
rect 28632 4558 28684 4564
rect 28172 4480 28224 4486
rect 28172 4422 28224 4428
rect 28540 4480 28592 4486
rect 28540 4422 28592 4428
rect 28184 3670 28212 4422
rect 28552 4214 28580 4422
rect 28644 4321 28672 4558
rect 28630 4312 28686 4321
rect 28828 4282 28856 4694
rect 28630 4247 28686 4256
rect 28816 4276 28868 4282
rect 28816 4218 28868 4224
rect 28540 4208 28592 4214
rect 28540 4150 28592 4156
rect 28920 4078 28948 5238
rect 30024 5234 30052 6054
rect 30300 5234 30328 6734
rect 33428 6458 33456 7375
rect 35452 7342 35480 7890
rect 35440 7336 35492 7342
rect 35438 7304 35440 7313
rect 35492 7304 35494 7313
rect 35438 7239 35494 7248
rect 34289 6556 34585 6576
rect 34345 6554 34369 6556
rect 34425 6554 34449 6556
rect 34505 6554 34529 6556
rect 34367 6502 34369 6554
rect 34431 6502 34443 6554
rect 34505 6502 34507 6554
rect 34345 6500 34369 6502
rect 34425 6500 34449 6502
rect 34505 6500 34529 6502
rect 34289 6480 34585 6500
rect 33416 6452 33468 6458
rect 33416 6394 33468 6400
rect 33232 6248 33284 6254
rect 33232 6190 33284 6196
rect 34610 6216 34666 6225
rect 30380 5568 30432 5574
rect 30380 5510 30432 5516
rect 30932 5568 30984 5574
rect 30932 5510 30984 5516
rect 30392 5370 30420 5510
rect 30380 5364 30432 5370
rect 30380 5306 30432 5312
rect 29644 5228 29696 5234
rect 29644 5170 29696 5176
rect 30012 5228 30064 5234
rect 30012 5170 30064 5176
rect 30288 5228 30340 5234
rect 30288 5170 30340 5176
rect 29368 5092 29420 5098
rect 29368 5034 29420 5040
rect 29460 5092 29512 5098
rect 29460 5034 29512 5040
rect 29380 4826 29408 5034
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 29472 4690 29500 5034
rect 29460 4684 29512 4690
rect 29460 4626 29512 4632
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 28908 4072 28960 4078
rect 28908 4014 28960 4020
rect 28172 3664 28224 3670
rect 28172 3606 28224 3612
rect 28920 3466 28948 4014
rect 29564 4010 29592 4422
rect 29656 4010 29684 5170
rect 29734 5128 29790 5137
rect 30944 5098 30972 5510
rect 31024 5364 31076 5370
rect 31024 5306 31076 5312
rect 31036 5098 31064 5306
rect 33244 5137 33272 6190
rect 34610 6151 34666 6160
rect 34289 5468 34585 5488
rect 34345 5466 34369 5468
rect 34425 5466 34449 5468
rect 34505 5466 34529 5468
rect 34367 5414 34369 5466
rect 34431 5414 34443 5466
rect 34505 5414 34507 5466
rect 34345 5412 34369 5414
rect 34425 5412 34449 5414
rect 34505 5412 34529 5414
rect 34289 5392 34585 5412
rect 33230 5128 33286 5137
rect 29734 5063 29790 5072
rect 30932 5092 30984 5098
rect 29552 4004 29604 4010
rect 29552 3946 29604 3952
rect 29644 4004 29696 4010
rect 29644 3946 29696 3952
rect 29000 3664 29052 3670
rect 29000 3606 29052 3612
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 29012 3194 29040 3606
rect 29748 3602 29776 5063
rect 30932 5034 30984 5040
rect 31024 5092 31076 5098
rect 33230 5063 33286 5072
rect 31024 5034 31076 5040
rect 30564 5024 30616 5030
rect 30564 4966 30616 4972
rect 29828 4820 29880 4826
rect 29828 4762 29880 4768
rect 29840 3738 29868 4762
rect 30576 4758 30604 4966
rect 30564 4752 30616 4758
rect 30564 4694 30616 4700
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30380 4548 30432 4554
rect 30380 4490 30432 4496
rect 30392 4434 30420 4490
rect 30300 4406 30420 4434
rect 30300 4078 30328 4406
rect 30378 4312 30434 4321
rect 30378 4247 30434 4256
rect 30392 4078 30420 4247
rect 30288 4072 30340 4078
rect 30288 4014 30340 4020
rect 30380 4072 30432 4078
rect 30380 4014 30432 4020
rect 30484 3738 30512 4558
rect 30576 4282 30604 4694
rect 30944 4622 30972 5034
rect 30932 4616 30984 4622
rect 34624 4593 34652 6151
rect 34702 4856 34758 4865
rect 34702 4791 34758 4800
rect 30932 4558 30984 4564
rect 34610 4584 34666 4593
rect 34610 4519 34666 4528
rect 34289 4380 34585 4400
rect 34345 4378 34369 4380
rect 34425 4378 34449 4380
rect 34505 4378 34529 4380
rect 34367 4326 34369 4378
rect 34431 4326 34443 4378
rect 34505 4326 34507 4378
rect 34345 4324 34369 4326
rect 34425 4324 34449 4326
rect 34505 4324 34529 4326
rect 34289 4304 34585 4324
rect 30564 4276 30616 4282
rect 30564 4218 30616 4224
rect 30840 4072 30892 4078
rect 30838 4040 30840 4049
rect 30892 4040 30894 4049
rect 30838 3975 30894 3984
rect 34716 3777 34744 4791
rect 37738 4040 37794 4049
rect 37738 3975 37794 3984
rect 31114 3768 31170 3777
rect 29828 3732 29880 3738
rect 29828 3674 29880 3680
rect 30472 3732 30524 3738
rect 31114 3703 31170 3712
rect 34702 3768 34758 3777
rect 34886 3768 34942 3777
rect 34702 3703 34758 3712
rect 34808 3726 34886 3754
rect 30472 3674 30524 3680
rect 31128 3602 31156 3703
rect 29736 3596 29788 3602
rect 31116 3596 31168 3602
rect 29788 3556 29868 3584
rect 29736 3538 29788 3544
rect 29552 3392 29604 3398
rect 29552 3334 29604 3340
rect 29000 3188 29052 3194
rect 29000 3130 29052 3136
rect 29564 2990 29592 3334
rect 29840 3194 29868 3556
rect 34808 3584 34836 3726
rect 34886 3703 34942 3712
rect 36818 3768 36874 3777
rect 36818 3703 36874 3712
rect 31116 3538 31168 3544
rect 34440 3556 34836 3584
rect 31128 3369 31156 3538
rect 34440 3505 34468 3556
rect 34426 3496 34482 3505
rect 34426 3431 34482 3440
rect 34610 3496 34666 3505
rect 34610 3431 34666 3440
rect 31114 3360 31170 3369
rect 31114 3295 31170 3304
rect 31128 3194 31156 3295
rect 34289 3292 34585 3312
rect 34345 3290 34369 3292
rect 34425 3290 34449 3292
rect 34505 3290 34529 3292
rect 34367 3238 34369 3290
rect 34431 3238 34443 3290
rect 34505 3238 34507 3290
rect 34345 3236 34369 3238
rect 34425 3236 34449 3238
rect 34505 3236 34529 3238
rect 32586 3224 32642 3233
rect 29828 3188 29880 3194
rect 29828 3130 29880 3136
rect 31116 3188 31168 3194
rect 34289 3216 34585 3236
rect 32586 3159 32642 3168
rect 31116 3130 31168 3136
rect 29736 3120 29788 3126
rect 29734 3088 29736 3097
rect 29788 3088 29790 3097
rect 29734 3023 29790 3032
rect 32218 3088 32274 3097
rect 32218 3023 32274 3032
rect 28080 2984 28132 2990
rect 29552 2984 29604 2990
rect 28080 2926 28132 2932
rect 28262 2952 28318 2961
rect 29552 2926 29604 2932
rect 30378 2952 30434 2961
rect 28262 2887 28318 2896
rect 28276 2854 28304 2887
rect 28264 2848 28316 2854
rect 28264 2790 28316 2796
rect 28722 2816 28778 2825
rect 28722 2751 28778 2760
rect 28736 2650 28764 2751
rect 23294 2615 23350 2624
rect 23388 2644 23440 2650
rect 22100 2586 22152 2592
rect 23308 2514 23336 2615
rect 23388 2586 23440 2592
rect 27988 2644 28040 2650
rect 27988 2586 28040 2592
rect 28724 2644 28776 2650
rect 28724 2586 28776 2592
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 21732 2508 21784 2514
rect 21732 2450 21784 2456
rect 23296 2508 23348 2514
rect 23296 2450 23348 2456
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 28540 2508 28592 2514
rect 28540 2450 28592 2456
rect 21744 2310 21772 2450
rect 21732 2304 21784 2310
rect 20442 2272 20498 2281
rect 21730 2272 21732 2281
rect 21784 2272 21786 2281
rect 20442 2207 20498 2216
rect 20456 1737 20484 2207
rect 20956 2204 21252 2224
rect 21730 2207 21786 2216
rect 21012 2202 21036 2204
rect 21092 2202 21116 2204
rect 21172 2202 21196 2204
rect 21034 2150 21036 2202
rect 21098 2150 21110 2202
rect 21172 2150 21174 2202
rect 21012 2148 21036 2150
rect 21092 2148 21116 2150
rect 21172 2148 21196 2150
rect 20956 2128 21252 2148
rect 23308 2009 23336 2450
rect 27632 2417 27660 2450
rect 27618 2408 27674 2417
rect 27618 2343 27674 2352
rect 28552 2281 28580 2450
rect 28538 2272 28594 2281
rect 28538 2207 28594 2216
rect 23294 2000 23350 2009
rect 23294 1935 23350 1944
rect 29564 1873 29592 2926
rect 30378 2887 30434 2896
rect 31574 2952 31630 2961
rect 31574 2887 31630 2896
rect 30286 2544 30342 2553
rect 30286 2479 30288 2488
rect 30340 2479 30342 2488
rect 30288 2450 30340 2456
rect 29550 1864 29606 1873
rect 29550 1799 29606 1808
rect 19154 1728 19210 1737
rect 19154 1663 19210 1672
rect 20442 1728 20498 1737
rect 20442 1663 20498 1672
rect 12438 1592 12494 1601
rect 12438 1527 12494 1536
rect 11886 1320 11942 1329
rect 11886 1255 11942 1264
rect 1398 776 1454 785
rect 1398 711 1454 720
rect 1858 0 1914 800
rect 2778 0 2834 800
rect 3698 0 3754 800
rect 4618 0 4674 800
rect 5538 0 5594 800
rect 6458 0 6514 800
rect 7378 0 7434 800
rect 8298 0 8354 800
rect 9218 0 9274 800
rect 10138 0 10194 800
rect 11058 0 11114 800
rect 19168 82 19196 1663
rect 30392 800 30420 2887
rect 31298 2816 31354 2825
rect 31298 2751 31354 2760
rect 31312 800 31340 2751
rect 31588 2650 31616 2887
rect 31576 2644 31628 2650
rect 31576 2586 31628 2592
rect 31392 2508 31444 2514
rect 31392 2450 31444 2456
rect 31404 1737 31432 2450
rect 31390 1728 31446 1737
rect 31390 1663 31446 1672
rect 32232 800 32260 3023
rect 32600 2514 32628 3159
rect 34058 2952 34114 2961
rect 34058 2887 34114 2896
rect 32770 2816 32826 2825
rect 32770 2751 32826 2760
rect 32784 2650 32812 2751
rect 32772 2644 32824 2650
rect 32772 2586 32824 2592
rect 32588 2508 32640 2514
rect 32588 2450 32640 2456
rect 33048 2440 33100 2446
rect 33100 2388 33180 2394
rect 33048 2382 33180 2388
rect 33060 2366 33180 2382
rect 33152 800 33180 2366
rect 34072 800 34100 2887
rect 34289 2204 34585 2224
rect 34345 2202 34369 2204
rect 34425 2202 34449 2204
rect 34505 2202 34529 2204
rect 34367 2150 34369 2202
rect 34431 2150 34443 2202
rect 34505 2150 34507 2202
rect 34345 2148 34369 2150
rect 34425 2148 34449 2150
rect 34505 2148 34529 2150
rect 34289 2128 34585 2148
rect 34624 2009 34652 3431
rect 35898 3088 35954 3097
rect 35898 3023 35954 3032
rect 34978 2816 35034 2825
rect 34978 2751 35034 2760
rect 34702 2136 34758 2145
rect 34702 2071 34758 2080
rect 34610 2000 34666 2009
rect 34610 1935 34666 1944
rect 34716 1193 34744 2071
rect 34702 1184 34758 1193
rect 34702 1119 34758 1128
rect 34992 800 35020 2751
rect 35912 800 35940 3023
rect 36832 800 36860 3703
rect 37752 800 37780 3975
rect 38658 3904 38714 3913
rect 38658 3839 38714 3848
rect 38672 800 38700 3839
rect 39578 2408 39634 2417
rect 39578 2343 39634 2352
rect 39592 800 39620 2343
rect 19246 96 19302 105
rect 19168 54 19246 82
rect 19246 31 19302 40
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 34058 0 34114 800
rect 34978 0 35034 800
rect 35898 0 35954 800
rect 36818 0 36874 800
rect 37738 0 37794 800
rect 38658 0 38714 800
rect 39578 0 39634 800
<< via2 >>
rect 3422 15680 3478 15736
rect 478 11600 534 11656
rect 14289 13626 14345 13628
rect 14369 13626 14425 13628
rect 14449 13626 14505 13628
rect 14529 13626 14585 13628
rect 14289 13574 14315 13626
rect 14315 13574 14345 13626
rect 14369 13574 14379 13626
rect 14379 13574 14425 13626
rect 14449 13574 14495 13626
rect 14495 13574 14505 13626
rect 14529 13574 14559 13626
rect 14559 13574 14585 13626
rect 14289 13572 14345 13574
rect 14369 13572 14425 13574
rect 14449 13572 14505 13574
rect 14529 13572 14585 13574
rect 7622 13082 7678 13084
rect 7702 13082 7758 13084
rect 7782 13082 7838 13084
rect 7862 13082 7918 13084
rect 7622 13030 7648 13082
rect 7648 13030 7678 13082
rect 7702 13030 7712 13082
rect 7712 13030 7758 13082
rect 7782 13030 7828 13082
rect 7828 13030 7838 13082
rect 7862 13030 7892 13082
rect 7892 13030 7918 13082
rect 7622 13028 7678 13030
rect 7702 13028 7758 13030
rect 7782 13028 7838 13030
rect 7862 13028 7918 13030
rect 14289 12538 14345 12540
rect 14369 12538 14425 12540
rect 14449 12538 14505 12540
rect 14529 12538 14585 12540
rect 14289 12486 14315 12538
rect 14315 12486 14345 12538
rect 14369 12486 14379 12538
rect 14379 12486 14425 12538
rect 14449 12486 14495 12538
rect 14495 12486 14505 12538
rect 14529 12486 14559 12538
rect 14559 12486 14585 12538
rect 14289 12484 14345 12486
rect 14369 12484 14425 12486
rect 14449 12484 14505 12486
rect 14529 12484 14585 12486
rect 7622 11994 7678 11996
rect 7702 11994 7758 11996
rect 7782 11994 7838 11996
rect 7862 11994 7918 11996
rect 7622 11942 7648 11994
rect 7648 11942 7678 11994
rect 7702 11942 7712 11994
rect 7712 11942 7758 11994
rect 7782 11942 7828 11994
rect 7828 11942 7838 11994
rect 7862 11942 7892 11994
rect 7892 11942 7918 11994
rect 7622 11940 7678 11942
rect 7702 11940 7758 11942
rect 7782 11940 7838 11942
rect 7862 11940 7918 11942
rect 15106 11600 15162 11656
rect 14289 11450 14345 11452
rect 14369 11450 14425 11452
rect 14449 11450 14505 11452
rect 14529 11450 14585 11452
rect 14289 11398 14315 11450
rect 14315 11398 14345 11450
rect 14369 11398 14379 11450
rect 14379 11398 14425 11450
rect 14449 11398 14495 11450
rect 14495 11398 14505 11450
rect 14529 11398 14559 11450
rect 14559 11398 14585 11450
rect 14289 11396 14345 11398
rect 14369 11396 14425 11398
rect 14449 11396 14505 11398
rect 14529 11396 14585 11398
rect 7622 10906 7678 10908
rect 7702 10906 7758 10908
rect 7782 10906 7838 10908
rect 7862 10906 7918 10908
rect 7622 10854 7648 10906
rect 7648 10854 7678 10906
rect 7702 10854 7712 10906
rect 7712 10854 7758 10906
rect 7782 10854 7828 10906
rect 7828 10854 7838 10906
rect 7862 10854 7892 10906
rect 7892 10854 7918 10906
rect 7622 10852 7678 10854
rect 7702 10852 7758 10854
rect 7782 10852 7838 10854
rect 7862 10852 7918 10854
rect 14289 10362 14345 10364
rect 14369 10362 14425 10364
rect 14449 10362 14505 10364
rect 14529 10362 14585 10364
rect 14289 10310 14315 10362
rect 14315 10310 14345 10362
rect 14369 10310 14379 10362
rect 14379 10310 14425 10362
rect 14449 10310 14495 10362
rect 14495 10310 14505 10362
rect 14529 10310 14559 10362
rect 14559 10310 14585 10362
rect 14289 10308 14345 10310
rect 14369 10308 14425 10310
rect 14449 10308 14505 10310
rect 14529 10308 14585 10310
rect 1582 10240 1638 10296
rect 7622 9818 7678 9820
rect 7702 9818 7758 9820
rect 7782 9818 7838 9820
rect 7862 9818 7918 9820
rect 7622 9766 7648 9818
rect 7648 9766 7678 9818
rect 7702 9766 7712 9818
rect 7712 9766 7758 9818
rect 7782 9766 7828 9818
rect 7828 9766 7838 9818
rect 7862 9766 7892 9818
rect 7892 9766 7918 9818
rect 7622 9764 7678 9766
rect 7702 9764 7758 9766
rect 7782 9764 7838 9766
rect 7862 9764 7918 9766
rect 14289 9274 14345 9276
rect 14369 9274 14425 9276
rect 14449 9274 14505 9276
rect 14529 9274 14585 9276
rect 14289 9222 14315 9274
rect 14315 9222 14345 9274
rect 14369 9222 14379 9274
rect 14379 9222 14425 9274
rect 14449 9222 14495 9274
rect 14495 9222 14505 9274
rect 14529 9222 14559 9274
rect 14559 9222 14585 9274
rect 14289 9220 14345 9222
rect 14369 9220 14425 9222
rect 14449 9220 14505 9222
rect 14529 9220 14585 9222
rect 1582 8880 1638 8936
rect 2318 8492 2374 8528
rect 2318 8472 2320 8492
rect 2320 8472 2372 8492
rect 2372 8472 2374 8492
rect 1950 8356 2006 8392
rect 1950 8336 1952 8356
rect 1952 8336 2004 8356
rect 2004 8336 2006 8356
rect 1582 7520 1638 7576
rect 18 3712 74 3768
rect 938 2760 994 2816
rect 2042 6060 2044 6080
rect 2044 6060 2096 6080
rect 2096 6060 2098 6080
rect 2042 6024 2098 6060
rect 2042 4936 2098 4992
rect 4158 6740 4160 6760
rect 4160 6740 4212 6760
rect 4212 6740 4214 6760
rect 4158 6704 4214 6740
rect 2502 5616 2558 5672
rect 3330 5364 3386 5400
rect 3330 5344 3332 5364
rect 3332 5344 3384 5364
rect 3384 5344 3386 5364
rect 3882 5228 3938 5264
rect 3882 5208 3884 5228
rect 3884 5208 3936 5228
rect 3936 5208 3938 5228
rect 2042 3304 2098 3360
rect 3054 2760 3110 2816
rect 3514 2388 3516 2408
rect 3516 2388 3568 2408
rect 3568 2388 3570 2408
rect 3514 2352 3570 2388
rect 2778 1944 2834 2000
rect 4526 5616 4582 5672
rect 5538 5344 5594 5400
rect 4710 3848 4766 3904
rect 4158 2896 4214 2952
rect 4342 2896 4398 2952
rect 5354 4528 5410 4584
rect 5262 4004 5318 4040
rect 5262 3984 5264 4004
rect 5264 3984 5316 4004
rect 5316 3984 5318 4004
rect 5538 3032 5594 3088
rect 4802 1672 4858 1728
rect 6182 5888 6238 5944
rect 15106 8880 15162 8936
rect 7622 8730 7678 8732
rect 7702 8730 7758 8732
rect 7782 8730 7838 8732
rect 7862 8730 7918 8732
rect 7622 8678 7648 8730
rect 7648 8678 7678 8730
rect 7702 8678 7712 8730
rect 7712 8678 7758 8730
rect 7782 8678 7828 8730
rect 7828 8678 7838 8730
rect 7862 8678 7892 8730
rect 7892 8678 7918 8730
rect 7622 8676 7678 8678
rect 7702 8676 7758 8678
rect 7782 8676 7838 8678
rect 7862 8676 7918 8678
rect 6550 7384 6606 7440
rect 6274 4664 6330 4720
rect 7102 8472 7158 8528
rect 13910 8336 13966 8392
rect 6826 7284 6828 7304
rect 6828 7284 6880 7304
rect 6880 7284 6882 7304
rect 6826 7248 6882 7284
rect 7102 3984 7158 4040
rect 6458 2760 6514 2816
rect 6090 2080 6146 2136
rect 6090 1536 6146 1592
rect 7622 7642 7678 7644
rect 7702 7642 7758 7644
rect 7782 7642 7838 7644
rect 7862 7642 7918 7644
rect 7622 7590 7648 7642
rect 7648 7590 7678 7642
rect 7702 7590 7712 7642
rect 7712 7590 7758 7642
rect 7782 7590 7828 7642
rect 7828 7590 7838 7642
rect 7862 7590 7892 7642
rect 7892 7590 7918 7642
rect 7622 7588 7678 7590
rect 7702 7588 7758 7590
rect 7782 7588 7838 7590
rect 7862 7588 7918 7590
rect 8206 7248 8262 7304
rect 7562 6740 7564 6760
rect 7564 6740 7616 6760
rect 7616 6740 7618 6760
rect 7562 6704 7618 6740
rect 7622 6554 7678 6556
rect 7702 6554 7758 6556
rect 7782 6554 7838 6556
rect 7862 6554 7918 6556
rect 7622 6502 7648 6554
rect 7648 6502 7678 6554
rect 7702 6502 7712 6554
rect 7712 6502 7758 6554
rect 7782 6502 7828 6554
rect 7828 6502 7838 6554
rect 7862 6502 7892 6554
rect 7892 6502 7918 6554
rect 7622 6500 7678 6502
rect 7702 6500 7758 6502
rect 7782 6500 7838 6502
rect 7862 6500 7918 6502
rect 7562 6296 7618 6352
rect 9126 6840 9182 6896
rect 11886 6840 11942 6896
rect 7286 4684 7342 4720
rect 7622 5466 7678 5468
rect 7702 5466 7758 5468
rect 7782 5466 7838 5468
rect 7862 5466 7918 5468
rect 7622 5414 7648 5466
rect 7648 5414 7678 5466
rect 7702 5414 7712 5466
rect 7712 5414 7758 5466
rect 7782 5414 7828 5466
rect 7828 5414 7838 5466
rect 7862 5414 7892 5466
rect 7892 5414 7918 5466
rect 7622 5412 7678 5414
rect 7702 5412 7758 5414
rect 7782 5412 7838 5414
rect 7862 5412 7918 5414
rect 7286 4664 7288 4684
rect 7288 4664 7340 4684
rect 7340 4664 7342 4684
rect 7622 4378 7678 4380
rect 7702 4378 7758 4380
rect 7782 4378 7838 4380
rect 7862 4378 7918 4380
rect 7622 4326 7648 4378
rect 7648 4326 7678 4378
rect 7702 4326 7712 4378
rect 7712 4326 7758 4378
rect 7782 4326 7828 4378
rect 7828 4326 7838 4378
rect 7862 4326 7892 4378
rect 7892 4326 7918 4378
rect 7622 4324 7678 4326
rect 7702 4324 7758 4326
rect 7782 4324 7838 4326
rect 7862 4324 7918 4326
rect 7378 2896 7434 2952
rect 7194 1672 7250 1728
rect 7622 3290 7678 3292
rect 7702 3290 7758 3292
rect 7782 3290 7838 3292
rect 7862 3290 7918 3292
rect 7622 3238 7648 3290
rect 7648 3238 7678 3290
rect 7702 3238 7712 3290
rect 7712 3238 7758 3290
rect 7782 3238 7828 3290
rect 7828 3238 7838 3290
rect 7862 3238 7892 3290
rect 7892 3238 7918 3290
rect 7622 3236 7678 3238
rect 7702 3236 7758 3238
rect 7782 3236 7838 3238
rect 7862 3236 7918 3238
rect 8574 3848 8630 3904
rect 9494 5072 9550 5128
rect 9126 4528 9182 4584
rect 8942 3712 8998 3768
rect 8942 3168 8998 3224
rect 7622 2202 7678 2204
rect 7702 2202 7758 2204
rect 7782 2202 7838 2204
rect 7862 2202 7918 2204
rect 7622 2150 7648 2202
rect 7648 2150 7678 2202
rect 7702 2150 7712 2202
rect 7712 2150 7758 2202
rect 7782 2150 7828 2202
rect 7828 2150 7838 2202
rect 7862 2150 7892 2202
rect 7892 2150 7918 2202
rect 7622 2148 7678 2150
rect 7702 2148 7758 2150
rect 7782 2148 7838 2150
rect 7862 2148 7918 2150
rect 8390 2252 8392 2272
rect 8392 2252 8444 2272
rect 8444 2252 8446 2272
rect 8390 2216 8446 2252
rect 10230 5072 10286 5128
rect 11334 6024 11390 6080
rect 9494 2932 9496 2952
rect 9496 2932 9548 2952
rect 9548 2932 9550 2952
rect 9494 2896 9550 2932
rect 10874 4936 10930 4992
rect 10874 4664 10930 4720
rect 11242 5108 11244 5128
rect 11244 5108 11296 5128
rect 11296 5108 11298 5128
rect 11242 5072 11298 5108
rect 9862 3304 9918 3360
rect 10322 3304 10378 3360
rect 12070 6840 12126 6896
rect 13542 7248 13598 7304
rect 12714 5888 12770 5944
rect 12990 5772 13046 5808
rect 12990 5752 12992 5772
rect 12992 5752 13044 5772
rect 13044 5752 13046 5772
rect 12806 5480 12862 5536
rect 10414 2508 10470 2544
rect 10414 2488 10416 2508
rect 10416 2488 10468 2508
rect 10468 2488 10470 2508
rect 12530 3848 12586 3904
rect 11886 3168 11942 3224
rect 11794 3052 11850 3088
rect 11794 3032 11796 3052
rect 11796 3032 11848 3052
rect 11848 3032 11850 3052
rect 12070 2080 12126 2136
rect 13634 6332 13636 6352
rect 13636 6332 13688 6352
rect 13688 6332 13690 6352
rect 13634 6296 13690 6332
rect 13542 2760 13598 2816
rect 14289 8186 14345 8188
rect 14369 8186 14425 8188
rect 14449 8186 14505 8188
rect 14529 8186 14585 8188
rect 14289 8134 14315 8186
rect 14315 8134 14345 8186
rect 14369 8134 14379 8186
rect 14379 8134 14425 8186
rect 14449 8134 14495 8186
rect 14495 8134 14505 8186
rect 14529 8134 14559 8186
rect 14559 8134 14585 8186
rect 14289 8132 14345 8134
rect 14369 8132 14425 8134
rect 14449 8132 14505 8134
rect 14529 8132 14585 8134
rect 15198 7928 15254 7984
rect 14738 7384 14794 7440
rect 14289 7098 14345 7100
rect 14369 7098 14425 7100
rect 14449 7098 14505 7100
rect 14529 7098 14585 7100
rect 14289 7046 14315 7098
rect 14315 7046 14345 7098
rect 14369 7046 14379 7098
rect 14379 7046 14425 7098
rect 14449 7046 14495 7098
rect 14495 7046 14505 7098
rect 14529 7046 14559 7098
rect 14559 7046 14585 7098
rect 14289 7044 14345 7046
rect 14369 7044 14425 7046
rect 14449 7044 14505 7046
rect 14529 7044 14585 7046
rect 14830 7112 14886 7168
rect 14094 4936 14150 4992
rect 14289 6010 14345 6012
rect 14369 6010 14425 6012
rect 14449 6010 14505 6012
rect 14529 6010 14585 6012
rect 14289 5958 14315 6010
rect 14315 5958 14345 6010
rect 14369 5958 14379 6010
rect 14379 5958 14425 6010
rect 14449 5958 14495 6010
rect 14495 5958 14505 6010
rect 14529 5958 14559 6010
rect 14559 5958 14585 6010
rect 14289 5956 14345 5958
rect 14369 5956 14425 5958
rect 14449 5956 14505 5958
rect 14529 5956 14585 5958
rect 15842 7112 15898 7168
rect 15750 6296 15806 6352
rect 14370 5208 14426 5264
rect 14289 4922 14345 4924
rect 14369 4922 14425 4924
rect 14449 4922 14505 4924
rect 14529 4922 14585 4924
rect 14289 4870 14315 4922
rect 14315 4870 14345 4922
rect 14369 4870 14379 4922
rect 14379 4870 14425 4922
rect 14449 4870 14495 4922
rect 14495 4870 14505 4922
rect 14529 4870 14559 4922
rect 14559 4870 14585 4922
rect 14289 4868 14345 4870
rect 14369 4868 14425 4870
rect 14449 4868 14505 4870
rect 14529 4868 14585 4870
rect 14289 3834 14345 3836
rect 14369 3834 14425 3836
rect 14449 3834 14505 3836
rect 14529 3834 14585 3836
rect 14289 3782 14315 3834
rect 14315 3782 14345 3834
rect 14369 3782 14379 3834
rect 14379 3782 14425 3834
rect 14449 3782 14495 3834
rect 14495 3782 14505 3834
rect 14529 3782 14559 3834
rect 14559 3782 14585 3834
rect 14289 3780 14345 3782
rect 14369 3780 14425 3782
rect 14449 3780 14505 3782
rect 14529 3780 14585 3782
rect 14186 3596 14242 3632
rect 14186 3576 14188 3596
rect 14188 3576 14240 3596
rect 14240 3576 14242 3596
rect 15106 3712 15162 3768
rect 16486 11056 16542 11112
rect 17038 10104 17094 10160
rect 18878 11056 18934 11112
rect 20956 13082 21012 13084
rect 21036 13082 21092 13084
rect 21116 13082 21172 13084
rect 21196 13082 21252 13084
rect 20956 13030 20982 13082
rect 20982 13030 21012 13082
rect 21036 13030 21046 13082
rect 21046 13030 21092 13082
rect 21116 13030 21162 13082
rect 21162 13030 21172 13082
rect 21196 13030 21226 13082
rect 21226 13030 21252 13082
rect 20956 13028 21012 13030
rect 21036 13028 21092 13030
rect 21116 13028 21172 13030
rect 21196 13028 21252 13030
rect 20956 11994 21012 11996
rect 21036 11994 21092 11996
rect 21116 11994 21172 11996
rect 21196 11994 21252 11996
rect 20956 11942 20982 11994
rect 20982 11942 21012 11994
rect 21036 11942 21046 11994
rect 21046 11942 21092 11994
rect 21116 11942 21162 11994
rect 21162 11942 21172 11994
rect 21196 11942 21226 11994
rect 21226 11942 21252 11994
rect 20956 11940 21012 11942
rect 21036 11940 21092 11942
rect 21116 11940 21172 11942
rect 21196 11940 21252 11942
rect 20956 10906 21012 10908
rect 21036 10906 21092 10908
rect 21116 10906 21172 10908
rect 21196 10906 21252 10908
rect 20956 10854 20982 10906
rect 20982 10854 21012 10906
rect 21036 10854 21046 10906
rect 21046 10854 21092 10906
rect 21116 10854 21162 10906
rect 21162 10854 21172 10906
rect 21196 10854 21226 10906
rect 21226 10854 21252 10906
rect 20956 10852 21012 10854
rect 21036 10852 21092 10854
rect 21116 10852 21172 10854
rect 21196 10852 21252 10854
rect 20956 9818 21012 9820
rect 21036 9818 21092 9820
rect 21116 9818 21172 9820
rect 21196 9818 21252 9820
rect 20956 9766 20982 9818
rect 20982 9766 21012 9818
rect 21036 9766 21046 9818
rect 21046 9766 21092 9818
rect 21116 9766 21162 9818
rect 21162 9766 21172 9818
rect 21196 9766 21226 9818
rect 21226 9766 21252 9818
rect 20956 9764 21012 9766
rect 21036 9764 21092 9766
rect 21116 9764 21172 9766
rect 21196 9764 21252 9766
rect 20956 8730 21012 8732
rect 21036 8730 21092 8732
rect 21116 8730 21172 8732
rect 21196 8730 21252 8732
rect 20956 8678 20982 8730
rect 20982 8678 21012 8730
rect 21036 8678 21046 8730
rect 21046 8678 21092 8730
rect 21116 8678 21162 8730
rect 21162 8678 21172 8730
rect 21196 8678 21226 8730
rect 21226 8678 21252 8730
rect 20956 8676 21012 8678
rect 21036 8676 21092 8678
rect 21116 8676 21172 8678
rect 21196 8676 21252 8678
rect 17130 7948 17186 7984
rect 17130 7928 17132 7948
rect 17132 7928 17184 7948
rect 17184 7928 17186 7948
rect 16946 6976 17002 7032
rect 17314 6296 17370 6352
rect 16394 6024 16450 6080
rect 16670 5752 16726 5808
rect 17222 5480 17278 5536
rect 17130 5228 17186 5264
rect 17130 5208 17132 5228
rect 17132 5208 17184 5228
rect 17184 5208 17186 5228
rect 19430 5752 19486 5808
rect 19706 6840 19762 6896
rect 20442 6296 20498 6352
rect 19798 6060 19800 6080
rect 19800 6060 19852 6080
rect 19852 6060 19854 6080
rect 19798 6024 19854 6060
rect 14738 2760 14794 2816
rect 14289 2746 14345 2748
rect 14369 2746 14425 2748
rect 14449 2746 14505 2748
rect 14529 2746 14585 2748
rect 14289 2694 14315 2746
rect 14315 2694 14345 2746
rect 14369 2694 14379 2746
rect 14379 2694 14425 2746
rect 14449 2694 14495 2746
rect 14495 2694 14505 2746
rect 14529 2694 14559 2746
rect 14559 2694 14585 2746
rect 14289 2692 14345 2694
rect 14369 2692 14425 2694
rect 14449 2692 14505 2694
rect 14529 2692 14585 2694
rect 15106 3168 15162 3224
rect 14922 2624 14978 2680
rect 17222 3712 17278 3768
rect 20956 7642 21012 7644
rect 21036 7642 21092 7644
rect 21116 7642 21172 7644
rect 21196 7642 21252 7644
rect 20956 7590 20982 7642
rect 20982 7590 21012 7642
rect 21036 7590 21046 7642
rect 21046 7590 21092 7642
rect 21116 7590 21162 7642
rect 21162 7590 21172 7642
rect 21196 7590 21226 7642
rect 21226 7590 21252 7642
rect 20956 7588 21012 7590
rect 21036 7588 21092 7590
rect 21116 7588 21172 7590
rect 21196 7588 21252 7590
rect 20956 6554 21012 6556
rect 21036 6554 21092 6556
rect 21116 6554 21172 6556
rect 21196 6554 21252 6556
rect 20956 6502 20982 6554
rect 20982 6502 21012 6554
rect 21036 6502 21046 6554
rect 21046 6502 21092 6554
rect 21116 6502 21162 6554
rect 21162 6502 21172 6554
rect 21196 6502 21226 6554
rect 21226 6502 21252 6554
rect 20956 6500 21012 6502
rect 21036 6500 21092 6502
rect 21116 6500 21172 6502
rect 21196 6500 21252 6502
rect 15474 3440 15530 3496
rect 15382 3304 15438 3360
rect 17406 3168 17462 3224
rect 15474 2896 15530 2952
rect 16670 2932 16672 2952
rect 16672 2932 16724 2952
rect 16724 2932 16726 2952
rect 16670 2896 16726 2932
rect 15198 2252 15200 2272
rect 15200 2252 15252 2272
rect 15252 2252 15254 2272
rect 15198 2216 15254 2252
rect 15382 2216 15438 2272
rect 16578 2080 16634 2136
rect 17038 2624 17094 2680
rect 17314 2488 17370 2544
rect 16670 1944 16726 2000
rect 12530 1808 12586 1864
rect 20718 5208 20774 5264
rect 24214 7384 24270 7440
rect 20956 5466 21012 5468
rect 21036 5466 21092 5468
rect 21116 5466 21172 5468
rect 21196 5466 21252 5468
rect 20956 5414 20982 5466
rect 20982 5414 21012 5466
rect 21036 5414 21046 5466
rect 21046 5414 21092 5466
rect 21116 5414 21162 5466
rect 21162 5414 21172 5466
rect 21196 5414 21226 5466
rect 21226 5414 21252 5466
rect 20956 5412 21012 5414
rect 21036 5412 21092 5414
rect 21116 5412 21172 5414
rect 21196 5412 21252 5414
rect 19706 3576 19762 3632
rect 20956 4378 21012 4380
rect 21036 4378 21092 4380
rect 21116 4378 21172 4380
rect 21196 4378 21252 4380
rect 20956 4326 20982 4378
rect 20982 4326 21012 4378
rect 21036 4326 21046 4378
rect 21046 4326 21092 4378
rect 21116 4326 21162 4378
rect 21162 4326 21172 4378
rect 21196 4326 21226 4378
rect 21226 4326 21252 4378
rect 20956 4324 21012 4326
rect 21036 4324 21092 4326
rect 21116 4324 21172 4326
rect 21196 4324 21252 4326
rect 21454 5616 21510 5672
rect 21822 5752 21878 5808
rect 22282 6160 22338 6216
rect 27622 13626 27678 13628
rect 27702 13626 27758 13628
rect 27782 13626 27838 13628
rect 27862 13626 27918 13628
rect 27622 13574 27648 13626
rect 27648 13574 27678 13626
rect 27702 13574 27712 13626
rect 27712 13574 27758 13626
rect 27782 13574 27828 13626
rect 27828 13574 27838 13626
rect 27862 13574 27892 13626
rect 27892 13574 27918 13626
rect 27622 13572 27678 13574
rect 27702 13572 27758 13574
rect 27782 13572 27838 13574
rect 27862 13572 27918 13574
rect 34289 13082 34345 13084
rect 34369 13082 34425 13084
rect 34449 13082 34505 13084
rect 34529 13082 34585 13084
rect 34289 13030 34315 13082
rect 34315 13030 34345 13082
rect 34369 13030 34379 13082
rect 34379 13030 34425 13082
rect 34449 13030 34495 13082
rect 34495 13030 34505 13082
rect 34529 13030 34559 13082
rect 34559 13030 34585 13082
rect 34289 13028 34345 13030
rect 34369 13028 34425 13030
rect 34449 13028 34505 13030
rect 34529 13028 34585 13030
rect 27622 12538 27678 12540
rect 27702 12538 27758 12540
rect 27782 12538 27838 12540
rect 27862 12538 27918 12540
rect 27622 12486 27648 12538
rect 27648 12486 27678 12538
rect 27702 12486 27712 12538
rect 27712 12486 27758 12538
rect 27782 12486 27828 12538
rect 27828 12486 27838 12538
rect 27862 12486 27892 12538
rect 27892 12486 27918 12538
rect 27622 12484 27678 12486
rect 27702 12484 27758 12486
rect 27782 12484 27838 12486
rect 27862 12484 27918 12486
rect 34289 11994 34345 11996
rect 34369 11994 34425 11996
rect 34449 11994 34505 11996
rect 34529 11994 34585 11996
rect 34289 11942 34315 11994
rect 34315 11942 34345 11994
rect 34369 11942 34379 11994
rect 34379 11942 34425 11994
rect 34449 11942 34495 11994
rect 34495 11942 34505 11994
rect 34529 11942 34559 11994
rect 34559 11942 34585 11994
rect 34289 11940 34345 11942
rect 34369 11940 34425 11942
rect 34449 11940 34505 11942
rect 34529 11940 34585 11942
rect 27622 11450 27678 11452
rect 27702 11450 27758 11452
rect 27782 11450 27838 11452
rect 27862 11450 27918 11452
rect 27622 11398 27648 11450
rect 27648 11398 27678 11450
rect 27702 11398 27712 11450
rect 27712 11398 27758 11450
rect 27782 11398 27828 11450
rect 27828 11398 27838 11450
rect 27862 11398 27892 11450
rect 27892 11398 27918 11450
rect 27622 11396 27678 11398
rect 27702 11396 27758 11398
rect 27782 11396 27838 11398
rect 27862 11396 27918 11398
rect 34289 10906 34345 10908
rect 34369 10906 34425 10908
rect 34449 10906 34505 10908
rect 34529 10906 34585 10908
rect 34289 10854 34315 10906
rect 34315 10854 34345 10906
rect 34369 10854 34379 10906
rect 34379 10854 34425 10906
rect 34449 10854 34495 10906
rect 34495 10854 34505 10906
rect 34529 10854 34559 10906
rect 34559 10854 34585 10906
rect 34289 10852 34345 10854
rect 34369 10852 34425 10854
rect 34449 10852 34505 10854
rect 34529 10852 34585 10854
rect 27622 10362 27678 10364
rect 27702 10362 27758 10364
rect 27782 10362 27838 10364
rect 27862 10362 27918 10364
rect 27622 10310 27648 10362
rect 27648 10310 27678 10362
rect 27702 10310 27712 10362
rect 27712 10310 27758 10362
rect 27782 10310 27828 10362
rect 27828 10310 27838 10362
rect 27862 10310 27892 10362
rect 27892 10310 27918 10362
rect 27622 10308 27678 10310
rect 27702 10308 27758 10310
rect 27782 10308 27838 10310
rect 27862 10308 27918 10310
rect 34289 9818 34345 9820
rect 34369 9818 34425 9820
rect 34449 9818 34505 9820
rect 34529 9818 34585 9820
rect 34289 9766 34315 9818
rect 34315 9766 34345 9818
rect 34369 9766 34379 9818
rect 34379 9766 34425 9818
rect 34449 9766 34495 9818
rect 34495 9766 34505 9818
rect 34529 9766 34559 9818
rect 34559 9766 34585 9818
rect 34289 9764 34345 9766
rect 34369 9764 34425 9766
rect 34449 9764 34505 9766
rect 34529 9764 34585 9766
rect 27622 9274 27678 9276
rect 27702 9274 27758 9276
rect 27782 9274 27838 9276
rect 27862 9274 27918 9276
rect 27622 9222 27648 9274
rect 27648 9222 27678 9274
rect 27702 9222 27712 9274
rect 27712 9222 27758 9274
rect 27782 9222 27828 9274
rect 27828 9222 27838 9274
rect 27862 9222 27892 9274
rect 27892 9222 27918 9274
rect 27622 9220 27678 9222
rect 27702 9220 27758 9222
rect 27782 9220 27838 9222
rect 27862 9220 27918 9222
rect 28998 8880 29054 8936
rect 35622 8880 35678 8936
rect 27622 8186 27678 8188
rect 27702 8186 27758 8188
rect 27782 8186 27838 8188
rect 27862 8186 27918 8188
rect 27622 8134 27648 8186
rect 27648 8134 27678 8186
rect 27702 8134 27712 8186
rect 27712 8134 27758 8186
rect 27782 8134 27828 8186
rect 27828 8134 27838 8186
rect 27862 8134 27892 8186
rect 27892 8134 27918 8186
rect 27622 8132 27678 8134
rect 27702 8132 27758 8134
rect 27782 8132 27838 8134
rect 27862 8132 27918 8134
rect 27158 7384 27214 7440
rect 24214 7112 24270 7168
rect 24306 6976 24362 7032
rect 24122 5772 24178 5808
rect 24122 5752 24124 5772
rect 24124 5752 24176 5772
rect 24176 5752 24178 5772
rect 23846 5616 23902 5672
rect 27622 7098 27678 7100
rect 27702 7098 27758 7100
rect 27782 7098 27838 7100
rect 27862 7098 27918 7100
rect 27622 7046 27648 7098
rect 27648 7046 27678 7098
rect 27702 7046 27712 7098
rect 27712 7046 27758 7098
rect 27782 7046 27828 7098
rect 27828 7046 27838 7098
rect 27862 7046 27892 7098
rect 27892 7046 27918 7098
rect 27622 7044 27678 7046
rect 27702 7044 27758 7046
rect 27782 7044 27838 7046
rect 27862 7044 27918 7046
rect 34289 8730 34345 8732
rect 34369 8730 34425 8732
rect 34449 8730 34505 8732
rect 34529 8730 34585 8732
rect 34289 8678 34315 8730
rect 34315 8678 34345 8730
rect 34369 8678 34379 8730
rect 34379 8678 34425 8730
rect 34449 8678 34495 8730
rect 34495 8678 34505 8730
rect 34529 8678 34559 8730
rect 34559 8678 34585 8730
rect 34289 8676 34345 8678
rect 34369 8676 34425 8678
rect 34449 8676 34505 8678
rect 34529 8676 34585 8678
rect 34289 7642 34345 7644
rect 34369 7642 34425 7644
rect 34449 7642 34505 7644
rect 34529 7642 34585 7644
rect 34289 7590 34315 7642
rect 34315 7590 34345 7642
rect 34369 7590 34379 7642
rect 34379 7590 34425 7642
rect 34449 7590 34495 7642
rect 34495 7590 34505 7642
rect 34529 7590 34559 7642
rect 34559 7590 34585 7642
rect 34289 7588 34345 7590
rect 34369 7588 34425 7590
rect 34449 7588 34505 7590
rect 34529 7588 34585 7590
rect 33414 7384 33470 7440
rect 25594 6196 25596 6216
rect 25596 6196 25648 6216
rect 25648 6196 25650 6216
rect 25594 6160 25650 6196
rect 25686 5244 25688 5264
rect 25688 5244 25740 5264
rect 25740 5244 25742 5264
rect 25686 5208 25742 5244
rect 20902 4120 20958 4176
rect 21270 4120 21326 4176
rect 20956 3290 21012 3292
rect 21036 3290 21092 3292
rect 21116 3290 21172 3292
rect 21196 3290 21252 3292
rect 20956 3238 20982 3290
rect 20982 3238 21012 3290
rect 21036 3238 21046 3290
rect 21046 3238 21092 3290
rect 21116 3238 21162 3290
rect 21162 3238 21172 3290
rect 21196 3238 21226 3290
rect 21226 3238 21252 3290
rect 20956 3236 21012 3238
rect 21036 3236 21092 3238
rect 21116 3236 21172 3238
rect 21196 3236 21252 3238
rect 24398 4548 24454 4584
rect 24398 4528 24400 4548
rect 24400 4528 24452 4548
rect 24452 4528 24454 4548
rect 23294 2932 23296 2952
rect 23296 2932 23348 2952
rect 23348 2932 23350 2952
rect 23294 2896 23350 2932
rect 23294 2624 23350 2680
rect 27710 6296 27766 6352
rect 27622 6010 27678 6012
rect 27702 6010 27758 6012
rect 27782 6010 27838 6012
rect 27862 6010 27918 6012
rect 27622 5958 27648 6010
rect 27648 5958 27678 6010
rect 27702 5958 27712 6010
rect 27712 5958 27758 6010
rect 27782 5958 27828 6010
rect 27828 5958 27838 6010
rect 27862 5958 27892 6010
rect 27892 5958 27918 6010
rect 27622 5956 27678 5958
rect 27702 5956 27758 5958
rect 27782 5956 27838 5958
rect 27862 5956 27918 5958
rect 27066 4392 27122 4448
rect 26606 4120 26662 4176
rect 27622 4922 27678 4924
rect 27702 4922 27758 4924
rect 27782 4922 27838 4924
rect 27862 4922 27918 4924
rect 27622 4870 27648 4922
rect 27648 4870 27678 4922
rect 27702 4870 27712 4922
rect 27712 4870 27758 4922
rect 27782 4870 27828 4922
rect 27828 4870 27838 4922
rect 27862 4870 27892 4922
rect 27892 4870 27918 4922
rect 27622 4868 27678 4870
rect 27702 4868 27758 4870
rect 27782 4868 27838 4870
rect 27862 4868 27918 4870
rect 27066 3168 27122 3224
rect 27622 3834 27678 3836
rect 27702 3834 27758 3836
rect 27782 3834 27838 3836
rect 27862 3834 27918 3836
rect 27622 3782 27648 3834
rect 27648 3782 27678 3834
rect 27702 3782 27712 3834
rect 27712 3782 27758 3834
rect 27782 3782 27828 3834
rect 27828 3782 27838 3834
rect 27862 3782 27892 3834
rect 27892 3782 27918 3834
rect 27622 3780 27678 3782
rect 27702 3780 27758 3782
rect 27782 3780 27838 3782
rect 27862 3780 27918 3782
rect 27622 2746 27678 2748
rect 27702 2746 27758 2748
rect 27782 2746 27838 2748
rect 27862 2746 27918 2748
rect 27622 2694 27648 2746
rect 27648 2694 27678 2746
rect 27702 2694 27712 2746
rect 27712 2694 27758 2746
rect 27782 2694 27828 2746
rect 27828 2694 27838 2746
rect 27862 2694 27892 2746
rect 27892 2694 27918 2746
rect 27622 2692 27678 2694
rect 27702 2692 27758 2694
rect 27782 2692 27838 2694
rect 27862 2692 27918 2694
rect 28630 4256 28686 4312
rect 35438 7284 35440 7304
rect 35440 7284 35492 7304
rect 35492 7284 35494 7304
rect 35438 7248 35494 7284
rect 34289 6554 34345 6556
rect 34369 6554 34425 6556
rect 34449 6554 34505 6556
rect 34529 6554 34585 6556
rect 34289 6502 34315 6554
rect 34315 6502 34345 6554
rect 34369 6502 34379 6554
rect 34379 6502 34425 6554
rect 34449 6502 34495 6554
rect 34495 6502 34505 6554
rect 34529 6502 34559 6554
rect 34559 6502 34585 6554
rect 34289 6500 34345 6502
rect 34369 6500 34425 6502
rect 34449 6500 34505 6502
rect 34529 6500 34585 6502
rect 29734 5072 29790 5128
rect 34610 6160 34666 6216
rect 34289 5466 34345 5468
rect 34369 5466 34425 5468
rect 34449 5466 34505 5468
rect 34529 5466 34585 5468
rect 34289 5414 34315 5466
rect 34315 5414 34345 5466
rect 34369 5414 34379 5466
rect 34379 5414 34425 5466
rect 34449 5414 34495 5466
rect 34495 5414 34505 5466
rect 34529 5414 34559 5466
rect 34559 5414 34585 5466
rect 34289 5412 34345 5414
rect 34369 5412 34425 5414
rect 34449 5412 34505 5414
rect 34529 5412 34585 5414
rect 33230 5072 33286 5128
rect 30378 4256 30434 4312
rect 34702 4800 34758 4856
rect 34610 4528 34666 4584
rect 34289 4378 34345 4380
rect 34369 4378 34425 4380
rect 34449 4378 34505 4380
rect 34529 4378 34585 4380
rect 34289 4326 34315 4378
rect 34315 4326 34345 4378
rect 34369 4326 34379 4378
rect 34379 4326 34425 4378
rect 34449 4326 34495 4378
rect 34495 4326 34505 4378
rect 34529 4326 34559 4378
rect 34559 4326 34585 4378
rect 34289 4324 34345 4326
rect 34369 4324 34425 4326
rect 34449 4324 34505 4326
rect 34529 4324 34585 4326
rect 30838 4020 30840 4040
rect 30840 4020 30892 4040
rect 30892 4020 30894 4040
rect 30838 3984 30894 4020
rect 37738 3984 37794 4040
rect 31114 3712 31170 3768
rect 34702 3712 34758 3768
rect 34886 3712 34942 3768
rect 36818 3712 36874 3768
rect 34426 3440 34482 3496
rect 34610 3440 34666 3496
rect 31114 3304 31170 3360
rect 34289 3290 34345 3292
rect 34369 3290 34425 3292
rect 34449 3290 34505 3292
rect 34529 3290 34585 3292
rect 34289 3238 34315 3290
rect 34315 3238 34345 3290
rect 34369 3238 34379 3290
rect 34379 3238 34425 3290
rect 34449 3238 34495 3290
rect 34495 3238 34505 3290
rect 34529 3238 34559 3290
rect 34559 3238 34585 3290
rect 34289 3236 34345 3238
rect 34369 3236 34425 3238
rect 34449 3236 34505 3238
rect 34529 3236 34585 3238
rect 32586 3168 32642 3224
rect 29734 3068 29736 3088
rect 29736 3068 29788 3088
rect 29788 3068 29790 3088
rect 29734 3032 29790 3068
rect 32218 3032 32274 3088
rect 28262 2896 28318 2952
rect 28722 2760 28778 2816
rect 20442 2216 20498 2272
rect 21730 2252 21732 2272
rect 21732 2252 21784 2272
rect 21784 2252 21786 2272
rect 21730 2216 21786 2252
rect 20956 2202 21012 2204
rect 21036 2202 21092 2204
rect 21116 2202 21172 2204
rect 21196 2202 21252 2204
rect 20956 2150 20982 2202
rect 20982 2150 21012 2202
rect 21036 2150 21046 2202
rect 21046 2150 21092 2202
rect 21116 2150 21162 2202
rect 21162 2150 21172 2202
rect 21196 2150 21226 2202
rect 21226 2150 21252 2202
rect 20956 2148 21012 2150
rect 21036 2148 21092 2150
rect 21116 2148 21172 2150
rect 21196 2148 21252 2150
rect 27618 2352 27674 2408
rect 28538 2216 28594 2272
rect 23294 1944 23350 2000
rect 30378 2896 30434 2952
rect 31574 2896 31630 2952
rect 30286 2508 30342 2544
rect 30286 2488 30288 2508
rect 30288 2488 30340 2508
rect 30340 2488 30342 2508
rect 29550 1808 29606 1864
rect 19154 1672 19210 1728
rect 20442 1672 20498 1728
rect 12438 1536 12494 1592
rect 11886 1264 11942 1320
rect 1398 720 1454 776
rect 31298 2760 31354 2816
rect 31390 1672 31446 1728
rect 34058 2896 34114 2952
rect 32770 2760 32826 2816
rect 34289 2202 34345 2204
rect 34369 2202 34425 2204
rect 34449 2202 34505 2204
rect 34529 2202 34585 2204
rect 34289 2150 34315 2202
rect 34315 2150 34345 2202
rect 34369 2150 34379 2202
rect 34379 2150 34425 2202
rect 34449 2150 34495 2202
rect 34495 2150 34505 2202
rect 34529 2150 34559 2202
rect 34559 2150 34585 2202
rect 34289 2148 34345 2150
rect 34369 2148 34425 2150
rect 34449 2148 34505 2150
rect 34529 2148 34585 2150
rect 35898 3032 35954 3088
rect 34978 2760 35034 2816
rect 34702 2080 34758 2136
rect 34610 1944 34666 2000
rect 34702 1128 34758 1184
rect 38658 3848 38714 3904
rect 39578 2352 39634 2408
rect 19246 40 19302 96
<< metal3 >>
rect 0 15738 800 15768
rect 3417 15738 3483 15741
rect 0 15736 3483 15738
rect 0 15680 3422 15736
rect 3478 15680 3483 15736
rect 0 15678 3483 15680
rect 0 15648 800 15678
rect 3417 15675 3483 15678
rect 14277 13632 14597 13633
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 13567 14597 13568
rect 27610 13632 27930 13633
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 13567 27930 13568
rect 7610 13088 7930 13089
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7930 13088
rect 7610 13023 7930 13024
rect 20944 13088 21264 13089
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 13023 21264 13024
rect 34277 13088 34597 13089
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 13023 34597 13024
rect 14277 12544 14597 12545
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 12479 14597 12480
rect 27610 12544 27930 12545
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 12479 27930 12480
rect 7610 12000 7930 12001
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7930 12000
rect 7610 11935 7930 11936
rect 20944 12000 21264 12001
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 11935 21264 11936
rect 34277 12000 34597 12001
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 11935 34597 11936
rect 473 11658 539 11661
rect 15101 11658 15167 11661
rect 473 11656 15167 11658
rect 473 11600 478 11656
rect 534 11600 15106 11656
rect 15162 11600 15167 11656
rect 473 11598 15167 11600
rect 473 11595 539 11598
rect 15101 11595 15167 11598
rect 14277 11456 14597 11457
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 11391 14597 11392
rect 27610 11456 27930 11457
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 11391 27930 11392
rect 16481 11114 16547 11117
rect 18873 11114 18939 11117
rect 16481 11112 18939 11114
rect 16481 11056 16486 11112
rect 16542 11056 18878 11112
rect 18934 11056 18939 11112
rect 16481 11054 18939 11056
rect 16481 11051 16547 11054
rect 18873 11051 18939 11054
rect 7610 10912 7930 10913
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7930 10912
rect 7610 10847 7930 10848
rect 20944 10912 21264 10913
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 10847 21264 10848
rect 34277 10912 34597 10913
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 10847 34597 10848
rect 28030 10374 39130 10434
rect 14277 10368 14597 10369
rect 0 10298 800 10328
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 10303 14597 10304
rect 27610 10368 27930 10369
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 10303 27930 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10208 800 10238
rect 1577 10235 1643 10238
rect 17033 10162 17099 10165
rect 28030 10162 28090 10374
rect 39070 10298 39130 10374
rect 39200 10298 40000 10328
rect 39070 10238 40000 10298
rect 39200 10208 40000 10238
rect 17033 10160 28090 10162
rect 17033 10104 17038 10160
rect 17094 10104 28090 10160
rect 17033 10102 28090 10104
rect 17033 10099 17099 10102
rect 7610 9824 7930 9825
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7930 9824
rect 7610 9759 7930 9760
rect 20944 9824 21264 9825
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 9759 21264 9760
rect 34277 9824 34597 9825
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 9759 34597 9760
rect 14277 9280 14597 9281
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 9215 14597 9216
rect 27610 9280 27930 9281
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 9215 27930 9216
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 15101 8938 15167 8941
rect 28993 8938 29059 8941
rect 15101 8936 29059 8938
rect 15101 8880 15106 8936
rect 15162 8880 28998 8936
rect 29054 8880 29059 8936
rect 15101 8878 29059 8880
rect 15101 8875 15167 8878
rect 28993 8875 29059 8878
rect 35617 8938 35683 8941
rect 39200 8938 40000 8968
rect 35617 8936 40000 8938
rect 35617 8880 35622 8936
rect 35678 8880 40000 8936
rect 35617 8878 40000 8880
rect 35617 8875 35683 8878
rect 39200 8848 40000 8878
rect 7610 8736 7930 8737
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7930 8736
rect 7610 8671 7930 8672
rect 20944 8736 21264 8737
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 8671 21264 8672
rect 34277 8736 34597 8737
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 8671 34597 8672
rect 2313 8530 2379 8533
rect 7097 8530 7163 8533
rect 2313 8528 7163 8530
rect 2313 8472 2318 8528
rect 2374 8472 7102 8528
rect 7158 8472 7163 8528
rect 2313 8470 7163 8472
rect 2313 8467 2379 8470
rect 7097 8467 7163 8470
rect 1945 8394 2011 8397
rect 13905 8394 13971 8397
rect 1945 8392 13971 8394
rect 1945 8336 1950 8392
rect 2006 8336 13910 8392
rect 13966 8336 13971 8392
rect 1945 8334 13971 8336
rect 1945 8331 2011 8334
rect 13905 8331 13971 8334
rect 14277 8192 14597 8193
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 8127 14597 8128
rect 27610 8192 27930 8193
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 8127 27930 8128
rect 15193 7986 15259 7989
rect 17125 7986 17191 7989
rect 15193 7984 17191 7986
rect 15193 7928 15198 7984
rect 15254 7928 17130 7984
rect 17186 7928 17191 7984
rect 15193 7926 17191 7928
rect 15193 7923 15259 7926
rect 17125 7923 17191 7926
rect 7610 7648 7930 7649
rect 0 7578 800 7608
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7930 7648
rect 7610 7583 7930 7584
rect 20944 7648 21264 7649
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 7583 21264 7584
rect 34277 7648 34597 7649
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 7583 34597 7584
rect 1577 7578 1643 7581
rect 39200 7578 40000 7608
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 34838 7518 40000 7578
rect 6545 7442 6611 7445
rect 14733 7442 14799 7445
rect 6545 7440 14799 7442
rect 6545 7384 6550 7440
rect 6606 7384 14738 7440
rect 14794 7384 14799 7440
rect 6545 7382 14799 7384
rect 6545 7379 6611 7382
rect 14733 7379 14799 7382
rect 24209 7442 24275 7445
rect 27153 7442 27219 7445
rect 24209 7440 27219 7442
rect 24209 7384 24214 7440
rect 24270 7384 27158 7440
rect 27214 7384 27219 7440
rect 24209 7382 27219 7384
rect 24209 7379 24275 7382
rect 27153 7379 27219 7382
rect 33409 7442 33475 7445
rect 34838 7442 34898 7518
rect 39200 7488 40000 7518
rect 33409 7440 34898 7442
rect 33409 7384 33414 7440
rect 33470 7384 34898 7440
rect 33409 7382 34898 7384
rect 33409 7379 33475 7382
rect 6821 7306 6887 7309
rect 8201 7306 8267 7309
rect 6821 7304 8267 7306
rect 6821 7248 6826 7304
rect 6882 7248 8206 7304
rect 8262 7248 8267 7304
rect 6821 7246 8267 7248
rect 6821 7243 6887 7246
rect 8201 7243 8267 7246
rect 13537 7306 13603 7309
rect 35433 7306 35499 7309
rect 13537 7304 35499 7306
rect 13537 7248 13542 7304
rect 13598 7248 35438 7304
rect 35494 7248 35499 7304
rect 13537 7246 35499 7248
rect 13537 7243 13603 7246
rect 35433 7243 35499 7246
rect 14825 7170 14891 7173
rect 15837 7170 15903 7173
rect 24209 7170 24275 7173
rect 14825 7168 24275 7170
rect 14825 7112 14830 7168
rect 14886 7112 15842 7168
rect 15898 7112 24214 7168
rect 24270 7112 24275 7168
rect 14825 7110 24275 7112
rect 14825 7107 14891 7110
rect 15837 7107 15903 7110
rect 24209 7107 24275 7110
rect 14277 7104 14597 7105
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 7039 14597 7040
rect 27610 7104 27930 7105
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 7039 27930 7040
rect 16941 7034 17007 7037
rect 24301 7034 24367 7037
rect 16941 7032 24367 7034
rect 16941 6976 16946 7032
rect 17002 6976 24306 7032
rect 24362 6976 24367 7032
rect 16941 6974 24367 6976
rect 16941 6971 17007 6974
rect 24301 6971 24367 6974
rect 9121 6898 9187 6901
rect 11881 6898 11947 6901
rect 9121 6896 11947 6898
rect 9121 6840 9126 6896
rect 9182 6840 11886 6896
rect 11942 6840 11947 6896
rect 9121 6838 11947 6840
rect 9121 6835 9187 6838
rect 11881 6835 11947 6838
rect 12065 6898 12131 6901
rect 19701 6898 19767 6901
rect 12065 6896 19767 6898
rect 12065 6840 12070 6896
rect 12126 6840 19706 6896
rect 19762 6840 19767 6896
rect 12065 6838 19767 6840
rect 12065 6835 12131 6838
rect 19701 6835 19767 6838
rect 4153 6762 4219 6765
rect 7557 6762 7623 6765
rect 4153 6760 7623 6762
rect 4153 6704 4158 6760
rect 4214 6704 7562 6760
rect 7618 6704 7623 6760
rect 4153 6702 7623 6704
rect 4153 6699 4219 6702
rect 7557 6699 7623 6702
rect 7610 6560 7930 6561
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7930 6560
rect 7610 6495 7930 6496
rect 20944 6560 21264 6561
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 6495 21264 6496
rect 34277 6560 34597 6561
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 6495 34597 6496
rect 7557 6354 7623 6357
rect 13629 6354 13695 6357
rect 15745 6354 15811 6357
rect 7557 6352 15811 6354
rect 7557 6296 7562 6352
rect 7618 6296 13634 6352
rect 13690 6296 15750 6352
rect 15806 6296 15811 6352
rect 7557 6294 15811 6296
rect 7557 6291 7623 6294
rect 13629 6291 13695 6294
rect 15745 6291 15811 6294
rect 17309 6354 17375 6357
rect 20437 6354 20503 6357
rect 27705 6354 27771 6357
rect 17309 6352 20503 6354
rect 17309 6296 17314 6352
rect 17370 6296 20442 6352
rect 20498 6296 20503 6352
rect 17309 6294 20503 6296
rect 17309 6291 17375 6294
rect 20437 6291 20503 6294
rect 20670 6352 27771 6354
rect 20670 6296 27710 6352
rect 27766 6296 27771 6352
rect 20670 6294 27771 6296
rect 0 6218 800 6248
rect 20670 6218 20730 6294
rect 27705 6291 27771 6294
rect 0 6158 20730 6218
rect 22277 6218 22343 6221
rect 25589 6218 25655 6221
rect 22277 6216 25655 6218
rect 22277 6160 22282 6216
rect 22338 6160 25594 6216
rect 25650 6160 25655 6216
rect 22277 6158 25655 6160
rect 0 6128 800 6158
rect 22277 6155 22343 6158
rect 25589 6155 25655 6158
rect 34605 6218 34671 6221
rect 39200 6218 40000 6248
rect 34605 6216 40000 6218
rect 34605 6160 34610 6216
rect 34666 6160 40000 6216
rect 34605 6158 40000 6160
rect 34605 6155 34671 6158
rect 39200 6128 40000 6158
rect 2037 6082 2103 6085
rect 11329 6082 11395 6085
rect 2037 6080 11395 6082
rect 2037 6024 2042 6080
rect 2098 6024 11334 6080
rect 11390 6024 11395 6080
rect 2037 6022 11395 6024
rect 2037 6019 2103 6022
rect 11329 6019 11395 6022
rect 16389 6082 16455 6085
rect 19793 6082 19859 6085
rect 16389 6080 19859 6082
rect 16389 6024 16394 6080
rect 16450 6024 19798 6080
rect 19854 6024 19859 6080
rect 16389 6022 19859 6024
rect 16389 6019 16455 6022
rect 19793 6019 19859 6022
rect 14277 6016 14597 6017
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 5951 14597 5952
rect 27610 6016 27930 6017
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 5951 27930 5952
rect 6177 5946 6243 5949
rect 12709 5946 12775 5949
rect 6177 5944 12775 5946
rect 6177 5888 6182 5944
rect 6238 5888 12714 5944
rect 12770 5888 12775 5944
rect 6177 5886 12775 5888
rect 6177 5883 6243 5886
rect 12709 5883 12775 5886
rect 12985 5810 13051 5813
rect 16665 5810 16731 5813
rect 19425 5810 19491 5813
rect 12985 5808 19491 5810
rect 12985 5752 12990 5808
rect 13046 5752 16670 5808
rect 16726 5752 19430 5808
rect 19486 5752 19491 5808
rect 12985 5750 19491 5752
rect 12985 5747 13051 5750
rect 16665 5747 16731 5750
rect 19425 5747 19491 5750
rect 21817 5810 21883 5813
rect 24117 5810 24183 5813
rect 21817 5808 24183 5810
rect 21817 5752 21822 5808
rect 21878 5752 24122 5808
rect 24178 5752 24183 5808
rect 21817 5750 24183 5752
rect 21817 5747 21883 5750
rect 24117 5747 24183 5750
rect 2497 5674 2563 5677
rect 4521 5674 4587 5677
rect 2497 5672 4587 5674
rect 2497 5616 2502 5672
rect 2558 5616 4526 5672
rect 4582 5616 4587 5672
rect 2497 5614 4587 5616
rect 2497 5611 2563 5614
rect 4521 5611 4587 5614
rect 21449 5674 21515 5677
rect 23841 5674 23907 5677
rect 21449 5672 23907 5674
rect 21449 5616 21454 5672
rect 21510 5616 23846 5672
rect 23902 5616 23907 5672
rect 21449 5614 23907 5616
rect 21449 5611 21515 5614
rect 23841 5611 23907 5614
rect 12801 5538 12867 5541
rect 17217 5538 17283 5541
rect 12801 5536 17283 5538
rect 12801 5480 12806 5536
rect 12862 5480 17222 5536
rect 17278 5480 17283 5536
rect 12801 5478 17283 5480
rect 12801 5475 12867 5478
rect 17217 5475 17283 5478
rect 7610 5472 7930 5473
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7930 5472
rect 7610 5407 7930 5408
rect 20944 5472 21264 5473
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 5407 21264 5408
rect 34277 5472 34597 5473
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 5407 34597 5408
rect 3325 5402 3391 5405
rect 5533 5402 5599 5405
rect 3325 5400 5599 5402
rect 3325 5344 3330 5400
rect 3386 5344 5538 5400
rect 5594 5344 5599 5400
rect 3325 5342 5599 5344
rect 3325 5339 3391 5342
rect 5533 5339 5599 5342
rect 3877 5266 3943 5269
rect 14365 5266 14431 5269
rect 17125 5266 17191 5269
rect 20713 5266 20779 5269
rect 25681 5266 25747 5269
rect 3877 5264 11530 5266
rect 3877 5208 3882 5264
rect 3938 5208 11530 5264
rect 3877 5206 11530 5208
rect 3877 5203 3943 5206
rect 9489 5130 9555 5133
rect 10225 5130 10291 5133
rect 11237 5130 11303 5133
rect 9489 5128 11303 5130
rect 9489 5072 9494 5128
rect 9550 5072 10230 5128
rect 10286 5072 11242 5128
rect 11298 5072 11303 5128
rect 9489 5070 11303 5072
rect 11470 5130 11530 5206
rect 14365 5264 25747 5266
rect 14365 5208 14370 5264
rect 14426 5208 17130 5264
rect 17186 5208 20718 5264
rect 20774 5208 25686 5264
rect 25742 5208 25747 5264
rect 14365 5206 25747 5208
rect 14365 5203 14431 5206
rect 17125 5203 17191 5206
rect 20713 5203 20779 5206
rect 25681 5203 25747 5206
rect 29729 5130 29795 5133
rect 33225 5130 33291 5133
rect 11470 5128 33291 5130
rect 11470 5072 29734 5128
rect 29790 5072 33230 5128
rect 33286 5072 33291 5128
rect 11470 5070 33291 5072
rect 9489 5067 9555 5070
rect 10225 5067 10291 5070
rect 11237 5067 11303 5070
rect 29729 5067 29795 5070
rect 33225 5067 33291 5070
rect 2037 4994 2103 4997
rect 10869 4994 10935 4997
rect 14089 4994 14155 4997
rect 2037 4992 7666 4994
rect 2037 4936 2042 4992
rect 2098 4936 7666 4992
rect 2037 4934 7666 4936
rect 2037 4931 2103 4934
rect 0 4858 800 4888
rect 7606 4858 7666 4934
rect 10869 4992 14155 4994
rect 10869 4936 10874 4992
rect 10930 4936 14094 4992
rect 14150 4936 14155 4992
rect 10869 4934 14155 4936
rect 10869 4931 10935 4934
rect 14089 4931 14155 4934
rect 14277 4928 14597 4929
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 4863 14597 4864
rect 27610 4928 27930 4929
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 4863 27930 4864
rect 34697 4858 34763 4861
rect 39200 4858 40000 4888
rect 0 4798 5274 4858
rect 7606 4798 14106 4858
rect 0 4768 800 4798
rect 5214 4178 5274 4798
rect 6269 4722 6335 4725
rect 7281 4722 7347 4725
rect 10869 4722 10935 4725
rect 6269 4720 10935 4722
rect 6269 4664 6274 4720
rect 6330 4664 7286 4720
rect 7342 4664 10874 4720
rect 10930 4664 10935 4720
rect 6269 4662 10935 4664
rect 6269 4659 6335 4662
rect 7281 4659 7347 4662
rect 10869 4659 10935 4662
rect 5349 4586 5415 4589
rect 9121 4586 9187 4589
rect 5349 4584 9187 4586
rect 5349 4528 5354 4584
rect 5410 4528 9126 4584
rect 9182 4528 9187 4584
rect 5349 4526 9187 4528
rect 14046 4586 14106 4798
rect 34697 4856 40000 4858
rect 34697 4800 34702 4856
rect 34758 4800 40000 4856
rect 34697 4798 40000 4800
rect 34697 4795 34763 4798
rect 39200 4768 40000 4798
rect 24393 4586 24459 4589
rect 34605 4586 34671 4589
rect 14046 4526 21466 4586
rect 5349 4523 5415 4526
rect 9121 4523 9187 4526
rect 21406 4450 21466 4526
rect 24393 4584 34671 4586
rect 24393 4528 24398 4584
rect 24454 4528 34610 4584
rect 34666 4528 34671 4584
rect 24393 4526 34671 4528
rect 24393 4523 24459 4526
rect 34605 4523 34671 4526
rect 27061 4450 27127 4453
rect 21406 4448 27127 4450
rect 21406 4392 27066 4448
rect 27122 4392 27127 4448
rect 21406 4390 27127 4392
rect 27061 4387 27127 4390
rect 7610 4384 7930 4385
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7930 4384
rect 7610 4319 7930 4320
rect 20944 4384 21264 4385
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 4319 21264 4320
rect 34277 4384 34597 4385
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 4319 34597 4320
rect 28625 4314 28691 4317
rect 30373 4314 30439 4317
rect 28625 4312 30439 4314
rect 28625 4256 28630 4312
rect 28686 4256 30378 4312
rect 30434 4256 30439 4312
rect 28625 4254 30439 4256
rect 28625 4251 28691 4254
rect 30373 4251 30439 4254
rect 20897 4178 20963 4181
rect 5214 4176 20963 4178
rect 5214 4120 20902 4176
rect 20958 4120 20963 4176
rect 5214 4118 20963 4120
rect 20897 4115 20963 4118
rect 21265 4178 21331 4181
rect 26601 4178 26667 4181
rect 21265 4176 26667 4178
rect 21265 4120 21270 4176
rect 21326 4120 26606 4176
rect 26662 4120 26667 4176
rect 21265 4118 26667 4120
rect 21265 4115 21331 4118
rect 26601 4115 26667 4118
rect 5257 4042 5323 4045
rect 7097 4042 7163 4045
rect 30833 4042 30899 4045
rect 37733 4042 37799 4045
rect 5257 4040 7163 4042
rect 5257 3984 5262 4040
rect 5318 3984 7102 4040
rect 7158 3984 7163 4040
rect 5257 3982 7163 3984
rect 5257 3979 5323 3982
rect 7097 3979 7163 3982
rect 14966 4040 37799 4042
rect 14966 3984 30838 4040
rect 30894 3984 37738 4040
rect 37794 3984 37799 4040
rect 14966 3982 37799 3984
rect 4705 3906 4771 3909
rect 8569 3906 8635 3909
rect 12525 3906 12591 3909
rect 4705 3904 12591 3906
rect 4705 3848 4710 3904
rect 4766 3848 8574 3904
rect 8630 3848 12530 3904
rect 12586 3848 12591 3904
rect 4705 3846 12591 3848
rect 4705 3843 4771 3846
rect 8569 3843 8635 3846
rect 12525 3843 12591 3846
rect 14277 3840 14597 3841
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 3775 14597 3776
rect 13 3770 79 3773
rect 8937 3770 9003 3773
rect 13 3768 9003 3770
rect 13 3712 18 3768
rect 74 3712 8942 3768
rect 8998 3712 9003 3768
rect 13 3710 9003 3712
rect 13 3707 79 3710
rect 8937 3707 9003 3710
rect 14181 3634 14247 3637
rect 798 3632 14247 3634
rect 798 3576 14186 3632
rect 14242 3576 14247 3632
rect 798 3574 14247 3576
rect 798 3528 858 3574
rect 14181 3571 14247 3574
rect 0 3438 858 3528
rect 14966 3498 15026 3982
rect 30833 3979 30899 3982
rect 37733 3979 37799 3982
rect 38653 3906 38719 3909
rect 30974 3904 38719 3906
rect 30974 3848 38658 3904
rect 38714 3848 38719 3904
rect 30974 3846 38719 3848
rect 27610 3840 27930 3841
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 3775 27930 3776
rect 15101 3770 15167 3773
rect 17217 3770 17283 3773
rect 15101 3768 17283 3770
rect 15101 3712 15106 3768
rect 15162 3712 17222 3768
rect 17278 3712 17283 3768
rect 15101 3710 17283 3712
rect 15101 3707 15167 3710
rect 17217 3707 17283 3710
rect 19701 3634 19767 3637
rect 30974 3634 31034 3846
rect 38653 3843 38719 3846
rect 31109 3770 31175 3773
rect 34697 3770 34763 3773
rect 31109 3768 34763 3770
rect 31109 3712 31114 3768
rect 31170 3712 34702 3768
rect 34758 3712 34763 3768
rect 31109 3710 34763 3712
rect 31109 3707 31175 3710
rect 34697 3707 34763 3710
rect 34881 3770 34947 3773
rect 36813 3770 36879 3773
rect 34881 3768 36879 3770
rect 34881 3712 34886 3768
rect 34942 3712 36818 3768
rect 36874 3712 36879 3768
rect 34881 3710 36879 3712
rect 34881 3707 34947 3710
rect 36813 3707 36879 3710
rect 19701 3632 31034 3634
rect 19701 3576 19706 3632
rect 19762 3576 31034 3632
rect 19701 3574 31034 3576
rect 19701 3571 19767 3574
rect 7422 3438 15026 3498
rect 15469 3498 15535 3501
rect 34421 3498 34487 3501
rect 15469 3496 34487 3498
rect 15469 3440 15474 3496
rect 15530 3440 34426 3496
rect 34482 3440 34487 3496
rect 15469 3438 34487 3440
rect 0 3408 800 3438
rect 2037 3362 2103 3365
rect 7422 3362 7482 3438
rect 15469 3435 15535 3438
rect 34421 3435 34487 3438
rect 34605 3498 34671 3501
rect 39200 3498 40000 3528
rect 34605 3496 40000 3498
rect 34605 3440 34610 3496
rect 34666 3440 40000 3496
rect 34605 3438 40000 3440
rect 34605 3435 34671 3438
rect 39200 3408 40000 3438
rect 2037 3360 7482 3362
rect 2037 3304 2042 3360
rect 2098 3304 7482 3360
rect 2037 3302 7482 3304
rect 9857 3362 9923 3365
rect 10317 3362 10383 3365
rect 15377 3362 15443 3365
rect 31109 3362 31175 3365
rect 9857 3360 15443 3362
rect 9857 3304 9862 3360
rect 9918 3304 10322 3360
rect 10378 3304 15382 3360
rect 15438 3304 15443 3360
rect 9857 3302 15443 3304
rect 2037 3299 2103 3302
rect 9857 3299 9923 3302
rect 10317 3299 10383 3302
rect 15377 3299 15443 3302
rect 26926 3360 31175 3362
rect 26926 3304 31114 3360
rect 31170 3304 31175 3360
rect 26926 3302 31175 3304
rect 7610 3296 7930 3297
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7930 3296
rect 7610 3231 7930 3232
rect 20944 3296 21264 3297
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 20944 3231 21264 3232
rect 8937 3226 9003 3229
rect 11881 3226 11947 3229
rect 8937 3224 11947 3226
rect 8937 3168 8942 3224
rect 8998 3168 11886 3224
rect 11942 3168 11947 3224
rect 8937 3166 11947 3168
rect 8937 3163 9003 3166
rect 11881 3163 11947 3166
rect 15101 3226 15167 3229
rect 17401 3226 17467 3229
rect 15101 3224 17467 3226
rect 15101 3168 15106 3224
rect 15162 3168 17406 3224
rect 17462 3168 17467 3224
rect 15101 3166 17467 3168
rect 15101 3163 15167 3166
rect 17401 3163 17467 3166
rect 5533 3090 5599 3093
rect 11789 3090 11855 3093
rect 26926 3090 26986 3302
rect 31109 3299 31175 3302
rect 34277 3296 34597 3297
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 3231 34597 3232
rect 27061 3226 27127 3229
rect 32581 3226 32647 3229
rect 27061 3224 32647 3226
rect 27061 3168 27066 3224
rect 27122 3168 32586 3224
rect 32642 3168 32647 3224
rect 27061 3166 32647 3168
rect 27061 3163 27127 3166
rect 32581 3163 32647 3166
rect 5533 3088 7666 3090
rect 5533 3032 5538 3088
rect 5594 3032 7666 3088
rect 5533 3030 7666 3032
rect 5533 3027 5599 3030
rect 4153 2954 4219 2957
rect 2822 2952 4219 2954
rect 2822 2896 4158 2952
rect 4214 2896 4219 2952
rect 2822 2894 4219 2896
rect 933 2818 999 2821
rect 2822 2818 2882 2894
rect 4153 2891 4219 2894
rect 4337 2954 4403 2957
rect 7373 2954 7439 2957
rect 4337 2952 7439 2954
rect 4337 2896 4342 2952
rect 4398 2896 7378 2952
rect 7434 2896 7439 2952
rect 4337 2894 7439 2896
rect 4337 2891 4403 2894
rect 7373 2891 7439 2894
rect 933 2816 2882 2818
rect 933 2760 938 2816
rect 994 2760 2882 2816
rect 933 2758 2882 2760
rect 3049 2818 3115 2821
rect 6453 2818 6519 2821
rect 3049 2816 6519 2818
rect 3049 2760 3054 2816
rect 3110 2760 6458 2816
rect 6514 2760 6519 2816
rect 3049 2758 6519 2760
rect 7606 2818 7666 3030
rect 11789 3088 26986 3090
rect 11789 3032 11794 3088
rect 11850 3032 26986 3088
rect 11789 3030 26986 3032
rect 29729 3090 29795 3093
rect 32213 3090 32279 3093
rect 29729 3088 32279 3090
rect 29729 3032 29734 3088
rect 29790 3032 32218 3088
rect 32274 3032 32279 3088
rect 29729 3030 32279 3032
rect 11789 3027 11855 3030
rect 29729 3027 29795 3030
rect 32213 3027 32279 3030
rect 35893 3092 35959 3093
rect 35893 3088 35940 3092
rect 36004 3090 36010 3092
rect 35893 3032 35898 3088
rect 35893 3028 35940 3032
rect 36004 3030 36050 3090
rect 36004 3028 36010 3030
rect 35893 3027 35959 3028
rect 9489 2954 9555 2957
rect 15469 2954 15535 2957
rect 9489 2952 15535 2954
rect 9489 2896 9494 2952
rect 9550 2896 15474 2952
rect 15530 2896 15535 2952
rect 9489 2894 15535 2896
rect 9489 2891 9555 2894
rect 15469 2891 15535 2894
rect 16665 2954 16731 2957
rect 23289 2954 23355 2957
rect 16665 2952 23355 2954
rect 16665 2896 16670 2952
rect 16726 2896 23294 2952
rect 23350 2896 23355 2952
rect 16665 2894 23355 2896
rect 16665 2891 16731 2894
rect 23289 2891 23355 2894
rect 28257 2954 28323 2957
rect 30373 2954 30439 2957
rect 28257 2952 30439 2954
rect 28257 2896 28262 2952
rect 28318 2896 30378 2952
rect 30434 2896 30439 2952
rect 28257 2894 30439 2896
rect 28257 2891 28323 2894
rect 30373 2891 30439 2894
rect 31569 2954 31635 2957
rect 34053 2954 34119 2957
rect 31569 2952 34119 2954
rect 31569 2896 31574 2952
rect 31630 2896 34058 2952
rect 34114 2896 34119 2952
rect 31569 2894 34119 2896
rect 31569 2891 31635 2894
rect 34053 2891 34119 2894
rect 13537 2818 13603 2821
rect 14733 2820 14799 2821
rect 14733 2818 14780 2820
rect 7606 2816 13603 2818
rect 7606 2760 13542 2816
rect 13598 2760 13603 2816
rect 7606 2758 13603 2760
rect 14688 2816 14780 2818
rect 14688 2760 14738 2816
rect 14688 2758 14780 2760
rect 933 2755 999 2758
rect 3049 2755 3115 2758
rect 6453 2755 6519 2758
rect 13537 2755 13603 2758
rect 14733 2756 14780 2758
rect 14844 2756 14850 2820
rect 28717 2818 28783 2821
rect 31293 2818 31359 2821
rect 28717 2816 31359 2818
rect 28717 2760 28722 2816
rect 28778 2760 31298 2816
rect 31354 2760 31359 2816
rect 28717 2758 31359 2760
rect 14733 2755 14799 2756
rect 28717 2755 28783 2758
rect 31293 2755 31359 2758
rect 32765 2818 32831 2821
rect 34973 2818 35039 2821
rect 32765 2816 35039 2818
rect 32765 2760 32770 2816
rect 32826 2760 34978 2816
rect 35034 2760 35039 2816
rect 32765 2758 35039 2760
rect 32765 2755 32831 2758
rect 34973 2755 35039 2758
rect 14277 2752 14597 2753
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2687 14597 2688
rect 27610 2752 27930 2753
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2687 27930 2688
rect 14917 2682 14983 2685
rect 17033 2682 17099 2685
rect 23289 2682 23355 2685
rect 14917 2680 17099 2682
rect 14917 2624 14922 2680
rect 14978 2624 17038 2680
rect 17094 2624 17099 2680
rect 14917 2622 17099 2624
rect 14917 2619 14983 2622
rect 17033 2619 17099 2622
rect 17174 2680 23355 2682
rect 17174 2624 23294 2680
rect 23350 2624 23355 2680
rect 17174 2622 23355 2624
rect 10409 2546 10475 2549
rect 17174 2546 17234 2622
rect 23289 2619 23355 2622
rect 10409 2544 17234 2546
rect 10409 2488 10414 2544
rect 10470 2488 17234 2544
rect 10409 2486 17234 2488
rect 17309 2546 17375 2549
rect 30281 2546 30347 2549
rect 17309 2544 30347 2546
rect 17309 2488 17314 2544
rect 17370 2488 30286 2544
rect 30342 2488 30347 2544
rect 17309 2486 30347 2488
rect 10409 2483 10475 2486
rect 17309 2483 17375 2486
rect 30281 2483 30347 2486
rect 3509 2410 3575 2413
rect 27613 2410 27679 2413
rect 39573 2410 39639 2413
rect 3509 2408 39639 2410
rect 3509 2352 3514 2408
rect 3570 2352 27618 2408
rect 27674 2352 39578 2408
rect 39634 2352 39639 2408
rect 3509 2350 39639 2352
rect 3509 2347 3575 2350
rect 27613 2347 27679 2350
rect 39573 2347 39639 2350
rect 8385 2274 8451 2277
rect 15193 2274 15259 2277
rect 8385 2272 15259 2274
rect 8385 2216 8390 2272
rect 8446 2216 15198 2272
rect 15254 2216 15259 2272
rect 8385 2214 15259 2216
rect 8385 2211 8451 2214
rect 15193 2211 15259 2214
rect 15377 2274 15443 2277
rect 20437 2274 20503 2277
rect 15377 2272 20503 2274
rect 15377 2216 15382 2272
rect 15438 2216 20442 2272
rect 20498 2216 20503 2272
rect 15377 2214 20503 2216
rect 15377 2211 15443 2214
rect 20437 2211 20503 2214
rect 21725 2274 21791 2277
rect 28533 2274 28599 2277
rect 21725 2272 28599 2274
rect 21725 2216 21730 2272
rect 21786 2216 28538 2272
rect 28594 2216 28599 2272
rect 21725 2214 28599 2216
rect 21725 2211 21791 2214
rect 28533 2211 28599 2214
rect 7610 2208 7930 2209
rect 0 2138 800 2168
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7930 2208
rect 7610 2143 7930 2144
rect 20944 2208 21264 2209
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2143 21264 2144
rect 34277 2208 34597 2209
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2143 34597 2144
rect 6085 2138 6151 2141
rect 0 2136 6151 2138
rect 0 2080 6090 2136
rect 6146 2080 6151 2136
rect 0 2078 6151 2080
rect 0 2048 800 2078
rect 6085 2075 6151 2078
rect 12065 2138 12131 2141
rect 16573 2138 16639 2141
rect 12065 2136 16639 2138
rect 12065 2080 12070 2136
rect 12126 2080 16578 2136
rect 16634 2080 16639 2136
rect 12065 2078 16639 2080
rect 12065 2075 12131 2078
rect 16573 2075 16639 2078
rect 34697 2138 34763 2141
rect 39200 2138 40000 2168
rect 34697 2136 40000 2138
rect 34697 2080 34702 2136
rect 34758 2080 40000 2136
rect 34697 2078 40000 2080
rect 34697 2075 34763 2078
rect 39200 2048 40000 2078
rect 2773 2002 2839 2005
rect 16665 2002 16731 2005
rect 2773 2000 16731 2002
rect 2773 1944 2778 2000
rect 2834 1944 16670 2000
rect 16726 1944 16731 2000
rect 2773 1942 16731 1944
rect 2773 1939 2839 1942
rect 16665 1939 16731 1942
rect 23289 2002 23355 2005
rect 34605 2002 34671 2005
rect 23289 2000 34671 2002
rect 23289 1944 23294 2000
rect 23350 1944 34610 2000
rect 34666 1944 34671 2000
rect 23289 1942 34671 1944
rect 23289 1939 23355 1942
rect 34605 1939 34671 1942
rect 12525 1866 12591 1869
rect 29545 1866 29611 1869
rect 12525 1864 29611 1866
rect 12525 1808 12530 1864
rect 12586 1808 29550 1864
rect 29606 1808 29611 1864
rect 12525 1806 29611 1808
rect 12525 1803 12591 1806
rect 29545 1803 29611 1806
rect 4797 1730 4863 1733
rect 7189 1730 7255 1733
rect 19149 1730 19215 1733
rect 4797 1728 19215 1730
rect 4797 1672 4802 1728
rect 4858 1672 7194 1728
rect 7250 1672 19154 1728
rect 19210 1672 19215 1728
rect 4797 1670 19215 1672
rect 4797 1667 4863 1670
rect 7189 1667 7255 1670
rect 19149 1667 19215 1670
rect 20437 1730 20503 1733
rect 31385 1730 31451 1733
rect 20437 1728 31451 1730
rect 20437 1672 20442 1728
rect 20498 1672 31390 1728
rect 31446 1672 31451 1728
rect 20437 1670 31451 1672
rect 20437 1667 20503 1670
rect 31385 1667 31451 1670
rect 6085 1594 6151 1597
rect 12433 1594 12499 1597
rect 6085 1592 12499 1594
rect 6085 1536 6090 1592
rect 6146 1536 12438 1592
rect 12494 1536 12499 1592
rect 6085 1534 12499 1536
rect 6085 1531 6151 1534
rect 12433 1531 12499 1534
rect 28942 1458 28948 1460
rect 22142 1398 28948 1458
rect 11881 1322 11947 1325
rect 22142 1322 22202 1398
rect 28942 1396 28948 1398
rect 29012 1396 29018 1460
rect 11881 1320 22202 1322
rect 11881 1264 11886 1320
rect 11942 1264 22202 1320
rect 11881 1262 22202 1264
rect 11881 1259 11947 1262
rect 28942 1124 28948 1188
rect 29012 1186 29018 1188
rect 34697 1186 34763 1189
rect 29012 1184 34763 1186
rect 29012 1128 34702 1184
rect 34758 1128 34763 1184
rect 29012 1126 34763 1128
rect 29012 1124 29018 1126
rect 34697 1123 34763 1126
rect 0 778 800 808
rect 1393 778 1459 781
rect 0 776 1459 778
rect 0 720 1398 776
rect 1454 720 1459 776
rect 0 718 1459 720
rect 0 688 800 718
rect 1393 715 1459 718
rect 28942 716 28948 780
rect 29012 778 29018 780
rect 39200 778 40000 808
rect 29012 718 40000 778
rect 29012 716 29018 718
rect 39200 688 40000 718
rect 28942 234 28948 236
rect 19244 174 28948 234
rect 19244 101 19304 174
rect 28942 172 28948 174
rect 29012 172 29018 236
rect 19241 96 19307 101
rect 19241 40 19246 96
rect 19302 40 19307 96
rect 19241 35 19307 40
<< via3 >>
rect 14285 13628 14349 13632
rect 14285 13572 14289 13628
rect 14289 13572 14345 13628
rect 14345 13572 14349 13628
rect 14285 13568 14349 13572
rect 14365 13628 14429 13632
rect 14365 13572 14369 13628
rect 14369 13572 14425 13628
rect 14425 13572 14429 13628
rect 14365 13568 14429 13572
rect 14445 13628 14509 13632
rect 14445 13572 14449 13628
rect 14449 13572 14505 13628
rect 14505 13572 14509 13628
rect 14445 13568 14509 13572
rect 14525 13628 14589 13632
rect 14525 13572 14529 13628
rect 14529 13572 14585 13628
rect 14585 13572 14589 13628
rect 14525 13568 14589 13572
rect 27618 13628 27682 13632
rect 27618 13572 27622 13628
rect 27622 13572 27678 13628
rect 27678 13572 27682 13628
rect 27618 13568 27682 13572
rect 27698 13628 27762 13632
rect 27698 13572 27702 13628
rect 27702 13572 27758 13628
rect 27758 13572 27762 13628
rect 27698 13568 27762 13572
rect 27778 13628 27842 13632
rect 27778 13572 27782 13628
rect 27782 13572 27838 13628
rect 27838 13572 27842 13628
rect 27778 13568 27842 13572
rect 27858 13628 27922 13632
rect 27858 13572 27862 13628
rect 27862 13572 27918 13628
rect 27918 13572 27922 13628
rect 27858 13568 27922 13572
rect 7618 13084 7682 13088
rect 7618 13028 7622 13084
rect 7622 13028 7678 13084
rect 7678 13028 7682 13084
rect 7618 13024 7682 13028
rect 7698 13084 7762 13088
rect 7698 13028 7702 13084
rect 7702 13028 7758 13084
rect 7758 13028 7762 13084
rect 7698 13024 7762 13028
rect 7778 13084 7842 13088
rect 7778 13028 7782 13084
rect 7782 13028 7838 13084
rect 7838 13028 7842 13084
rect 7778 13024 7842 13028
rect 7858 13084 7922 13088
rect 7858 13028 7862 13084
rect 7862 13028 7918 13084
rect 7918 13028 7922 13084
rect 7858 13024 7922 13028
rect 20952 13084 21016 13088
rect 20952 13028 20956 13084
rect 20956 13028 21012 13084
rect 21012 13028 21016 13084
rect 20952 13024 21016 13028
rect 21032 13084 21096 13088
rect 21032 13028 21036 13084
rect 21036 13028 21092 13084
rect 21092 13028 21096 13084
rect 21032 13024 21096 13028
rect 21112 13084 21176 13088
rect 21112 13028 21116 13084
rect 21116 13028 21172 13084
rect 21172 13028 21176 13084
rect 21112 13024 21176 13028
rect 21192 13084 21256 13088
rect 21192 13028 21196 13084
rect 21196 13028 21252 13084
rect 21252 13028 21256 13084
rect 21192 13024 21256 13028
rect 34285 13084 34349 13088
rect 34285 13028 34289 13084
rect 34289 13028 34345 13084
rect 34345 13028 34349 13084
rect 34285 13024 34349 13028
rect 34365 13084 34429 13088
rect 34365 13028 34369 13084
rect 34369 13028 34425 13084
rect 34425 13028 34429 13084
rect 34365 13024 34429 13028
rect 34445 13084 34509 13088
rect 34445 13028 34449 13084
rect 34449 13028 34505 13084
rect 34505 13028 34509 13084
rect 34445 13024 34509 13028
rect 34525 13084 34589 13088
rect 34525 13028 34529 13084
rect 34529 13028 34585 13084
rect 34585 13028 34589 13084
rect 34525 13024 34589 13028
rect 14285 12540 14349 12544
rect 14285 12484 14289 12540
rect 14289 12484 14345 12540
rect 14345 12484 14349 12540
rect 14285 12480 14349 12484
rect 14365 12540 14429 12544
rect 14365 12484 14369 12540
rect 14369 12484 14425 12540
rect 14425 12484 14429 12540
rect 14365 12480 14429 12484
rect 14445 12540 14509 12544
rect 14445 12484 14449 12540
rect 14449 12484 14505 12540
rect 14505 12484 14509 12540
rect 14445 12480 14509 12484
rect 14525 12540 14589 12544
rect 14525 12484 14529 12540
rect 14529 12484 14585 12540
rect 14585 12484 14589 12540
rect 14525 12480 14589 12484
rect 27618 12540 27682 12544
rect 27618 12484 27622 12540
rect 27622 12484 27678 12540
rect 27678 12484 27682 12540
rect 27618 12480 27682 12484
rect 27698 12540 27762 12544
rect 27698 12484 27702 12540
rect 27702 12484 27758 12540
rect 27758 12484 27762 12540
rect 27698 12480 27762 12484
rect 27778 12540 27842 12544
rect 27778 12484 27782 12540
rect 27782 12484 27838 12540
rect 27838 12484 27842 12540
rect 27778 12480 27842 12484
rect 27858 12540 27922 12544
rect 27858 12484 27862 12540
rect 27862 12484 27918 12540
rect 27918 12484 27922 12540
rect 27858 12480 27922 12484
rect 7618 11996 7682 12000
rect 7618 11940 7622 11996
rect 7622 11940 7678 11996
rect 7678 11940 7682 11996
rect 7618 11936 7682 11940
rect 7698 11996 7762 12000
rect 7698 11940 7702 11996
rect 7702 11940 7758 11996
rect 7758 11940 7762 11996
rect 7698 11936 7762 11940
rect 7778 11996 7842 12000
rect 7778 11940 7782 11996
rect 7782 11940 7838 11996
rect 7838 11940 7842 11996
rect 7778 11936 7842 11940
rect 7858 11996 7922 12000
rect 7858 11940 7862 11996
rect 7862 11940 7918 11996
rect 7918 11940 7922 11996
rect 7858 11936 7922 11940
rect 20952 11996 21016 12000
rect 20952 11940 20956 11996
rect 20956 11940 21012 11996
rect 21012 11940 21016 11996
rect 20952 11936 21016 11940
rect 21032 11996 21096 12000
rect 21032 11940 21036 11996
rect 21036 11940 21092 11996
rect 21092 11940 21096 11996
rect 21032 11936 21096 11940
rect 21112 11996 21176 12000
rect 21112 11940 21116 11996
rect 21116 11940 21172 11996
rect 21172 11940 21176 11996
rect 21112 11936 21176 11940
rect 21192 11996 21256 12000
rect 21192 11940 21196 11996
rect 21196 11940 21252 11996
rect 21252 11940 21256 11996
rect 21192 11936 21256 11940
rect 34285 11996 34349 12000
rect 34285 11940 34289 11996
rect 34289 11940 34345 11996
rect 34345 11940 34349 11996
rect 34285 11936 34349 11940
rect 34365 11996 34429 12000
rect 34365 11940 34369 11996
rect 34369 11940 34425 11996
rect 34425 11940 34429 11996
rect 34365 11936 34429 11940
rect 34445 11996 34509 12000
rect 34445 11940 34449 11996
rect 34449 11940 34505 11996
rect 34505 11940 34509 11996
rect 34445 11936 34509 11940
rect 34525 11996 34589 12000
rect 34525 11940 34529 11996
rect 34529 11940 34585 11996
rect 34585 11940 34589 11996
rect 34525 11936 34589 11940
rect 14285 11452 14349 11456
rect 14285 11396 14289 11452
rect 14289 11396 14345 11452
rect 14345 11396 14349 11452
rect 14285 11392 14349 11396
rect 14365 11452 14429 11456
rect 14365 11396 14369 11452
rect 14369 11396 14425 11452
rect 14425 11396 14429 11452
rect 14365 11392 14429 11396
rect 14445 11452 14509 11456
rect 14445 11396 14449 11452
rect 14449 11396 14505 11452
rect 14505 11396 14509 11452
rect 14445 11392 14509 11396
rect 14525 11452 14589 11456
rect 14525 11396 14529 11452
rect 14529 11396 14585 11452
rect 14585 11396 14589 11452
rect 14525 11392 14589 11396
rect 27618 11452 27682 11456
rect 27618 11396 27622 11452
rect 27622 11396 27678 11452
rect 27678 11396 27682 11452
rect 27618 11392 27682 11396
rect 27698 11452 27762 11456
rect 27698 11396 27702 11452
rect 27702 11396 27758 11452
rect 27758 11396 27762 11452
rect 27698 11392 27762 11396
rect 27778 11452 27842 11456
rect 27778 11396 27782 11452
rect 27782 11396 27838 11452
rect 27838 11396 27842 11452
rect 27778 11392 27842 11396
rect 27858 11452 27922 11456
rect 27858 11396 27862 11452
rect 27862 11396 27918 11452
rect 27918 11396 27922 11452
rect 27858 11392 27922 11396
rect 7618 10908 7682 10912
rect 7618 10852 7622 10908
rect 7622 10852 7678 10908
rect 7678 10852 7682 10908
rect 7618 10848 7682 10852
rect 7698 10908 7762 10912
rect 7698 10852 7702 10908
rect 7702 10852 7758 10908
rect 7758 10852 7762 10908
rect 7698 10848 7762 10852
rect 7778 10908 7842 10912
rect 7778 10852 7782 10908
rect 7782 10852 7838 10908
rect 7838 10852 7842 10908
rect 7778 10848 7842 10852
rect 7858 10908 7922 10912
rect 7858 10852 7862 10908
rect 7862 10852 7918 10908
rect 7918 10852 7922 10908
rect 7858 10848 7922 10852
rect 20952 10908 21016 10912
rect 20952 10852 20956 10908
rect 20956 10852 21012 10908
rect 21012 10852 21016 10908
rect 20952 10848 21016 10852
rect 21032 10908 21096 10912
rect 21032 10852 21036 10908
rect 21036 10852 21092 10908
rect 21092 10852 21096 10908
rect 21032 10848 21096 10852
rect 21112 10908 21176 10912
rect 21112 10852 21116 10908
rect 21116 10852 21172 10908
rect 21172 10852 21176 10908
rect 21112 10848 21176 10852
rect 21192 10908 21256 10912
rect 21192 10852 21196 10908
rect 21196 10852 21252 10908
rect 21252 10852 21256 10908
rect 21192 10848 21256 10852
rect 34285 10908 34349 10912
rect 34285 10852 34289 10908
rect 34289 10852 34345 10908
rect 34345 10852 34349 10908
rect 34285 10848 34349 10852
rect 34365 10908 34429 10912
rect 34365 10852 34369 10908
rect 34369 10852 34425 10908
rect 34425 10852 34429 10908
rect 34365 10848 34429 10852
rect 34445 10908 34509 10912
rect 34445 10852 34449 10908
rect 34449 10852 34505 10908
rect 34505 10852 34509 10908
rect 34445 10848 34509 10852
rect 34525 10908 34589 10912
rect 34525 10852 34529 10908
rect 34529 10852 34585 10908
rect 34585 10852 34589 10908
rect 34525 10848 34589 10852
rect 14285 10364 14349 10368
rect 14285 10308 14289 10364
rect 14289 10308 14345 10364
rect 14345 10308 14349 10364
rect 14285 10304 14349 10308
rect 14365 10364 14429 10368
rect 14365 10308 14369 10364
rect 14369 10308 14425 10364
rect 14425 10308 14429 10364
rect 14365 10304 14429 10308
rect 14445 10364 14509 10368
rect 14445 10308 14449 10364
rect 14449 10308 14505 10364
rect 14505 10308 14509 10364
rect 14445 10304 14509 10308
rect 14525 10364 14589 10368
rect 14525 10308 14529 10364
rect 14529 10308 14585 10364
rect 14585 10308 14589 10364
rect 14525 10304 14589 10308
rect 27618 10364 27682 10368
rect 27618 10308 27622 10364
rect 27622 10308 27678 10364
rect 27678 10308 27682 10364
rect 27618 10304 27682 10308
rect 27698 10364 27762 10368
rect 27698 10308 27702 10364
rect 27702 10308 27758 10364
rect 27758 10308 27762 10364
rect 27698 10304 27762 10308
rect 27778 10364 27842 10368
rect 27778 10308 27782 10364
rect 27782 10308 27838 10364
rect 27838 10308 27842 10364
rect 27778 10304 27842 10308
rect 27858 10364 27922 10368
rect 27858 10308 27862 10364
rect 27862 10308 27918 10364
rect 27918 10308 27922 10364
rect 27858 10304 27922 10308
rect 7618 9820 7682 9824
rect 7618 9764 7622 9820
rect 7622 9764 7678 9820
rect 7678 9764 7682 9820
rect 7618 9760 7682 9764
rect 7698 9820 7762 9824
rect 7698 9764 7702 9820
rect 7702 9764 7758 9820
rect 7758 9764 7762 9820
rect 7698 9760 7762 9764
rect 7778 9820 7842 9824
rect 7778 9764 7782 9820
rect 7782 9764 7838 9820
rect 7838 9764 7842 9820
rect 7778 9760 7842 9764
rect 7858 9820 7922 9824
rect 7858 9764 7862 9820
rect 7862 9764 7918 9820
rect 7918 9764 7922 9820
rect 7858 9760 7922 9764
rect 20952 9820 21016 9824
rect 20952 9764 20956 9820
rect 20956 9764 21012 9820
rect 21012 9764 21016 9820
rect 20952 9760 21016 9764
rect 21032 9820 21096 9824
rect 21032 9764 21036 9820
rect 21036 9764 21092 9820
rect 21092 9764 21096 9820
rect 21032 9760 21096 9764
rect 21112 9820 21176 9824
rect 21112 9764 21116 9820
rect 21116 9764 21172 9820
rect 21172 9764 21176 9820
rect 21112 9760 21176 9764
rect 21192 9820 21256 9824
rect 21192 9764 21196 9820
rect 21196 9764 21252 9820
rect 21252 9764 21256 9820
rect 21192 9760 21256 9764
rect 34285 9820 34349 9824
rect 34285 9764 34289 9820
rect 34289 9764 34345 9820
rect 34345 9764 34349 9820
rect 34285 9760 34349 9764
rect 34365 9820 34429 9824
rect 34365 9764 34369 9820
rect 34369 9764 34425 9820
rect 34425 9764 34429 9820
rect 34365 9760 34429 9764
rect 34445 9820 34509 9824
rect 34445 9764 34449 9820
rect 34449 9764 34505 9820
rect 34505 9764 34509 9820
rect 34445 9760 34509 9764
rect 34525 9820 34589 9824
rect 34525 9764 34529 9820
rect 34529 9764 34585 9820
rect 34585 9764 34589 9820
rect 34525 9760 34589 9764
rect 14285 9276 14349 9280
rect 14285 9220 14289 9276
rect 14289 9220 14345 9276
rect 14345 9220 14349 9276
rect 14285 9216 14349 9220
rect 14365 9276 14429 9280
rect 14365 9220 14369 9276
rect 14369 9220 14425 9276
rect 14425 9220 14429 9276
rect 14365 9216 14429 9220
rect 14445 9276 14509 9280
rect 14445 9220 14449 9276
rect 14449 9220 14505 9276
rect 14505 9220 14509 9276
rect 14445 9216 14509 9220
rect 14525 9276 14589 9280
rect 14525 9220 14529 9276
rect 14529 9220 14585 9276
rect 14585 9220 14589 9276
rect 14525 9216 14589 9220
rect 27618 9276 27682 9280
rect 27618 9220 27622 9276
rect 27622 9220 27678 9276
rect 27678 9220 27682 9276
rect 27618 9216 27682 9220
rect 27698 9276 27762 9280
rect 27698 9220 27702 9276
rect 27702 9220 27758 9276
rect 27758 9220 27762 9276
rect 27698 9216 27762 9220
rect 27778 9276 27842 9280
rect 27778 9220 27782 9276
rect 27782 9220 27838 9276
rect 27838 9220 27842 9276
rect 27778 9216 27842 9220
rect 27858 9276 27922 9280
rect 27858 9220 27862 9276
rect 27862 9220 27918 9276
rect 27918 9220 27922 9276
rect 27858 9216 27922 9220
rect 7618 8732 7682 8736
rect 7618 8676 7622 8732
rect 7622 8676 7678 8732
rect 7678 8676 7682 8732
rect 7618 8672 7682 8676
rect 7698 8732 7762 8736
rect 7698 8676 7702 8732
rect 7702 8676 7758 8732
rect 7758 8676 7762 8732
rect 7698 8672 7762 8676
rect 7778 8732 7842 8736
rect 7778 8676 7782 8732
rect 7782 8676 7838 8732
rect 7838 8676 7842 8732
rect 7778 8672 7842 8676
rect 7858 8732 7922 8736
rect 7858 8676 7862 8732
rect 7862 8676 7918 8732
rect 7918 8676 7922 8732
rect 7858 8672 7922 8676
rect 20952 8732 21016 8736
rect 20952 8676 20956 8732
rect 20956 8676 21012 8732
rect 21012 8676 21016 8732
rect 20952 8672 21016 8676
rect 21032 8732 21096 8736
rect 21032 8676 21036 8732
rect 21036 8676 21092 8732
rect 21092 8676 21096 8732
rect 21032 8672 21096 8676
rect 21112 8732 21176 8736
rect 21112 8676 21116 8732
rect 21116 8676 21172 8732
rect 21172 8676 21176 8732
rect 21112 8672 21176 8676
rect 21192 8732 21256 8736
rect 21192 8676 21196 8732
rect 21196 8676 21252 8732
rect 21252 8676 21256 8732
rect 21192 8672 21256 8676
rect 34285 8732 34349 8736
rect 34285 8676 34289 8732
rect 34289 8676 34345 8732
rect 34345 8676 34349 8732
rect 34285 8672 34349 8676
rect 34365 8732 34429 8736
rect 34365 8676 34369 8732
rect 34369 8676 34425 8732
rect 34425 8676 34429 8732
rect 34365 8672 34429 8676
rect 34445 8732 34509 8736
rect 34445 8676 34449 8732
rect 34449 8676 34505 8732
rect 34505 8676 34509 8732
rect 34445 8672 34509 8676
rect 34525 8732 34589 8736
rect 34525 8676 34529 8732
rect 34529 8676 34585 8732
rect 34585 8676 34589 8732
rect 34525 8672 34589 8676
rect 14285 8188 14349 8192
rect 14285 8132 14289 8188
rect 14289 8132 14345 8188
rect 14345 8132 14349 8188
rect 14285 8128 14349 8132
rect 14365 8188 14429 8192
rect 14365 8132 14369 8188
rect 14369 8132 14425 8188
rect 14425 8132 14429 8188
rect 14365 8128 14429 8132
rect 14445 8188 14509 8192
rect 14445 8132 14449 8188
rect 14449 8132 14505 8188
rect 14505 8132 14509 8188
rect 14445 8128 14509 8132
rect 14525 8188 14589 8192
rect 14525 8132 14529 8188
rect 14529 8132 14585 8188
rect 14585 8132 14589 8188
rect 14525 8128 14589 8132
rect 27618 8188 27682 8192
rect 27618 8132 27622 8188
rect 27622 8132 27678 8188
rect 27678 8132 27682 8188
rect 27618 8128 27682 8132
rect 27698 8188 27762 8192
rect 27698 8132 27702 8188
rect 27702 8132 27758 8188
rect 27758 8132 27762 8188
rect 27698 8128 27762 8132
rect 27778 8188 27842 8192
rect 27778 8132 27782 8188
rect 27782 8132 27838 8188
rect 27838 8132 27842 8188
rect 27778 8128 27842 8132
rect 27858 8188 27922 8192
rect 27858 8132 27862 8188
rect 27862 8132 27918 8188
rect 27918 8132 27922 8188
rect 27858 8128 27922 8132
rect 7618 7644 7682 7648
rect 7618 7588 7622 7644
rect 7622 7588 7678 7644
rect 7678 7588 7682 7644
rect 7618 7584 7682 7588
rect 7698 7644 7762 7648
rect 7698 7588 7702 7644
rect 7702 7588 7758 7644
rect 7758 7588 7762 7644
rect 7698 7584 7762 7588
rect 7778 7644 7842 7648
rect 7778 7588 7782 7644
rect 7782 7588 7838 7644
rect 7838 7588 7842 7644
rect 7778 7584 7842 7588
rect 7858 7644 7922 7648
rect 7858 7588 7862 7644
rect 7862 7588 7918 7644
rect 7918 7588 7922 7644
rect 7858 7584 7922 7588
rect 20952 7644 21016 7648
rect 20952 7588 20956 7644
rect 20956 7588 21012 7644
rect 21012 7588 21016 7644
rect 20952 7584 21016 7588
rect 21032 7644 21096 7648
rect 21032 7588 21036 7644
rect 21036 7588 21092 7644
rect 21092 7588 21096 7644
rect 21032 7584 21096 7588
rect 21112 7644 21176 7648
rect 21112 7588 21116 7644
rect 21116 7588 21172 7644
rect 21172 7588 21176 7644
rect 21112 7584 21176 7588
rect 21192 7644 21256 7648
rect 21192 7588 21196 7644
rect 21196 7588 21252 7644
rect 21252 7588 21256 7644
rect 21192 7584 21256 7588
rect 34285 7644 34349 7648
rect 34285 7588 34289 7644
rect 34289 7588 34345 7644
rect 34345 7588 34349 7644
rect 34285 7584 34349 7588
rect 34365 7644 34429 7648
rect 34365 7588 34369 7644
rect 34369 7588 34425 7644
rect 34425 7588 34429 7644
rect 34365 7584 34429 7588
rect 34445 7644 34509 7648
rect 34445 7588 34449 7644
rect 34449 7588 34505 7644
rect 34505 7588 34509 7644
rect 34445 7584 34509 7588
rect 34525 7644 34589 7648
rect 34525 7588 34529 7644
rect 34529 7588 34585 7644
rect 34585 7588 34589 7644
rect 34525 7584 34589 7588
rect 14285 7100 14349 7104
rect 14285 7044 14289 7100
rect 14289 7044 14345 7100
rect 14345 7044 14349 7100
rect 14285 7040 14349 7044
rect 14365 7100 14429 7104
rect 14365 7044 14369 7100
rect 14369 7044 14425 7100
rect 14425 7044 14429 7100
rect 14365 7040 14429 7044
rect 14445 7100 14509 7104
rect 14445 7044 14449 7100
rect 14449 7044 14505 7100
rect 14505 7044 14509 7100
rect 14445 7040 14509 7044
rect 14525 7100 14589 7104
rect 14525 7044 14529 7100
rect 14529 7044 14585 7100
rect 14585 7044 14589 7100
rect 14525 7040 14589 7044
rect 27618 7100 27682 7104
rect 27618 7044 27622 7100
rect 27622 7044 27678 7100
rect 27678 7044 27682 7100
rect 27618 7040 27682 7044
rect 27698 7100 27762 7104
rect 27698 7044 27702 7100
rect 27702 7044 27758 7100
rect 27758 7044 27762 7100
rect 27698 7040 27762 7044
rect 27778 7100 27842 7104
rect 27778 7044 27782 7100
rect 27782 7044 27838 7100
rect 27838 7044 27842 7100
rect 27778 7040 27842 7044
rect 27858 7100 27922 7104
rect 27858 7044 27862 7100
rect 27862 7044 27918 7100
rect 27918 7044 27922 7100
rect 27858 7040 27922 7044
rect 7618 6556 7682 6560
rect 7618 6500 7622 6556
rect 7622 6500 7678 6556
rect 7678 6500 7682 6556
rect 7618 6496 7682 6500
rect 7698 6556 7762 6560
rect 7698 6500 7702 6556
rect 7702 6500 7758 6556
rect 7758 6500 7762 6556
rect 7698 6496 7762 6500
rect 7778 6556 7842 6560
rect 7778 6500 7782 6556
rect 7782 6500 7838 6556
rect 7838 6500 7842 6556
rect 7778 6496 7842 6500
rect 7858 6556 7922 6560
rect 7858 6500 7862 6556
rect 7862 6500 7918 6556
rect 7918 6500 7922 6556
rect 7858 6496 7922 6500
rect 20952 6556 21016 6560
rect 20952 6500 20956 6556
rect 20956 6500 21012 6556
rect 21012 6500 21016 6556
rect 20952 6496 21016 6500
rect 21032 6556 21096 6560
rect 21032 6500 21036 6556
rect 21036 6500 21092 6556
rect 21092 6500 21096 6556
rect 21032 6496 21096 6500
rect 21112 6556 21176 6560
rect 21112 6500 21116 6556
rect 21116 6500 21172 6556
rect 21172 6500 21176 6556
rect 21112 6496 21176 6500
rect 21192 6556 21256 6560
rect 21192 6500 21196 6556
rect 21196 6500 21252 6556
rect 21252 6500 21256 6556
rect 21192 6496 21256 6500
rect 34285 6556 34349 6560
rect 34285 6500 34289 6556
rect 34289 6500 34345 6556
rect 34345 6500 34349 6556
rect 34285 6496 34349 6500
rect 34365 6556 34429 6560
rect 34365 6500 34369 6556
rect 34369 6500 34425 6556
rect 34425 6500 34429 6556
rect 34365 6496 34429 6500
rect 34445 6556 34509 6560
rect 34445 6500 34449 6556
rect 34449 6500 34505 6556
rect 34505 6500 34509 6556
rect 34445 6496 34509 6500
rect 34525 6556 34589 6560
rect 34525 6500 34529 6556
rect 34529 6500 34585 6556
rect 34585 6500 34589 6556
rect 34525 6496 34589 6500
rect 14285 6012 14349 6016
rect 14285 5956 14289 6012
rect 14289 5956 14345 6012
rect 14345 5956 14349 6012
rect 14285 5952 14349 5956
rect 14365 6012 14429 6016
rect 14365 5956 14369 6012
rect 14369 5956 14425 6012
rect 14425 5956 14429 6012
rect 14365 5952 14429 5956
rect 14445 6012 14509 6016
rect 14445 5956 14449 6012
rect 14449 5956 14505 6012
rect 14505 5956 14509 6012
rect 14445 5952 14509 5956
rect 14525 6012 14589 6016
rect 14525 5956 14529 6012
rect 14529 5956 14585 6012
rect 14585 5956 14589 6012
rect 14525 5952 14589 5956
rect 27618 6012 27682 6016
rect 27618 5956 27622 6012
rect 27622 5956 27678 6012
rect 27678 5956 27682 6012
rect 27618 5952 27682 5956
rect 27698 6012 27762 6016
rect 27698 5956 27702 6012
rect 27702 5956 27758 6012
rect 27758 5956 27762 6012
rect 27698 5952 27762 5956
rect 27778 6012 27842 6016
rect 27778 5956 27782 6012
rect 27782 5956 27838 6012
rect 27838 5956 27842 6012
rect 27778 5952 27842 5956
rect 27858 6012 27922 6016
rect 27858 5956 27862 6012
rect 27862 5956 27918 6012
rect 27918 5956 27922 6012
rect 27858 5952 27922 5956
rect 7618 5468 7682 5472
rect 7618 5412 7622 5468
rect 7622 5412 7678 5468
rect 7678 5412 7682 5468
rect 7618 5408 7682 5412
rect 7698 5468 7762 5472
rect 7698 5412 7702 5468
rect 7702 5412 7758 5468
rect 7758 5412 7762 5468
rect 7698 5408 7762 5412
rect 7778 5468 7842 5472
rect 7778 5412 7782 5468
rect 7782 5412 7838 5468
rect 7838 5412 7842 5468
rect 7778 5408 7842 5412
rect 7858 5468 7922 5472
rect 7858 5412 7862 5468
rect 7862 5412 7918 5468
rect 7918 5412 7922 5468
rect 7858 5408 7922 5412
rect 20952 5468 21016 5472
rect 20952 5412 20956 5468
rect 20956 5412 21012 5468
rect 21012 5412 21016 5468
rect 20952 5408 21016 5412
rect 21032 5468 21096 5472
rect 21032 5412 21036 5468
rect 21036 5412 21092 5468
rect 21092 5412 21096 5468
rect 21032 5408 21096 5412
rect 21112 5468 21176 5472
rect 21112 5412 21116 5468
rect 21116 5412 21172 5468
rect 21172 5412 21176 5468
rect 21112 5408 21176 5412
rect 21192 5468 21256 5472
rect 21192 5412 21196 5468
rect 21196 5412 21252 5468
rect 21252 5412 21256 5468
rect 21192 5408 21256 5412
rect 34285 5468 34349 5472
rect 34285 5412 34289 5468
rect 34289 5412 34345 5468
rect 34345 5412 34349 5468
rect 34285 5408 34349 5412
rect 34365 5468 34429 5472
rect 34365 5412 34369 5468
rect 34369 5412 34425 5468
rect 34425 5412 34429 5468
rect 34365 5408 34429 5412
rect 34445 5468 34509 5472
rect 34445 5412 34449 5468
rect 34449 5412 34505 5468
rect 34505 5412 34509 5468
rect 34445 5408 34509 5412
rect 34525 5468 34589 5472
rect 34525 5412 34529 5468
rect 34529 5412 34585 5468
rect 34585 5412 34589 5468
rect 34525 5408 34589 5412
rect 14285 4924 14349 4928
rect 14285 4868 14289 4924
rect 14289 4868 14345 4924
rect 14345 4868 14349 4924
rect 14285 4864 14349 4868
rect 14365 4924 14429 4928
rect 14365 4868 14369 4924
rect 14369 4868 14425 4924
rect 14425 4868 14429 4924
rect 14365 4864 14429 4868
rect 14445 4924 14509 4928
rect 14445 4868 14449 4924
rect 14449 4868 14505 4924
rect 14505 4868 14509 4924
rect 14445 4864 14509 4868
rect 14525 4924 14589 4928
rect 14525 4868 14529 4924
rect 14529 4868 14585 4924
rect 14585 4868 14589 4924
rect 14525 4864 14589 4868
rect 27618 4924 27682 4928
rect 27618 4868 27622 4924
rect 27622 4868 27678 4924
rect 27678 4868 27682 4924
rect 27618 4864 27682 4868
rect 27698 4924 27762 4928
rect 27698 4868 27702 4924
rect 27702 4868 27758 4924
rect 27758 4868 27762 4924
rect 27698 4864 27762 4868
rect 27778 4924 27842 4928
rect 27778 4868 27782 4924
rect 27782 4868 27838 4924
rect 27838 4868 27842 4924
rect 27778 4864 27842 4868
rect 27858 4924 27922 4928
rect 27858 4868 27862 4924
rect 27862 4868 27918 4924
rect 27918 4868 27922 4924
rect 27858 4864 27922 4868
rect 7618 4380 7682 4384
rect 7618 4324 7622 4380
rect 7622 4324 7678 4380
rect 7678 4324 7682 4380
rect 7618 4320 7682 4324
rect 7698 4380 7762 4384
rect 7698 4324 7702 4380
rect 7702 4324 7758 4380
rect 7758 4324 7762 4380
rect 7698 4320 7762 4324
rect 7778 4380 7842 4384
rect 7778 4324 7782 4380
rect 7782 4324 7838 4380
rect 7838 4324 7842 4380
rect 7778 4320 7842 4324
rect 7858 4380 7922 4384
rect 7858 4324 7862 4380
rect 7862 4324 7918 4380
rect 7918 4324 7922 4380
rect 7858 4320 7922 4324
rect 20952 4380 21016 4384
rect 20952 4324 20956 4380
rect 20956 4324 21012 4380
rect 21012 4324 21016 4380
rect 20952 4320 21016 4324
rect 21032 4380 21096 4384
rect 21032 4324 21036 4380
rect 21036 4324 21092 4380
rect 21092 4324 21096 4380
rect 21032 4320 21096 4324
rect 21112 4380 21176 4384
rect 21112 4324 21116 4380
rect 21116 4324 21172 4380
rect 21172 4324 21176 4380
rect 21112 4320 21176 4324
rect 21192 4380 21256 4384
rect 21192 4324 21196 4380
rect 21196 4324 21252 4380
rect 21252 4324 21256 4380
rect 21192 4320 21256 4324
rect 34285 4380 34349 4384
rect 34285 4324 34289 4380
rect 34289 4324 34345 4380
rect 34345 4324 34349 4380
rect 34285 4320 34349 4324
rect 34365 4380 34429 4384
rect 34365 4324 34369 4380
rect 34369 4324 34425 4380
rect 34425 4324 34429 4380
rect 34365 4320 34429 4324
rect 34445 4380 34509 4384
rect 34445 4324 34449 4380
rect 34449 4324 34505 4380
rect 34505 4324 34509 4380
rect 34445 4320 34509 4324
rect 34525 4380 34589 4384
rect 34525 4324 34529 4380
rect 34529 4324 34585 4380
rect 34585 4324 34589 4380
rect 34525 4320 34589 4324
rect 14285 3836 14349 3840
rect 14285 3780 14289 3836
rect 14289 3780 14345 3836
rect 14345 3780 14349 3836
rect 14285 3776 14349 3780
rect 14365 3836 14429 3840
rect 14365 3780 14369 3836
rect 14369 3780 14425 3836
rect 14425 3780 14429 3836
rect 14365 3776 14429 3780
rect 14445 3836 14509 3840
rect 14445 3780 14449 3836
rect 14449 3780 14505 3836
rect 14505 3780 14509 3836
rect 14445 3776 14509 3780
rect 14525 3836 14589 3840
rect 14525 3780 14529 3836
rect 14529 3780 14585 3836
rect 14585 3780 14589 3836
rect 14525 3776 14589 3780
rect 27618 3836 27682 3840
rect 27618 3780 27622 3836
rect 27622 3780 27678 3836
rect 27678 3780 27682 3836
rect 27618 3776 27682 3780
rect 27698 3836 27762 3840
rect 27698 3780 27702 3836
rect 27702 3780 27758 3836
rect 27758 3780 27762 3836
rect 27698 3776 27762 3780
rect 27778 3836 27842 3840
rect 27778 3780 27782 3836
rect 27782 3780 27838 3836
rect 27838 3780 27842 3836
rect 27778 3776 27842 3780
rect 27858 3836 27922 3840
rect 27858 3780 27862 3836
rect 27862 3780 27918 3836
rect 27918 3780 27922 3836
rect 27858 3776 27922 3780
rect 7618 3292 7682 3296
rect 7618 3236 7622 3292
rect 7622 3236 7678 3292
rect 7678 3236 7682 3292
rect 7618 3232 7682 3236
rect 7698 3292 7762 3296
rect 7698 3236 7702 3292
rect 7702 3236 7758 3292
rect 7758 3236 7762 3292
rect 7698 3232 7762 3236
rect 7778 3292 7842 3296
rect 7778 3236 7782 3292
rect 7782 3236 7838 3292
rect 7838 3236 7842 3292
rect 7778 3232 7842 3236
rect 7858 3292 7922 3296
rect 7858 3236 7862 3292
rect 7862 3236 7918 3292
rect 7918 3236 7922 3292
rect 7858 3232 7922 3236
rect 20952 3292 21016 3296
rect 20952 3236 20956 3292
rect 20956 3236 21012 3292
rect 21012 3236 21016 3292
rect 20952 3232 21016 3236
rect 21032 3292 21096 3296
rect 21032 3236 21036 3292
rect 21036 3236 21092 3292
rect 21092 3236 21096 3292
rect 21032 3232 21096 3236
rect 21112 3292 21176 3296
rect 21112 3236 21116 3292
rect 21116 3236 21172 3292
rect 21172 3236 21176 3292
rect 21112 3232 21176 3236
rect 21192 3292 21256 3296
rect 21192 3236 21196 3292
rect 21196 3236 21252 3292
rect 21252 3236 21256 3292
rect 21192 3232 21256 3236
rect 34285 3292 34349 3296
rect 34285 3236 34289 3292
rect 34289 3236 34345 3292
rect 34345 3236 34349 3292
rect 34285 3232 34349 3236
rect 34365 3292 34429 3296
rect 34365 3236 34369 3292
rect 34369 3236 34425 3292
rect 34425 3236 34429 3292
rect 34365 3232 34429 3236
rect 34445 3292 34509 3296
rect 34445 3236 34449 3292
rect 34449 3236 34505 3292
rect 34505 3236 34509 3292
rect 34445 3232 34509 3236
rect 34525 3292 34589 3296
rect 34525 3236 34529 3292
rect 34529 3236 34585 3292
rect 34585 3236 34589 3292
rect 34525 3232 34589 3236
rect 35940 3088 36004 3092
rect 35940 3032 35954 3088
rect 35954 3032 36004 3088
rect 35940 3028 36004 3032
rect 14780 2816 14844 2820
rect 14780 2760 14794 2816
rect 14794 2760 14844 2816
rect 14780 2756 14844 2760
rect 14285 2748 14349 2752
rect 14285 2692 14289 2748
rect 14289 2692 14345 2748
rect 14345 2692 14349 2748
rect 14285 2688 14349 2692
rect 14365 2748 14429 2752
rect 14365 2692 14369 2748
rect 14369 2692 14425 2748
rect 14425 2692 14429 2748
rect 14365 2688 14429 2692
rect 14445 2748 14509 2752
rect 14445 2692 14449 2748
rect 14449 2692 14505 2748
rect 14505 2692 14509 2748
rect 14445 2688 14509 2692
rect 14525 2748 14589 2752
rect 14525 2692 14529 2748
rect 14529 2692 14585 2748
rect 14585 2692 14589 2748
rect 14525 2688 14589 2692
rect 27618 2748 27682 2752
rect 27618 2692 27622 2748
rect 27622 2692 27678 2748
rect 27678 2692 27682 2748
rect 27618 2688 27682 2692
rect 27698 2748 27762 2752
rect 27698 2692 27702 2748
rect 27702 2692 27758 2748
rect 27758 2692 27762 2748
rect 27698 2688 27762 2692
rect 27778 2748 27842 2752
rect 27778 2692 27782 2748
rect 27782 2692 27838 2748
rect 27838 2692 27842 2748
rect 27778 2688 27842 2692
rect 27858 2748 27922 2752
rect 27858 2692 27862 2748
rect 27862 2692 27918 2748
rect 27918 2692 27922 2748
rect 27858 2688 27922 2692
rect 7618 2204 7682 2208
rect 7618 2148 7622 2204
rect 7622 2148 7678 2204
rect 7678 2148 7682 2204
rect 7618 2144 7682 2148
rect 7698 2204 7762 2208
rect 7698 2148 7702 2204
rect 7702 2148 7758 2204
rect 7758 2148 7762 2204
rect 7698 2144 7762 2148
rect 7778 2204 7842 2208
rect 7778 2148 7782 2204
rect 7782 2148 7838 2204
rect 7838 2148 7842 2204
rect 7778 2144 7842 2148
rect 7858 2204 7922 2208
rect 7858 2148 7862 2204
rect 7862 2148 7918 2204
rect 7918 2148 7922 2204
rect 7858 2144 7922 2148
rect 20952 2204 21016 2208
rect 20952 2148 20956 2204
rect 20956 2148 21012 2204
rect 21012 2148 21016 2204
rect 20952 2144 21016 2148
rect 21032 2204 21096 2208
rect 21032 2148 21036 2204
rect 21036 2148 21092 2204
rect 21092 2148 21096 2204
rect 21032 2144 21096 2148
rect 21112 2204 21176 2208
rect 21112 2148 21116 2204
rect 21116 2148 21172 2204
rect 21172 2148 21176 2204
rect 21112 2144 21176 2148
rect 21192 2204 21256 2208
rect 21192 2148 21196 2204
rect 21196 2148 21252 2204
rect 21252 2148 21256 2204
rect 21192 2144 21256 2148
rect 34285 2204 34349 2208
rect 34285 2148 34289 2204
rect 34289 2148 34345 2204
rect 34345 2148 34349 2204
rect 34285 2144 34349 2148
rect 34365 2204 34429 2208
rect 34365 2148 34369 2204
rect 34369 2148 34425 2204
rect 34425 2148 34429 2204
rect 34365 2144 34429 2148
rect 34445 2204 34509 2208
rect 34445 2148 34449 2204
rect 34449 2148 34505 2204
rect 34505 2148 34509 2204
rect 34445 2144 34509 2148
rect 34525 2204 34589 2208
rect 34525 2148 34529 2204
rect 34529 2148 34585 2204
rect 34585 2148 34589 2204
rect 34525 2144 34589 2148
rect 28948 1396 29012 1460
rect 28948 1124 29012 1188
rect 28948 716 29012 780
rect 28948 172 29012 236
<< metal4 >>
rect 7610 13088 7931 13648
rect 7610 13024 7618 13088
rect 7682 13024 7698 13088
rect 7762 13024 7778 13088
rect 7842 13024 7858 13088
rect 7922 13024 7931 13088
rect 7610 12000 7931 13024
rect 7610 11936 7618 12000
rect 7682 11936 7698 12000
rect 7762 11936 7778 12000
rect 7842 11936 7858 12000
rect 7922 11936 7931 12000
rect 7610 10912 7931 11936
rect 7610 10848 7618 10912
rect 7682 10848 7698 10912
rect 7762 10848 7778 10912
rect 7842 10848 7858 10912
rect 7922 10848 7931 10912
rect 7610 9824 7931 10848
rect 7610 9760 7618 9824
rect 7682 9760 7698 9824
rect 7762 9760 7778 9824
rect 7842 9760 7858 9824
rect 7922 9760 7931 9824
rect 7610 8736 7931 9760
rect 7610 8672 7618 8736
rect 7682 8672 7698 8736
rect 7762 8672 7778 8736
rect 7842 8672 7858 8736
rect 7922 8672 7931 8736
rect 7610 7648 7931 8672
rect 7610 7584 7618 7648
rect 7682 7584 7698 7648
rect 7762 7584 7778 7648
rect 7842 7584 7858 7648
rect 7922 7584 7931 7648
rect 7610 6560 7931 7584
rect 7610 6496 7618 6560
rect 7682 6496 7698 6560
rect 7762 6496 7778 6560
rect 7842 6496 7858 6560
rect 7922 6496 7931 6560
rect 7610 5472 7931 6496
rect 7610 5408 7618 5472
rect 7682 5408 7698 5472
rect 7762 5408 7778 5472
rect 7842 5408 7858 5472
rect 7922 5408 7931 5472
rect 7610 4384 7931 5408
rect 7610 4320 7618 4384
rect 7682 4320 7698 4384
rect 7762 4320 7778 4384
rect 7842 4320 7858 4384
rect 7922 4320 7931 4384
rect 7610 3296 7931 4320
rect 7610 3232 7618 3296
rect 7682 3232 7698 3296
rect 7762 3232 7778 3296
rect 7842 3232 7858 3296
rect 7922 3232 7931 3296
rect 7610 2208 7931 3232
rect 7610 2144 7618 2208
rect 7682 2144 7698 2208
rect 7762 2144 7778 2208
rect 7842 2144 7858 2208
rect 7922 2144 7931 2208
rect 7610 2128 7931 2144
rect 14277 13632 14597 13648
rect 14277 13568 14285 13632
rect 14349 13568 14365 13632
rect 14429 13568 14445 13632
rect 14509 13568 14525 13632
rect 14589 13568 14597 13632
rect 14277 12544 14597 13568
rect 14277 12480 14285 12544
rect 14349 12480 14365 12544
rect 14429 12480 14445 12544
rect 14509 12480 14525 12544
rect 14589 12480 14597 12544
rect 14277 11456 14597 12480
rect 14277 11392 14285 11456
rect 14349 11392 14365 11456
rect 14429 11392 14445 11456
rect 14509 11392 14525 11456
rect 14589 11392 14597 11456
rect 14277 10368 14597 11392
rect 14277 10304 14285 10368
rect 14349 10304 14365 10368
rect 14429 10304 14445 10368
rect 14509 10304 14525 10368
rect 14589 10304 14597 10368
rect 14277 9280 14597 10304
rect 14277 9216 14285 9280
rect 14349 9216 14365 9280
rect 14429 9216 14445 9280
rect 14509 9216 14525 9280
rect 14589 9216 14597 9280
rect 14277 8192 14597 9216
rect 14277 8128 14285 8192
rect 14349 8128 14365 8192
rect 14429 8128 14445 8192
rect 14509 8128 14525 8192
rect 14589 8128 14597 8192
rect 14277 7104 14597 8128
rect 14277 7040 14285 7104
rect 14349 7040 14365 7104
rect 14429 7040 14445 7104
rect 14509 7040 14525 7104
rect 14589 7040 14597 7104
rect 14277 6016 14597 7040
rect 14277 5952 14285 6016
rect 14349 5952 14365 6016
rect 14429 5952 14445 6016
rect 14509 5952 14525 6016
rect 14589 5952 14597 6016
rect 14277 4928 14597 5952
rect 14277 4864 14285 4928
rect 14349 4864 14365 4928
rect 14429 4864 14445 4928
rect 14509 4864 14525 4928
rect 14589 4864 14597 4928
rect 14277 3840 14597 4864
rect 14277 3776 14285 3840
rect 14349 3776 14365 3840
rect 14429 3776 14445 3840
rect 14509 3776 14525 3840
rect 14589 3776 14597 3840
rect 14277 2752 14597 3776
rect 20944 13088 21264 13648
rect 20944 13024 20952 13088
rect 21016 13024 21032 13088
rect 21096 13024 21112 13088
rect 21176 13024 21192 13088
rect 21256 13024 21264 13088
rect 20944 12000 21264 13024
rect 20944 11936 20952 12000
rect 21016 11936 21032 12000
rect 21096 11936 21112 12000
rect 21176 11936 21192 12000
rect 21256 11936 21264 12000
rect 20944 10912 21264 11936
rect 20944 10848 20952 10912
rect 21016 10848 21032 10912
rect 21096 10848 21112 10912
rect 21176 10848 21192 10912
rect 21256 10848 21264 10912
rect 20944 9824 21264 10848
rect 20944 9760 20952 9824
rect 21016 9760 21032 9824
rect 21096 9760 21112 9824
rect 21176 9760 21192 9824
rect 21256 9760 21264 9824
rect 20944 8736 21264 9760
rect 20944 8672 20952 8736
rect 21016 8672 21032 8736
rect 21096 8672 21112 8736
rect 21176 8672 21192 8736
rect 21256 8672 21264 8736
rect 20944 7648 21264 8672
rect 20944 7584 20952 7648
rect 21016 7584 21032 7648
rect 21096 7584 21112 7648
rect 21176 7584 21192 7648
rect 21256 7584 21264 7648
rect 20944 6560 21264 7584
rect 20944 6496 20952 6560
rect 21016 6496 21032 6560
rect 21096 6496 21112 6560
rect 21176 6496 21192 6560
rect 21256 6496 21264 6560
rect 20944 5472 21264 6496
rect 20944 5408 20952 5472
rect 21016 5408 21032 5472
rect 21096 5408 21112 5472
rect 21176 5408 21192 5472
rect 21256 5408 21264 5472
rect 20944 4384 21264 5408
rect 20944 4320 20952 4384
rect 21016 4320 21032 4384
rect 21096 4320 21112 4384
rect 21176 4320 21192 4384
rect 21256 4320 21264 4384
rect 20944 3296 21264 4320
rect 20944 3232 20952 3296
rect 21016 3232 21032 3296
rect 21096 3232 21112 3296
rect 21176 3232 21192 3296
rect 21256 3232 21264 3296
rect 14782 2821 14842 2942
rect 14779 2820 14845 2821
rect 14779 2756 14780 2820
rect 14844 2756 14845 2820
rect 14779 2755 14845 2756
rect 14277 2688 14285 2752
rect 14349 2688 14365 2752
rect 14429 2688 14445 2752
rect 14509 2688 14525 2752
rect 14589 2688 14597 2752
rect 14277 2128 14597 2688
rect 20944 2208 21264 3232
rect 20944 2144 20952 2208
rect 21016 2144 21032 2208
rect 21096 2144 21112 2208
rect 21176 2144 21192 2208
rect 21256 2144 21264 2208
rect 20944 2128 21264 2144
rect 27610 13632 27930 13648
rect 27610 13568 27618 13632
rect 27682 13568 27698 13632
rect 27762 13568 27778 13632
rect 27842 13568 27858 13632
rect 27922 13568 27930 13632
rect 27610 12544 27930 13568
rect 27610 12480 27618 12544
rect 27682 12480 27698 12544
rect 27762 12480 27778 12544
rect 27842 12480 27858 12544
rect 27922 12480 27930 12544
rect 27610 11456 27930 12480
rect 27610 11392 27618 11456
rect 27682 11392 27698 11456
rect 27762 11392 27778 11456
rect 27842 11392 27858 11456
rect 27922 11392 27930 11456
rect 27610 10368 27930 11392
rect 27610 10304 27618 10368
rect 27682 10304 27698 10368
rect 27762 10304 27778 10368
rect 27842 10304 27858 10368
rect 27922 10304 27930 10368
rect 27610 9280 27930 10304
rect 27610 9216 27618 9280
rect 27682 9216 27698 9280
rect 27762 9216 27778 9280
rect 27842 9216 27858 9280
rect 27922 9216 27930 9280
rect 27610 8192 27930 9216
rect 27610 8128 27618 8192
rect 27682 8128 27698 8192
rect 27762 8128 27778 8192
rect 27842 8128 27858 8192
rect 27922 8128 27930 8192
rect 27610 7104 27930 8128
rect 27610 7040 27618 7104
rect 27682 7040 27698 7104
rect 27762 7040 27778 7104
rect 27842 7040 27858 7104
rect 27922 7040 27930 7104
rect 27610 6016 27930 7040
rect 27610 5952 27618 6016
rect 27682 5952 27698 6016
rect 27762 5952 27778 6016
rect 27842 5952 27858 6016
rect 27922 5952 27930 6016
rect 27610 4928 27930 5952
rect 27610 4864 27618 4928
rect 27682 4864 27698 4928
rect 27762 4864 27778 4928
rect 27842 4864 27858 4928
rect 27922 4864 27930 4928
rect 27610 3840 27930 4864
rect 27610 3776 27618 3840
rect 27682 3776 27698 3840
rect 27762 3776 27778 3840
rect 27842 3776 27858 3840
rect 27922 3776 27930 3840
rect 27610 2752 27930 3776
rect 27610 2688 27618 2752
rect 27682 2688 27698 2752
rect 27762 2688 27778 2752
rect 27842 2688 27858 2752
rect 27922 2688 27930 2752
rect 27610 2128 27930 2688
rect 34277 13088 34597 13648
rect 34277 13024 34285 13088
rect 34349 13024 34365 13088
rect 34429 13024 34445 13088
rect 34509 13024 34525 13088
rect 34589 13024 34597 13088
rect 34277 12000 34597 13024
rect 34277 11936 34285 12000
rect 34349 11936 34365 12000
rect 34429 11936 34445 12000
rect 34509 11936 34525 12000
rect 34589 11936 34597 12000
rect 34277 10912 34597 11936
rect 34277 10848 34285 10912
rect 34349 10848 34365 10912
rect 34429 10848 34445 10912
rect 34509 10848 34525 10912
rect 34589 10848 34597 10912
rect 34277 9824 34597 10848
rect 34277 9760 34285 9824
rect 34349 9760 34365 9824
rect 34429 9760 34445 9824
rect 34509 9760 34525 9824
rect 34589 9760 34597 9824
rect 34277 8736 34597 9760
rect 34277 8672 34285 8736
rect 34349 8672 34365 8736
rect 34429 8672 34445 8736
rect 34509 8672 34525 8736
rect 34589 8672 34597 8736
rect 34277 7648 34597 8672
rect 34277 7584 34285 7648
rect 34349 7584 34365 7648
rect 34429 7584 34445 7648
rect 34509 7584 34525 7648
rect 34589 7584 34597 7648
rect 34277 6560 34597 7584
rect 34277 6496 34285 6560
rect 34349 6496 34365 6560
rect 34429 6496 34445 6560
rect 34509 6496 34525 6560
rect 34589 6496 34597 6560
rect 34277 5472 34597 6496
rect 34277 5408 34285 5472
rect 34349 5408 34365 5472
rect 34429 5408 34445 5472
rect 34509 5408 34525 5472
rect 34589 5408 34597 5472
rect 34277 4384 34597 5408
rect 34277 4320 34285 4384
rect 34349 4320 34365 4384
rect 34429 4320 34445 4384
rect 34509 4320 34525 4384
rect 34589 4320 34597 4384
rect 34277 3296 34597 4320
rect 34277 3232 34285 3296
rect 34349 3232 34365 3296
rect 34429 3232 34445 3296
rect 34509 3232 34525 3296
rect 34589 3232 34597 3296
rect 34277 2208 34597 3232
rect 34277 2144 34285 2208
rect 34349 2144 34365 2208
rect 34429 2144 34445 2208
rect 34509 2144 34525 2208
rect 34589 2144 34597 2208
rect 34277 2128 34597 2144
rect 28947 1460 29013 1461
rect 28947 1396 28948 1460
rect 29012 1396 29013 1460
rect 28947 1395 29013 1396
rect 28950 1189 29010 1395
rect 28947 1188 29013 1189
rect 28947 1124 28948 1188
rect 29012 1124 29013 1188
rect 28947 1123 29013 1124
rect 28947 780 29013 781
rect 28947 716 28948 780
rect 29012 716 29013 780
rect 28947 715 29013 716
rect 28950 237 29010 715
rect 28947 236 29013 237
rect 28947 172 28948 236
rect 29012 172 29013 236
rect 28947 171 29013 172
<< via4 >>
rect 14694 2942 14930 3178
rect 35854 3092 36090 3178
rect 35854 3028 35940 3092
rect 35940 3028 36004 3092
rect 36004 3028 36090 3092
rect 35854 2942 36090 3028
<< metal5 >>
rect 14652 3178 36132 3220
rect 14652 2942 14694 3178
rect 14930 2942 35854 3178
rect 36090 2942 36132 3178
rect 14652 2900 36132 2942
use scs8hd_fill_1  FILLER_1_3 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1380 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_7 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1748 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_3
timestamp 1586364061
transform 1 0 1380 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_3  PHY_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_0
timestamp 1586364061
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_17
timestamp 1586364061
transform 1 0 2668 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_13
timestamp 1586364061
transform 1 0 2300 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_15 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2484 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_11
timestamp 1586364061
transform 1 0 2116 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 1932 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_8  _088_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 1472 0 1 2720
box -38 -48 866 592
use scs8hd_decap_4  FILLER_1_21
timestamp 1586364061
transform 1 0 3036 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_23
timestamp 1586364061
transform 1 0 3220 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__090__A
timestamp 1586364061
transform 1 0 3404 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__088__A
timestamp 1586364061
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__106__A
timestamp 1586364061
transform 1 0 3404 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _106_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 2852 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_0_32
timestamp 1586364061
transform 1 0 4048 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_0_27
timestamp 1586364061
transform 1 0 3588 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_42 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _105_
timestamp 1586364061
transform 1 0 4140 0 -1 2720
box -38 -48 406 592
use scs8hd_inv_8  _090_
timestamp 1586364061
transform 1 0 3588 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_40
timestamp 1586364061
transform 1 0 4784 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_36
timestamp 1586364061
transform 1 0 4416 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_41
timestamp 1586364061
transform 1 0 4876 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_37
timestamp 1586364061
transform 1 0 4508 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__091__A
timestamp 1586364061
transform 1 0 5060 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 4600 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__105__A
timestamp 1586364061
transform 1 0 4692 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_53
timestamp 1586364061
transform 1 0 5980 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5152 0 1 2720
box -38 -48 866 592
use scs8hd_inv_8  _091_
timestamp 1586364061
transform 1 0 5244 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_57
timestamp 1586364061
transform 1 0 6348 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_58
timestamp 1586364061
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_54
timestamp 1586364061
transform 1 0 6072 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_55
timestamp 1586364061
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_43
timestamp 1586364061
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_71
timestamp 1586364061
transform 1 0 7636 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_63
timestamp 1586364061
transform 1 0 6900 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7176 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_75
timestamp 1586364061
transform 1 0 8004 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_75
timestamp 1586364061
transform 1 0 8004 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7820 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _103_
timestamp 1586364061
transform 1 0 8372 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_1_87
timestamp 1586364061
transform 1 0 9108 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_83
timestamp 1586364061
transform 1 0 8740 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__103__A
timestamp 1586364061
transform 1 0 8924 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_79 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 8372 0 -1 2720
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_0_98
timestamp 1586364061
transform 1 0 10120 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 9476 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__101__A
timestamp 1586364061
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_44
timestamp 1586364061
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _100_
timestamp 1586364061
transform 1 0 9752 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_105
timestamp 1586364061
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_101
timestamp 1586364061
transform 1 0 10396 0 1 2720
box -38 -48 406 592
use scs8hd_decap_3  FILLER_0_102
timestamp 1586364061
transform 1 0 10488 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 10764 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 10856 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__100__A
timestamp 1586364061
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 9568 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 10948 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_108
timestamp 1586364061
transform 1 0 11040 0 1 2720
box -38 -48 130 592
use scs8hd_buf_2  _098_
timestamp 1586364061
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_113
timestamp 1586364061
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_116
timestamp 1586364061
transform 1 0 11776 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__098__A
timestamp 1586364061
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_121
timestamp 1586364061
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_117
timestamp 1586364061
transform 1 0 11868 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_120
timestamp 1586364061
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12052 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_56
timestamp 1586364061
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_45
timestamp 1586364061
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_130
timestamp 1586364061
transform 1 0 13064 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_126
timestamp 1586364061
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13248 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 12880 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_138
timestamp 1586364061
transform 1 0 13800 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_134
timestamp 1586364061
transform 1 0 13432 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 13432 0 1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_147
timestamp 1586364061
transform 1 0 14628 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_143
timestamp 1586364061
transform 1 0 14260 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_149
timestamp 1586364061
transform 1 0 14812 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_145
timestamp 1586364061
transform 1 0 14444 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14812 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14628 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 14444 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_160
timestamp 1586364061
transform 1 0 15824 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_159
timestamp 1586364061
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_153
timestamp 1586364061
transform 1 0 15180 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_46
timestamp 1586364061
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 15456 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 14996 0 1 2720
box -38 -48 866 592
use scs8hd_fill_2  FILLER_1_164
timestamp 1586364061
transform 1 0 16192 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 16008 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 15916 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 16560 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_175
timestamp 1586364061
transform 1 0 17204 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_171
timestamp 1586364061
transform 1 0 16836 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_175 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 17204 0 -1 2720
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 17388 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 17020 0 1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_163
timestamp 1586364061
transform 1 0 16100 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_184
timestamp 1586364061
transform 1 0 18032 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_179
timestamp 1586364061
transform 1 0 17572 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_0_183
timestamp 1586364061
transform 1 0 17940 0 -1 2720
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 17756 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_57
timestamp 1586364061
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use scs8hd_fill_1  FILLER_1_188
timestamp 1586364061
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_187 tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 18308 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18492 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_47
timestamp 1586364061
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 18676 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_194
timestamp 1586364061
transform 1 0 18952 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_196
timestamp 1586364061
transform 1 0 19136 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_193
timestamp 1586364061
transform 1 0 18860 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 18952 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19504 0 -1 2720
box -38 -48 866 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19688 0 1 2720
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19504 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 20700 0 1 2720
box -38 -48 222 592
use scs8hd_decap_8  FILLER_0_209
timestamp 1586364061
transform 1 0 20332 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_1_198
timestamp 1586364061
transform 1 0 19320 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_211
timestamp 1586364061
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_1_215
timestamp 1586364061
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_221
timestamp 1586364061
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 21068 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_48
timestamp 1586364061
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 21160 0 -1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_228
timestamp 1586364061
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_225
timestamp 1586364061
transform 1 0 21804 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21988 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22264 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 21620 0 -1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 22172 0 -1 2720
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21252 0 1 2720
box -38 -48 866 592
use scs8hd_fill_1  FILLER_1_240
timestamp 1586364061
transform 1 0 23184 0 1 2720
box -38 -48 130 592
use scs8hd_decap_4  FILLER_1_236
timestamp 1586364061
transform 1 0 22816 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_232
timestamp 1586364061
transform 1 0 22448 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_232
timestamp 1586364061
transform 1 0 22448 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22632 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 22632 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_243
timestamp 1586364061
transform 1 0 23460 0 1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 23276 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_58
timestamp 1586364061
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_49
timestamp 1586364061
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_245
timestamp 1586364061
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_249
timestamp 1586364061
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_236
timestamp 1586364061
transform 1 0 22816 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_261
timestamp 1586364061
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_257
timestamp 1586364061
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_1_269
timestamp 1586364061
transform 1 0 25852 0 1 2720
box -38 -48 590 592
use scs8hd_decap_6  FILLER_0_273
timestamp 1586364061
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_1_278
timestamp 1586364061
transform 1 0 26680 0 1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_1_275
timestamp 1586364061
transform 1 0 26404 0 1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_280
timestamp 1586364061
transform 1 0 26864 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26864 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 26496 0 1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_50
timestamp 1586364061
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use scs8hd_fill_2  FILLER_1_285
timestamp 1586364061
transform 1 0 27324 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27048 0 1 2720
box -38 -48 314 592
use scs8hd_fill_2  FILLER_1_289
timestamp 1586364061
transform 1 0 27692 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_290
timestamp 1586364061
transform 1 0 27784 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_1  FILLER_0_286
timestamp 1586364061
transform 1 0 27416 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27508 0 1 2720
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27508 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_294
timestamp 1586364061
transform 1 0 28152 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 27876 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 27968 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _107_
timestamp 1586364061
transform 1 0 28060 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_297
timestamp 1586364061
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__107__A
timestamp 1586364061
transform 1 0 28612 0 1 2720
box -38 -48 222 592
use scs8hd_buf_2  _109_
timestamp 1586364061
transform 1 0 28520 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_301
timestamp 1586364061
transform 1 0 28796 0 1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_302
timestamp 1586364061
transform 1 0 28888 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 2720
box -38 -48 222 592
use scs8hd_decap_3  FILLER_1_306
timestamp 1586364061
transform 1 0 29256 0 1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_0_306
timestamp 1586364061
transform 1 0 29256 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__109__A
timestamp 1586364061
transform 1 0 29072 0 -1 2720
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_59
timestamp 1586364061
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_51
timestamp 1586364061
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use scs8hd_buf_2  _110_
timestamp 1586364061
transform 1 0 29532 0 1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_1_313
timestamp 1586364061
transform 1 0 29900 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_0_311
timestamp 1586364061
transform 1 0 29716 0 -1 2720
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30084 0 1 2720
box -38 -48 222 592
use scs8hd_decap_6  FILLER_1_317
timestamp 1586364061
transform 1 0 30268 0 1 2720
box -38 -48 590 592
use scs8hd_fill_2  FILLER_0_321
timestamp 1586364061
transform 1 0 30636 0 -1 2720
box -38 -48 222 592
use scs8hd_buf_2  _112_
timestamp 1586364061
transform 1 0 30268 0 -1 2720
box -38 -48 406 592
use scs8hd_buf_2  _114_
timestamp 1586364061
transform 1 0 31372 0 -1 2720
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__114__A
timestamp 1586364061
transform 1 0 31924 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__112__A
timestamp 1586364061
transform 1 0 30820 0 -1 2720
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 30820 0 1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_325
timestamp 1586364061
transform 1 0 31004 0 -1 2720
box -38 -48 406 592
use scs8hd_fill_2  FILLER_0_333
timestamp 1586364061
transform 1 0 31740 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_4  FILLER_0_337
timestamp 1586364061
transform 1 0 32108 0 -1 2720
box -38 -48 406 592
use scs8hd_decap_12  FILLER_1_325
timestamp 1586364061
transform 1 0 31004 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_337
timestamp 1586364061
transform 1 0 32108 0 1 2720
box -38 -48 1142 592
use scs8hd_buf_2  _115_
timestamp 1586364061
transform 1 0 32568 0 -1 2720
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_52
timestamp 1586364061
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__115__A
timestamp 1586364061
transform 1 0 33120 0 -1 2720
box -38 -48 222 592
use scs8hd_fill_2  FILLER_0_346
timestamp 1586364061
transform 1 0 32936 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_350
timestamp 1586364061
transform 1 0 33304 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_349
timestamp 1586364061
transform 1 0 33212 0 1 2720
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_53
timestamp 1586364061
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_60
timestamp 1586364061
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use scs8hd_decap_8  FILLER_0_362
timestamp 1586364061
transform 1 0 34408 0 -1 2720
box -38 -48 774 592
use scs8hd_fill_2  FILLER_0_370
timestamp 1586364061
transform 1 0 35144 0 -1 2720
box -38 -48 222 592
use scs8hd_decap_12  FILLER_0_373
timestamp 1586364061
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_1_361
timestamp 1586364061
transform 1 0 34316 0 1 2720
box -38 -48 406 592
use scs8hd_fill_1  FILLER_1_365
timestamp 1586364061
transform 1 0 34684 0 1 2720
box -38 -48 130 592
use scs8hd_decap_12  FILLER_1_367
timestamp 1586364061
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_0_385
timestamp 1586364061
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_379
timestamp 1586364061
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_1_391
timestamp 1586364061
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use scs8hd_decap_3  PHY_1
timestamp 1586364061
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_3  PHY_3
timestamp 1586364061
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_54
timestamp 1586364061
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use scs8hd_decap_6  FILLER_0_397
timestamp 1586364061
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use scs8hd_decap_3  FILLER_0_404
timestamp 1586364061
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use scs8hd_decap_4  FILLER_1_403
timestamp 1586364061
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1472 0 -1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_4
timestamp 1586364061
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 2484 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_3
timestamp 1586364061
transform 1 0 1380 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_13
timestamp 1586364061
transform 1 0 2300 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_17
timestamp 1586364061
transform 1 0 2668 0 -1 3808
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_61
timestamp 1586364061
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__089__A
timestamp 1586364061
transform 1 0 4232 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3772 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 3312 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2852 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_21
timestamp 1586364061
transform 1 0 3036 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_26
timestamp 1586364061
transform 1 0 3496 0 -1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_2_32
timestamp 1586364061
transform 1 0 4048 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_1_.latch tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 5520 0 -1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 4508 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__085__C
timestamp 1586364061
transform 1 0 5336 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__B
timestamp 1586364061
transform 1 0 4968 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_36
timestamp 1586364061
transform 1 0 4416 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_40
timestamp 1586364061
transform 1 0 4784 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_44
timestamp 1586364061
transform 1 0 5152 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_2.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7268 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 6808 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_59
timestamp 1586364061
transform 1 0 6532 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_64
timestamp 1586364061
transform 1 0 6992 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_76
timestamp 1586364061
transform 1 0 8096 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_8  FILLER_2_80
timestamp 1586364061
transform 1 0 8464 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_88
timestamp 1586364061
transform 1 0 9200 0 -1 3808
box -38 -48 222 592
use scs8hd_buf_2  _101_
timestamp 1586364061
transform 1 0 9660 0 -1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 10856 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_62
timestamp 1586364061
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__074__D
timestamp 1586364061
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__C
timestamp 1586364061
transform 1 0 10580 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_97
timestamp 1586364061
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_101
timestamp 1586364061
transform 1 0 10396 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_2_105
timestamp 1586364061
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 12052 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_117
timestamp 1586364061
transform 1 0 11868 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_121
timestamp 1586364061
transform 1 0 12236 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 14168 0 -1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12604 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 13616 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 13984 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_134
timestamp 1586364061
transform 1 0 13432 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_138
timestamp 1586364061
transform 1 0 13800 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 15272 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_63
timestamp 1586364061
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 14628 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 14996 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_145
timestamp 1586364061
transform 1 0 14444 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_149
timestamp 1586364061
transform 1 0 14812 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 17020 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__A
timestamp 1586364061
transform 1 0 16744 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_165
timestamp 1586364061
transform 1 0 16284 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_169
timestamp 1586364061
transform 1 0 16652 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_172
timestamp 1586364061
transform 1 0 16928 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18124 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_2_182
timestamp 1586364061
transform 1 0 17848 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_8  FILLER_2_187
timestamp 1586364061
transform 1 0 18308 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_195
timestamp 1586364061
transform 1 0 19044 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_64
timestamp 1586364061
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 20240 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_206
timestamp 1586364061
transform 1 0 20056 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_210
timestamp 1586364061
transform 1 0 20424 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21712 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 21252 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_215
timestamp 1586364061
transform 1 0 20884 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_3  FILLER_2_221
timestamp 1586364061
transform 1 0 21436 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 23276 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 22724 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_233
timestamp 1586364061
transform 1 0 22540 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_237
timestamp 1586364061
transform 1 0 22908 0 -1 3808
box -38 -48 406 592
use scs8hd_decap_12  FILLER_2_244
timestamp 1586364061
transform 1 0 23552 0 -1 3808
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__050__C
timestamp 1586364061
transform 1 0 25300 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__A
timestamp 1586364061
transform 1 0 25668 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_6  FILLER_2_256
timestamp 1586364061
transform 1 0 24656 0 -1 3808
box -38 -48 590 592
use scs8hd_fill_1  FILLER_2_262
timestamp 1586364061
transform 1 0 25208 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_2_265
timestamp 1586364061
transform 1 0 25484 0 -1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 26496 0 -1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_65
timestamp 1586364061
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__050__B
timestamp 1586364061
transform 1 0 26036 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_269
timestamp 1586364061
transform 1 0 25852 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_273
timestamp 1586364061
transform 1 0 26220 0 -1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28244 0 -1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 27692 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28060 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_287
timestamp 1586364061
transform 1 0 27508 0 -1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_2_291
timestamp 1586364061
transform 1 0 27876 0 -1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_2_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29808 0 -1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__110__A
timestamp 1586364061
transform 1 0 29532 0 -1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30360 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_2_304
timestamp 1586364061
transform 1 0 29072 0 -1 3808
box -38 -48 406 592
use scs8hd_fill_1  FILLER_2_308
timestamp 1586364061
transform 1 0 29440 0 -1 3808
box -38 -48 130 592
use scs8hd_fill_1  FILLER_2_311
timestamp 1586364061
transform 1 0 29716 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_3  FILLER_2_315
timestamp 1586364061
transform 1 0 30084 0 -1 3808
box -38 -48 314 592
use scs8hd_decap_3  FILLER_2_320
timestamp 1586364061
transform 1 0 30544 0 -1 3808
box -38 -48 314 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_5_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_66
timestamp 1586364061
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_326
timestamp 1586364061
transform 1 0 31096 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_2  FILLER_2_334
timestamp 1586364061
transform 1 0 31832 0 -1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_2_337
timestamp 1586364061
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_349
timestamp 1586364061
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_361
timestamp 1586364061
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_373
timestamp 1586364061
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_2_385
timestamp 1586364061
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_5
timestamp 1586364061
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_67
timestamp 1586364061
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use scs8hd_decap_8  FILLER_2_398
timestamp 1586364061
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use scs8hd_fill_1  FILLER_2_406
timestamp 1586364061
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1748 0 1 3808
box -38 -48 866 592
use scs8hd_decap_3  PHY_6
timestamp 1586364061
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 1564 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_3
timestamp 1586364061
transform 1 0 1380 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_16
timestamp 1586364061
transform 1 0 2576 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 3312 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 3128 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_20
timestamp 1586364061
transform 1 0 2944 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_33
timestamp 1586364061
transform 1 0 4140 0 1 3808
box -38 -48 314 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 5152 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 4968 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__C
timestamp 1586364061
transform 1 0 4416 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_38
timestamp 1586364061
transform 1 0 4600 0 1 3808
box -38 -48 406 592
use scs8hd_fill_2  FILLER_3_53
timestamp 1586364061
transform 1 0 5980 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_68
timestamp 1586364061
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__085__D
timestamp 1586364061
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_57
timestamp 1586364061
transform 1 0 6348 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 9200 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8832 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8372 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_73
timestamp 1586364061
transform 1 0 7820 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_77
timestamp 1586364061
transform 1 0 8188 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_81
timestamp 1586364061
transform 1 0 8556 0 1 3808
box -38 -48 314 592
use scs8hd_fill_2  FILLER_3_86
timestamp 1586364061
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 9384 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__074__A
timestamp 1586364061
transform 1 0 10580 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__074__B
timestamp 1586364061
transform 1 0 10948 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_101
timestamp 1586364061
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_105
timestamp 1586364061
transform 1 0 10764 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_1_.latch
timestamp 1586364061
transform 1 0 12420 0 1 3808
box -38 -48 1050 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 3808
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_69
timestamp 1586364061
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 12144 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_109
timestamp 1586364061
transform 1 0 11132 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_114
timestamp 1586364061
transform 1 0 11592 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_118
timestamp 1586364061
transform 1 0 11960 0 1 3808
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 14168 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 13616 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 13984 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_134
timestamp 1586364061
transform 1 0 13432 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_138
timestamp 1586364061
transform 1 0 13800 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__064__A
timestamp 1586364061
transform 1 0 15364 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__B
timestamp 1586364061
transform 1 0 15732 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_153
timestamp 1586364061
transform 1 0 15180 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_157
timestamp 1586364061
transform 1 0 15548 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 15916 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__062__C
timestamp 1586364061
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__062__D
timestamp 1586364061
transform 1 0 17296 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_170
timestamp 1586364061
transform 1 0 16744 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_174
timestamp 1586364061
transform 1 0 17112 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_178
timestamp 1586364061
transform 1 0 17480 0 1 3808
box -38 -48 314 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_0_.latch
timestamp 1586364061
transform 1 0 18124 0 1 3808
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_70
timestamp 1586364061
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use scs8hd_fill_1  FILLER_3_184
timestamp 1586364061
transform 1 0 18032 0 1 3808
box -38 -48 130 592
use scs8hd_fill_2  FILLER_3_196
timestamp 1586364061
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19872 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20332 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 19688 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_200
timestamp 1586364061
transform 1 0 19504 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_207
timestamp 1586364061
transform 1 0 20148 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_211
timestamp 1586364061
transform 1 0 20516 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_2_.latch
timestamp 1586364061
transform 1 0 21252 0 1 3808
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 20884 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_217
timestamp 1586364061
transform 1 0 21068 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_230
timestamp 1586364061
transform 1 0 22264 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 23644 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_71
timestamp 1586364061
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 23368 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_2_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22448 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22816 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_234
timestamp 1586364061
transform 1 0 22632 0 1 3808
box -38 -48 222 592
use scs8hd_decap_4  FILLER_3_238
timestamp 1586364061
transform 1 0 23000 0 1 3808
box -38 -48 406 592
use scs8hd_nor4_4  _050_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 25300 0 1 3808
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__113__A
timestamp 1586364061
transform 1 0 24656 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__050__D
timestamp 1586364061
transform 1 0 25116 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_254
timestamp 1586364061
transform 1 0 24472 0 1 3808
box -38 -48 222 592
use scs8hd_decap_3  FILLER_3_258
timestamp 1586364061
transform 1 0 24840 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_2_.latch_D
timestamp 1586364061
transform 1 0 27048 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_280
timestamp 1586364061
transform 1 0 26864 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_284
timestamp 1586364061
transform 1 0 27232 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 3808
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 28612 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28980 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 27416 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_297
timestamp 1586364061
transform 1 0 28428 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_301
timestamp 1586364061
transform 1 0 28796 0 1 3808
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 3808
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_72
timestamp 1586364061
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30268 0 1 3808
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30636 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_315
timestamp 1586364061
transform 1 0 30084 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_319
timestamp 1586364061
transform 1 0 30452 0 1 3808
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 30820 0 1 3808
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 31280 0 1 3808
box -38 -48 222 592
use scs8hd_fill_2  FILLER_3_326
timestamp 1586364061
transform 1 0 31096 0 1 3808
box -38 -48 222 592
use scs8hd_decap_12  FILLER_3_330
timestamp 1586364061
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_342
timestamp 1586364061
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_354
timestamp 1586364061
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_73
timestamp 1586364061
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use scs8hd_decap_12  FILLER_3_367
timestamp 1586364061
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_379
timestamp 1586364061
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_3_391
timestamp 1586364061
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use scs8hd_decap_3  PHY_7
timestamp 1586364061
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use scs8hd_decap_4  FILLER_3_403
timestamp 1586364061
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 1472 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_8
timestamp 1586364061
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 2668 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_4_3
timestamp 1586364061
transform 1 0 1380 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_4_15
timestamp 1586364061
transform 1 0 2484 0 -1 4896
box -38 -48 222 592
use scs8hd_inv_8  _089_
timestamp 1586364061
transform 1 0 4048 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_74
timestamp 1586364061
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__084__B
timestamp 1586364061
transform 1 0 3772 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_8  FILLER_4_19
timestamp 1586364061
transform 1 0 2852 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_2  FILLER_4_27
timestamp 1586364061
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _085_
timestamp 1586364061
transform 1 0 5704 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__085__A
timestamp 1586364061
transform 1 0 5520 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__084__A
timestamp 1586364061
transform 1 0 5060 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_41
timestamp 1586364061
transform 1 0 4876 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_45
timestamp 1586364061
transform 1 0 5244 0 -1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__079__A
timestamp 1586364061
transform 1 0 7452 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_67
timestamp 1586364061
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_71
timestamp 1586364061
transform 1 0 7636 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 8004 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 7820 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_84
timestamp 1586364061
transform 1 0 8832 0 -1 4896
box -38 -48 590 592
use scs8hd_nor4_4  _074_
timestamp 1586364061
transform 1 0 10212 0 -1 4896
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_75
timestamp 1586364061
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__073__A
timestamp 1586364061
transform 1 0 10028 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__D
timestamp 1586364061
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_93
timestamp 1586364061
transform 1 0 9660 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__070__A
timestamp 1586364061
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__C
timestamp 1586364061
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_116
timestamp 1586364061
transform 1 0 11776 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_122
timestamp 1586364061
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 13432 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__071__D
timestamp 1586364061
transform 1 0 13248 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__070__D
timestamp 1586364061
transform 1 0 12880 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_126
timestamp 1586364061
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_130
timestamp 1586364061
transform 1 0 13064 0 -1 4896
box -38 -48 222 592
use scs8hd_buf_1  _064_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 15272 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_76
timestamp 1586364061
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__071__C
timestamp 1586364061
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 14996 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 15824 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_145
timestamp 1586364061
transform 1 0 14444 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_149
timestamp 1586364061
transform 1 0 14812 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_4_157
timestamp 1586364061
transform 1 0 15548 0 -1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _062_
timestamp 1586364061
transform 1 0 16744 0 -1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__063__A
timestamp 1586364061
transform 1 0 16560 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__B
timestamp 1586364061
transform 1 0 16192 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_162
timestamp 1586364061
transform 1 0 16008 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_166
timestamp 1586364061
transform 1 0 16376 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 18492 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_187
timestamp 1586364061
transform 1 0 18308 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_4_191
timestamp 1586364061
transform 1 0 18676 0 -1 4896
box -38 -48 590 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 19228 0 -1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_77
timestamp 1586364061
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__C
timestamp 1586364061
transform 1 0 20516 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_206
timestamp 1586364061
transform 1 0 20056 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_4_210
timestamp 1586364061
transform 1 0 20424 0 -1 4896
box -38 -48 130 592
use scs8hd_fill_1  FILLER_4_213
timestamp 1586364061
transform 1 0 20700 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_3_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 4896
box -38 -48 1050 592
use scs8hd_decap_8  FILLER_4_226
timestamp 1586364061
transform 1 0 21896 0 -1 4896
box -38 -48 774 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 22632 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 23644 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_243
timestamp 1586364061
transform 1 0 23460 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_247
timestamp 1586364061
transform 1 0 23828 0 -1 4896
box -38 -48 406 592
use scs8hd_buf_2  _113_
timestamp 1586364061
transform 1 0 24196 0 -1 4896
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__052__D
timestamp 1586364061
transform 1 0 25300 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__C
timestamp 1586364061
transform 1 0 25668 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__C
timestamp 1586364061
transform 1 0 24748 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_255
timestamp 1586364061
transform 1 0 24564 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_259
timestamp 1586364061
transform 1 0 24932 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_265
timestamp 1586364061
transform 1 0 25484 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_2_.latch
timestamp 1586364061
transform 1 0 26864 0 -1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_78
timestamp 1586364061
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__D
timestamp 1586364061
transform 1 0 26680 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__B
timestamp 1586364061
transform 1 0 26220 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_269
timestamp 1586364061
transform 1 0 25852 0 -1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_4_276
timestamp 1586364061
transform 1 0 26496 0 -1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_0_.latch
timestamp 1586364061
transform 1 0 28612 0 -1 4896
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28060 0 -1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_291
timestamp 1586364061
transform 1 0 27876 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_295
timestamp 1586364061
transform 1 0 28244 0 -1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30360 0 -1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 29808 0 -1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_4_310
timestamp 1586364061
transform 1 0 29624 0 -1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_4_314
timestamp 1586364061
transform 1 0 29992 0 -1 4896
box -38 -48 406 592
use scs8hd_tapvpwrvgnd_1  PHY_79
timestamp 1586364061
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_327
timestamp 1586364061
transform 1 0 31188 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_335
timestamp 1586364061
transform 1 0 31924 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_12  FILLER_4_337
timestamp 1586364061
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_349
timestamp 1586364061
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_361
timestamp 1586364061
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_373
timestamp 1586364061
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_4_385
timestamp 1586364061
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_9
timestamp 1586364061
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_80
timestamp 1586364061
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use scs8hd_decap_8  FILLER_4_398
timestamp 1586364061
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use scs8hd_fill_1  FILLER_4_406
timestamp 1586364061
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use scs8hd_lpflow_inputisolatch_1  mem_top_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 1564 0 1 4896
box -38 -48 1050 592
use scs8hd_decap_3  PHY_10
timestamp 1586364061
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_3
timestamp 1586364061
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_16
timestamp 1586364061
transform 1 0 2576 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 3312 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__080__A
timestamp 1586364061
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 3772 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 2760 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_SLEEPB
timestamp 1586364061
transform 1 0 3128 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_20
timestamp 1586364061
transform 1 0 2944 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_27
timestamp 1586364061
transform 1 0 3588 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_31
timestamp 1586364061
transform 1 0 3956 0 1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _084_
timestamp 1586364061
transform 1 0 4416 0 1 4896
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_5_53
timestamp 1586364061
transform 1 0 5980 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_0_.latch
timestamp 1586364061
transform 1 0 6808 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_81
timestamp 1586364061
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__079__B
timestamp 1586364061
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_57
timestamp 1586364061
transform 1 0 6348 0 1 4896
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 9016 0 1 4896
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8464 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__C
timestamp 1586364061
transform 1 0 8004 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 8832 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_73
timestamp 1586364061
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_77
timestamp 1586364061
transform 1 0 8188 0 1 4896
box -38 -48 314 592
use scs8hd_fill_2  FILLER_5_82
timestamp 1586364061
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_89
timestamp 1586364061
transform 1 0 9292 0 1 4896
box -38 -48 222 592
use scs8hd_nor4_4  _073_
timestamp 1586364061
transform 1 0 10028 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__068__B
timestamp 1586364061
transform 1 0 9844 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__A
timestamp 1586364061
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_93
timestamp 1586364061
transform 1 0 9660 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 12512 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_82
timestamp 1586364061
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__070__B
timestamp 1586364061
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__B
timestamp 1586364061
transform 1 0 11776 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_114
timestamp 1586364061
transform 1 0 11592 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_118
timestamp 1586364061
transform 1 0 11960 0 1 4896
box -38 -48 222 592
use scs8hd_fill_1  FILLER_5_123
timestamp 1586364061
transform 1 0 12420 0 1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _071_
timestamp 1586364061
transform 1 0 14076 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__071__A
timestamp 1586364061
transform 1 0 13892 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__071__B
timestamp 1586364061
transform 1 0 13524 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_133
timestamp 1586364061
transform 1 0 13340 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_137
timestamp 1586364061
transform 1 0 13708 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__039__A
timestamp 1586364061
transform 1 0 15824 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_158
timestamp 1586364061
transform 1 0 15640 0 1 4896
box -38 -48 222 592
use scs8hd_inv_8  _047_
timestamp 1586364061
transform 1 0 16376 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__047__A
timestamp 1586364061
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__063__C
timestamp 1586364061
transform 1 0 17388 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_162
timestamp 1586364061
transform 1 0 16008 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_175
timestamp 1586364061
transform 1 0 17204 0 1 4896
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_1_.latch
timestamp 1586364061
transform 1 0 18032 0 1 4896
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_83
timestamp 1586364061
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 17756 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_179
timestamp 1586364061
transform 1 0 17572 0 1 4896
box -38 -48 222 592
use scs8hd_decap_3  FILLER_5_195
timestamp 1586364061
transform 1 0 19044 0 1 4896
box -38 -48 314 592
use scs8hd_nor4_4  _059_
timestamp 1586364061
transform 1 0 20516 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 19688 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 20332 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__D
timestamp 1586364061
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_200
timestamp 1586364061
transform 1 0 19504 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_204
timestamp 1586364061
transform 1 0 19872 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_208
timestamp 1586364061
transform 1 0 20240 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__059__B
timestamp 1586364061
transform 1 0 22264 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_228
timestamp 1586364061
transform 1 0 22080 0 1 4896
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_84
timestamp 1586364061
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__046__D
timestamp 1586364061
transform 1 0 23368 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 22632 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_232
timestamp 1586364061
transform 1 0 22448 0 1 4896
box -38 -48 222 592
use scs8hd_decap_6  FILLER_5_236
timestamp 1586364061
transform 1 0 22816 0 1 4896
box -38 -48 590 592
use scs8hd_decap_4  FILLER_5_245
timestamp 1586364061
transform 1 0 23644 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_249
timestamp 1586364061
transform 1 0 24012 0 1 4896
box -38 -48 130 592
use scs8hd_nor4_4  _052_
timestamp 1586364061
transform 1 0 25300 0 1 4896
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__052__A
timestamp 1586364061
transform 1 0 25116 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__A
timestamp 1586364061
transform 1 0 24104 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__046__B
timestamp 1586364061
transform 1 0 24472 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_252
timestamp 1586364061
transform 1 0 24288 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_256
timestamp 1586364061
transform 1 0 24656 0 1 4896
box -38 -48 406 592
use scs8hd_fill_1  FILLER_5_260
timestamp 1586364061
transform 1 0 25024 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__049__C
timestamp 1586364061
transform 1 0 27048 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_280
timestamp 1586364061
transform 1 0 26864 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_284
timestamp 1586364061
transform 1 0 27232 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 27600 0 1 4896
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_D
timestamp 1586364061
transform 1 0 28796 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__049__A
timestamp 1586364061
transform 1 0 27416 0 1 4896
box -38 -48 222 592
use scs8hd_decap_4  FILLER_5_297
timestamp 1586364061
transform 1 0 28428 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_5_303
timestamp 1586364061
transform 1 0 28980 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29256 0 1 4896
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_85
timestamp 1586364061
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 30636 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_315
timestamp 1586364061
transform 1 0 30084 0 1 4896
box -38 -48 222 592
use scs8hd_fill_2  FILLER_5_319
timestamp 1586364061
transform 1 0 30452 0 1 4896
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 30820 0 1 4896
box -38 -48 866 592
use scs8hd_decap_12  FILLER_5_332
timestamp 1586364061
transform 1 0 31648 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_344
timestamp 1586364061
transform 1 0 32752 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_5_356
timestamp 1586364061
transform 1 0 33856 0 1 4896
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_86
timestamp 1586364061
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use scs8hd_fill_2  FILLER_5_364
timestamp 1586364061
transform 1 0 34592 0 1 4896
box -38 -48 222 592
use scs8hd_decap_12  FILLER_5_367
timestamp 1586364061
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_379
timestamp 1586364061
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_5_391
timestamp 1586364061
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use scs8hd_decap_3  PHY_11
timestamp 1586364061
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use scs8hd_decap_4  FILLER_5_403
timestamp 1586364061
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_7
timestamp 1586364061
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_7
timestamp 1586364061
transform 1 0 1748 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_3
timestamp 1586364061
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_top_ipin_1.LATCH_0_.latch_D
timestamp 1586364061
transform 1 0 1564 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  PHY_14
timestamp 1586364061
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_12
timestamp 1586364061
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use scs8hd_buf_2  _104_
timestamp 1586364061
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use scs8hd_decap_8  FILLER_7_15
timestamp 1586364061
transform 1 0 2484 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_11
timestamp 1586364061
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__104__A
timestamp 1586364061
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use scs8hd_ebufn_2  mux_top_ipin_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 1932 0 -1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_23
timestamp 1586364061
transform 1 0 3220 0 1 5984
box -38 -48 222 592
use scs8hd_conb_1  _097_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 3404 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_32
timestamp 1586364061
transform 1 0 4048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_28
timestamp 1586364061
transform 1 0 3680 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_32
timestamp 1586364061
transform 1 0 4048 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_1  FILLER_6_30
timestamp 1586364061
transform 1 0 3864 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__082__A
timestamp 1586364061
transform 1 0 3864 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__D
timestamp 1586364061
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_87
timestamp 1586364061
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_18
timestamp 1586364061
transform 1 0 2760 0 -1 5984
box -38 -48 1142 592
use scs8hd_inv_8  _080_
timestamp 1586364061
transform 1 0 4600 0 -1 5984
box -38 -48 866 592
use scs8hd_nor4_4  _082_
timestamp 1586364061
transform 1 0 4416 0 1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__084__D
timestamp 1586364061
transform 1 0 4416 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__D
timestamp 1586364061
transform 1 0 5612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__079__D
timestamp 1586364061
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_47
timestamp 1586364061
transform 1 0 5428 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_51
timestamp 1586364061
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_53
timestamp 1586364061
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _078_
timestamp 1586364061
transform 1 0 6808 0 1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _079_
timestamp 1586364061
transform 1 0 6164 0 -1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_94
timestamp 1586364061
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__078__B
timestamp 1586364061
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__083__A
timestamp 1586364061
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_57
timestamp 1586364061
transform 1 0 6348 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_79
timestamp 1586364061
transform 1 0 8372 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_76
timestamp 1586364061
transform 1 0 8096 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_72
timestamp 1586364061
transform 1 0 7728 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 8280 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 7912 0 -1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_2.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 8464 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_83
timestamp 1586364061
transform 1 0 8740 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_89
timestamp 1586364061
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_6  FILLER_6_83
timestamp 1586364061
transform 1 0 8740 0 -1 5984
box -38 -48 590 592
use scs8hd_diode_2  ANTENNA__087__A
timestamp 1586364061
transform 1 0 8924 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__C
timestamp 1586364061
transform 1 0 8556 0 1 5984
box -38 -48 222 592
use scs8hd_inv_8  _087_
timestamp 1586364061
transform 1 0 9108 0 1 5984
box -38 -48 866 592
use scs8hd_fill_2  FILLER_7_96
timestamp 1586364061
transform 1 0 9936 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_93
timestamp 1586364061
transform 1 0 9660 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__068__D
timestamp 1586364061
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__068__C
timestamp 1586364061
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__073__C
timestamp 1586364061
transform 1 0 9936 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_88
timestamp 1586364061
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_7_107
timestamp 1586364061
transform 1 0 10948 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_104
timestamp 1586364061
transform 1 0 10672 0 1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_100
timestamp 1586364061
transform 1 0 10304 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 10764 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _068_
timestamp 1586364061
transform 1 0 10120 0 -1 5984
box -38 -48 1602 592
use scs8hd_fill_2  FILLER_7_114
timestamp 1586364061
transform 1 0 11592 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_115
timestamp 1586364061
transform 1 0 11684 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__B
timestamp 1586364061
transform 1 0 11132 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 11316 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_118
timestamp 1586364061
transform 1 0 11960 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_119
timestamp 1586364061
transform 1 0 12052 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__066__C
timestamp 1586364061
transform 1 0 12328 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__076__A
timestamp 1586364061
transform 1 0 11868 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__081__B
timestamp 1586364061
transform 1 0 12144 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_top_ipin_0.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 11776 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_95
timestamp 1586364061
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use scs8hd_or2_4  _081_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12420 0 1 5984
box -38 -48 682 592
use scs8hd_nor4_4  _070_
timestamp 1586364061
transform 1 0 12512 0 -1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _072_
timestamp 1586364061
transform 1 0 13892 0 1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__081__A
timestamp 1586364061
transform 1 0 13248 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__066__B
timestamp 1586364061
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_141
timestamp 1586364061
transform 1 0 14076 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_130
timestamp 1586364061
transform 1 0 13064 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_134
timestamp 1586364061
transform 1 0 13432 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_7_138
timestamp 1586364061
transform 1 0 13800 0 1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_149
timestamp 1586364061
transform 1 0 14812 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_145
timestamp 1586364061
transform 1 0 14444 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__D
timestamp 1586364061
transform 1 0 14628 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__B
timestamp 1586364061
transform 1 0 14260 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__B
timestamp 1586364061
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_160
timestamp 1586364061
transform 1 0 15824 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_156
timestamp 1586364061
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__A
timestamp 1586364061
transform 1 0 15640 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_89
timestamp 1586364061
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use scs8hd_inv_8  _039_
timestamp 1586364061
transform 1 0 15272 0 -1 5984
box -38 -48 866 592
use scs8hd_decap_4  FILLER_6_167
timestamp 1586364061
transform 1 0 16468 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_6_163
timestamp 1586364061
transform 1 0 16100 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__D
timestamp 1586364061
transform 1 0 16284 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__038__A
timestamp 1586364061
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use scs8hd_decap_6  FILLER_7_177
timestamp 1586364061
transform 1 0 17388 0 1 5984
box -38 -48 590 592
use scs8hd_fill_2  FILLER_7_173
timestamp 1586364061
transform 1 0 17020 0 1 5984
box -38 -48 222 592
use scs8hd_fill_1  FILLER_6_171
timestamp 1586364061
transform 1 0 16836 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__063__D
timestamp 1586364061
transform 1 0 16928 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__061__A
timestamp 1586364061
transform 1 0 17204 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _063_
timestamp 1586364061
transform 1 0 17112 0 -1 5984
box -38 -48 1602 592
use scs8hd_inv_8  _038_
timestamp 1586364061
transform 1 0 16192 0 1 5984
box -38 -48 866 592
use scs8hd_buf_1  _060_
timestamp 1586364061
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_96
timestamp 1586364061
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__060__A
timestamp 1586364061
transform 1 0 18492 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__055__A
timestamp 1586364061
transform 1 0 18860 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_191
timestamp 1586364061
transform 1 0 18676 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_187
timestamp 1586364061
transform 1 0 18308 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_191
timestamp 1586364061
transform 1 0 18676 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_7_195
timestamp 1586364061
transform 1 0 19044 0 1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_201
timestamp 1586364061
transform 1 0 19596 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_205
timestamp 1586364061
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_6_199
timestamp 1586364061
transform 1 0 19412 0 -1 5984
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__058__A
timestamp 1586364061
transform 1 0 19412 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__C
timestamp 1586364061
transform 1 0 19780 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_2.INVTX1_3_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 19688 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_1  FILLER_6_213
timestamp 1586364061
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use scs8hd_fill_2  FILLER_6_209
timestamp 1586364061
transform 1 0 20332 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__B
timestamp 1586364061
transform 1 0 20148 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__059__A
timestamp 1586364061
transform 1 0 20516 0 -1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_90
timestamp 1586364061
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use scs8hd_nor4_4  _058_
timestamp 1586364061
transform 1 0 19964 0 1 5984
box -38 -48 1602 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_4_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 5984
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA__056__A
timestamp 1586364061
transform 1 0 21712 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__B
timestamp 1586364061
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_226
timestamp 1586364061
transform 1 0 21896 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_222
timestamp 1586364061
transform 1 0 21528 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_226
timestamp 1586364061
transform 1 0 21896 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_230
timestamp 1586364061
transform 1 0 22264 0 1 5984
box -38 -48 222 592
use scs8hd_buf_1  _045_
timestamp 1586364061
transform 1 0 23644 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_97
timestamp 1586364061
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__056__C
timestamp 1586364061
transform 1 0 22448 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_238
timestamp 1586364061
transform 1 0 23000 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_234
timestamp 1586364061
transform 1 0 22632 0 1 5984
box -38 -48 774 592
use scs8hd_fill_2  FILLER_7_242
timestamp 1586364061
transform 1 0 23368 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_248
timestamp 1586364061
transform 1 0 23920 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _046_
timestamp 1586364061
transform 1 0 24104 0 -1 5984
box -38 -48 1602 592
use scs8hd_nor4_4  _051_
timestamp 1586364061
transform 1 0 25116 0 1 5984
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__045__A
timestamp 1586364061
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__A
timestamp 1586364061
transform 1 0 24932 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__C
timestamp 1586364061
transform 1 0 24564 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_6_267
timestamp 1586364061
transform 1 0 25668 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_252
timestamp 1586364061
transform 1 0 24288 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_257
timestamp 1586364061
transform 1 0 24748 0 1 5984
box -38 -48 222 592
use scs8hd_nor4_4  _049_
timestamp 1586364061
transform 1 0 26496 0 -1 5984
box -38 -48 1602 592
use scs8hd_tapvpwrvgnd_1  PHY_91
timestamp 1586364061
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 27232 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__052__B
timestamp 1586364061
transform 1 0 25852 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 26864 0 1 5984
box -38 -48 222 592
use scs8hd_decap_4  FILLER_6_271
timestamp 1586364061
transform 1 0 26036 0 -1 5984
box -38 -48 406 592
use scs8hd_fill_2  FILLER_7_278
timestamp 1586364061
transform 1 0 26680 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_282
timestamp 1586364061
transform 1 0 27048 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_292
timestamp 1586364061
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_286
timestamp 1586364061
transform 1 0 27416 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_293
timestamp 1586364061
transform 1 0 28060 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 28152 0 1 5984
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.INVTX1_4_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 27692 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_301
timestamp 1586364061
transform 1 0 28796 0 1 5984
box -38 -48 222 592
use scs8hd_decap_3  FILLER_7_296
timestamp 1586364061
transform 1 0 28336 0 1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_6_297
timestamp 1586364061
transform 1 0 28428 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28244 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_4_.latch_SLEEPB
timestamp 1586364061
transform 1 0 28612 0 -1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28612 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_D
timestamp 1586364061
transform 1 0 28980 0 1 5984
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_4_.latch
timestamp 1586364061
transform 1 0 28796 0 -1 5984
box -38 -48 1050 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_3_.latch
timestamp 1586364061
transform 1 0 29256 0 1 5984
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_98
timestamp 1586364061
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_0.LATCH_3_.latch_SLEEPB
timestamp 1586364061
transform 1 0 30452 0 1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_312
timestamp 1586364061
transform 1 0 29808 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_320
timestamp 1586364061
transform 1 0 30544 0 -1 5984
box -38 -48 314 592
use scs8hd_fill_2  FILLER_7_317
timestamp 1586364061
transform 1 0 30268 0 1 5984
box -38 -48 222 592
use scs8hd_fill_2  FILLER_7_321
timestamp 1586364061
transform 1 0 30636 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_92
timestamp 1586364061
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 1 5984
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 30820 0 -1 5984
box -38 -48 222 592
use scs8hd_decap_8  FILLER_6_325
timestamp 1586364061
transform 1 0 31004 0 -1 5984
box -38 -48 774 592
use scs8hd_decap_3  FILLER_6_333
timestamp 1586364061
transform 1 0 31740 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_12  FILLER_6_337
timestamp 1586364061
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_325
timestamp 1586364061
transform 1 0 31004 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_337
timestamp 1586364061
transform 1 0 32108 0 1 5984
box -38 -48 1142 592
use scs8hd_buf_2  _111_
timestamp 1586364061
transform 1 0 33212 0 1 5984
box -38 -48 406 592
use scs8hd_diode_2  ANTENNA__111__A
timestamp 1586364061
transform 1 0 33764 0 1 5984
box -38 -48 222 592
use scs8hd_decap_12  FILLER_6_349
timestamp 1586364061
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_7_353
timestamp 1586364061
transform 1 0 33580 0 1 5984
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_99
timestamp 1586364061
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_6_361
timestamp 1586364061
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_373
timestamp 1586364061
transform 1 0 35420 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_7_357
timestamp 1586364061
transform 1 0 33948 0 1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_7_365
timestamp 1586364061
transform 1 0 34684 0 1 5984
box -38 -48 130 592
use scs8hd_decap_12  FILLER_7_367
timestamp 1586364061
transform 1 0 34868 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_6_385
timestamp 1586364061
transform 1 0 36524 0 -1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_379
timestamp 1586364061
transform 1 0 35972 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_7_391
timestamp 1586364061
transform 1 0 37076 0 1 5984
box -38 -48 1142 592
use scs8hd_decap_3  PHY_13
timestamp 1586364061
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use scs8hd_decap_3  PHY_15
timestamp 1586364061
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_93
timestamp 1586364061
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_8  FILLER_6_398
timestamp 1586364061
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use scs8hd_fill_1  FILLER_6_406
timestamp 1586364061
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use scs8hd_decap_4  FILLER_7_403
timestamp 1586364061
transform 1 0 38180 0 1 5984
box -38 -48 406 592
use scs8hd_inv_1  mux_top_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_16
timestamp 1586364061
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_6
timestamp 1586364061
transform 1 0 1656 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _093_
timestamp 1586364061
transform 1 0 4140 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_100
timestamp 1586364061
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_12  FILLER_8_18
timestamp 1586364061
transform 1 0 2760 0 -1 7072
box -38 -48 1142 592
use scs8hd_fill_1  FILLER_8_30
timestamp 1586364061
transform 1 0 3864 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_1  FILLER_8_32
timestamp 1586364061
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use scs8hd_nor4_4  _083_
timestamp 1586364061
transform 1 0 5152 0 -1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__083__B
timestamp 1586364061
transform 1 0 4968 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__B
timestamp 1586364061
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_36
timestamp 1586364061
transform 1 0 4416 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_40
timestamp 1586364061
transform 1 0 4784 0 -1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 7452 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__078__D
timestamp 1586364061
transform 1 0 6900 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__078__A
timestamp 1586364061
transform 1 0 7268 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_61
timestamp 1586364061
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_65
timestamp 1586364061
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_78
timestamp 1586364061
transform 1 0 8280 0 -1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _095_
timestamp 1586364061
transform 1 0 9660 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_101
timestamp 1586364061
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_90
timestamp 1586364061
transform 1 0 9384 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_8_96
timestamp 1586364061
transform 1 0 9936 0 -1 7072
box -38 -48 1142 592
use scs8hd_or2_4  _076_
timestamp 1586364061
transform 1 0 11592 0 -1 7072
box -38 -48 682 592
use scs8hd_diode_2  ANTENNA__066__A
timestamp 1586364061
transform 1 0 12420 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_8_108
timestamp 1586364061
transform 1 0 11040 0 -1 7072
box -38 -48 590 592
use scs8hd_fill_2  FILLER_8_121
timestamp 1586364061
transform 1 0 12236 0 -1 7072
box -38 -48 222 592
use scs8hd_or4_4  _066_ tech/SW/EFS8A/libs.ref/mag/scs8hd
timestamp 1586364061
transform 1 0 12972 0 -1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__066__D
timestamp 1586364061
transform 1 0 12788 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__A
timestamp 1586364061
transform 1 0 13984 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_125
timestamp 1586364061
transform 1 0 12604 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_138
timestamp 1586364061
transform 1 0 13800 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_142
timestamp 1586364061
transform 1 0 14168 0 -1 7072
box -38 -48 406 592
use scs8hd_or4_4  _054_
timestamp 1586364061
transform 1 0 15640 0 -1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_102
timestamp 1586364061
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__053__A
timestamp 1586364061
transform 1 0 14628 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__040__A
timestamp 1586364061
transform 1 0 15456 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__054__C
timestamp 1586364061
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_8_146
timestamp 1586364061
transform 1 0 14536 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_149
timestamp 1586364061
transform 1 0 14812 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_154
timestamp 1586364061
transform 1 0 15272 0 -1 7072
box -38 -48 222 592
use scs8hd_buf_1  _061_
timestamp 1586364061
transform 1 0 17204 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_167
timestamp 1586364061
transform 1 0 16468 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_178
timestamp 1586364061
transform 1 0 17480 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _055_
timestamp 1586364061
transform 1 0 18216 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_189
timestamp 1586364061
transform 1 0 18492 0 -1 7072
box -38 -48 774 592
use scs8hd_conb_1  _094_
timestamp 1586364061
transform 1 0 19780 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_103
timestamp 1586364061
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__B
timestamp 1586364061
transform 1 0 19504 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__058__D
timestamp 1586364061
transform 1 0 20240 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__056__D
timestamp 1586364061
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_197
timestamp 1586364061
transform 1 0 19228 0 -1 7072
box -38 -48 314 592
use scs8hd_fill_1  FILLER_8_202
timestamp 1586364061
transform 1 0 19688 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_206
timestamp 1586364061
transform 1 0 20056 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_210
timestamp 1586364061
transform 1 0 20424 0 -1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _056_
timestamp 1586364061
transform 1 0 20884 0 -1 7072
box -38 -48 1602 592
use scs8hd_decap_12  FILLER_8_232
timestamp 1586364061
transform 1 0 22448 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_8_244
timestamp 1586364061
transform 1 0 23552 0 -1 7072
box -38 -48 774 592
use scs8hd_buf_1  _043_
timestamp 1586364061
transform 1 0 24472 0 -1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__044__B
timestamp 1586364061
transform 1 0 25208 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__043__A
timestamp 1586364061
transform 1 0 24288 0 -1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__051__D
timestamp 1586364061
transform 1 0 25576 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_8_257
timestamp 1586364061
transform 1 0 24748 0 -1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_8_261
timestamp 1586364061
transform 1 0 25116 0 -1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_8_264
timestamp 1586364061
transform 1 0 25392 0 -1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_0.LATCH_5_.latch
timestamp 1586364061
transform 1 0 27232 0 -1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_104
timestamp 1586364061
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__051__B
timestamp 1586364061
transform 1 0 25944 0 -1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_8_268
timestamp 1586364061
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_8_272
timestamp 1586364061
transform 1 0 26128 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_8_276
timestamp 1586364061
transform 1 0 26496 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_8  FILLER_8_295
timestamp 1586364061
transform 1 0 28244 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_303
timestamp 1586364061
transform 1 0 28980 0 -1 7072
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 29072 0 -1 7072
box -38 -48 866 592
use scs8hd_decap_12  FILLER_8_313
timestamp 1586364061
transform 1 0 29900 0 -1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_105
timestamp 1586364061
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_325
timestamp 1586364061
transform 1 0 31004 0 -1 7072
box -38 -48 774 592
use scs8hd_decap_3  FILLER_8_333
timestamp 1586364061
transform 1 0 31740 0 -1 7072
box -38 -48 314 592
use scs8hd_decap_12  FILLER_8_337
timestamp 1586364061
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_349
timestamp 1586364061
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_361
timestamp 1586364061
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_373
timestamp 1586364061
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_8_385
timestamp 1586364061
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_17
timestamp 1586364061
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_106
timestamp 1586364061
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_8_398
timestamp 1586364061
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use scs8hd_fill_1  FILLER_8_406
timestamp 1586364061
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use scs8hd_conb_1  _096_
timestamp 1586364061
transform 1 0 1380 0 1 7072
box -38 -48 314 592
use scs8hd_decap_3  PHY_18
timestamp 1586364061
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__102__A
timestamp 1586364061
transform 1 0 1840 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_6
timestamp 1586364061
transform 1 0 1656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_10
timestamp 1586364061
transform 1 0 2024 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_22
timestamp 1586364061
transform 1 0 3128 0 1 7072
box -38 -48 1142 592
use scs8hd_fill_2  FILLER_9_34
timestamp 1586364061
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _086_
timestamp 1586364061
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__083__C
timestamp 1586364061
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__082__C
timestamp 1586364061
transform 1 0 4416 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_38
timestamp 1586364061
transform 1 0 4600 0 1 7072
box -38 -48 406 592
use scs8hd_fill_2  FILLER_9_53
timestamp 1586364061
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_1.LATCH_1_.latch
timestamp 1586364061
transform 1 0 6808 0 1 7072
box -38 -48 1050 592
use scs8hd_tapvpwrvgnd_1  PHY_107
timestamp 1586364061
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_D
timestamp 1586364061
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_57
timestamp 1586364061
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use scs8hd_buf_1  _077_
timestamp 1586364061
transform 1 0 8556 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__077__A
timestamp 1586364061
transform 1 0 9016 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_1.LATCH_1_.latch_SLEEPB
timestamp 1586364061
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_73
timestamp 1586364061
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_77
timestamp 1586364061
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_84
timestamp 1586364061
transform 1 0 8832 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_88
timestamp 1586364061
transform 1 0 9200 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_100
timestamp 1586364061
transform 1 0 10304 0 1 7072
box -38 -48 1142 592
use scs8hd_inv_8  _065_
timestamp 1586364061
transform 1 0 12420 0 1 7072
box -38 -48 866 592
use scs8hd_tapvpwrvgnd_1  PHY_108
timestamp 1586364061
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__065__A
timestamp 1586364061
transform 1 0 12144 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_112
timestamp 1586364061
transform 1 0 11408 0 1 7072
box -38 -48 774 592
use scs8hd_diode_2  ANTENNA__069__A
timestamp 1586364061
transform 1 0 14168 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__067__A
timestamp 1586364061
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__072__C
timestamp 1586364061
transform 1 0 13800 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_132
timestamp 1586364061
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_136
timestamp 1586364061
transform 1 0 13616 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_140
timestamp 1586364061
transform 1 0 13984 0 1 7072
box -38 -48 222 592
use scs8hd_inv_8  _053_
timestamp 1586364061
transform 1 0 14628 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__042__B
timestamp 1586364061
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_144
timestamp 1586364061
transform 1 0 14352 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_156
timestamp 1586364061
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_160
timestamp 1586364061
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use scs8hd_or4_4  _042_
timestamp 1586364061
transform 1 0 16192 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__048__A
timestamp 1586364061
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__C
timestamp 1586364061
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_173
timestamp 1586364061
transform 1 0 17020 0 1 7072
box -38 -48 222 592
use scs8hd_decap_6  FILLER_9_177
timestamp 1586364061
transform 1 0 17388 0 1 7072
box -38 -48 590 592
use scs8hd_buf_1  _037_
timestamp 1586364061
transform 1 0 18032 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_109
timestamp 1586364061
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__037__A
timestamp 1586364061
transform 1 0 18492 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__057__D
timestamp 1586364061
transform 1 0 18952 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_187
timestamp 1586364061
transform 1 0 18308 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_191
timestamp 1586364061
transform 1 0 18676 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_196
timestamp 1586364061
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use scs8hd_nor4_4  _057_
timestamp 1586364061
transform 1 0 19504 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__057__A
timestamp 1586364061
transform 1 0 19320 0 1 7072
box -38 -48 222 592
use scs8hd_ebufn_2  mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 21804 0 1 7072
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_D
timestamp 1586364061
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_217
timestamp 1586364061
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_221
timestamp 1586364061
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use scs8hd_tapvpwrvgnd_1  PHY_110
timestamp 1586364061
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use scs8hd_decap_8  FILLER_9_234
timestamp 1586364061
transform 1 0 22632 0 1 7072
box -38 -48 774 592
use scs8hd_fill_2  FILLER_9_242
timestamp 1586364061
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use scs8hd_decap_8  FILLER_9_245
timestamp 1586364061
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use scs8hd_nor4_4  _044_
timestamp 1586364061
transform 1 0 25208 0 1 7072
box -38 -48 1602 592
use scs8hd_diode_2  ANTENNA__044__A
timestamp 1586364061
transform 1 0 25024 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__044__D
timestamp 1586364061
transform 1 0 24656 0 1 7072
box -38 -48 222 592
use scs8hd_decap_3  FILLER_9_253
timestamp 1586364061
transform 1 0 24380 0 1 7072
box -38 -48 314 592
use scs8hd_fill_2  FILLER_9_258
timestamp 1586364061
transform 1 0 24840 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_279
timestamp 1586364061
transform 1 0 26772 0 1 7072
box -38 -48 1142 592
use scs8hd_conb_1  _092_
timestamp 1586364061
transform 1 0 27968 0 1 7072
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 28428 0 1 7072
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 28796 0 1 7072
box -38 -48 222 592
use scs8hd_fill_1  FILLER_9_291
timestamp 1586364061
transform 1 0 27876 0 1 7072
box -38 -48 130 592
use scs8hd_fill_2  FILLER_9_295
timestamp 1586364061
transform 1 0 28244 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_299
timestamp 1586364061
transform 1 0 28612 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_303
timestamp 1586364061
transform 1 0 28980 0 1 7072
box -38 -48 222 592
use scs8hd_inv_1  mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 29256 0 1 7072
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_111
timestamp 1586364061
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_0.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 29716 0 1 7072
box -38 -48 222 592
use scs8hd_fill_2  FILLER_9_309
timestamp 1586364061
transform 1 0 29532 0 1 7072
box -38 -48 222 592
use scs8hd_decap_12  FILLER_9_313
timestamp 1586364061
transform 1 0 29900 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_325
timestamp 1586364061
transform 1 0 31004 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_337
timestamp 1586364061
transform 1 0 32108 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_349
timestamp 1586364061
transform 1 0 33212 0 1 7072
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_112
timestamp 1586364061
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__108__A
timestamp 1586364061
transform 1 0 35420 0 1 7072
box -38 -48 222 592
use scs8hd_decap_4  FILLER_9_361
timestamp 1586364061
transform 1 0 34316 0 1 7072
box -38 -48 406 592
use scs8hd_fill_1  FILLER_9_365
timestamp 1586364061
transform 1 0 34684 0 1 7072
box -38 -48 130 592
use scs8hd_decap_6  FILLER_9_367
timestamp 1586364061
transform 1 0 34868 0 1 7072
box -38 -48 590 592
use scs8hd_decap_12  FILLER_9_375
timestamp 1586364061
transform 1 0 35604 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_9_387
timestamp 1586364061
transform 1 0 36708 0 1 7072
box -38 -48 1142 592
use scs8hd_decap_3  PHY_19
timestamp 1586364061
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use scs8hd_decap_8  FILLER_9_399
timestamp 1586364061
transform 1 0 37812 0 1 7072
box -38 -48 774 592
use scs8hd_buf_2  _102_
timestamp 1586364061
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_3  PHY_20
timestamp 1586364061
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_7
timestamp 1586364061
transform 1 0 1748 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_113
timestamp 1586364061
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_19
timestamp 1586364061
transform 1 0 2852 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_32
timestamp 1586364061
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 5796 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__086__A
timestamp 1586364061
transform 1 0 5152 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_46
timestamp 1586364061
transform 1 0 5336 0 -1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_10_50
timestamp 1586364061
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use scs8hd_ebufn_2  mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 6808 0 -1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A
timestamp 1586364061
transform 1 0 6624 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_6  FILLER_10_54
timestamp 1586364061
transform 1 0 6072 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_71
timestamp 1586364061
transform 1 0 7636 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_83
timestamp 1586364061
transform 1 0 8740 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_114
timestamp 1586364061
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use scs8hd_fill_1  FILLER_10_91
timestamp 1586364061
transform 1 0 9476 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_93
timestamp 1586364061
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_105
timestamp 1586364061
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_117
timestamp 1586364061
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_1  _067_
timestamp 1586364061
transform 1 0 13156 0 -1 8160
box -38 -48 314 592
use scs8hd_buf_1  _069_
timestamp 1586364061
transform 1 0 14168 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_129
timestamp 1586364061
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_134
timestamp 1586364061
transform 1 0 13432 0 -1 8160
box -38 -48 774 592
use scs8hd_buf_1  _040_
timestamp 1586364061
transform 1 0 15640 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_115
timestamp 1586364061
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_145
timestamp 1586364061
transform 1 0 14444 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_4  FILLER_10_154
timestamp 1586364061
transform 1 0 15272 0 -1 8160
box -38 -48 406 592
use scs8hd_buf_1  _048_
timestamp 1586364061
transform 1 0 17112 0 -1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__042__A
timestamp 1586364061
transform 1 0 16192 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA__042__D
timestamp 1586364061
transform 1 0 16560 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_161
timestamp 1586364061
transform 1 0 15916 0 -1 8160
box -38 -48 314 592
use scs8hd_fill_2  FILLER_10_166
timestamp 1586364061
transform 1 0 16376 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_4  FILLER_10_170
timestamp 1586364061
transform 1 0 16744 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_177
timestamp 1586364061
transform 1 0 17388 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_189
timestamp 1586364061
transform 1 0 18492 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_116
timestamp 1586364061
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__057__C
timestamp 1586364061
transform 1 0 19504 0 -1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mem_bottom_ipin_2.LATCH_5_.latch_SLEEPB
timestamp 1586364061
transform 1 0 20608 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_3  FILLER_10_197
timestamp 1586364061
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_8  FILLER_10_202
timestamp 1586364061
transform 1 0 19688 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_2  FILLER_10_210
timestamp 1586364061
transform 1 0 20424 0 -1 8160
box -38 -48 222 592
use scs8hd_lpflow_inputisolatch_1  mem_bottom_ipin_2.LATCH_5_.latch
timestamp 1586364061
transform 1 0 20884 0 -1 8160
box -38 -48 1050 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB
timestamp 1586364061
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_10_226
timestamp 1586364061
transform 1 0 21896 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_10_230
timestamp 1586364061
transform 1 0 22264 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_242
timestamp 1586364061
transform 1 0 23368 0 -1 8160
box -38 -48 1142 592
use scs8hd_diode_2  ANTENNA__044__C
timestamp 1586364061
transform 1 0 25208 0 -1 8160
box -38 -48 222 592
use scs8hd_decap_8  FILLER_10_254
timestamp 1586364061
transform 1 0 24472 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_8  FILLER_10_264
timestamp 1586364061
transform 1 0 25392 0 -1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_117
timestamp 1586364061
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_3  FILLER_10_272
timestamp 1586364061
transform 1 0 26128 0 -1 8160
box -38 -48 314 592
use scs8hd_decap_12  FILLER_10_276
timestamp 1586364061
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use scs8hd_ebufn_2  mux_bottom_ipin_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2
timestamp 1586364061
transform 1 0 28152 0 -1 8160
box -38 -48 866 592
use scs8hd_decap_6  FILLER_10_288
timestamp 1586364061
transform 1 0 27600 0 -1 8160
box -38 -48 590 592
use scs8hd_decap_12  FILLER_10_303
timestamp 1586364061
transform 1 0 28980 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_315
timestamp 1586364061
transform 1 0 30084 0 -1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_118
timestamp 1586364061
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_327
timestamp 1586364061
transform 1 0 31188 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_335
timestamp 1586364061
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_10_337
timestamp 1586364061
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_349
timestamp 1586364061
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use scs8hd_buf_2  _108_
timestamp 1586364061
transform 1 0 35420 0 -1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_10_361
timestamp 1586364061
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_10_377
timestamp 1586364061
transform 1 0 35788 0 -1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_10_389
timestamp 1586364061
transform 1 0 36892 0 -1 8160
box -38 -48 774 592
use scs8hd_decap_3  PHY_21
timestamp 1586364061
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_119
timestamp 1586364061
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_10_398
timestamp 1586364061
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use scs8hd_fill_1  FILLER_10_406
timestamp 1586364061
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use scs8hd_inv_1  mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 1380 0 1 8160
box -38 -48 314 592
use scs8hd_decap_3  PHY_22
timestamp 1586364061
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA__099__A
timestamp 1586364061
transform 1 0 1840 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 2208 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_6
timestamp 1586364061
transform 1 0 1656 0 1 8160
box -38 -48 222 592
use scs8hd_fill_2  FILLER_11_10
timestamp 1586364061
transform 1 0 2024 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_14
timestamp 1586364061
transform 1 0 2392 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_26
timestamp 1586364061
transform 1 0 3496 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_38
timestamp 1586364061
transform 1 0 4600 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_11_50
timestamp 1586364061
transform 1 0 5704 0 1 8160
box -38 -48 774 592
use scs8hd_inv_1  mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 6808 0 1 8160
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_120
timestamp 1586364061
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use scs8hd_diode_2  ANTENNA__075__A
timestamp 1586364061
transform 1 0 6440 0 1 8160
box -38 -48 222 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_1.INVTX1_1_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_60
timestamp 1586364061
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_65
timestamp 1586364061
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_69
timestamp 1586364061
transform 1 0 7452 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_81
timestamp 1586364061
transform 1 0 8556 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_93
timestamp 1586364061
transform 1 0 9660 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_105
timestamp 1586364061
transform 1 0 10764 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_121
timestamp 1586364061
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_117
timestamp 1586364061
transform 1 0 11868 0 1 8160
box -38 -48 406 592
use scs8hd_fill_1  FILLER_11_121
timestamp 1586364061
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_123
timestamp 1586364061
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_135
timestamp 1586364061
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_147
timestamp 1586364061
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_11_159
timestamp 1586364061
transform 1 0 15732 0 1 8160
box -38 -48 406 592
use scs8hd_inv_8  _041_
timestamp 1586364061
transform 1 0 16376 0 1 8160
box -38 -48 866 592
use scs8hd_diode_2  ANTENNA__041__A
timestamp 1586364061
transform 1 0 16192 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_163
timestamp 1586364061
transform 1 0 16100 0 1 8160
box -38 -48 130 592
use scs8hd_decap_8  FILLER_11_175
timestamp 1586364061
transform 1 0 17204 0 1 8160
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_122
timestamp 1586364061
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_184
timestamp 1586364061
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_196
timestamp 1586364061
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use scs8hd_inv_1  mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1
timestamp 1586364061
transform 1 0 20332 0 1 8160
box -38 -48 314 592
use scs8hd_diode_2  ANTENNA_mux_bottom_ipin_2.tap_buf4_0_.scs8hd_inv_1_A
timestamp 1586364061
transform 1 0 20792 0 1 8160
box -38 -48 222 592
use scs8hd_fill_1  FILLER_11_208
timestamp 1586364061
transform 1 0 20240 0 1 8160
box -38 -48 130 592
use scs8hd_fill_2  FILLER_11_212
timestamp 1586364061
transform 1 0 20608 0 1 8160
box -38 -48 222 592
use scs8hd_decap_12  FILLER_11_216
timestamp 1586364061
transform 1 0 20976 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_228
timestamp 1586364061
transform 1 0 22080 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_123
timestamp 1586364061
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use scs8hd_decap_4  FILLER_11_240
timestamp 1586364061
transform 1 0 23184 0 1 8160
box -38 -48 406 592
use scs8hd_decap_12  FILLER_11_245
timestamp 1586364061
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_257
timestamp 1586364061
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_269
timestamp 1586364061
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_281
timestamp 1586364061
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_293
timestamp 1586364061
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_124
timestamp 1586364061
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_306
timestamp 1586364061
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_318
timestamp 1586364061
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_330
timestamp 1586364061
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_342
timestamp 1586364061
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_354
timestamp 1586364061
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_125
timestamp 1586364061
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use scs8hd_decap_12  FILLER_11_367
timestamp 1586364061
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_379
timestamp 1586364061
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_11_391
timestamp 1586364061
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use scs8hd_decap_3  PHY_23
timestamp 1586364061
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use scs8hd_decap_4  FILLER_11_403
timestamp 1586364061
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use scs8hd_buf_2  _099_
timestamp 1586364061
transform 1 0 1380 0 -1 9248
box -38 -48 406 592
use scs8hd_decap_3  PHY_24
timestamp 1586364061
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use scs8hd_decap_12  FILLER_12_7
timestamp 1586364061
transform 1 0 1748 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_126
timestamp 1586364061
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_19
timestamp 1586364061
transform 1 0 2852 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_32
timestamp 1586364061
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_44
timestamp 1586364061
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use scs8hd_buf_1  _075_
timestamp 1586364061
transform 1 0 6440 0 -1 9248
box -38 -48 314 592
use scs8hd_fill_2  FILLER_12_56
timestamp 1586364061
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_12_61
timestamp 1586364061
transform 1 0 6716 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_73
timestamp 1586364061
transform 1 0 7820 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_12_85
timestamp 1586364061
transform 1 0 8924 0 -1 9248
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_127
timestamp 1586364061
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use scs8hd_fill_1  FILLER_12_91
timestamp 1586364061
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_93
timestamp 1586364061
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_105
timestamp 1586364061
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_117
timestamp 1586364061
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_129
timestamp 1586364061
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_141
timestamp 1586364061
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_128
timestamp 1586364061
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_154
timestamp 1586364061
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_166
timestamp 1586364061
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_178
timestamp 1586364061
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_190
timestamp 1586364061
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_129
timestamp 1586364061
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_202
timestamp 1586364061
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_215
timestamp 1586364061
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_227
timestamp 1586364061
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_239
timestamp 1586364061
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_251
timestamp 1586364061
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_263
timestamp 1586364061
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_130
timestamp 1586364061
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_276
timestamp 1586364061
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_288
timestamp 1586364061
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_300
timestamp 1586364061
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_312
timestamp 1586364061
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_131
timestamp 1586364061
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_12_324
timestamp 1586364061
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_337
timestamp 1586364061
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_349
timestamp 1586364061
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_361
timestamp 1586364061
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_373
timestamp 1586364061
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_12_385
timestamp 1586364061
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use scs8hd_decap_3  PHY_25
timestamp 1586364061
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_132
timestamp 1586364061
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_8  FILLER_12_398
timestamp 1586364061
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use scs8hd_fill_1  FILLER_12_406
timestamp 1586364061
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use scs8hd_decap_3  PHY_26
timestamp 1586364061
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_28
timestamp 1586364061
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_13_3
timestamp 1586364061
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_15
timestamp 1586364061
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_3
timestamp 1586364061
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_15
timestamp 1586364061
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_139
timestamp 1586364061
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_27
timestamp 1586364061
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_14_27
timestamp 1586364061
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use scs8hd_decap_12  FILLER_14_32
timestamp 1586364061
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_39
timestamp 1586364061
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_13_51
timestamp 1586364061
transform 1 0 5796 0 1 9248
box -38 -48 774 592
use scs8hd_decap_12  FILLER_14_44
timestamp 1586364061
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_133
timestamp 1586364061
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use scs8hd_fill_2  FILLER_13_59
timestamp 1586364061
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use scs8hd_decap_12  FILLER_13_62
timestamp 1586364061
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_56
timestamp 1586364061
transform 1 0 6256 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_68
timestamp 1586364061
transform 1 0 7360 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_74
timestamp 1586364061
transform 1 0 7912 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_86
timestamp 1586364061
transform 1 0 9016 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_80
timestamp 1586364061
transform 1 0 8464 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_140
timestamp 1586364061
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_98
timestamp 1586364061
transform 1 0 10120 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_93
timestamp 1586364061
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_105
timestamp 1586364061
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_134
timestamp 1586364061
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_110
timestamp 1586364061
transform 1 0 11224 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_123
timestamp 1586364061
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_117
timestamp 1586364061
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_135
timestamp 1586364061
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_129
timestamp 1586364061
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_141
timestamp 1586364061
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_141
timestamp 1586364061
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_147
timestamp 1586364061
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_159
timestamp 1586364061
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_154
timestamp 1586364061
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_171
timestamp 1586364061
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_166
timestamp 1586364061
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_178
timestamp 1586364061
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_135
timestamp 1586364061
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_184
timestamp 1586364061
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_196
timestamp 1586364061
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_190
timestamp 1586364061
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_142
timestamp 1586364061
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_208
timestamp 1586364061
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_202
timestamp 1586364061
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_220
timestamp 1586364061
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_215
timestamp 1586364061
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_227
timestamp 1586364061
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_136
timestamp 1586364061
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_232
timestamp 1586364061
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_245
timestamp 1586364061
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_239
timestamp 1586364061
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_257
timestamp 1586364061
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_251
timestamp 1586364061
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_263
timestamp 1586364061
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_143
timestamp 1586364061
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_269
timestamp 1586364061
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_281
timestamp 1586364061
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_276
timestamp 1586364061
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_293
timestamp 1586364061
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_288
timestamp 1586364061
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_300
timestamp 1586364061
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_137
timestamp 1586364061
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_306
timestamp 1586364061
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_318
timestamp 1586364061
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_312
timestamp 1586364061
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_144
timestamp 1586364061
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_330
timestamp 1586364061
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_324
timestamp 1586364061
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_337
timestamp 1586364061
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_342
timestamp 1586364061
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_354
timestamp 1586364061
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_349
timestamp 1586364061
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_138
timestamp 1586364061
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use scs8hd_decap_12  FILLER_13_367
timestamp 1586364061
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_361
timestamp 1586364061
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_373
timestamp 1586364061
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_379
timestamp 1586364061
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_13_391
timestamp 1586364061
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_14_385
timestamp 1586364061
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_27
timestamp 1586364061
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use scs8hd_decap_3  PHY_29
timestamp 1586364061
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_145
timestamp 1586364061
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_4  FILLER_13_403
timestamp 1586364061
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use scs8hd_decap_8  FILLER_14_398
timestamp 1586364061
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use scs8hd_fill_1  FILLER_14_406
timestamp 1586364061
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use scs8hd_decap_3  PHY_30
timestamp 1586364061
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use scs8hd_decap_12  FILLER_15_3
timestamp 1586364061
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_15
timestamp 1586364061
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_27
timestamp 1586364061
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_39
timestamp 1586364061
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_15_51
timestamp 1586364061
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_146
timestamp 1586364061
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use scs8hd_fill_2  FILLER_15_59
timestamp 1586364061
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use scs8hd_decap_12  FILLER_15_62
timestamp 1586364061
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_74
timestamp 1586364061
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_86
timestamp 1586364061
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_98
timestamp 1586364061
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_147
timestamp 1586364061
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_110
timestamp 1586364061
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_123
timestamp 1586364061
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_135
timestamp 1586364061
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_147
timestamp 1586364061
transform 1 0 14628 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_159
timestamp 1586364061
transform 1 0 15732 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_171
timestamp 1586364061
transform 1 0 16836 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_148
timestamp 1586364061
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_184
timestamp 1586364061
transform 1 0 18032 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_196
timestamp 1586364061
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_208
timestamp 1586364061
transform 1 0 20240 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_220
timestamp 1586364061
transform 1 0 21344 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_149
timestamp 1586364061
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_232
timestamp 1586364061
transform 1 0 22448 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_245
timestamp 1586364061
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_257
timestamp 1586364061
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_269
timestamp 1586364061
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_281
timestamp 1586364061
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_293
timestamp 1586364061
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_150
timestamp 1586364061
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_306
timestamp 1586364061
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_318
timestamp 1586364061
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_330
timestamp 1586364061
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_342
timestamp 1586364061
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_354
timestamp 1586364061
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_151
timestamp 1586364061
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use scs8hd_decap_12  FILLER_15_367
timestamp 1586364061
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_379
timestamp 1586364061
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_15_391
timestamp 1586364061
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use scs8hd_decap_3  PHY_31
timestamp 1586364061
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use scs8hd_decap_4  FILLER_15_403
timestamp 1586364061
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use scs8hd_decap_3  PHY_32
timestamp 1586364061
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_16_3
timestamp 1586364061
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_15
timestamp 1586364061
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_152
timestamp 1586364061
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_4  FILLER_16_27
timestamp 1586364061
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use scs8hd_decap_12  FILLER_16_32
timestamp 1586364061
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_44
timestamp 1586364061
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_56
timestamp 1586364061
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_68
timestamp 1586364061
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_80
timestamp 1586364061
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_153
timestamp 1586364061
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_93
timestamp 1586364061
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_105
timestamp 1586364061
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_117
timestamp 1586364061
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_129
timestamp 1586364061
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_141
timestamp 1586364061
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_154
timestamp 1586364061
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_154
timestamp 1586364061
transform 1 0 15272 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_166
timestamp 1586364061
transform 1 0 16376 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_178
timestamp 1586364061
transform 1 0 17480 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_190
timestamp 1586364061
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_155
timestamp 1586364061
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_202
timestamp 1586364061
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_215
timestamp 1586364061
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_227
timestamp 1586364061
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_239
timestamp 1586364061
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_251
timestamp 1586364061
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_263
timestamp 1586364061
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_156
timestamp 1586364061
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_276
timestamp 1586364061
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_288
timestamp 1586364061
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_300
timestamp 1586364061
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_312
timestamp 1586364061
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_157
timestamp 1586364061
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_16_324
timestamp 1586364061
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_337
timestamp 1586364061
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_349
timestamp 1586364061
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_361
timestamp 1586364061
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_373
timestamp 1586364061
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_16_385
timestamp 1586364061
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_33
timestamp 1586364061
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_158
timestamp 1586364061
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_8  FILLER_16_398
timestamp 1586364061
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use scs8hd_fill_1  FILLER_16_406
timestamp 1586364061
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use scs8hd_decap_3  PHY_34
timestamp 1586364061
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use scs8hd_decap_12  FILLER_17_3
timestamp 1586364061
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_15
timestamp 1586364061
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_27
timestamp 1586364061
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_39
timestamp 1586364061
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_17_51
timestamp 1586364061
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use scs8hd_tapvpwrvgnd_1  PHY_159
timestamp 1586364061
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use scs8hd_fill_2  FILLER_17_59
timestamp 1586364061
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use scs8hd_decap_12  FILLER_17_62
timestamp 1586364061
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_74
timestamp 1586364061
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_86
timestamp 1586364061
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_98
timestamp 1586364061
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_160
timestamp 1586364061
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_110
timestamp 1586364061
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_123
timestamp 1586364061
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_135
timestamp 1586364061
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_147
timestamp 1586364061
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_159
timestamp 1586364061
transform 1 0 15732 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_171
timestamp 1586364061
transform 1 0 16836 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_161
timestamp 1586364061
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_184
timestamp 1586364061
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_196
timestamp 1586364061
transform 1 0 19136 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_208
timestamp 1586364061
transform 1 0 20240 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_220
timestamp 1586364061
transform 1 0 21344 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_162
timestamp 1586364061
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_232
timestamp 1586364061
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_245
timestamp 1586364061
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_257
timestamp 1586364061
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_269
timestamp 1586364061
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_281
timestamp 1586364061
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_293
timestamp 1586364061
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_163
timestamp 1586364061
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_306
timestamp 1586364061
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_318
timestamp 1586364061
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_330
timestamp 1586364061
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_342
timestamp 1586364061
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_354
timestamp 1586364061
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_164
timestamp 1586364061
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use scs8hd_decap_12  FILLER_17_367
timestamp 1586364061
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_379
timestamp 1586364061
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_17_391
timestamp 1586364061
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use scs8hd_decap_3  PHY_35
timestamp 1586364061
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use scs8hd_decap_4  FILLER_17_403
timestamp 1586364061
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use scs8hd_decap_3  PHY_36
timestamp 1586364061
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use scs8hd_decap_12  FILLER_18_3
timestamp 1586364061
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_15
timestamp 1586364061
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_165
timestamp 1586364061
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_4  FILLER_18_27
timestamp 1586364061
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use scs8hd_decap_12  FILLER_18_32
timestamp 1586364061
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_44
timestamp 1586364061
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_56
timestamp 1586364061
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_68
timestamp 1586364061
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_80
timestamp 1586364061
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_166
timestamp 1586364061
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_93
timestamp 1586364061
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_105
timestamp 1586364061
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_117
timestamp 1586364061
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_129
timestamp 1586364061
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_141
timestamp 1586364061
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_167
timestamp 1586364061
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_154
timestamp 1586364061
transform 1 0 15272 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_166
timestamp 1586364061
transform 1 0 16376 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_178
timestamp 1586364061
transform 1 0 17480 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_190
timestamp 1586364061
transform 1 0 18584 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_168
timestamp 1586364061
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_202
timestamp 1586364061
transform 1 0 19688 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_215
timestamp 1586364061
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_227
timestamp 1586364061
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_239
timestamp 1586364061
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_251
timestamp 1586364061
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_263
timestamp 1586364061
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_169
timestamp 1586364061
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_276
timestamp 1586364061
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_288
timestamp 1586364061
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_300
timestamp 1586364061
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_312
timestamp 1586364061
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_170
timestamp 1586364061
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_12  FILLER_18_324
timestamp 1586364061
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_337
timestamp 1586364061
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_349
timestamp 1586364061
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_361
timestamp 1586364061
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_373
timestamp 1586364061
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_18_385
timestamp 1586364061
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use scs8hd_decap_3  PHY_37
timestamp 1586364061
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_171
timestamp 1586364061
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_8  FILLER_18_398
timestamp 1586364061
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use scs8hd_fill_1  FILLER_18_406
timestamp 1586364061
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use scs8hd_decap_3  PHY_38
timestamp 1586364061
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_40
timestamp 1586364061
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use scs8hd_decap_12  FILLER_19_3
timestamp 1586364061
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_15
timestamp 1586364061
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_3
timestamp 1586364061
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_15
timestamp 1586364061
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_178
timestamp 1586364061
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_27
timestamp 1586364061
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_4  FILLER_20_27
timestamp 1586364061
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use scs8hd_decap_12  FILLER_20_32
timestamp 1586364061
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_39
timestamp 1586364061
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_8  FILLER_19_51
timestamp 1586364061
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use scs8hd_decap_12  FILLER_20_44
timestamp 1586364061
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_172
timestamp 1586364061
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_179
timestamp 1586364061
transform 1 0 6808 0 -1 13600
box -38 -48 130 592
use scs8hd_fill_2  FILLER_19_59
timestamp 1586364061
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use scs8hd_decap_12  FILLER_19_62
timestamp 1586364061
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_56
timestamp 1586364061
transform 1 0 6256 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_63
timestamp 1586364061
transform 1 0 6900 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_74
timestamp 1586364061
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_86
timestamp 1586364061
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_75
timestamp 1586364061
transform 1 0 8004 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_87
timestamp 1586364061
transform 1 0 9108 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_180
timestamp 1586364061
transform 1 0 9660 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_98
timestamp 1586364061
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_94
timestamp 1586364061
transform 1 0 9752 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_106
timestamp 1586364061
transform 1 0 10856 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_173
timestamp 1586364061
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_181
timestamp 1586364061
transform 1 0 12512 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_110
timestamp 1586364061
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_123
timestamp 1586364061
transform 1 0 12420 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_118
timestamp 1586364061
transform 1 0 11960 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_19_135
timestamp 1586364061
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_125
timestamp 1586364061
transform 1 0 12604 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_137
timestamp 1586364061
transform 1 0 13708 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_182
timestamp 1586364061
transform 1 0 15364 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_147
timestamp 1586364061
transform 1 0 14628 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_159
timestamp 1586364061
transform 1 0 15732 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_149
timestamp 1586364061
transform 1 0 14812 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_156
timestamp 1586364061
transform 1 0 15456 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_171
timestamp 1586364061
transform 1 0 16836 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_168
timestamp 1586364061
transform 1 0 16560 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_174
timestamp 1586364061
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_183
timestamp 1586364061
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_184
timestamp 1586364061
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_196
timestamp 1586364061
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_180
timestamp 1586364061
transform 1 0 17664 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_187
timestamp 1586364061
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_208
timestamp 1586364061
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_199
timestamp 1586364061
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_211
timestamp 1586364061
transform 1 0 20516 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_184
timestamp 1586364061
transform 1 0 21068 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_220
timestamp 1586364061
transform 1 0 21344 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_218
timestamp 1586364061
transform 1 0 21160 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_230
timestamp 1586364061
transform 1 0 22264 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_175
timestamp 1586364061
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_185
timestamp 1586364061
transform 1 0 23920 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_232
timestamp 1586364061
transform 1 0 22448 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_245
timestamp 1586364061
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_242
timestamp 1586364061
transform 1 0 23368 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_249
timestamp 1586364061
transform 1 0 24012 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_257
timestamp 1586364061
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_261
timestamp 1586364061
transform 1 0 25116 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_186
timestamp 1586364061
transform 1 0 26772 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_269
timestamp 1586364061
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_281
timestamp 1586364061
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_273
timestamp 1586364061
transform 1 0 26220 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_280
timestamp 1586364061
transform 1 0 26864 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_293
timestamp 1586364061
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_292
timestamp 1586364061
transform 1 0 27968 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_176
timestamp 1586364061
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_187
timestamp 1586364061
transform 1 0 29624 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_306
timestamp 1586364061
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_318
timestamp 1586364061
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_304
timestamp 1586364061
transform 1 0 29072 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_311
timestamp 1586364061
transform 1 0 29716 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_330
timestamp 1586364061
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_323
timestamp 1586364061
transform 1 0 30820 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_335
timestamp 1586364061
transform 1 0 31924 0 -1 13600
box -38 -48 590 592
use scs8hd_tapvpwrvgnd_1  PHY_188
timestamp 1586364061
transform 1 0 32476 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_342
timestamp 1586364061
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_354
timestamp 1586364061
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_342
timestamp 1586364061
transform 1 0 32568 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_354
timestamp 1586364061
transform 1 0 33672 0 -1 13600
box -38 -48 1142 592
use scs8hd_tapvpwrvgnd_1  PHY_177
timestamp 1586364061
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use scs8hd_tapvpwrvgnd_1  PHY_189
timestamp 1586364061
transform 1 0 35328 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_12  FILLER_19_367
timestamp 1586364061
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_6  FILLER_20_366
timestamp 1586364061
transform 1 0 34776 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_12  FILLER_20_373
timestamp 1586364061
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_379
timestamp 1586364061
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_19_391
timestamp 1586364061
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use scs8hd_decap_12  FILLER_20_385
timestamp 1586364061
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use scs8hd_decap_3  PHY_39
timestamp 1586364061
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use scs8hd_decap_3  PHY_41
timestamp 1586364061
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use scs8hd_tapvpwrvgnd_1  PHY_190
timestamp 1586364061
transform 1 0 38180 0 -1 13600
box -38 -48 130 592
use scs8hd_decap_4  FILLER_19_403
timestamp 1586364061
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use scs8hd_decap_6  FILLER_20_397
timestamp 1586364061
transform 1 0 37628 0 -1 13600
box -38 -48 590 592
use scs8hd_decap_3  FILLER_20_404
timestamp 1586364061
transform 1 0 38272 0 -1 13600
box -38 -48 314 592
<< labels >>
rlabel metal2 s 27158 15200 27214 16000 6 address[0]
port 0 nsew default input
rlabel metal2 s 15198 15200 15254 16000 6 address[1]
port 1 nsew default input
rlabel metal2 s 16118 15200 16174 16000 6 address[2]
port 2 nsew default input
rlabel metal2 s 17038 15200 17094 16000 6 address[3]
port 3 nsew default input
rlabel metal2 s 17958 15200 18014 16000 6 address[4]
port 4 nsew default input
rlabel metal2 s 18878 15200 18934 16000 6 address[5]
port 5 nsew default input
rlabel metal2 s 18 0 74 800 6 bottom_grid_pin_0_
port 6 nsew default tristate
rlabel metal3 s 0 688 800 808 6 bottom_grid_pin_4_
port 7 nsew default tristate
rlabel metal2 s 938 0 994 800 6 bottom_grid_pin_8_
port 8 nsew default tristate
rlabel metal2 s 1858 0 1914 800 6 chanx_left_in[0]
port 9 nsew default input
rlabel metal3 s 0 2048 800 2168 6 chanx_left_in[1]
port 10 nsew default input
rlabel metal2 s 2778 0 2834 800 6 chanx_left_in[2]
port 11 nsew default input
rlabel metal3 s 0 3408 800 3528 6 chanx_left_in[3]
port 12 nsew default input
rlabel metal2 s 3698 0 3754 800 6 chanx_left_in[4]
port 13 nsew default input
rlabel metal2 s 4618 0 4674 800 6 chanx_left_in[5]
port 14 nsew default input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[6]
port 15 nsew default input
rlabel metal2 s 5538 0 5594 800 6 chanx_left_in[7]
port 16 nsew default input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[8]
port 17 nsew default input
rlabel metal2 s 6458 0 6514 800 6 chanx_left_out[0]
port 18 nsew default tristate
rlabel metal2 s 7378 0 7434 800 6 chanx_left_out[1]
port 19 nsew default tristate
rlabel metal3 s 0 7488 800 7608 6 chanx_left_out[2]
port 20 nsew default tristate
rlabel metal2 s 8298 0 8354 800 6 chanx_left_out[3]
port 21 nsew default tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_out[4]
port 22 nsew default tristate
rlabel metal2 s 9218 0 9274 800 6 chanx_left_out[5]
port 23 nsew default tristate
rlabel metal2 s 10138 0 10194 800 6 chanx_left_out[6]
port 24 nsew default tristate
rlabel metal3 s 0 10208 800 10328 6 chanx_left_out[7]
port 25 nsew default tristate
rlabel metal2 s 11058 0 11114 800 6 chanx_left_out[8]
port 26 nsew default tristate
rlabel metal2 s 39578 0 39634 800 6 chanx_right_in[0]
port 27 nsew default input
rlabel metal3 s 39200 688 40000 808 6 chanx_right_in[1]
port 28 nsew default input
rlabel metal2 s 38658 0 38714 800 6 chanx_right_in[2]
port 29 nsew default input
rlabel metal3 s 39200 2048 40000 2168 6 chanx_right_in[3]
port 30 nsew default input
rlabel metal2 s 37738 0 37794 800 6 chanx_right_in[4]
port 31 nsew default input
rlabel metal2 s 36818 0 36874 800 6 chanx_right_in[5]
port 32 nsew default input
rlabel metal3 s 39200 3408 40000 3528 6 chanx_right_in[6]
port 33 nsew default input
rlabel metal2 s 35898 0 35954 800 6 chanx_right_in[7]
port 34 nsew default input
rlabel metal3 s 39200 4768 40000 4888 6 chanx_right_in[8]
port 35 nsew default input
rlabel metal2 s 34978 0 35034 800 6 chanx_right_out[0]
port 36 nsew default tristate
rlabel metal2 s 34058 0 34114 800 6 chanx_right_out[1]
port 37 nsew default tristate
rlabel metal3 s 39200 6128 40000 6248 6 chanx_right_out[2]
port 38 nsew default tristate
rlabel metal2 s 33138 0 33194 800 6 chanx_right_out[3]
port 39 nsew default tristate
rlabel metal3 s 39200 7488 40000 7608 6 chanx_right_out[4]
port 40 nsew default tristate
rlabel metal2 s 32218 0 32274 800 6 chanx_right_out[5]
port 41 nsew default tristate
rlabel metal2 s 31298 0 31354 800 6 chanx_right_out[6]
port 42 nsew default tristate
rlabel metal3 s 39200 8848 40000 8968 6 chanx_right_out[7]
port 43 nsew default tristate
rlabel metal2 s 30378 0 30434 800 6 chanx_right_out[8]
port 44 nsew default tristate
rlabel metal2 s 19798 15200 19854 16000 6 data_in
port 45 nsew default input
rlabel metal3 s 39200 10208 40000 10328 6 enable
port 46 nsew default input
rlabel metal3 s 0 15648 800 15768 6 top_grid_pin_14_
port 47 nsew default tristate
rlabel metal2 s 478 15200 534 16000 6 top_grid_pin_2_
port 48 nsew default tristate
rlabel metal2 s 1398 15200 1454 16000 6 top_grid_pin_6_
port 49 nsew default tristate
rlabel metal4 s 7611 2128 7931 13648 6 vpwr
port 50 nsew default input
rlabel metal4 s 14277 2128 14597 13648 6 vgnd
port 51 nsew default input
<< properties >>
string FIXED_BBOX 0 0 40000 16000
<< end >>
