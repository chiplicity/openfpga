* NGSPICE file created from sb_1__1_.ext - technology: EFS8A

* Black-box entry subcircuit for scs8hd_fill_2 abstract view
.subckt scs8hd_fill_2 vpwr vgnd
.ends

* Black-box entry subcircuit for scs8hd_inv_1 abstract view
.subckt scs8hd_inv_1 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_diode_2 abstract view
.subckt scs8hd_diode_2 DIODE vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_lpflow_inputisolatch_1 abstract view
.subckt scs8hd_lpflow_inputisolatch_1 D Q SLEEPB vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_fill_1 abstract view
.subckt scs8hd_fill_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_ebufn_2 abstract view
.subckt scs8hd_ebufn_2 A TEB Z vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_buf_2 abstract view
.subckt scs8hd_buf_2 A X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nor2_4 abstract view
.subckt scs8hd_nor2_4 A B Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_3 abstract view
.subckt scs8hd_decap_3 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or4_4 abstract view
.subckt scs8hd_or4_4 A B C D X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_inv_8 abstract view
.subckt scs8hd_inv_8 A Y vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_4 abstract view
.subckt scs8hd_decap_4 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_12 abstract view
.subckt scs8hd_decap_12 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_8 abstract view
.subckt scs8hd_decap_8 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_tapvpwrvgnd_1 abstract view
.subckt scs8hd_tapvpwrvgnd_1 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or3_4 abstract view
.subckt scs8hd_or3_4 A B C X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_or2_4 abstract view
.subckt scs8hd_or2_4 A B X vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_conb_1 abstract view
.subckt scs8hd_conb_1 HI LO vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_decap_6 abstract view
.subckt scs8hd_decap_6 vgnd vpwr
.ends

* Black-box entry subcircuit for scs8hd_nand2_4 abstract view
.subckt scs8hd_nand2_4 A B Y vgnd vpwr
.ends

.subckt sb_1__1_ address[0] address[1] address[2] address[6] bottom_left_grid_pin_13_
+ bottom_right_grid_pin_11_ chanx_left_in[1] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7]
+ chanx_left_in[8] chanx_left_out[0] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_right_in[0] chanx_right_in[1] chanx_right_in[2] chanx_right_in[3] chanx_right_in[4]
+ chanx_right_in[6] chanx_right_in[7] chanx_right_in[8] chanx_right_out[0] chanx_right_out[1]
+ chanx_right_out[2] chanx_right_out[3] chanx_right_out[4] chanx_right_out[5] chanx_right_out[6]
+ chanx_right_out[7] chanx_right_out[8] vgnd chany_bottom_in[1] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_out[0]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_top_in[0] chany_top_in[1] chany_top_in[3] chany_top_in[4] chany_top_in[5]
+ chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_out[0] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] enable left_bottom_grid_pin_12_ left_top_grid_pin_10_
+ right_bottom_grid_pin_12_ right_top_grid_pin_10_ top_left_grid_pin_13_ top_right_grid_pin_11_
+ vgnd
XFILLER_22_166 vgnd vgnd scs8hd_fill_2
XFILLER_22_100 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[4] mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_26_41 vgnd vgnd scs8hd_fill_2
XFILLER_13_155 vgnd vgnd scs8hd_fill_2
XANTENNA__113__B _045_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_0_.scs8hd_inv_1 top_right_grid_pin_11_ mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmem_left_track_1.LATCH_6_.latch vgnd mem_left_track_1.LATCH_6_.latch/Q _116_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_27_214 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_10_147 vgnd vgnd scs8hd_fill_2
XFILLER_10_158 vgnd vgnd scs8hd_fill_2
XFILLER_12_32 vgnd vgnd scs8hd_fill_2
XFILLER_12_54 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_SLEEPB _138_/Y vgnd vgnd scs8hd_diode_2
XFILLER_12_87 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__108__B _110_/B vgnd vgnd scs8hd_diode_2
XANTENNA__124__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB chany_bottom_in[1]
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _161_/HI mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_4_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_23_20 vgnd vgnd scs8hd_fill_2
X_200_ chany_bottom_in[6] chany_top_out[7] vgnd vgnd scs8hd_buf_2
XFILLER_15_217 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_right_track_16.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
X_062_ _056_/B vgnd _062_/Y vgnd vgnd scs8hd_nor2_4
X_131_ vgnd _124_/B _131_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_23_53 vgnd vgnd scs8hd_decap_3
XFILLER_2_198 vgnd vgnd scs8hd_fill_2
XFILLER_2_154 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__119__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_9_77 vgnd vgnd scs8hd_fill_2
XFILLER_9_99 vgnd vgnd scs8hd_fill_2
Xmem_bottom_track_17.LATCH_2_.latch vgnd mem_bottom_track_17.LATCH_2_.latch/Q _150_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ _194_/A vgnd vgnd scs8hd_inv_1
XFILLER_12_209 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_18_64 vgnd vgnd scs8hd_fill_2
XFILLER_18_97 vgnd vgnd scs8hd_fill_1
XFILLER_34_63 vgnd vgnd scs8hd_fill_2
X_114_ vgnd vgnd vgnd chanx_right_in[2] _114_/X vgnd vgnd scs8hd_or4_4
X_045_ address[6] _045_/Y vgnd vgnd scs8hd_inv_8
XANTENNA_mem_top_track_0.LATCH_2_.latch_SLEEPB _062_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__121__B _114_/X vgnd vgnd scs8hd_diode_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ chany_bottom_in[1] vgnd vgnd vgnd scs8hd_ebufn_2
Xmux_bottom_track_9.INVTX1_6_.scs8hd_inv_1 vgnd mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[1] mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ mem_top_track_0.LATCH_5_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_205 vgnd vgnd scs8hd_fill_2
XFILLER_20_32 vgnd vgnd scs8hd_fill_1
XFILLER_29_96 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_20_87 vgnd vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[7] mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__116__B _114_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA__132__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_19_150 vgnd vgnd scs8hd_decap_4
XFILLER_34_197 vgnd vgnd scs8hd_decap_12
XFILLER_34_142 vgnd vgnd scs8hd_decap_8
Xmem_right_track_8.LATCH_1_.latch vgnd mem_right_track_8.LATCH_1_.latch/Q _093_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__042__A address[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_25_153 vgnd vgnd scs8hd_fill_1
XFILLER_25_197 vgnd vgnd scs8hd_fill_2
XFILLER_15_98 vgnd vgnd scs8hd_fill_2
XFILLER_0_230 vgnd vgnd scs8hd_decap_3
XFILLER_31_112 vgnd vgnd scs8hd_fill_2
XPHY_170 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA__127__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_16_120 vgnd vgnd scs8hd_fill_2
XFILLER_16_186 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_4_.latch_SLEEPB _127_/Y vgnd vgnd scs8hd_diode_2
XPHY_192 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_181 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA_mem_top_track_8.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _161_/HI vgnd
+ vgnd scs8hd_diode_2
XFILLER_22_145 vgnd vgnd scs8hd_fill_2
XFILLER_22_134 vgnd vgnd scs8hd_decap_4
XFILLER_13_123 vgnd vgnd scs8hd_decap_3
XFILLER_9_138 vgnd vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_6_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
Xmux_top_track_0.INVTX1_3_.scs8hd_inv_1 chanx_right_in[7] mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_27_226 vgnd vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_10_104 vgnd vgnd scs8hd_fill_2
XFILLER_10_115 vgnd vgnd scs8hd_fill_2
XFILLER_10_126 vgnd vgnd scs8hd_fill_2
XFILLER_12_22 vgnd vgnd scs8hd_fill_2
XFILLER_33_218 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_204 vgnd vgnd scs8hd_fill_2
XANTENNA__124__B _124_/B vgnd vgnd scs8hd_diode_2
XFILLER_5_174 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__140__A _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.INVTX1_0_.scs8hd_inv_1_A top_left_grid_pin_13_ vgnd vgnd
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_4_.scs8hd_inv_1 vgnd mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_right_track_8.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA__050__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmem_top_track_8.LATCH_6_.latch vgnd mem_top_track_8.LATCH_6_.latch/Q _069_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.INVTX1_0_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
Xmem_right_track_0.LATCH_6_.latch vgnd mem_right_track_0.LATCH_6_.latch/Q _078_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _171_/HI mem_top_track_8.LATCH_7_.latch/Q
+ mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
X_130_ vgnd _124_/B _130_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_23_43 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_061_ address[2] _043_/Y address[0] vgnd vgnd vgnd scs8hd_or3_4
XFILLER_23_76 vgnd vgnd scs8hd_fill_2
XFILLER_2_100 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ chany_bottom_in[1] mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__119__B _114_/X vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
XFILLER_9_56 vgnd vgnd scs8hd_fill_2
XANTENNA__135__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_20_232 vgnd vgnd scs8hd_fill_1
XFILLER_20_210 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_SLEEPB _097_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__045__A address[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_54 vgnd vgnd scs8hd_fill_1
XFILLER_7_214 vgnd vgnd scs8hd_fill_1
XFILLER_7_225 vgnd vgnd scs8hd_fill_2
X_113_ vgnd _045_/Y chanx_right_in[2] vgnd vgnd scs8hd_or2_4
XFILLER_11_210 vgnd vgnd scs8hd_decap_4
XFILLER_11_221 vgnd vgnd scs8hd_fill_2
X_044_ address[0] _063_/C vgnd vgnd scs8hd_inv_8
XANTENNA_mem_left_track_1.LATCH_0_.latch_SLEEPB _122_/Y vgnd vgnd scs8hd_diode_2
XFILLER_15_7 vgnd vgnd scs8hd_fill_2
Xmux_left_track_1.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[6] mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1_A bottom_right_grid_pin_11_ vgnd
+ vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_4_228 vgnd vgnd scs8hd_fill_2
XFILLER_20_55 vgnd vgnd scs8hd_fill_2
XFILLER_20_66 vgnd vgnd scs8hd_decap_3
XFILLER_29_75 vgnd vgnd scs8hd_fill_2
XFILLER_29_53 vgnd vgnd scs8hd_fill_2
XFILLER_28_140 vgnd vgnd scs8hd_fill_2
XANTENNA__132__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_SLEEPB _145_/Y vgnd vgnd scs8hd_diode_2
XFILLER_19_173 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd scs8hd_diode_2
XFILLER_25_132 vgnd vgnd scs8hd_fill_2
XFILLER_25_110 vgnd vgnd scs8hd_fill_2
XFILLER_15_11 vgnd vgnd scs8hd_fill_2
XFILLER_15_22 vgnd vgnd scs8hd_fill_2
XFILLER_15_55 vgnd vgnd scs8hd_fill_2
XFILLER_31_87 vgnd vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XPHY_193 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_left_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XPHY_182 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_171 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_160 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA__127__B _124_/B vgnd vgnd scs8hd_diode_2
XFILLER_16_154 vgnd vgnd scs8hd_fill_2
XFILLER_16_198 vgnd vgnd scs8hd_decap_3
Xmux_right_track_16.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__143__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_22_179 vgnd vgnd scs8hd_decap_4
XANTENNA__053__A _055_/A vgnd vgnd scs8hd_diode_2
XFILLER_7_9 vgnd vgnd scs8hd_fill_2
XFILLER_26_32 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_13_102 vgnd vgnd scs8hd_fill_2
XFILLER_13_113 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_5_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ _190_/A vgnd vgnd scs8hd_inv_1
XANTENNA__138__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_8_161 vgnd vgnd scs8hd_decap_4
Xmem_left_track_9.LATCH_7_.latch vgnd mem_left_track_9.LATCH_7_.latch/Q _124_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_8_183 vgnd vgnd scs8hd_decap_3
XANTENNA__048__A enable vgnd vgnd scs8hd_diode_2
XFILLER_12_67 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_33_208 vgnd vgnd scs8hd_decap_4
XFILLER_5_164 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__140__B _141_/B vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.INVTX1_7_.scs8hd_inv_1 vgnd mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_4_90 vgnd vgnd scs8hd_fill_2
XANTENNA__050__B address[6] vgnd vgnd scs8hd_diode_2
XFILLER_15_208 vgnd vgnd scs8hd_decap_3
XFILLER_23_11 vgnd vgnd scs8hd_fill_2
X_060_ _056_/B chanx_right_in[2] _060_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_3_3 vgnd vgnd scs8hd_fill_1
XFILLER_2_123 vgnd vgnd scs8hd_fill_2
XFILLER_2_112 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_2_167 vgnd vgnd scs8hd_fill_2
XANTENNA__135__B vgnd vgnd vgnd scs8hd_diode_2
X_189_ _189_/A chanx_right_out[0] vgnd vgnd scs8hd_buf_2
XANTENNA__151__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__061__A address[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vgnd scs8hd_diode_2
XFILLER_18_11 vgnd vgnd scs8hd_fill_2
XFILLER_18_22 vgnd vgnd scs8hd_fill_2
XFILLER_34_32 vgnd vgnd scs8hd_decap_3
XFILLER_34_21 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_88 vgnd vgnd scs8hd_fill_2
X_043_ address[1] _043_/Y vgnd vgnd scs8hd_inv_8
X_112_ vgnd _110_/B _112_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA__146__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_29_108 vgnd vgnd scs8hd_fill_2
XANTENNA__056__A _056_/B vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_6_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_29_32 vgnd vgnd scs8hd_fill_2
XFILLER_28_163 vgnd vgnd scs8hd_fill_2
XFILLER_28_152 vgnd vgnd scs8hd_fill_1
XANTENNA__132__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_19_130 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_25_177 vgnd vgnd scs8hd_decap_4
XFILLER_25_166 vgnd vgnd scs8hd_decap_4
XFILLER_31_66 vgnd vgnd scs8hd_fill_2
XFILLER_31_44 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _160_/HI vgnd vgnd
+ scs8hd_diode_2
XFILLER_16_133 vgnd vgnd scs8hd_fill_2
XFILLER_16_144 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XPHY_194 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_31_136 vgnd vgnd scs8hd_fill_2
XPHY_183 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_172 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_161 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_150 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA_mem_right_track_8.LATCH_5_.latch_SLEEPB _089_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__143__B _141_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__053__B _043_/Y vgnd vgnd scs8hd_diode_2
XFILLER_30_191 vgnd vgnd scs8hd_fill_2
XFILLER_30_180 vgnd vgnd scs8hd_decap_4
XFILLER_26_11 vgnd vgnd scs8hd_fill_2
XFILLER_26_88 vgnd vgnd scs8hd_fill_2
XFILLER_9_118 vgnd vgnd scs8hd_fill_2
XFILLER_13_136 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vgnd scs8hd_diode_2
XFILLER_3_59 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[8] mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__138__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__154__A _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_27_217 vgnd vgnd scs8hd_fill_1
XANTENNA__064__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_12_79 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_18_228 vgnd vgnd scs8hd_fill_2
XFILLER_5_187 vgnd vgnd scs8hd_fill_2
XFILLER_5_143 vgnd vgnd scs8hd_fill_2
XFILLER_5_132 vgnd vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_0_.latch vgnd mem_top_track_0.LATCH_0_.latch/Q _066_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__149__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_24_209 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_32_231 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 vgnd mem_bottom_track_17.LATCH_3_.latch/Q
+ mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
Xmem_right_track_8.LATCH_7_.latch vgnd mem_right_track_8.LATCH_7_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__059__A address[2] vgnd vgnd scs8hd_diode_2
XFILLER_2_146 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[7] vgnd vgnd scs8hd_diode_2
XFILLER_9_36 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmem_left_track_17.LATCH_3_.latch vgnd mem_left_track_17.LATCH_3_.latch/Q _156_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
X_188_ vgnd chanx_right_out[1] vgnd vgnd scs8hd_buf_2
XANTENNA__151__B _152_/B vgnd vgnd scs8hd_diode_2
XFILLER_20_201 vgnd vgnd scs8hd_fill_1
XANTENNA__061__B _043_/Y vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y vgnd vgnd scs8hd_ebufn_2
XFILLER_34_88 vgnd vgnd scs8hd_fill_2
X_111_ vgnd _110_/B _111_/Y vgnd vgnd scs8hd_nor2_4
X_042_ address[2] _055_/A vgnd vgnd scs8hd_inv_8
XANTENNA_mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[0] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_SLEEPB _083_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__146__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__056__B _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA__072__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_20_24 vgnd vgnd scs8hd_fill_2
XFILLER_29_88 vgnd vgnd scs8hd_fill_2
XFILLER_28_197 vgnd vgnd scs8hd_fill_2
XFILLER_28_186 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_6_26 vgnd vgnd scs8hd_fill_2
XANTENNA__132__D _067_/D vgnd vgnd scs8hd_diode_2
XFILLER_10_90 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_7 vgnd vgnd scs8hd_fill_2
XFILLER_34_123 vgnd vgnd scs8hd_fill_2
XANTENNA__157__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_19_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_1.LATCH_2_.latch vgnd mem_bottom_track_1.LATCH_2_.latch/Q _101_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_SLEEPB _072_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__067__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_25_156 vgnd vgnd scs8hd_fill_1
XFILLER_15_79 vgnd vgnd scs8hd_fill_2
XFILLER_31_56 vgnd vgnd scs8hd_fill_2
XFILLER_31_23 vgnd vgnd scs8hd_fill_2
XFILLER_31_12 vgnd vgnd scs8hd_fill_2
XFILLER_0_222 vgnd vgnd scs8hd_fill_2
XFILLER_0_200 vgnd vgnd scs8hd_fill_2
XFILLER_31_104 vgnd vgnd scs8hd_fill_2
XFILLER_16_101 vgnd vgnd scs8hd_fill_2
XPHY_195 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_184 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_173 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_162 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_151 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_140 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_22_115 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__053__C address[0] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_left_track_1.LATCH_1_.latch vgnd mem_left_track_1.LATCH_1_.latch/Q _121_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_26_67 vgnd vgnd scs8hd_fill_2
XFILLER_26_56 vgnd vgnd scs8hd_fill_2
XFILLER_26_23 vgnd vgnd scs8hd_decap_4
XFILLER_13_159 vgnd vgnd scs8hd_fill_2
XANTENNA__154__B _159_/B vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_12_181 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__064__B vgnd vgnd vgnd scs8hd_diode_2
Xmem_right_track_16.LATCH_2_.latch vgnd chany_bottom_in[1] _143_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_12_36 vgnd vgnd scs8hd_decap_3
XANTENNA__080__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__149__B _152_/B vgnd vgnd scs8hd_diode_2
XANTENNA__059__B _043_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_23_221 vgnd vgnd scs8hd_fill_2
XFILLER_23_210 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__075__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_24 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_2_158 vgnd vgnd scs8hd_fill_2
XFILLER_9_48 vgnd vgnd scs8hd_fill_2
XFILLER_14_232 vgnd vgnd scs8hd_fill_1
X_187_ chanx_left_in[1] chanx_right_out[2] vgnd vgnd scs8hd_buf_2
XFILLER_20_224 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_3_.scs8hd_inv_1 chanx_right_in[3] mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_9.INVTX1_0_.scs8hd_inv_1 vgnd mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__061__C address[0] vgnd vgnd scs8hd_diode_2
XFILLER_18_46 vgnd vgnd scs8hd_fill_2
XFILLER_18_68 vgnd vgnd scs8hd_fill_2
XFILLER_34_67 vgnd vgnd scs8hd_fill_2
X_110_ vgnd _110_/B vgnd vgnd vgnd scs8hd_nor2_4
XFILLER_7_217 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__146__C vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] vgnd vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__072__B _067_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_209 vgnd vgnd scs8hd_fill_2
XFILLER_20_36 vgnd vgnd scs8hd_decap_4
XFILLER_29_12 vgnd vgnd scs8hd_decap_4
XFILLER_28_110 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_7_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XFILLER_34_102 vgnd vgnd scs8hd_fill_2
XANTENNA__157__B _159_/B vgnd vgnd scs8hd_diode_2
XANTENNA__173__A chanx_right_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_SLEEPB _130_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__067__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__083__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_15_36 vgnd vgnd scs8hd_fill_2
XFILLER_0_212 vgnd vgnd scs8hd_fill_2
XFILLER_31_149 vgnd vgnd scs8hd_fill_2
XFILLER_31_116 vgnd vgnd scs8hd_decap_4
XPHY_152 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XPHY_130 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_141 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_196 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_185 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_174 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_163 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA_mem_left_track_17.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_22_149 vgnd vgnd scs8hd_fill_2
XFILLER_22_138 vgnd vgnd scs8hd_fill_1
Xmux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.INVTX1_0_.scs8hd_inv_1 top_left_grid_pin_13_ mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__078__A _053_/X vgnd vgnd scs8hd_diode_2
XFILLER_21_193 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_8_131 vgnd vgnd scs8hd_fill_2
XFILLER_8_197 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_10_119 vgnd vgnd scs8hd_fill_2
XFILLER_12_26 vgnd vgnd scs8hd_fill_2
XANTENNA__080__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_18_208 vgnd vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_1_.latch vgnd mem_right_track_0.LATCH_1_.latch/Q _083_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmem_top_track_8.LATCH_1_.latch vgnd mem_top_track_8.LATCH_1_.latch/Q _074_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_5_178 vgnd vgnd scs8hd_decap_3
XFILLER_5_156 vgnd vgnd scs8hd_fill_2
XFILLER_5_123 vgnd vgnd scs8hd_fill_2
XFILLER_5_101 vgnd vgnd scs8hd_fill_2
XFILLER_32_211 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_17_230 vgnd vgnd scs8hd_decap_3
XANTENNA__181__A _181_/A vgnd vgnd scs8hd_diode_2
XANTENNA__059__C _063_/C vgnd vgnd scs8hd_diode_2
XANTENNA__075__B _067_/X vgnd vgnd scs8hd_diode_2
XANTENNA__091__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_23_58 vgnd vgnd scs8hd_decap_3
XFILLER_23_47 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_SLEEPB _100_/Y vgnd vgnd scs8hd_diode_2
XFILLER_0_29 vgnd vgnd scs8hd_fill_2
XFILLER_14_200 vgnd vgnd scs8hd_fill_2
XFILLER_9_16 vgnd vgnd scs8hd_fill_2
XFILLER_13_91 vgnd vgnd scs8hd_fill_2
X_186_ vgnd chanx_right_out[3] vgnd vgnd scs8hd_buf_2
XANTENNA__176__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_6_.scs8hd_inv_1 chanx_left_in[1] vgnd vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.INVTX1_3_.scs8hd_inv_1 chanx_right_in[0] mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_34_13 vgnd vgnd scs8hd_fill_2
XANTENNA__086__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_34_46 vgnd vgnd scs8hd_fill_2
XFILLER_7_229 vgnd vgnd scs8hd_fill_2
XFILLER_11_214 vgnd vgnd scs8hd_fill_1
XFILLER_11_225 vgnd vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_5_.scs8hd_inv_1 vgnd mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_169_ _169_/HI _169_/LO vgnd vgnd scs8hd_conb_1
XANTENNA__146__D chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_34_3 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_right_track_8.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_59 vgnd vgnd scs8hd_fill_2
XFILLER_29_57 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_28_144 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_3_221 vgnd vgnd scs8hd_fill_2
XFILLER_3_210 vgnd vgnd scs8hd_decap_4
Xmux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_34_136 vgnd vgnd scs8hd_decap_4
Xmem_top_track_0.LATCH_6_.latch vgnd mem_top_track_0.LATCH_6_.latch/Q _054_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_3_.latch vgnd mem_bottom_track_9.LATCH_3_.latch/Q _109_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__067__C vgnd vgnd vgnd scs8hd_diode_2
XFILLER_25_136 vgnd vgnd scs8hd_fill_2
XFILLER_25_114 vgnd vgnd scs8hd_fill_2
XFILLER_25_103 vgnd vgnd scs8hd_fill_2
XFILLER_15_26 vgnd vgnd scs8hd_fill_2
XANTENNA__083__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_15_59 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XPHY_175 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_164 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_24_180 vgnd vgnd scs8hd_decap_4
XPHY_153 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_120 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_131 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_16_158 vgnd vgnd scs8hd_fill_1
XPHY_142 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_197 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_186 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_91 vgnd vgnd scs8hd_fill_2
XFILLER_21_80 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_4_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XPHY_0 vgnd vgnd scs8hd_decap_3
XANTENNA__184__A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_15_180 vgnd vgnd scs8hd_decap_3
Xmem_left_track_9.LATCH_2_.latch vgnd mem_left_track_9.LATCH_2_.latch/Q _129_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA__078__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__094__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_13_106 vgnd vgnd scs8hd_fill_2
XFILLER_13_117 vgnd vgnd scs8hd_fill_2
XFILLER_13_128 vgnd vgnd scs8hd_fill_2
XFILLER_21_161 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_top_track_0.LATCH_7_.latch_SLEEPB _052_/Y vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.INVTX1_8_.scs8hd_inv_1 left_bottom_grid_pin_12_ mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_8_110 vgnd vgnd scs8hd_fill_2
XFILLER_12_150 vgnd vgnd scs8hd_decap_3
XFILLER_12_161 vgnd vgnd scs8hd_fill_2
XFILLER_12_194 vgnd vgnd scs8hd_fill_2
XANTENNA__179__A chanx_right_in[0] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_SLEEPB _148_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__089__A _056_/B vgnd vgnd scs8hd_diode_2
Xmem_top_track_16.LATCH_3_.latch vgnd mem_top_track_16.LATCH_3_.latch/Q _135_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_5_168 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_left_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_23_15 vgnd vgnd scs8hd_fill_2
XANTENNA__091__B _086_/X vgnd vgnd scs8hd_diode_2
XFILLER_2_127 vgnd vgnd scs8hd_fill_2
XFILLER_2_116 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_14_212 vgnd vgnd scs8hd_fill_2
X_185_ vgnd chanx_right_out[4] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_left_track_9.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vgnd scs8hd_diode_2
XFILLER_1_160 vgnd vgnd scs8hd_fill_2
XFILLER_1_193 vgnd vgnd scs8hd_fill_2
XANTENNA__192__A chany_top_in[5] vgnd vgnd scs8hd_diode_2
XFILLER_18_26 vgnd vgnd scs8hd_fill_2
XANTENNA__086__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_34_25 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_top_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vgnd scs8hd_diode_2
Xmem_left_track_1.LATCH_7_.latch vgnd mem_left_track_1.LATCH_7_.latch/Q _115_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_top_track_0.INVTX1_8_.scs8hd_inv_1 chany_bottom_in[1] vgnd vgnd vgnd scs8hd_inv_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_168_ _168_/HI _168_/LO vgnd vgnd scs8hd_conb_1
XFILLER_24_91 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_left_track_9.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
X_099_ vgnd vgnd _099_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA__187__A chanx_left_in[1] vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_6_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_29_36 vgnd vgnd scs8hd_fill_2
XFILLER_28_123 vgnd vgnd scs8hd_fill_2
XANTENNA__097__A _053_/X vgnd vgnd scs8hd_diode_2
XFILLER_28_167 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_10_71 vgnd vgnd scs8hd_fill_2
XFILLER_10_82 vgnd vgnd scs8hd_fill_2
XFILLER_19_156 vgnd vgnd scs8hd_fill_2
XFILLER_19_134 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_right_track_8.LATCH_2_.latch_SLEEPB _092_/Y vgnd vgnd scs8hd_diode_2
XFILLER_33_170 vgnd vgnd scs8hd_fill_1
XANTENNA__067__D _067_/D vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_17.LATCH_3_.latch vgnd mem_bottom_track_17.LATCH_3_.latch/Q _149_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_16_137 vgnd vgnd scs8hd_fill_2
XFILLER_16_148 vgnd vgnd scs8hd_fill_2
XPHY_198 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_187 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_176 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_165 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_154 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_110 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_121 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_132 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_143 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_1 vgnd vgnd scs8hd_decap_3
XFILLER_30_195 vgnd vgnd scs8hd_decap_4
XFILLER_7_83 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_26_37 vgnd vgnd scs8hd_fill_2
XFILLER_26_15 vgnd vgnd scs8hd_fill_2
XANTENNA__094__B _086_/X vgnd vgnd scs8hd_diode_2
XFILLER_21_173 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_SLEEPB _117_/Y vgnd vgnd scs8hd_diode_2
XFILLER_35_221 vgnd vgnd scs8hd_fill_2
XANTENNA__195__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_left_track_1.LATCH_5_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA__089__B _086_/X vgnd vgnd scs8hd_diode_2
XFILLER_26_232 vgnd vgnd scs8hd_fill_1
Xmem_right_track_8.LATCH_2_.latch vgnd mem_right_track_8.LATCH_2_.latch/Q _092_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_5_114 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_SLEEPB _140_/Y vgnd vgnd scs8hd_diode_2
XFILLER_17_210 vgnd vgnd scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_2_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_17.INVTX1_6_.scs8hd_inv_1 vgnd mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_14_224 vgnd vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[8] mux_right_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_184_ chany_bottom_in[1] chanx_right_out[5] vgnd vgnd scs8hd_buf_2
Xmux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_right_track_16.LATCH_5_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_13_71 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 vgnd mem_top_track_0.LATCH_6_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
Xmux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__086__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
X_098_ _056_/B vgnd vgnd vgnd vgnd scs8hd_nor2_4
X_167_ _167_/HI _167_/LO vgnd vgnd scs8hd_conb_1
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_20_28 vgnd vgnd scs8hd_decap_3
XANTENNA__097__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_0_.latch_SLEEPB _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A _067_/X vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_SLEEPB _156_/Y vgnd vgnd scs8hd_diode_2
XFILLER_10_50 vgnd vgnd scs8hd_fill_2
Xmem_right_track_0.LATCH_7_.latch vgnd mem_right_track_0.LATCH_7_.latch/Q _077_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_19_102 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_17.tap_buf4_0_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_19_179 vgnd vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_7_.latch vgnd mem_top_track_8.LATCH_7_.latch/Q _068_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_19_81 vgnd vgnd scs8hd_fill_2
XFILLER_35_80 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__198__A _198_/A vgnd vgnd scs8hd_diode_2
XFILLER_33_193 vgnd vgnd scs8hd_fill_2
XFILLER_25_149 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB chany_bottom_in[1]
+ vgnd vgnd scs8hd_diode_2
XFILLER_31_27 vgnd vgnd scs8hd_fill_2
XFILLER_31_16 vgnd vgnd scs8hd_fill_2
XFILLER_0_226 vgnd vgnd scs8hd_fill_2
XPHY_100 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_16_105 vgnd vgnd scs8hd_fill_2
XFILLER_16_116 vgnd vgnd scs8hd_fill_2
XPHY_199 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_188 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_177 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_166 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_155 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_144 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _170_/HI mem_top_track_16.LATCH_2_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XPHY_111 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_122 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_133 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _165_/HI mem_left_track_9.LATCH_7_.latch/Q
+ mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XFILLER_22_119 vgnd vgnd scs8hd_fill_2
XPHY_2 vgnd vgnd scs8hd_decap_3
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_15_193 vgnd vgnd scs8hd_fill_2
XFILLER_30_163 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_5_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 vgnd vgnd mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_16_60 vgnd vgnd scs8hd_fill_2
XFILLER_32_70 vgnd vgnd scs8hd_fill_1
XFILLER_8_145 vgnd vgnd scs8hd_fill_2
XFILLER_8_178 vgnd vgnd scs8hd_decap_3
XFILLER_35_211 vgnd vgnd scs8hd_decap_6
XFILLER_35_200 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_12_18 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.tap_buf4_0_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_17_222 vgnd vgnd scs8hd_fill_2
XFILLER_32_203 vgnd vgnd scs8hd_decap_8
XFILLER_27_92 vgnd vgnd scs8hd_decap_4
Xmux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.tap_buf4_0_.scs8hd_inv_1 mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _180_/A vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_8.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[8] vgnd vgnd scs8hd_diode_2
XFILLER_23_225 vgnd vgnd scs8hd_fill_2
XFILLER_23_214 vgnd vgnd scs8hd_fill_1
XFILLER_23_39 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A _124_/Y vgnd vgnd
+ scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_183_ chanx_left_in[5] chanx_right_out[6] vgnd vgnd scs8hd_buf_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_228 vgnd vgnd scs8hd_fill_2
XFILLER_20_206 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA__086__D _086_/D vgnd vgnd scs8hd_diode_2
XFILLER_11_217 vgnd vgnd scs8hd_fill_1
Xmux_top_track_16.INVTX1_1_.scs8hd_inv_1 chanx_right_in[3] mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_097_ _053_/X vgnd _097_/Y vgnd vgnd scs8hd_nor2_4
X_166_ _166_/HI _166_/LO vgnd vgnd scs8hd_conb_1
XFILLER_6_232 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_left_track_17.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_SLEEPB _110_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[8] vgnd vgnd scs8hd_diode_2
XFILLER_29_49 vgnd vgnd scs8hd_fill_2
XFILLER_29_16 vgnd vgnd scs8hd_fill_1
XFILLER_19_114 vgnd vgnd scs8hd_fill_2
XFILLER_34_106 vgnd vgnd scs8hd_fill_2
XFILLER_19_169 vgnd vgnd scs8hd_fill_2
X_149_ chanx_right_in[2] _152_/B _149_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_180 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_0_216 vgnd vgnd scs8hd_fill_1
XFILLER_24_150 vgnd vgnd scs8hd_fill_1
XPHY_101 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_112 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_123 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_134 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_189 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_178 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_167 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_156 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_145 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XPHY_3 vgnd vgnd scs8hd_decap_3
XFILLER_15_161 vgnd vgnd scs8hd_fill_1
XFILLER_30_186 vgnd vgnd scs8hd_fill_2
XFILLER_7_96 vgnd vgnd scs8hd_fill_2
XFILLER_21_197 vgnd vgnd scs8hd_fill_2
XFILLER_21_153 vgnd vgnd scs8hd_fill_2
XFILLER_21_142 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_6_.latch_SLEEPB _078_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_8_102 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_16_72 vgnd vgnd scs8hd_fill_1
XFILLER_8_135 vgnd vgnd scs8hd_fill_1
XFILLER_8_157 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_26_201 vgnd vgnd scs8hd_decap_12
XFILLER_5_105 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XFILLER_27_71 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_SLEEPB _103_/Y vgnd vgnd scs8hd_diode_2
XFILLER_4_86 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_3_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_14_204 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_3_.scs8hd_inv_1 vgnd mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_182_ chanx_left_in[6] chanx_right_out[7] vgnd vgnd scs8hd_buf_2
Xmux_left_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mem_left_track_1.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_13_95 vgnd vgnd scs8hd_fill_2
XFILLER_1_130 vgnd vgnd scs8hd_fill_2
XANTENNA__100__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_2_.scs8hd_inv_1 chanx_right_in[6] mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_18_18 vgnd vgnd scs8hd_fill_2
XFILLER_34_17 vgnd vgnd scs8hd_fill_2
XFILLER_11_229 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _160_/HI mem_bottom_track_1.LATCH_7_.latch/Q
+ mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
X_165_ _165_/HI _165_/LO vgnd vgnd scs8hd_conb_1
XFILLER_24_83 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_SLEEPB _136_/Y vgnd vgnd scs8hd_diode_2
X_096_ vgnd vgnd vgnd vgnd vgnd scs8hd_nor2_4
Xmem_top_track_0.LATCH_1_.latch vgnd vgnd vgnd vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_28_148 vgnd vgnd scs8hd_fill_2
XFILLER_3_225 vgnd vgnd scs8hd_fill_2
XFILLER_3_214 vgnd vgnd scs8hd_fill_1
XFILLER_10_96 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.INVTX1_0_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_19_94 vgnd vgnd scs8hd_fill_2
XFILLER_19_126 vgnd vgnd scs8hd_fill_2
XFILLER_27_170 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_148_ vgnd _152_/B _148_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_079_ _056_/B vgnd _079_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_25_118 vgnd vgnd scs8hd_fill_2
XFILLER_33_173 vgnd vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_4_.latch vgnd mem_left_track_17.LATCH_4_.latch/Q _155_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XPHY_157 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_102 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_113 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_124 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_135 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_146 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_179 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_168 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_62 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vgnd scs8hd_diode_2
XFILLER_21_95 vgnd vgnd scs8hd_fill_2
XFILLER_21_84 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_SLEEPB _058_/Y vgnd vgnd scs8hd_diode_2
XFILLER_11_9 vgnd vgnd scs8hd_fill_2
XFILLER_30_121 vgnd vgnd scs8hd_fill_2
XPHY_4 vgnd vgnd scs8hd_decap_3
Xmux_bottom_track_9.INVTX1_8_.scs8hd_inv_1 chanx_left_in[8] mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_15_140 vgnd vgnd scs8hd_fill_1
XFILLER_15_173 vgnd vgnd scs8hd_decap_4
Xmux_left_track_9.INVTX1_5_.scs8hd_inv_1 vgnd mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_7_53 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_26_29 vgnd vgnd scs8hd_fill_2
XFILLER_21_110 vgnd vgnd scs8hd_fill_2
XFILLER_29_221 vgnd vgnd scs8hd_fill_2
XFILLER_29_210 vgnd vgnd scs8hd_decap_4
XFILLER_8_114 vgnd vgnd scs8hd_fill_2
XFILLER_12_121 vgnd vgnd scs8hd_fill_2
XFILLER_12_143 vgnd vgnd scs8hd_fill_1
XFILLER_12_165 vgnd vgnd scs8hd_fill_1
XFILLER_16_84 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_SLEEPB _151_/Y vgnd vgnd scs8hd_diode_2
XFILLER_12_198 vgnd vgnd scs8hd_fill_2
XANTENNA__103__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_bottom_track_17.LATCH_4_.latch/Q mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_26_224 vgnd vgnd scs8hd_decap_8
XFILLER_26_213 vgnd vgnd scs8hd_fill_1
XFILLER_5_139 vgnd vgnd scs8hd_fill_2
XFILLER_5_128 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[4] vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_1.LATCH_3_.latch vgnd vgnd _100_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_4_194 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_SLEEPB _125_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
X_181_ _181_/A chanx_right_out[8] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[3] vgnd vgnd scs8hd_diode_2
XANTENNA__100__B vgnd vgnd vgnd scs8hd_diode_2
Xmem_left_track_1.LATCH_2_.latch vgnd mem_left_track_1.LATCH_2_.latch/Q _120_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_1_164 vgnd vgnd scs8hd_decap_4
XFILLER_1_175 vgnd vgnd scs8hd_fill_2
XFILLER_1_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_9_231 vgnd vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[4] mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__201__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_24_51 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmem_right_track_16.LATCH_3_.latch vgnd mem_right_track_16.LATCH_3_.latch/Q _142_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
X_095_ vgnd _086_/D chany_top_in[1] vgnd vgnd vgnd vgnd scs8hd_or4_4
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_24_73 vgnd vgnd scs8hd_fill_1
X_164_ vgnd _164_/LO vgnd vgnd scs8hd_conb_1
XFILLER_6_201 vgnd vgnd scs8hd_fill_2
XANTENNA__111__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_28_127 vgnd vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[4] mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_10_86 vgnd vgnd scs8hd_fill_2
XFILLER_34_119 vgnd vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_19_62 vgnd vgnd scs8hd_fill_2
XFILLER_35_72 vgnd vgnd scs8hd_fill_2
XFILLER_27_193 vgnd vgnd scs8hd_fill_2
XANTENNA__106__A _053_/X vgnd vgnd scs8hd_diode_2
X_147_ _056_/B _152_/B _147_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
X_078_ _053_/X vgnd _078_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_18_3 vgnd vgnd scs8hd_fill_1
XFILLER_18_171 vgnd vgnd scs8hd_fill_2
XFILLER_18_193 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XPHY_169 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_24_163 vgnd vgnd scs8hd_fill_2
XPHY_158 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_103 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_114 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_125 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_136 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_147 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_30 vgnd vgnd scs8hd_decap_4
Xmux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_top_track_16.LATCH_3_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_SLEEPB _120_/Y vgnd vgnd scs8hd_diode_2
XPHY_5 vgnd vgnd scs8hd_decap_3
XFILLER_7_43 vgnd vgnd scs8hd_fill_1
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 _067_/X mem_bottom_track_17.LATCH_2_.latch/Q
+ mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_8_.scs8hd_inv_1 left_top_grid_pin_10_ mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_7_65 vgnd vgnd scs8hd_decap_3
XFILLER_26_19 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_21_177 vgnd vgnd scs8hd_decap_4
XFILLER_32_73 vgnd vgnd scs8hd_fill_2
XFILLER_32_62 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 vgnd mem_left_track_17.LATCH_3_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_12_177 vgnd vgnd scs8hd_fill_2
XFILLER_32_84 vgnd vgnd scs8hd_fill_2
XANTENNA__103__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_35_225 vgnd vgnd scs8hd_decap_8
XANTENNA_mem_right_track_16.LATCH_2_.latch_SLEEPB _143_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__204__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_5_118 vgnd vgnd scs8hd_fill_2
XFILLER_27_40 vgnd vgnd scs8hd_fill_2
XFILLER_17_214 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__114__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_16.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_4_162 vgnd vgnd scs8hd_fill_2
XFILLER_4_140 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[2] mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_217 vgnd vgnd scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_2_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_228 vgnd vgnd scs8hd_fill_2
X_180_ _180_/A chanx_left_out[0] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_13_53 vgnd vgnd scs8hd_fill_2
XFILLER_13_75 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A _124_/B vgnd vgnd
+ scs8hd_diode_2
XFILLER_1_143 vgnd vgnd scs8hd_fill_2
XANTENNA__109__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _163_/HI vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_094_ vgnd _086_/X _094_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_213 vgnd vgnd scs8hd_fill_1
XFILLER_6_224 vgnd vgnd scs8hd_fill_2
X_163_ _163_/HI _163_/LO vgnd vgnd scs8hd_conb_1
XANTENNA__111__B _110_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_SLEEPB _159_/Y vgnd vgnd scs8hd_diode_2
Xmem_top_track_8.LATCH_2_.latch vgnd mem_top_track_8.LATCH_2_.latch/Q _073_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmem_right_track_0.LATCH_2_.latch vgnd mem_right_track_0.LATCH_2_.latch/Q _082_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_29_19 vgnd vgnd scs8hd_fill_2
XFILLER_28_106 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_10_32 vgnd vgnd scs8hd_fill_2
XFILLER_10_54 vgnd vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 vgnd mem_top_track_16.LATCH_1_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XANTENNA__106__B _110_/B vgnd vgnd scs8hd_diode_2
X_146_ vgnd vgnd vgnd chanx_right_in[2] _152_/B vgnd vgnd scs8hd_or4_4
XANTENNA__122__A vgnd vgnd vgnd scs8hd_diode_2
X_077_ vgnd vgnd _077_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_32_6 vgnd vgnd scs8hd_fill_2
XFILLER_33_197 vgnd vgnd scs8hd_fill_2
XFILLER_33_153 vgnd vgnd scs8hd_fill_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_1_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vgnd scs8hd_diode_2
XFILLER_0_208 vgnd vgnd scs8hd_fill_2
XANTENNA__207__A _207_/A vgnd vgnd scs8hd_diode_2
XFILLER_24_197 vgnd vgnd scs8hd_fill_2
XFILLER_24_186 vgnd vgnd scs8hd_fill_2
XFILLER_24_142 vgnd vgnd scs8hd_fill_2
XPHY_159 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_148 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_104 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_115 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_126 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_137 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_53 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_30_101 vgnd vgnd scs8hd_fill_2
XPHY_6 vgnd vgnd scs8hd_decap_3
XFILLER_30_167 vgnd vgnd scs8hd_decap_4
XFILLER_30_145 vgnd vgnd scs8hd_fill_2
XFILLER_30_134 vgnd vgnd scs8hd_fill_2
XANTENNA__117__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_15_197 vgnd vgnd scs8hd_fill_2
XFILLER_30_3 vgnd vgnd scs8hd_fill_2
X_129_ vgnd _124_/B _129_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_top_track_16.INVTX1_3_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_21_123 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ chany_bottom_in[1] mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_12_101 vgnd vgnd scs8hd_fill_2
XFILLER_16_64 vgnd vgnd scs8hd_fill_2
XFILLER_8_127 vgnd vgnd scs8hd_fill_2
XFILLER_8_149 vgnd vgnd scs8hd_fill_2
XFILLER_16_97 vgnd vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_right_track_0.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_7_193 vgnd vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_7_.latch vgnd mem_top_track_0.LATCH_7_.latch/Q _052_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_4_.latch vgnd vgnd _110_/B vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_17_226 vgnd vgnd scs8hd_fill_2
XFILLER_27_96 vgnd vgnd scs8hd_fill_1
XANTENNA__114__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__130__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_4_152 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_229 vgnd vgnd scs8hd_decap_4
XFILLER_13_32 vgnd vgnd scs8hd_fill_2
XFILLER_8_3 vgnd vgnd scs8hd_fill_1
Xmem_left_track_9.LATCH_3_.latch vgnd mem_left_track_9.LATCH_3_.latch/Q _128_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__109__B _110_/B vgnd vgnd scs8hd_diode_2
XFILLER_9_211 vgnd vgnd scs8hd_decap_4
XANTENNA__125__A _053_/X vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_6_.scs8hd_inv_1 vgnd mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_SLEEPB _111_/Y vgnd vgnd scs8hd_diode_2
XFILLER_24_42 vgnd vgnd scs8hd_decap_3
X_162_ _162_/HI _162_/LO vgnd vgnd scs8hd_conb_1
XFILLER_10_232 vgnd vgnd scs8hd_fill_1
Xmux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_3_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
X_093_ vgnd _086_/X _093_/Y vgnd vgnd scs8hd_nor2_4
Xmem_top_track_16.LATCH_4_.latch vgnd mem_top_track_16.LATCH_4_.latch/Q _134_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_3_217 vgnd vgnd scs8hd_fill_1
XFILLER_19_53 vgnd vgnd scs8hd_fill_2
XFILLER_19_118 vgnd vgnd scs8hd_fill_2
XFILLER_35_85 vgnd vgnd scs8hd_fill_2
XFILLER_35_52 vgnd vgnd scs8hd_decap_4
XFILLER_35_41 vgnd vgnd scs8hd_fill_2
XFILLER_27_173 vgnd vgnd scs8hd_fill_2
X_145_ vgnd _141_/B _145_/Y vgnd vgnd scs8hd_nor2_4
Xmux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ mem_right_track_0.LATCH_5_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA__122__B _114_/X vgnd vgnd scs8hd_diode_2
X_076_ chany_top_in[1] vgnd vgnd _067_/D vgnd vgnd vgnd scs8hd_or4_4
XFILLER_33_132 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_1_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XPHY_105 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_116 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_149 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_10 vgnd vgnd scs8hd_fill_2
XPHY_127 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_138 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_7 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_right_track_0.LATCH_3_.latch_SLEEPB _081_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_15_132 vgnd vgnd scs8hd_fill_2
XFILLER_15_143 vgnd vgnd scs8hd_fill_2
XFILLER_15_154 vgnd vgnd scs8hd_decap_4
XANTENNA__117__B _114_/X vgnd vgnd scs8hd_diode_2
XANTENNA__133__A _056_/B vgnd vgnd scs8hd_diode_2
X_128_ chanx_right_in[2] _124_/B _128_/Y vgnd vgnd scs8hd_nor2_4
X_059_ address[2] _043_/Y _063_/C chanx_right_in[2] vgnd vgnd scs8hd_or3_4
Xmux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XFILLER_21_157 vgnd vgnd scs8hd_fill_2
XFILLER_21_146 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__043__A address[1] vgnd vgnd scs8hd_diode_2
XFILLER_12_135 vgnd vgnd scs8hd_fill_2
XFILLER_16_32 vgnd vgnd scs8hd_fill_2
XFILLER_16_43 vgnd vgnd scs8hd_fill_2
XFILLER_8_106 vgnd vgnd scs8hd_fill_2
XFILLER_12_146 vgnd vgnd scs8hd_fill_2
XFILLER_12_157 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.INVTX1_5_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__128__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_5_109 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_SLEEPB _070_/Y vgnd vgnd scs8hd_diode_2
XFILLER_27_75 vgnd vgnd scs8hd_fill_2
XFILLER_27_53 vgnd vgnd scs8hd_fill_2
XFILLER_27_20 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_top_track_0.INVTX1_7_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_32_219 vgnd vgnd scs8hd_decap_12
XANTENNA__114__C vgnd vgnd vgnd scs8hd_diode_2
XFILLER_4_175 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA__130__B _124_/B vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmem_bottom_track_17.LATCH_4_.latch vgnd mem_bottom_track_17.LATCH_4_.latch/Q _148_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_13_22 vgnd vgnd scs8hd_decap_3
XFILLER_14_208 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__125__B _124_/B vgnd vgnd scs8hd_diode_2
XFILLER_9_223 vgnd vgnd scs8hd_fill_2
XFILLER_13_230 vgnd vgnd scs8hd_decap_3
XANTENNA__141__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _168_/HI mem_right_track_8.LATCH_7_.latch/Q
+ mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XANTENNA__051__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_24_87 vgnd vgnd scs8hd_fill_2
XFILLER_24_65 vgnd vgnd scs8hd_fill_2
XFILLER_24_32 vgnd vgnd scs8hd_decap_3
XFILLER_24_21 vgnd vgnd scs8hd_fill_2
X_161_ _161_/HI _161_/LO vgnd vgnd scs8hd_conb_1
XFILLER_10_211 vgnd vgnd scs8hd_fill_1
X_092_ vgnd _086_/X _092_/Y vgnd vgnd scs8hd_nor2_4
Xmux_right_track_0.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmem_right_track_8.LATCH_3_.latch vgnd mem_right_track_8.LATCH_3_.latch/Q _091_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__136__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__046__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_3_229 vgnd vgnd scs8hd_fill_2
XFILLER_10_67 vgnd vgnd scs8hd_fill_2
XFILLER_10_78 vgnd vgnd scs8hd_fill_2
XFILLER_19_10 vgnd vgnd scs8hd_fill_2
XFILLER_19_98 vgnd vgnd scs8hd_decap_4
X_075_ vgnd _067_/X _056_/B vgnd vgnd scs8hd_nor2_4
X_144_ vgnd _141_/B _144_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_25_7 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_141 vgnd vgnd scs8hd_fill_1
XFILLER_18_163 vgnd vgnd scs8hd_fill_2
XFILLER_33_177 vgnd vgnd scs8hd_decap_4
XFILLER_33_166 vgnd vgnd scs8hd_decap_4
XANTENNA_mem_top_track_0.LATCH_1_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_2_90 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_5_.scs8hd_inv_1 bottom_left_grid_pin_13_ mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XPHY_106 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_117 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_128 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_139 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_21_22 vgnd vgnd scs8hd_fill_2
XFILLER_21_66 vgnd vgnd scs8hd_fill_1
XPHY_8 vgnd vgnd scs8hd_decap_3
XFILLER_15_177 vgnd vgnd scs8hd_fill_1
X_058_ _056_/B vgnd _058_/Y vgnd vgnd scs8hd_nor2_4
X_127_ vgnd _124_/B _127_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_7_79 vgnd vgnd scs8hd_fill_2
XANTENNA__133__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_16_3 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1 mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ _198_/A vgnd vgnd scs8hd_inv_1
XFILLER_21_114 vgnd vgnd scs8hd_fill_2
Xmux_top_track_16.INVTX1_6_.scs8hd_inv_1 chanx_left_in[5] vgnd vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_6_.latch/Q mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_29_225 vgnd vgnd scs8hd_fill_2
XFILLER_29_214 vgnd vgnd scs8hd_fill_1
XFILLER_16_11 vgnd vgnd scs8hd_fill_1
XFILLER_32_10 vgnd vgnd scs8hd_fill_2
XFILLER_12_125 vgnd vgnd scs8hd_fill_1
XFILLER_16_88 vgnd vgnd scs8hd_fill_2
XFILLER_32_32 vgnd vgnd scs8hd_fill_2
XFILLER_20_180 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__144__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__128__B _124_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
XANTENNA__054__A _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_3_.latch_SLEEPB _128_/Y vgnd vgnd scs8hd_diode_2
XFILLER_17_217 vgnd vgnd scs8hd_fill_1
XANTENNA__114__D chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XFILLER_4_198 vgnd vgnd scs8hd_fill_2
XFILLER_4_154 vgnd vgnd scs8hd_fill_2
XFILLER_4_110 vgnd vgnd scs8hd_fill_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _169_/HI mem_top_track_0.LATCH_7_.latch/Q
+ mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XANTENNA__139__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__049__A _055_/A vgnd vgnd scs8hd_diode_2
XFILLER_13_45 vgnd vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_2_.scs8hd_inv_1 vgnd mux_top_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_1_168 vgnd vgnd scs8hd_fill_1
XFILLER_1_179 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__141__B _141_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__051__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_24_11 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _169_/HI vgnd vgnd
+ scs8hd_diode_2
Xmux_right_track_8.INVTX1_3_.scs8hd_inv_1 right_bottom_grid_pin_12_ mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_091_ chanx_right_in[2] _086_/X _091_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_24_55 vgnd vgnd scs8hd_fill_1
X_160_ _160_/HI _160_/LO vgnd vgnd scs8hd_conb_1
XFILLER_6_205 vgnd vgnd scs8hd_fill_2
XANTENNA__136__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__152__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__062__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_27_153 vgnd vgnd scs8hd_fill_2
XFILLER_19_77 vgnd vgnd scs8hd_fill_2
XFILLER_35_76 vgnd vgnd scs8hd_fill_2
XFILLER_35_10 vgnd vgnd scs8hd_fill_2
XFILLER_27_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_5_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
X_143_ vgnd _141_/B _143_/Y vgnd vgnd scs8hd_nor2_4
X_074_ vgnd _067_/X _074_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_1_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_18_7 vgnd vgnd scs8hd_fill_2
XFILLER_18_197 vgnd vgnd scs8hd_fill_2
XANTENNA__147__A _056_/B vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vgnd scs8hd_diode_2
XFILLER_24_167 vgnd vgnd scs8hd_fill_2
XANTENNA__057__A _055_/A vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_8_.scs8hd_inv_1 chanx_left_in[7] mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.INVTX1_5_.scs8hd_inv_1 vgnd mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XPHY_107 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_118 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_129 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_9 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_057_ _055_/A address[1] address[0] vgnd vgnd vgnd scs8hd_or3_4
X_126_ _056_/B _124_/B vgnd vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_top_track_0.INVTX1_2_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[5] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _166_/HI vgnd vgnd
+ scs8hd_diode_2
XFILLER_16_23 vgnd vgnd scs8hd_fill_2
XFILLER_32_88 vgnd vgnd scs8hd_fill_2
XFILLER_32_66 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_35_207 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA__144__B _141_/B vgnd vgnd scs8hd_diode_2
XFILLER_7_141 vgnd vgnd scs8hd_decap_4
XFILLER_7_163 vgnd vgnd scs8hd_decap_4
XFILLER_7_174 vgnd vgnd scs8hd_fill_2
X_109_ chanx_right_in[2] _110_/B _109_/Y vgnd vgnd scs8hd_nor2_4
Xmux_left_track_17.INVTX1_0_.scs8hd_inv_1 chany_top_in[1] vgnd vgnd vgnd scs8hd_inv_1
XANTENNA__054__B _053_/X vgnd vgnd scs8hd_diode_2
XANTENNA__070__A _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_27_99 vgnd vgnd scs8hd_decap_4
XFILLER_27_88 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_144 vgnd vgnd scs8hd_fill_2
XANTENNA__155__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_31_221 vgnd vgnd scs8hd_fill_2
XFILLER_31_210 vgnd vgnd scs8hd_decap_4
XANTENNA__139__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[5] vgnd vgnd scs8hd_diode_2
XANTENNA__049__B _043_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__065__A address[2] vgnd vgnd scs8hd_diode_2
XFILLER_22_232 vgnd vgnd scs8hd_fill_1
XFILLER_13_57 vgnd vgnd scs8hd_fill_2
XFILLER_13_79 vgnd vgnd scs8hd_fill_1
XFILLER_1_147 vgnd vgnd scs8hd_fill_2
XANTENNA__051__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_6_228 vgnd vgnd scs8hd_fill_2
XFILLER_10_224 vgnd vgnd scs8hd_fill_2
X_090_ vgnd _086_/X _090_/Y vgnd vgnd scs8hd_nor2_4
Xmux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_0_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmux_right_track_0.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[7] mux_right_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__152__B _152_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__062__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_10_36 vgnd vgnd scs8hd_decap_3
XFILLER_27_132 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 vgnd mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_19_23 vgnd vgnd scs8hd_fill_2
XFILLER_19_34 vgnd vgnd scs8hd_fill_2
X_142_ chanx_right_in[2] _141_/B _142_/Y vgnd vgnd scs8hd_nor2_4
X_073_ vgnd _067_/X _073_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_bottom_track_17.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_33_102 vgnd vgnd scs8hd_fill_2
XANTENNA__147__B _152_/B vgnd vgnd scs8hd_diode_2
XFILLER_18_121 vgnd vgnd scs8hd_fill_2
XFILLER_18_132 vgnd vgnd scs8hd_fill_2
XFILLER_18_176 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_24_102 vgnd vgnd scs8hd_fill_2
XFILLER_24_146 vgnd vgnd scs8hd_decap_4
XANTENNA__057__B address[1] vgnd vgnd scs8hd_diode_2
XPHY_108 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_119 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA__073__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_21_57 vgnd vgnd scs8hd_fill_2
XFILLER_15_102 vgnd vgnd scs8hd_decap_4
XFILLER_15_113 vgnd vgnd scs8hd_decap_3
X_125_ _053_/X _124_/B _125_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_30_149 vgnd vgnd scs8hd_fill_2
XFILLER_30_138 vgnd vgnd scs8hd_fill_2
XFILLER_30_105 vgnd vgnd scs8hd_decap_3
XFILLER_7_59 vgnd vgnd scs8hd_fill_2
X_056_ _056_/B _056_/B vgnd vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__158__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_21_127 vgnd vgnd scs8hd_fill_2
XANTENNA__068__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_16_68 vgnd vgnd scs8hd_fill_2
XFILLER_32_45 vgnd vgnd scs8hd_fill_2
XFILLER_32_23 vgnd vgnd scs8hd_fill_2
XFILLER_20_193 vgnd vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_2_.latch vgnd vgnd _062_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_12_105 vgnd vgnd scs8hd_fill_1
X_108_ vgnd _110_/B _110_/B vgnd vgnd scs8hd_nor2_4
XFILLER_7_197 vgnd vgnd scs8hd_fill_2
XFILLER_11_193 vgnd vgnd scs8hd_fill_2
XFILLER_21_3 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vgnd
+ scs8hd_diode_2
Xmux_top_track_8.tap_buf4_0_.scs8hd_inv_1 mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ _203_/A vgnd vgnd scs8hd_inv_1
XANTENNA__070__B _067_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_4_.latch_SLEEPB _090_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_27_12 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_left_track_17.LATCH_5_.latch vgnd mem_left_track_17.LATCH_5_.latch/Q _154_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_123 vgnd vgnd scs8hd_fill_2
XANTENNA__139__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__155__B _159_/B vgnd vgnd scs8hd_diode_2
XANTENNA__049__C _063_/C vgnd vgnd scs8hd_diode_2
XFILLER_22_211 vgnd vgnd scs8hd_decap_3
XFILLER_22_200 vgnd vgnd scs8hd_fill_1
XANTENNA__065__B address[1] vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_3_.scs8hd_inv_1 chanx_right_in[6] mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_13_14 vgnd vgnd scs8hd_fill_2
XFILLER_1_126 vgnd vgnd scs8hd_fill_2
XANTENNA__081__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_7_.latch_SLEEPB _115_/Y vgnd vgnd scs8hd_diode_2
XFILLER_13_222 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_0_181 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__051__D _067_/D vgnd vgnd scs8hd_diode_2
XFILLER_10_203 vgnd vgnd scs8hd_fill_2
XANTENNA__076__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_1_.scs8hd_inv_1_A chany_top_in[6] vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_1.LATCH_4_.latch vgnd mem_bottom_track_1.LATCH_4_.latch/Q _099_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_0_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_35_45 vgnd vgnd scs8hd_fill_2
XFILLER_35_23 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_3_.scs8hd_inv_1_A right_bottom_grid_pin_12_ vgnd
+ vgnd scs8hd_diode_2
XFILLER_27_177 vgnd vgnd scs8hd_decap_4
XFILLER_27_166 vgnd vgnd scs8hd_decap_4
XFILLER_19_57 vgnd vgnd scs8hd_fill_2
XFILLER_35_89 vgnd vgnd scs8hd_fill_2
X_141_ vgnd _141_/B _141_/Y vgnd vgnd scs8hd_nor2_4
X_072_ chanx_right_in[2] _067_/X _072_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_2_232 vgnd vgnd scs8hd_fill_1
Xmux_right_track_16.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XFILLER_33_136 vgnd vgnd scs8hd_fill_2
XFILLER_33_114 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_0_.latch_SLEEPB _084_/Y vgnd vgnd scs8hd_diode_2
Xmem_left_track_1.LATCH_3_.latch vgnd mem_left_track_1.LATCH_3_.latch/Q _119_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_24_125 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_32_180 vgnd vgnd scs8hd_decap_4
XFILLER_24_136 vgnd vgnd scs8hd_decap_4
XANTENNA__057__C address[0] vgnd vgnd scs8hd_diode_2
XPHY_109 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA__073__B _067_/X vgnd vgnd scs8hd_diode_2
XFILLER_21_36 vgnd vgnd scs8hd_fill_2
XFILLER_21_14 vgnd vgnd scs8hd_fill_2
XFILLER_30_117 vgnd vgnd scs8hd_fill_2
XFILLER_15_136 vgnd vgnd scs8hd_decap_4
XFILLER_15_158 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
X_055_ _055_/A address[1] _063_/C _056_/B vgnd vgnd scs8hd_or3_4
X_124_ vgnd _124_/B _124_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_left_track_17.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[7] vgnd vgnd scs8hd_diode_2
XFILLER_23_7 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_11_91 vgnd vgnd scs8hd_fill_2
XANTENNA__158__B _159_/B vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 vgnd mem_bottom_track_17.LATCH_5_.latch/Q
+ mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
Xmem_right_track_16.LATCH_4_.latch vgnd chany_bottom_in[1] _141_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__174__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_29_217 vgnd vgnd scs8hd_fill_1
XANTENNA__068__B _067_/X vgnd vgnd scs8hd_diode_2
XFILLER_12_117 vgnd vgnd scs8hd_fill_2
XFILLER_16_47 vgnd vgnd scs8hd_fill_2
XANTENNA__084__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_161 vgnd vgnd scs8hd_fill_2
XFILLER_12_139 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_SLEEPB _073_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_SLEEPB _154_/Y vgnd vgnd scs8hd_diode_2
X_107_ _056_/B _110_/B _107_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_27_57 vgnd vgnd scs8hd_fill_2
XFILLER_27_24 vgnd vgnd scs8hd_fill_1
XANTENNA__079__A _056_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[4] vgnd vgnd scs8hd_diode_2
XFILLER_4_102 vgnd vgnd scs8hd_fill_2
XFILLER_4_179 vgnd vgnd scs8hd_fill_2
XANTENNA__139__D _086_/D vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 vgnd mem_left_track_9.LATCH_0_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__065__C address[0] vgnd vgnd scs8hd_diode_2
XANTENNA__081__B vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_1_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_9_227 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.INVTX1_2_.scs8hd_inv_1_A chanx_right_in[2] vgnd vgnd
+ scs8hd_diode_2
XANTENNA__182__A chanx_left_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_5_71 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_24_69 vgnd vgnd scs8hd_fill_2
XFILLER_24_47 vgnd vgnd scs8hd_fill_2
XFILLER_24_25 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__076__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__092__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_1_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_14_91 vgnd vgnd scs8hd_fill_1
XANTENNA__177__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA__087__A vgnd vgnd vgnd scs8hd_diode_2
X_071_ vgnd _067_/X vgnd vgnd vgnd scs8hd_nor2_4
X_140_ _056_/B _141_/B _140_/Y vgnd vgnd scs8hd_nor2_4
Xmux_bottom_track_9.INVTX1_2_.scs8hd_inv_1 chanx_right_in[0] mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_4_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_18_145 vgnd vgnd scs8hd_fill_2
XFILLER_18_167 vgnd vgnd scs8hd_fill_2
XPHY_90 vgnd vgnd scs8hd_tapvpwrvgnd_1
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_21_26 vgnd vgnd scs8hd_fill_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_4_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
Xmux_top_track_16.INVTX1_3_.scs8hd_inv_1 vgnd mux_top_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_123_ chany_top_in[1] vgnd vgnd chanx_right_in[2] _124_/B vgnd vgnd scs8hd_or4_4
X_054_ _056_/B _053_/X _054_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_11_70 vgnd vgnd scs8hd_decap_4
XFILLER_16_7 vgnd vgnd scs8hd_fill_2
XFILLER_21_118 vgnd vgnd scs8hd_fill_2
XFILLER_14_170 vgnd vgnd scs8hd_fill_2
XANTENNA__190__A _190_/A vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_6_.latch_SLEEPB _106_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_29_229 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmem_right_track_0.LATCH_3_.latch vgnd mem_right_track_0.LATCH_3_.latch/Q _081_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_3_.latch vgnd mem_top_track_8.LATCH_3_.latch/Q _072_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__084__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_20_140 vgnd vgnd scs8hd_decap_4
XFILLER_7_100 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_0_.latch_SLEEPB _131_/Y vgnd vgnd scs8hd_diode_2
X_106_ _053_/X _110_/B _106_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_22_91 vgnd vgnd scs8hd_fill_1
XFILLER_34_232 vgnd vgnd scs8hd_fill_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_3_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA__185__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_27_36 vgnd vgnd scs8hd_fill_2
XFILLER_25_221 vgnd vgnd scs8hd_fill_2
XFILLER_25_210 vgnd vgnd scs8hd_decap_4
XANTENNA__079__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__095__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_4_158 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_16_232 vgnd vgnd scs8hd_fill_1
XFILLER_22_224 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_13_49 vgnd vgnd scs8hd_fill_2
XFILLER_13_213 vgnd vgnd scs8hd_fill_2
XFILLER_9_217 vgnd vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_0_.scs8hd_inv_1 chany_top_in[0] mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_6_209 vgnd vgnd scs8hd_fill_2
XANTENNA__076__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__092__B _086_/X vgnd vgnd scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_9.LATCH_5_.latch vgnd mem_bottom_track_9.LATCH_5_.latch/Q _107_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_bottom_track_1.LATCH_2_.latch_SLEEPB _101_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__193__A chany_top_in[4] vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_2_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_2_.scs8hd_inv_1_A chany_top_in[7] vgnd vgnd scs8hd_diode_2
XFILLER_10_28 vgnd vgnd scs8hd_decap_3
XFILLER_35_58 vgnd vgnd scs8hd_fill_2
XANTENNA__087__B _086_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_070_ _056_/B _067_/X _070_/Y vgnd vgnd scs8hd_nor2_4
Xmux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 _180_/A vgnd mux_left_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_left_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_bottom_track_1.INVTX1_5_.scs8hd_inv_1 bottom_right_grid_pin_11_ mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_18_113 vgnd vgnd scs8hd_fill_2
XFILLER_33_149 vgnd vgnd scs8hd_fill_2
XPHY_91 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_80 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_199_ _199_/A chany_top_out[8] vgnd vgnd scs8hd_buf_2
Xmem_left_track_9.LATCH_4_.latch vgnd mem_left_track_9.LATCH_4_.latch/Q _127_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.INVTX1_4_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA__188__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 vgnd mem_bottom_track_9.LATCH_5_.latch/Q
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
Xmux_top_track_8.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[1] mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_21_49 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__098__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_23_193 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_ebufn_2
X_053_ _055_/A _043_/Y address[0] _053_/X vgnd vgnd scs8hd_or3_4
X_122_ vgnd _114_/X _122_/Y vgnd vgnd scs8hd_nor2_4
Xmux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_3_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_4_.latch_SLEEPB _134_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _162_/HI vgnd vgnd
+ scs8hd_diode_2
Xmem_top_track_16.LATCH_5_.latch vgnd mem_top_track_16.LATCH_5_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_16_27 vgnd vgnd scs8hd_fill_2
X_105_ vgnd _110_/B vgnd vgnd vgnd scs8hd_nor2_4
XFILLER_7_123 vgnd vgnd scs8hd_fill_2
XFILLER_7_145 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_7_178 vgnd vgnd scs8hd_decap_3
XFILLER_19_230 vgnd vgnd scs8hd_decap_3
XFILLER_8_61 vgnd vgnd scs8hd_fill_2
XANTENNA__095__B _086_/D vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_148 vgnd vgnd scs8hd_fill_2
XFILLER_31_225 vgnd vgnd scs8hd_decap_8
XFILLER_31_214 vgnd vgnd scs8hd_fill_1
XFILLER_16_211 vgnd vgnd scs8hd_decap_3
XFILLER_17_92 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_6_.latch_SLEEPB _054_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__196__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[4] mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_22_203 vgnd vgnd scs8hd_fill_2
XFILLER_13_28 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_0_173 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_3_.latch_SLEEPB _149_/Y vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.INVTX1_3_.scs8hd_inv_1 right_top_grid_pin_10_ mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_5_84 vgnd vgnd scs8hd_fill_2
XFILLER_24_38 vgnd vgnd scs8hd_fill_2
XANTENNA__076__D _067_/D vgnd vgnd scs8hd_diode_2
XFILLER_10_228 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_60 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_6_.latch/Q mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_5_210 vgnd vgnd scs8hd_decap_4
XFILLER_5_221 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
Xmem_bottom_track_17.LATCH_5_.latch vgnd mem_bottom_track_17.LATCH_5_.latch/Q _147_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_27_136 vgnd vgnd scs8hd_fill_2
XFILLER_27_114 vgnd vgnd scs8hd_fill_2
XFILLER_19_27 vgnd vgnd scs8hd_fill_2
XFILLER_19_38 vgnd vgnd scs8hd_fill_2
XFILLER_2_213 vgnd vgnd scs8hd_fill_1
XFILLER_2_224 vgnd vgnd scs8hd_fill_2
XFILLER_33_106 vgnd vgnd scs8hd_fill_2
XFILLER_26_180 vgnd vgnd scs8hd_fill_2
XFILLER_18_136 vgnd vgnd scs8hd_decap_3
XPHY_70 vgnd vgnd scs8hd_decap_3
XPHY_92 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_81 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_198_ _198_/A chany_bottom_out[0] vgnd vgnd scs8hd_buf_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_2_96 vgnd vgnd scs8hd_fill_1
XFILLER_32_150 vgnd vgnd scs8hd_fill_1
XFILLER_24_106 vgnd vgnd scs8hd_fill_2
XFILLER_17_180 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.INVTX1_7_.scs8hd_inv_1 vgnd mux_top_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA__098__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_15_106 vgnd vgnd scs8hd_fill_1
X_121_ vgnd _114_/X _121_/Y vgnd vgnd scs8hd_nor2_4
X_052_ vgnd _056_/B _052_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_left_track_1.INVTX1_6_.scs8hd_inv_1_A chany_bottom_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_183 vgnd vgnd scs8hd_fill_2
XANTENNA__199__A _199_/A vgnd vgnd scs8hd_diode_2
Xmem_right_track_8.LATCH_4_.latch vgnd mem_right_track_8.LATCH_4_.latch/Q _090_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_32_49 vgnd vgnd scs8hd_fill_2
XFILLER_32_27 vgnd vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_8_.scs8hd_inv_1 chanx_left_in[5] mux_right_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_0.INVTX1_8_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_20_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_1_.latch_SLEEPB _093_/Y vgnd vgnd scs8hd_diode_2
X_104_ chany_top_in[1] vgnd vgnd _086_/D _110_/B vgnd vgnd scs8hd_or4_4
XFILLER_22_60 vgnd vgnd scs8hd_fill_2
Xmem_left_track_17.LATCH_0_.latch vgnd mem_left_track_17.LATCH_0_.latch/Q _159_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_11_164 vgnd vgnd scs8hd_fill_2
XFILLER_11_175 vgnd vgnd scs8hd_fill_2
XFILLER_11_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_8_.scs8hd_inv_1_A left_bottom_grid_pin_12_ vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_8_84 vgnd vgnd scs8hd_fill_2
XFILLER_27_16 vgnd vgnd scs8hd_fill_2
XANTENNA__095__C chany_top_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_4_127 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_0_.scs8hd_inv_1 vgnd mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_3_193 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_SLEEPB _118_/Y vgnd vgnd scs8hd_diode_2
XFILLER_13_18 vgnd vgnd scs8hd_fill_2
XFILLER_13_204 vgnd vgnd scs8hd_fill_2
XFILLER_13_226 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_7_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_0_185 vgnd vgnd scs8hd_fill_1
XFILLER_0_196 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_4_.latch_SLEEPB _141_/Y vgnd vgnd scs8hd_diode_2
XFILLER_10_207 vgnd vgnd scs8hd_decap_4
XFILLER_14_83 vgnd vgnd scs8hd_fill_2
XFILLER_30_93 vgnd vgnd scs8hd_fill_1
Xmux_left_track_17.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[1] _180_/A vgnd vgnd scs8hd_inv_1
Xmux_right_track_16.INVTX1_4_.scs8hd_inv_1 chany_bottom_in[6] mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_35_27 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XPHY_71 vgnd vgnd scs8hd_decap_3
XFILLER_33_118 vgnd vgnd scs8hd_fill_2
XPHY_60 vgnd vgnd scs8hd_decap_3
XPHY_82 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_197_ chany_top_in[0] chany_bottom_out[1] vgnd vgnd scs8hd_buf_2
XFILLER_25_82 vgnd vgnd scs8hd_fill_2
XPHY_93 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_top_track_16.tap_buf4_0_.scs8hd_inv_1 mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A
+ _199_/A vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _163_/HI mem_left_track_1.LATCH_7_.latch/Q
+ mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XFILLER_21_18 vgnd vgnd scs8hd_fill_1
XFILLER_15_118 vgnd vgnd scs8hd_fill_2
X_051_ vgnd vgnd vgnd _067_/D _056_/B vgnd vgnd scs8hd_or4_4
X_120_ vgnd _114_/X _120_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_23_173 vgnd vgnd scs8hd_fill_2
XFILLER_11_95 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd scs8hd_diode_2
XFILLER_14_151 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_17.LATCH_2_.latch_SLEEPB _157_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_176 vgnd vgnd scs8hd_fill_2
XFILLER_20_165 vgnd vgnd scs8hd_fill_2
XFILLER_20_121 vgnd vgnd scs8hd_fill_2
XFILLER_28_232 vgnd vgnd scs8hd_fill_1
XFILLER_11_132 vgnd vgnd scs8hd_fill_2
X_103_ vgnd vgnd _103_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_22_83 vgnd vgnd scs8hd_fill_2
XFILLER_7_114 vgnd vgnd scs8hd_fill_2
XFILLER_7_169 vgnd vgnd scs8hd_fill_2
XFILLER_11_143 vgnd vgnd scs8hd_decap_4
XFILLER_34_224 vgnd vgnd scs8hd_decap_8
XFILLER_34_213 vgnd vgnd scs8hd_fill_1
XFILLER_19_210 vgnd vgnd scs8hd_decap_4
XFILLER_8_30 vgnd vgnd scs8hd_fill_1
XANTENNA__095__D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_4_106 vgnd vgnd scs8hd_fill_2
XFILLER_16_224 vgnd vgnd scs8hd_fill_2
XFILLER_33_60 vgnd vgnd scs8hd_fill_1
XFILLER_3_172 vgnd vgnd scs8hd_decap_4
Xmux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_0_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_0_153 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_17.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_28_93 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_24_29 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.tap_buf4_0_.scs8hd_inv_1 mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd vgnd scs8hd_inv_1
XFILLER_30_83 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 vgnd mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA__101__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_7_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_1_.scs8hd_inv_1_A chany_top_in[3] vgnd vgnd scs8hd_diode_2
XFILLER_35_182 vgnd vgnd scs8hd_fill_2
XFILLER_27_149 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_18_149 vgnd vgnd scs8hd_fill_2
XPHY_61 vgnd vgnd scs8hd_decap_3
XPHY_50 vgnd vgnd scs8hd_decap_3
XPHY_94 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_83 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_72 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_196_ chany_top_in[1] chany_bottom_out[2] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_top_track_0.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[7] vgnd vgnd scs8hd_diode_2
Xmux_top_track_16.INVTX1_0_.scs8hd_inv_1 chanx_right_in[0] mux_top_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_2_32 vgnd vgnd scs8hd_fill_1
XFILLER_24_119 vgnd vgnd scs8hd_decap_4
XFILLER_32_163 vgnd vgnd scs8hd_decap_8
XANTENNA_mux_left_track_9.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_17_193 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_152 vgnd vgnd scs8hd_fill_2
XFILLER_23_130 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
X_050_ vgnd address[6] _067_/D vgnd vgnd scs8hd_or2_4
XANTENNA_mem_bottom_track_9.LATCH_3_.latch_SLEEPB _109_/Y vgnd vgnd scs8hd_diode_2
XFILLER_11_74 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_top_track_8.INVTX1_5_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_141 vgnd vgnd scs8hd_decap_4
XFILLER_14_174 vgnd vgnd scs8hd_fill_2
X_179_ chanx_right_in[0] chanx_left_out[1] vgnd vgnd scs8hd_buf_2
XFILLER_20_144 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_7_104 vgnd vgnd scs8hd_fill_1
X_102_ vgnd vgnd _102_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_7_137 vgnd vgnd scs8hd_fill_2
XFILLER_7_148 vgnd vgnd scs8hd_fill_2
XFILLER_19_222 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1_A chanx_left_in[7] vgnd vgnd scs8hd_diode_2
XFILLER_25_214 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_25_225 vgnd vgnd scs8hd_fill_2
XFILLER_31_217 vgnd vgnd scs8hd_fill_1
XFILLER_16_203 vgnd vgnd scs8hd_fill_2
XFILLER_17_73 vgnd vgnd scs8hd_fill_2
XFILLER_33_72 vgnd vgnd scs8hd_fill_2
XANTENNA__104__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_3_151 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_right_track_0.LATCH_5_.latch_SLEEPB _079_/Y vgnd vgnd scs8hd_diode_2
XFILLER_22_228 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_1_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_13_217 vgnd vgnd scs8hd_fill_1
XFILLER_28_72 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_8_232 vgnd vgnd scs8hd_fill_1
Xmem_top_track_0.LATCH_3_.latch vgnd mem_top_track_0.LATCH_3_.latch/Q _060_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmem_bottom_track_9.LATCH_0_.latch vgnd mem_bottom_track_9.LATCH_0_.latch/Q _112_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_1_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_top_track_8.LATCH_7_.latch_SLEEPB _068_/Y vgnd vgnd scs8hd_diode_2
XFILLER_14_30 vgnd vgnd scs8hd_fill_1
XFILLER_14_41 vgnd vgnd scs8hd_fill_2
XFILLER_14_96 vgnd vgnd scs8hd_fill_2
XFILLER_30_62 vgnd vgnd scs8hd_fill_2
XANTENNA__101__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_1.INVTX1_2_.scs8hd_inv_1 chanx_right_in[1] mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_2_205 vgnd vgnd scs8hd_fill_2
XANTENNA__202__A chany_bottom_in[4] vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_1_.scs8hd_inv_1 chanx_right_in[2] _124_/B vgnd vgnd scs8hd_inv_1
XFILLER_18_117 vgnd vgnd scs8hd_fill_2
XPHY_62 vgnd vgnd scs8hd_decap_3
XFILLER_26_150 vgnd vgnd scs8hd_fill_1
XPHY_51 vgnd vgnd scs8hd_decap_3
XPHY_95 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_84 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_73 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_40 vgnd vgnd scs8hd_decap_3
X_195_ vgnd chany_bottom_out[3] vgnd vgnd scs8hd_buf_2
XANTENNA__112__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_17_172 vgnd vgnd scs8hd_fill_2
XFILLER_32_197 vgnd vgnd scs8hd_decap_4
XFILLER_32_186 vgnd vgnd scs8hd_fill_2
XFILLER_32_142 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_1_.latch_SLEEPB _137_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_197 vgnd vgnd scs8hd_fill_2
XFILLER_23_120 vgnd vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_0_.latch vgnd mem_top_track_16.LATCH_0_.latch/Q _138_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_15_109 vgnd vgnd scs8hd_fill_2
XFILLER_11_20 vgnd vgnd scs8hd_fill_2
XFILLER_11_53 vgnd vgnd scs8hd_fill_2
XANTENNA__107__A _056_/B vgnd vgnd scs8hd_diode_2
X_178_ chanx_right_in[1] chanx_left_out[2] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_bottom_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vgnd
+ scs8hd_diode_2
Xmem_bottom_track_1.LATCH_5_.latch vgnd mem_bottom_track_1.LATCH_5_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_28_201 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_101_ vgnd vgnd _101_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_22_41 vgnd vgnd scs8hd_fill_2
XFILLER_22_30 vgnd vgnd scs8hd_fill_1
XFILLER_7_127 vgnd vgnd scs8hd_fill_1
XFILLER_22_96 vgnd vgnd scs8hd_fill_2
XFILLER_8_32 vgnd vgnd scs8hd_fill_1
XFILLER_8_65 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_6_182 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_3_.latch_SLEEPB _060_/Y vgnd vgnd scs8hd_diode_2
Xmem_left_track_1.LATCH_4_.latch vgnd mem_left_track_1.LATCH_4_.latch/Q _118_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_bottom_track_9.INVTX1_7_.scs8hd_inv_1 chanx_left_in[6] mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_9.INVTX1_4_.scs8hd_inv_1 vgnd vgnd vgnd vgnd scs8hd_inv_1
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_17_96 vgnd vgnd scs8hd_fill_2
XFILLER_33_62 vgnd vgnd scs8hd_fill_1
XANTENNA__104__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_3_130 vgnd vgnd scs8hd_fill_2
XANTENNA__120__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_22_207 vgnd vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_left_track_9.LATCH_4_.latch/Q mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA_mem_bottom_track_17.LATCH_0_.latch_SLEEPB _152_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_right_track_16.LATCH_5_.latch vgnd mem_right_track_16.LATCH_5_.latch/Q _140_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_0.INVTX1_0_.scs8hd_inv_1 vgnd mux_right_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_right_track_0.INVTX1_2_.scs8hd_inv_1_A chany_top_in[8] vgnd vgnd scs8hd_diode_2
XANTENNA__205__A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_28_84 vgnd vgnd scs8hd_fill_2
XFILLER_28_51 vgnd vgnd scs8hd_fill_2
XFILLER_0_177 vgnd vgnd scs8hd_fill_2
XANTENNA__115__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_5_88 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 mem_bottom_track_9.LATCH_1_.latch/Q
+ mem_bottom_track_9.LATCH_1_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_17.LATCH_0_.latch vgnd mem_bottom_track_17.LATCH_0_.latch/Q _152_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_8.INVTX1_4_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_5_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ mem_top_track_8.LATCH_5_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_30_41 vgnd vgnd scs8hd_fill_2
XFILLER_5_214 vgnd vgnd scs8hd_fill_1
XFILLER_5_225 vgnd vgnd scs8hd_fill_2
XFILLER_14_64 vgnd vgnd scs8hd_fill_2
XFILLER_29_170 vgnd vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_27_118 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_0_.scs8hd_inv_1_A top_right_grid_pin_11_ vgnd vgnd
+ scs8hd_diode_2
XFILLER_35_151 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_2_228 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_6_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.INVTX1_4_.scs8hd_inv_1 vgnd mux_top_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XPHY_30 vgnd vgnd scs8hd_decap_3
XPHY_63 vgnd vgnd scs8hd_decap_3
XFILLER_26_184 vgnd vgnd scs8hd_fill_2
XPHY_52 vgnd vgnd scs8hd_decap_3
XPHY_41 vgnd vgnd scs8hd_decap_3
XPHY_85 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_74 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_96 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_194_ _194_/A chany_bottom_out[4] vgnd vgnd scs8hd_buf_2
XANTENNA__112__B _110_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_165 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.INVTX1_3_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_11_43 vgnd vgnd scs8hd_fill_1
XFILLER_11_87 vgnd vgnd scs8hd_fill_2
Xmux_right_track_8.INVTX1_5_.scs8hd_inv_1 chany_bottom_in[3] mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_14_154 vgnd vgnd scs8hd_decap_3
XANTENNA__107__B _110_/B vgnd vgnd scs8hd_diode_2
X_177_ chanx_right_in[2] chanx_left_out[3] vgnd vgnd scs8hd_buf_2
XFILLER_14_187 vgnd vgnd scs8hd_fill_2
XANTENNA__123__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_20_157 vgnd vgnd scs8hd_fill_2
XFILLER_28_213 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1_A bottom_left_grid_pin_13_ vgnd
+ vgnd scs8hd_diode_2
XFILLER_28_224 vgnd vgnd scs8hd_decap_8
X_100_ chanx_right_in[2] vgnd _100_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_22_64 vgnd vgnd scs8hd_decap_3
XFILLER_11_113 vgnd vgnd scs8hd_fill_2
XFILLER_11_168 vgnd vgnd scs8hd_fill_2
XFILLER_11_179 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__118__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_8_44 vgnd vgnd scs8hd_fill_2
XFILLER_8_88 vgnd vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_1_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_SLEEPB _121_/Y vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_2_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmux_left_track_1.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[8] mux_left_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_17_20 vgnd vgnd scs8hd_fill_2
XFILLER_17_31 vgnd vgnd scs8hd_fill_2
XPHY_200 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_33_52 vgnd vgnd scs8hd_fill_2
XFILLER_17_53 vgnd vgnd scs8hd_fill_2
XFILLER_33_85 vgnd vgnd scs8hd_fill_2
XANTENNA__104__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_3_197 vgnd vgnd scs8hd_fill_2
XANTENNA__120__B _114_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[6] vgnd vgnd
+ scs8hd_diode_2
XFILLER_21_230 vgnd vgnd scs8hd_decap_3
XFILLER_13_208 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mem_top_track_8.LATCH_2_.latch/Q
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_0_134 vgnd vgnd scs8hd_fill_2
XFILLER_0_145 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_0_156 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_SLEEPB _144_/Y vgnd vgnd scs8hd_diode_2
Xmem_right_track_0.LATCH_4_.latch vgnd mem_right_track_0.LATCH_4_.latch/Q _080_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_8_201 vgnd vgnd scs8hd_fill_1
XFILLER_8_212 vgnd vgnd scs8hd_fill_2
Xmem_top_track_8.LATCH_4_.latch vgnd vgnd vgnd vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__115__B _114_/X vgnd vgnd scs8hd_diode_2
XANTENNA__131__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_17.INVTX1_2_.scs8hd_inv_1 chany_top_in[7] mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_right_track_16.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_14_32 vgnd vgnd scs8hd_fill_2
XFILLER_14_87 vgnd vgnd scs8hd_fill_2
XFILLER_30_97 vgnd vgnd scs8hd_fill_2
XFILLER_30_75 vgnd vgnd scs8hd_fill_2
XFILLER_30_20 vgnd vgnd scs8hd_decap_3
Xmux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A
+ mem_top_track_16.LATCH_5_.latch/Q mux_top_track_16.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XFILLER_29_193 vgnd vgnd scs8hd_fill_2
XANTENNA__126__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_35_196 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_diode_2
XPHY_64 vgnd vgnd scs8hd_decap_3
XPHY_53 vgnd vgnd scs8hd_decap_3
XFILLER_26_163 vgnd vgnd scs8hd_fill_2
XFILLER_25_53 vgnd vgnd scs8hd_fill_2
XFILLER_25_42 vgnd vgnd scs8hd_fill_2
XPHY_42 vgnd vgnd scs8hd_decap_3
XPHY_20 vgnd vgnd scs8hd_decap_3
XPHY_31 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_16.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vgnd scs8hd_diode_2
Xmux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_left_track_17.LATCH_5_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_25_86 vgnd vgnd scs8hd_fill_2
X_193_ chany_top_in[4] chany_bottom_out[5] vgnd vgnd scs8hd_buf_2
XPHY_86 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_75 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_97 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_17_141 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_23_177 vgnd vgnd scs8hd_decap_4
XFILLER_11_66 vgnd vgnd scs8hd_fill_2
XFILLER_11_77 vgnd vgnd scs8hd_fill_1
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_bottom_track_1.LATCH_4_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_14_100 vgnd vgnd scs8hd_fill_2
XFILLER_14_111 vgnd vgnd scs8hd_fill_2
XFILLER_14_122 vgnd vgnd scs8hd_fill_2
XFILLER_14_166 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.INVTX1_8_.scs8hd_inv_1 chany_bottom_in[1] mux_right_track_0.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_176_ vgnd chanx_left_out[4] vgnd vgnd scs8hd_buf_2
XFILLER_35_6 vgnd vgnd scs8hd_fill_2
XANTENNA__123__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_20_147 vgnd vgnd scs8hd_decap_4
Xmem_bottom_track_9.LATCH_6_.latch vgnd mem_bottom_track_9.LATCH_6_.latch/Q _106_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_20_125 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_22_87 vgnd vgnd scs8hd_fill_2
XFILLER_22_32 vgnd vgnd scs8hd_fill_2
XFILLER_22_10 vgnd vgnd scs8hd_fill_2
XFILLER_7_118 vgnd vgnd scs8hd_fill_2
XFILLER_11_136 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_19_214 vgnd vgnd scs8hd_fill_1
XANTENNA__118__B _114_/X vgnd vgnd scs8hd_diode_2
X_159_ vgnd _159_/B _159_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_140 vgnd vgnd scs8hd_fill_2
XANTENNA__134__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_25_217 vgnd vgnd scs8hd_fill_1
XANTENNA__044__A address[0] vgnd vgnd scs8hd_diode_2
Xmem_left_track_9.LATCH_5_.latch vgnd vgnd vgnd vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_16_228 vgnd vgnd scs8hd_fill_2
XFILLER_17_43 vgnd vgnd scs8hd_fill_2
XPHY_201 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_33_31 vgnd vgnd scs8hd_fill_2
XANTENNA__104__D _086_/D vgnd vgnd scs8hd_diode_2
XFILLER_3_143 vgnd vgnd scs8hd_fill_2
XFILLER_3_176 vgnd vgnd scs8hd_fill_1
XANTENNA__129__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1_A mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_8_224 vgnd vgnd scs8hd_fill_2
XANTENNA__131__B _124_/B vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_3_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_3_.latch/Q mux_left_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_17.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mem_right_track_8.LATCH_6_.latch_SLEEPB _088_/Y vgnd vgnd scs8hd_diode_2
XFILLER_14_22 vgnd vgnd scs8hd_fill_2
XFILLER_30_87 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_5_.scs8hd_inv_1_A chanx_left_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA__126__B _124_/B vgnd vgnd scs8hd_diode_2
XANTENNA__142__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_35_142 vgnd vgnd scs8hd_fill_1
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_8_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_6_.latch/Q mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_top_track_16.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__052__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_5_.scs8hd_inv_1 vgnd _067_/X vgnd vgnd scs8hd_inv_1
XFILLER_18_109 vgnd vgnd scs8hd_fill_2
XPHY_65 vgnd vgnd scs8hd_decap_3
XFILLER_26_197 vgnd vgnd scs8hd_fill_2
XFILLER_26_142 vgnd vgnd scs8hd_fill_2
XPHY_54 vgnd vgnd scs8hd_decap_3
XFILLER_25_65 vgnd vgnd scs8hd_fill_2
XPHY_43 vgnd vgnd scs8hd_decap_3
XPHY_10 vgnd vgnd scs8hd_decap_3
XPHY_87 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_5_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_1_.latch/Q mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_ebufn_2
XPHY_76 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_98 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_21 vgnd vgnd scs8hd_decap_3
XPHY_32 vgnd vgnd scs8hd_decap_3
X_192_ chany_top_in[5] chany_bottom_out[6] vgnd vgnd scs8hd_buf_2
XFILLER_1_230 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_bottom_track_9.INVTX1_0_.scs8hd_inv_1_A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_0_.latch_SLEEPB _112_/Y vgnd vgnd scs8hd_diode_2
XFILLER_17_153 vgnd vgnd scs8hd_fill_2
XANTENNA__137__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_17_197 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB chany_bottom_in[1]
+ vgnd vgnd scs8hd_diode_2
XFILLER_23_134 vgnd vgnd scs8hd_fill_2
XFILLER_23_112 vgnd vgnd scs8hd_fill_2
XANTENNA__047__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_178 vgnd vgnd scs8hd_fill_2
XANTENNA__123__C vgnd vgnd vgnd scs8hd_diode_2
X_175_ chanx_right_in[4] chanx_left_out[5] vgnd vgnd scs8hd_buf_2
XFILLER_28_6 vgnd vgnd scs8hd_fill_2
XFILLER_9_160 vgnd vgnd scs8hd_fill_2
XFILLER_20_104 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_19_226 vgnd vgnd scs8hd_fill_2
X_158_ vgnd _159_/B vgnd vgnd vgnd scs8hd_nor2_4
X_089_ _056_/B _086_/X _089_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_152 vgnd vgnd scs8hd_fill_1
XANTENNA__134__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_10_192 vgnd vgnd scs8hd_fill_2
XANTENNA__150__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_25_229 vgnd vgnd scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_2_.latch_SLEEPB _082_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__060__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_16_207 vgnd vgnd scs8hd_fill_2
XFILLER_17_77 vgnd vgnd scs8hd_fill_2
XPHY_202 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_33_76 vgnd vgnd scs8hd_decap_4
XFILLER_3_155 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__129__B _124_/B vgnd vgnd scs8hd_diode_2
XFILLER_30_232 vgnd vgnd scs8hd_fill_1
XANTENNA__145__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__055__A _055_/A vgnd vgnd scs8hd_diode_2
XFILLER_21_210 vgnd vgnd scs8hd_decap_4
XFILLER_28_32 vgnd vgnd scs8hd_fill_2
XFILLER_28_10 vgnd vgnd scs8hd_fill_2
XFILLER_0_169 vgnd vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_5_.latch vgnd mem_right_track_8.LATCH_5_.latch/Q _089_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_28_76 vgnd vgnd scs8hd_decap_3
Xmux_right_track_0.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _166_/HI mem_right_track_0.LATCH_7_.latch/Q
+ mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XFILLER_12_232 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_3_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
Xmem_left_track_17.LATCH_1_.latch vgnd mem_left_track_17.LATCH_1_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_5_206 vgnd vgnd scs8hd_fill_2
XFILLER_5_217 vgnd vgnd scs8hd_fill_1
XFILLER_14_45 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA__142__B _141_/B vgnd vgnd scs8hd_diode_2
Xmux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2 _167_/HI chany_bottom_in[1]
+ mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XFILLER_35_176 vgnd vgnd scs8hd_decap_4
XFILLER_35_165 vgnd vgnd scs8hd_fill_2
XANTENNA__052__B _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_2_209 vgnd vgnd scs8hd_fill_2
XPHY_66 vgnd vgnd scs8hd_decap_3
XPHY_55 vgnd vgnd scs8hd_decap_3
XFILLER_25_99 vgnd vgnd scs8hd_fill_2
XFILLER_25_11 vgnd vgnd scs8hd_decap_3
XPHY_44 vgnd vgnd scs8hd_decap_3
XPHY_88 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_77 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_11 vgnd vgnd scs8hd_decap_3
XPHY_99 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_22 vgnd vgnd scs8hd_decap_3
XPHY_33 vgnd vgnd scs8hd_decap_3
X_191_ chany_top_in[6] chany_bottom_out[7] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_left_track_1.INVTX1_7_.scs8hd_inv_1_A chany_bottom_in[8] vgnd vgnd scs8hd_diode_2
XFILLER_32_102 vgnd vgnd scs8hd_fill_2
XFILLER_17_176 vgnd vgnd scs8hd_decap_4
XFILLER_32_146 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA__137__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__153__A chany_top_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__063__A address[2] vgnd vgnd scs8hd_diode_2
XFILLER_11_24 vgnd vgnd scs8hd_fill_2
XFILLER_11_35 vgnd vgnd scs8hd_fill_2
XFILLER_11_57 vgnd vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_0_.latch vgnd mem_bottom_track_1.LATCH_0_.latch/Q _103_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__123__D chanx_right_in[2] vgnd vgnd scs8hd_diode_2
X_174_ vgnd chanx_left_out[6] vgnd vgnd scs8hd_buf_2
XANTENNA__148__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_9_194 vgnd vgnd scs8hd_fill_2
XFILLER_28_205 vgnd vgnd scs8hd_decap_8
XANTENNA__058__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_22_23 vgnd vgnd scs8hd_decap_4
XFILLER_11_149 vgnd vgnd scs8hd_fill_2
XFILLER_22_78 vgnd vgnd scs8hd_decap_3
XFILLER_22_56 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_0_.latch_SLEEPB _066_/Y vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_9.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_bottom_track_9.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
X_157_ vgnd _159_/B _157_/Y vgnd vgnd scs8hd_nor2_4
Xmux_left_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[6] _124_/Y vgnd vgnd scs8hd_inv_1
XFILLER_8_69 vgnd vgnd scs8hd_fill_2
XANTENNA__150__B _152_/B vgnd vgnd scs8hd_diode_2
X_088_ _053_/X _086_/X _088_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_186 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__060__B chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XPHY_203 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_33_44 vgnd vgnd scs8hd_fill_2
XFILLER_33_11 vgnd vgnd scs8hd_decap_4
Xmem_right_track_16.LATCH_0_.latch vgnd vgnd _145_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_top_track_16.INVTX1_5_.scs8hd_inv_1 chanx_left_in[1] mux_top_track_16.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_15_230 vgnd vgnd scs8hd_decap_3
XANTENNA__145__B _141_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.tap_buf4_0_.scs8hd_inv_1_A mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_0_92 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__055__B address[1] vgnd vgnd scs8hd_diode_2
XFILLER_21_222 vgnd vgnd scs8hd_fill_2
XANTENNA__071__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.INVTX1_0_.scs8hd_inv_1_A chanx_right_in[0] vgnd vgnd scs8hd_diode_2
XFILLER_28_88 vgnd vgnd scs8hd_fill_2
XFILLER_28_55 vgnd vgnd scs8hd_fill_2
XFILLER_8_204 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_9.LATCH_2_.latch_SLEEPB _129_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A vgnd vgnd vgnd
+ scs8hd_diode_2
XANTENNA__156__A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA__066__A _056_/B vgnd vgnd scs8hd_diode_2
XFILLER_30_45 vgnd vgnd scs8hd_fill_2
XFILLER_5_229 vgnd vgnd scs8hd_fill_2
XFILLER_14_79 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _165_/HI vgnd vgnd
+ scs8hd_diode_2
XFILLER_29_174 vgnd vgnd scs8hd_fill_2
Xmux_top_track_0.INVTX1_1_.scs8hd_inv_1 chanx_right_in[1] mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XPHY_12 vgnd vgnd scs8hd_decap_3
XPHY_67 vgnd vgnd scs8hd_decap_3
XPHY_56 vgnd vgnd scs8hd_decap_3
XPHY_45 vgnd vgnd scs8hd_decap_3
XPHY_89 vgnd vgnd scs8hd_tapvpwrvgnd_1
XPHY_78 vgnd vgnd scs8hd_tapvpwrvgnd_1
X_190_ _190_/A chany_bottom_out[8] vgnd vgnd scs8hd_buf_2
XPHY_23 vgnd vgnd scs8hd_decap_3
XPHY_34 vgnd vgnd scs8hd_decap_3
XFILLER_1_210 vgnd vgnd scs8hd_fill_2
XFILLER_32_136 vgnd vgnd scs8hd_decap_4
XFILLER_32_125 vgnd vgnd scs8hd_fill_2
XFILLER_17_100 vgnd vgnd scs8hd_decap_3
XANTENNA__153__B vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_8.INVTX1_2_.scs8hd_inv_1 chany_top_in[4] mux_right_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_23_169 vgnd vgnd scs8hd_fill_2
XANTENNA__063__B address[1] vgnd vgnd scs8hd_diode_2
X_173_ chanx_right_in[6] chanx_left_out[7] vgnd vgnd scs8hd_buf_2
XFILLER_14_147 vgnd vgnd scs8hd_fill_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_0_.latch/Q mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA__148__B _152_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_4_.latch_SLEEPB _099_/Y vgnd vgnd scs8hd_diode_2
XFILLER_9_184 vgnd vgnd scs8hd_fill_1
XANTENNA__058__B vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__074__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_11_117 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_left_track_9.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_19_217 vgnd vgnd scs8hd_fill_1
XFILLER_34_209 vgnd vgnd scs8hd_decap_4
X_087_ vgnd _086_/X vgnd vgnd vgnd scs8hd_nor2_4
X_156_ chanx_right_in[2] _159_/B _156_/Y vgnd vgnd scs8hd_nor2_4
Xmux_bottom_track_1.INVTX1_7_.scs8hd_inv_1 chanx_left_in[5] mux_bottom_track_1.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[4] mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_6_110 vgnd vgnd scs8hd_fill_2
XFILLER_6_154 vgnd vgnd scs8hd_fill_2
XFILLER_6_165 vgnd vgnd scs8hd_fill_2
XFILLER_8_48 vgnd vgnd scs8hd_fill_2
XANTENNA__159__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__069__A _053_/X vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.INVTX1_6_.scs8hd_inv_1 vgnd mem_top_track_8.LATCH_2_.latch/Q vgnd
+ vgnd scs8hd_inv_1
XPHY_204 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_17_24 vgnd vgnd scs8hd_fill_2
XFILLER_17_35 vgnd vgnd scs8hd_fill_2
XFILLER_17_57 vgnd vgnd scs8hd_fill_2
XFILLER_33_89 vgnd vgnd scs8hd_fill_2
XFILLER_33_56 vgnd vgnd scs8hd_fill_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 _124_/B mem_top_track_8.LATCH_1_.latch/Q
+ mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
XFILLER_3_179 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_139_ vgnd vgnd vgnd _086_/D _141_/B vgnd vgnd scs8hd_or4_4
XANTENNA__055__C _063_/C vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_9_91 vgnd vgnd scs8hd_fill_2
XANTENNA__071__B _067_/X vgnd vgnd scs8hd_diode_2
XFILLER_0_138 vgnd vgnd scs8hd_fill_2
XFILLER_0_149 vgnd vgnd scs8hd_fill_2
XFILLER_28_23 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_1.tap_buf4_0_.scs8hd_inv_1_A mux_left_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XANTENNA__156__B _159_/B vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.INVTX1_8_.scs8hd_inv_1_A chany_bottom_in[1] vgnd vgnd scs8hd_diode_2
XANTENNA__172__A _172_/A vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_2_.scs8hd_inv_1_A chany_top_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA__066__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_14_14 vgnd vgnd scs8hd_fill_2
XFILLER_14_36 vgnd vgnd scs8hd_fill_2
XANTENNA__082__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_30_79 vgnd vgnd scs8hd_fill_2
XFILLER_29_197 vgnd vgnd scs8hd_fill_2
XFILLER_29_153 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_4_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB chany_bottom_in[1]
+ vgnd vgnd scs8hd_diode_2
XFILLER_35_134 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_9.INVTX1_4_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_26_167 vgnd vgnd scs8hd_fill_2
XPHY_46 vgnd vgnd scs8hd_decap_3
XPHY_13 vgnd vgnd scs8hd_decap_3
XPHY_24 vgnd vgnd scs8hd_decap_3
XANTENNA__077__A vgnd vgnd vgnd scs8hd_diode_2
XPHY_35 vgnd vgnd scs8hd_decap_3
XPHY_68 vgnd vgnd scs8hd_decap_3
XPHY_57 vgnd vgnd scs8hd_decap_3
XFILLER_25_57 vgnd vgnd scs8hd_fill_2
XFILLER_25_46 vgnd vgnd scs8hd_fill_2
XPHY_79 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_1_222 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_17_112 vgnd vgnd scs8hd_decap_4
XFILLER_17_123 vgnd vgnd scs8hd_decap_4
XFILLER_17_145 vgnd vgnd scs8hd_decap_3
XANTENNA__153__C vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_5_.latch_SLEEPB _147_/Y vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.INVTX1_5_.scs8hd_inv_1 vgnd mux_right_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_31_170 vgnd vgnd scs8hd_fill_1
XFILLER_23_148 vgnd vgnd scs8hd_fill_2
XFILLER_23_126 vgnd vgnd scs8hd_fill_2
Xmem_top_track_0.LATCH_4_.latch vgnd mem_top_track_0.LATCH_4_.latch/Q _058_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__063__C _063_/C vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_9.LATCH_1_.latch vgnd mem_bottom_track_9.LATCH_1_.latch/Q _111_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_4_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_9.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_14_137 vgnd vgnd scs8hd_fill_2
XFILLER_14_159 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_0.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
X_172_ _172_/A chanx_left_out[8] vgnd vgnd scs8hd_buf_2
XANTENNA_mem_bottom_track_9.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__180__A _180_/A vgnd vgnd scs8hd_diode_2
XANTENNA__074__B _067_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_9.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_left_track_9.LATCH_0_.latch vgnd mem_left_track_9.LATCH_0_.latch/Q _131_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__090__A vgnd vgnd vgnd scs8hd_diode_2
X_086_ vgnd vgnd vgnd _086_/D _086_/X vgnd vgnd scs8hd_or4_4
X_155_ vgnd _159_/B _155_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_144 vgnd vgnd scs8hd_fill_2
XFILLER_10_151 vgnd vgnd scs8hd_fill_2
XFILLER_10_173 vgnd vgnd scs8hd_fill_2
XFILLER_12_91 vgnd vgnd scs8hd_fill_1
XFILLER_33_7 vgnd vgnd scs8hd_fill_2
XFILLER_33_232 vgnd vgnd scs8hd_fill_1
XANTENNA__159__B _159_/B vgnd vgnd scs8hd_diode_2
XANTENNA__175__A chanx_right_in[4] vgnd vgnd scs8hd_diode_2
XANTENNA__069__B _067_/X vgnd vgnd scs8hd_diode_2
XFILLER_24_232 vgnd vgnd scs8hd_fill_1
XANTENNA__085__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_16.LATCH_2_.latch/Q mux_top_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_3_114 vgnd vgnd scs8hd_fill_2
XFILLER_3_147 vgnd vgnd scs8hd_fill_2
Xmem_top_track_16.LATCH_1_.latch vgnd mem_top_track_16.LATCH_1_.latch/Q _137_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_30_224 vgnd vgnd scs8hd_decap_8
XFILLER_30_202 vgnd vgnd scs8hd_decap_12
X_207_ _207_/A chany_top_out[0] vgnd vgnd scs8hd_buf_2
XFILLER_23_90 vgnd vgnd scs8hd_decap_3
X_069_ _053_/X _067_/X _069_/Y vgnd vgnd scs8hd_nor2_4
X_138_ vgnd vgnd _138_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_24_3 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_17.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_16.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_2_.TGATE_1_.scs8hd_ebufn_2 vgnd mem_bottom_track_17.LATCH_1_.latch/Q
+ vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_9_81 vgnd vgnd scs8hd_fill_1
Xmux_left_track_17.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_28_68 vgnd vgnd scs8hd_fill_2
XFILLER_8_228 vgnd vgnd scs8hd_fill_2
XFILLER_12_213 vgnd vgnd scs8hd_fill_1
XFILLER_12_224 vgnd vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_6_.latch vgnd mem_bottom_track_1.LATCH_6_.latch/Q _097_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_right_track_8.LATCH_3_.latch_SLEEPB _091_/Y vgnd vgnd scs8hd_diode_2
XFILLER_10_9 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_TEB mem_bottom_track_17.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_8.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_14_26 vgnd vgnd scs8hd_fill_2
XANTENNA__082__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_30_58 vgnd vgnd scs8hd_fill_2
XFILLER_30_25 vgnd vgnd scs8hd_decap_4
Xmux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_0_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_0_.latch/Q mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_29_132 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.INVTX1_2_.scs8hd_inv_1 chanx_right_in[2] vgnd vgnd vgnd scs8hd_inv_1
Xmem_left_track_1.LATCH_5_.latch vgnd mem_left_track_1.LATCH_5_.latch/Q _117_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_20_91 vgnd vgnd scs8hd_fill_1
Xmux_right_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ mem_right_track_16.LATCH_3_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XANTENNA__183__A chanx_left_in[5] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_6_.latch_SLEEPB _116_/Y vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ mem_top_track_0.LATCH_4_.latch/Q mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.tap_buf4_0_.scs8hd_inv_1 mux_top_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _207_/A vgnd vgnd scs8hd_inv_1
XPHY_69 vgnd vgnd scs8hd_decap_3
XPHY_58 vgnd vgnd scs8hd_decap_3
XFILLER_26_146 vgnd vgnd scs8hd_decap_4
XFILLER_26_102 vgnd vgnd scs8hd_fill_2
XFILLER_25_69 vgnd vgnd scs8hd_fill_2
XFILLER_25_25 vgnd vgnd scs8hd_fill_2
XPHY_47 vgnd vgnd scs8hd_decap_3
XPHY_14 vgnd vgnd scs8hd_decap_3
Xmux_right_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_5_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_1_.latch/Q mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XPHY_25 vgnd vgnd scs8hd_decap_3
XANTENNA__077__B vgnd vgnd vgnd scs8hd_diode_2
XPHY_36 vgnd vgnd scs8hd_decap_3
XANTENNA__093__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_17_157 vgnd vgnd scs8hd_fill_2
XANTENNA__153__D chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_23_138 vgnd vgnd scs8hd_fill_1
XFILLER_23_116 vgnd vgnd scs8hd_fill_2
XANTENNA__178__A chanx_right_in[1] vgnd vgnd scs8hd_diode_2
XFILLER_31_193 vgnd vgnd scs8hd_fill_2
XANTENNA__088__A _053_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_17.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_A mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
X_171_ _171_/HI _171_/LO vgnd vgnd scs8hd_conb_1
Xmem_bottom_track_17.LATCH_1_.latch vgnd mem_bottom_track_17.LATCH_1_.latch/Q _151_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_9_142 vgnd vgnd scs8hd_decap_3
XFILLER_9_164 vgnd vgnd scs8hd_fill_2
XFILLER_9_175 vgnd vgnd scs8hd_fill_2
XFILLER_13_182 vgnd vgnd scs8hd_fill_1
XFILLER_13_193 vgnd vgnd scs8hd_fill_2
XFILLER_20_108 vgnd vgnd scs8hd_fill_2
Xmux_right_track_16.INVTX1_6_.scs8hd_inv_1 vgnd mux_right_track_16.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_17.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[7] mux_left_track_17.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_22_37 vgnd vgnd scs8hd_fill_2
XANTENNA__090__B _086_/X vgnd vgnd scs8hd_diode_2
XFILLER_27_230 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_left_track_17.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_10_130 vgnd vgnd scs8hd_fill_2
X_154_ _056_/B _159_/B _154_/Y vgnd vgnd scs8hd_nor2_4
X_085_ vgnd _045_/Y _086_/D vgnd vgnd scs8hd_nand2_4
XFILLER_6_123 vgnd vgnd scs8hd_fill_2
XFILLER_10_196 vgnd vgnd scs8hd_fill_2
XFILLER_26_7 vgnd vgnd scs8hd_fill_2
Xmux_top_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 vgnd mem_top_track_16.LATCH_0_.latch/Q
+ mux_top_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XFILLER_19_6 vgnd vgnd scs8hd_fill_2
XFILLER_33_222 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 vgnd vgnd mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA__191__A chany_top_in[6] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__085__B _045_/Y vgnd vgnd scs8hd_diode_2
Xmux_left_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_left_track_1.LATCH_0_.latch/Q mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_0.INVTX1_3_.scs8hd_inv_1_A right_top_grid_pin_10_ vgnd vgnd
+ scs8hd_diode_2
XFILLER_3_159 vgnd vgnd scs8hd_fill_2
XFILLER_3_126 vgnd vgnd scs8hd_fill_2
Xmem_right_track_8.LATCH_0_.latch vgnd mem_right_track_8.LATCH_0_.latch/Q _094_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_15_222 vgnd vgnd scs8hd_fill_2
XFILLER_23_80 vgnd vgnd scs8hd_fill_1
X_206_ vgnd chany_top_out[1] vgnd vgnd scs8hd_buf_2
X_137_ vgnd vgnd _137_/Y vgnd vgnd scs8hd_nor2_4
Xmux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2 mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_17.LATCH_0_.latch/Q mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
X_068_ vgnd _067_/X _068_/Y vgnd vgnd scs8hd_nor2_4
Xmux_bottom_track_9.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_bottom_track_9.INVTX1_2_.scs8hd_inv_1/Y
+ mem_bottom_track_9.LATCH_2_.latch/Q mux_bottom_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_17_3 vgnd vgnd scs8hd_decap_4
XFILLER_21_214 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_top_track_8.LATCH_1_.latch_SLEEPB _074_/Y vgnd vgnd scs8hd_diode_2
XFILLER_9_60 vgnd vgnd scs8hd_fill_1
XANTENNA__186__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_4_.latch_SLEEPB _155_/Y vgnd vgnd scs8hd_diode_2
Xmux_left_track_17.tap_buf4_0_.scs8hd_inv_1 vgnd _172_/A vgnd vgnd scs8hd_inv_1
XFILLER_28_36 vgnd vgnd scs8hd_decap_4
XANTENNA_mux_right_track_8.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[3] vgnd vgnd scs8hd_diode_2
XANTENNA__096__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_8_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_6_.latch/Q mux_top_track_8.tap_buf4_0_.scs8hd_inv_1/A vgnd
+ vgnd scs8hd_ebufn_2
Xmux_right_track_16.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_16.LATCH_1_.latch/Q mux_right_track_16.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
Xmux_top_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_5_.scs8hd_inv_1/Y
+ vgnd mux_top_track_0.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_top_track_8.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[2] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_17.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XFILLER_29_166 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _171_/HI vgnd vgnd
+ scs8hd_diode_2
XFILLER_4_232 vgnd vgnd scs8hd_fill_1
XFILLER_35_169 vgnd vgnd scs8hd_fill_2
XFILLER_35_147 vgnd vgnd scs8hd_fill_2
XFILLER_35_103 vgnd vgnd scs8hd_fill_2
Xmux_left_track_9.tap_buf4_0_.scs8hd_inv_1 mux_left_track_9.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd vgnd scs8hd_inv_1
XFILLER_34_180 vgnd vgnd scs8hd_decap_8
XPHY_59 vgnd vgnd scs8hd_decap_3
XFILLER_26_136 vgnd vgnd scs8hd_decap_4
XFILLER_26_125 vgnd vgnd scs8hd_fill_2
XPHY_48 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[7] vgnd vgnd scs8hd_diode_2
XPHY_15 vgnd vgnd scs8hd_decap_3
XPHY_26 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_bottom_track_9.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XPHY_37 vgnd vgnd scs8hd_decap_3
XANTENNA__093__B _086_/X vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_32_106 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_2_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
Xmem_top_track_8.LATCH_5_.latch vgnd mem_top_track_8.LATCH_5_.latch/Q _070_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__194__A _194_/A vgnd vgnd scs8hd_diode_2
Xmem_right_track_0.LATCH_5_.latch vgnd mem_right_track_0.LATCH_5_.latch/Q _079_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd
+ scs8hd_diode_2
XFILLER_11_39 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_9.INVTX1_6_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__088__B _086_/X vgnd vgnd scs8hd_diode_2
XFILLER_22_183 vgnd vgnd scs8hd_fill_1
X_170_ _170_/HI _170_/LO vgnd vgnd scs8hd_conb_1
Xmux_left_track_9.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ mem_left_track_9.LATCH_2_.latch/Q vgnd vgnd vgnd scs8hd_ebufn_2
XFILLER_9_154 vgnd vgnd scs8hd_decap_4
XFILLER_9_198 vgnd vgnd scs8hd_fill_2
XFILLER_13_172 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_9.INVTX1_1_.scs8hd_inv_1 chany_top_in[5] mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_inv_1
XANTENNA__189__A _189_/A vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_11_109 vgnd vgnd scs8hd_fill_2
XFILLER_22_27 vgnd vgnd scs8hd_fill_1
XANTENNA__099__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_3_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_3_.latch/Q mux_right_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
X_153_ chany_top_in[1] vgnd vgnd chanx_right_in[2] _159_/B vgnd vgnd scs8hd_or4_4
XFILLER_6_102 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_A _168_/HI vgnd vgnd
+ scs8hd_diode_2
X_084_ vgnd vgnd _084_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_12_71 vgnd vgnd scs8hd_fill_2
XFILLER_33_212 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_bottom_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[8] vgnd vgnd
+ scs8hd_diode_2
Xmux_top_track_16.INVTX1_2_.scs8hd_inv_1 chanx_right_in[4] mux_top_track_16.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_24_201 vgnd vgnd scs8hd_fill_2
XFILLER_17_49 vgnd vgnd scs8hd_fill_2
XFILLER_33_48 vgnd vgnd scs8hd_fill_2
XFILLER_33_15 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_right_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _167_/HI vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_3_.latch/Q mux_top_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mem_bottom_track_9.LATCH_5_.latch_SLEEPB _107_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_205_ chany_bottom_in[1] chany_top_out[2] vgnd vgnd scs8hd_buf_2
X_136_ vgnd vgnd _136_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB vgnd vgnd vgnd scs8hd_diode_2
X_067_ vgnd vgnd vgnd _067_/D _067_/X vgnd vgnd scs8hd_or4_4
XFILLER_2_182 vgnd vgnd scs8hd_fill_2
XFILLER_21_226 vgnd vgnd scs8hd_fill_2
XANTENNA__096__B vgnd vgnd vgnd scs8hd_diode_2
Xmem_bottom_track_9.LATCH_7_.latch vgnd mem_bottom_track_9.LATCH_7_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_8_208 vgnd vgnd scs8hd_fill_2
XFILLER_34_80 vgnd vgnd scs8hd_fill_2
X_119_ chanx_right_in[2] _114_/X _119_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA__197__A chany_top_in[0] vgnd vgnd scs8hd_diode_2
XFILLER_30_16 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vgnd scs8hd_diode_2
XFILLER_29_178 vgnd vgnd scs8hd_decap_3
XFILLER_29_112 vgnd vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_6_.latch vgnd mem_left_track_9.LATCH_6_.latch/Q _125_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_20_71 vgnd vgnd scs8hd_decap_3
XFILLER_35_115 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_0.LATCH_7_.latch_SLEEPB _077_/Y vgnd vgnd scs8hd_diode_2
XFILLER_6_73 vgnd vgnd scs8hd_fill_2
XFILLER_6_84 vgnd vgnd scs8hd_fill_2
XPHY_49 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_right_track_0.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XPHY_16 vgnd vgnd scs8hd_decap_3
XPHY_27 vgnd vgnd scs8hd_decap_3
XPHY_38 vgnd vgnd scs8hd_decap_3
XANTENNA_mem_bottom_track_1.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_1_214 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ mem_bottom_track_1.LATCH_5_.latch/Q mux_bottom_track_1.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_25_170 vgnd vgnd scs8hd_fill_1
XFILLER_15_71 vgnd vgnd scs8hd_fill_2
XFILLER_31_70 vgnd vgnd scs8hd_fill_2
XFILLER_23_107 vgnd vgnd scs8hd_decap_3
XFILLER_16_170 vgnd vgnd scs8hd_fill_2
XFILLER_16_181 vgnd vgnd scs8hd_decap_3
XFILLER_31_173 vgnd vgnd scs8hd_fill_2
XFILLER_14_107 vgnd vgnd scs8hd_fill_2
XFILLER_14_118 vgnd vgnd scs8hd_fill_2
XFILLER_22_162 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_bottom_track_1.LATCH_1_.latch_SLEEPB _102_/Y vgnd vgnd scs8hd_diode_2
XFILLER_13_140 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_left_track_17.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A _180_/A vgnd vgnd
+ scs8hd_diode_2
XFILLER_3_41 vgnd vgnd scs8hd_fill_1
Xmux_bottom_track_1.INVTX1_4_.scs8hd_inv_1 chanx_right_in[7] mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_left_track_1.INVTX1_1_.scs8hd_inv_1 chany_top_in[3] mux_left_track_1.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_top_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA__099__B vgnd vgnd vgnd scs8hd_diode_2
XFILLER_27_210 vgnd vgnd scs8hd_decap_4
X_152_ vgnd _152_/B _152_/Y vgnd vgnd scs8hd_nor2_4
X_083_ vgnd vgnd _083_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_10_143 vgnd vgnd scs8hd_fill_2
XFILLER_10_154 vgnd vgnd scs8hd_fill_2
Xmux_top_track_8.INVTX1_3_.scs8hd_inv_1 chanx_right_in[8] mux_top_track_8.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_12_50 vgnd vgnd scs8hd_fill_2
XFILLER_6_169 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_8.INVTX1_0_.scs8hd_inv_1_A chany_top_in[0] vgnd vgnd scs8hd_diode_2
XFILLER_12_83 vgnd vgnd scs8hd_fill_2
XFILLER_18_232 vgnd vgnd scs8hd_fill_1
XFILLER_5_191 vgnd vgnd scs8hd_fill_2
XFILLER_24_224 vgnd vgnd scs8hd_decap_8
XFILLER_24_213 vgnd vgnd scs8hd_fill_1
XANTENNA_mem_top_track_16.LATCH_3_.latch_SLEEPB _135_/Y vgnd vgnd scs8hd_diode_2
XFILLER_17_39 vgnd vgnd scs8hd_fill_2
XFILLER_33_27 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_right_track_16.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_16.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_204_ vgnd chany_top_out[3] vgnd vgnd scs8hd_buf_2
XFILLER_15_213 vgnd vgnd scs8hd_fill_2
X_066_ _056_/B vgnd _066_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_23_71 vgnd vgnd scs8hd_decap_3
X_135_ chanx_right_in[2] vgnd _135_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mem_top_track_0.LATCH_0_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_2_194 vgnd vgnd scs8hd_fill_2
XFILLER_2_150 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_left_track_17.INVTX1_4_.scs8hd_inv_1_A chanx_right_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_9_73 vgnd vgnd scs8hd_fill_2
XFILLER_9_95 vgnd vgnd scs8hd_fill_2
XFILLER_28_27 vgnd vgnd scs8hd_fill_2
XFILLER_12_205 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_93 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_6_.scs8hd_inv_1_A chanx_left_in[5] vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_049_ _055_/A _043_/Y _063_/C vgnd vgnd vgnd scs8hd_or3_4
X_118_ vgnd _114_/X _118_/Y vgnd vgnd scs8hd_nor2_4
Xmux_bottom_track_9.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2 _162_/HI mem_bottom_track_9.LATCH_7_.latch/Q
+ mux_bottom_track_9.tap_buf4_0_.scs8hd_inv_1/A vgnd vgnd scs8hd_ebufn_2
XFILLER_14_18 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2 vgnd mem_bottom_track_1.LATCH_2_.latch/Q
+ mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_3_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_16.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_top_track_0.LATCH_5_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.INVTX1_6_.scs8hd_inv_1 chany_bottom_in[3] mux_left_track_9.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mux_bottom_track_9.INVTX1_1_.scs8hd_inv_1_A chany_top_in[5] vgnd vgnd scs8hd_diode_2
XFILLER_20_83 vgnd vgnd scs8hd_fill_2
XFILLER_29_92 vgnd vgnd scs8hd_fill_2
XFILLER_35_138 vgnd vgnd scs8hd_decap_4
XANTENNA_mem_bottom_track_9.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_6_63 vgnd vgnd scs8hd_fill_1
XPHY_17 vgnd vgnd scs8hd_decap_3
XPHY_28 vgnd vgnd scs8hd_decap_3
XPHY_39 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_3_.scs8hd_ebufn_2_TEB mem_left_track_1.LATCH_7_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_17.LATCH_2_.latch_SLEEPB _150_/Y vgnd vgnd scs8hd_diode_2
Xmux_right_track_0.INVTX1_2_.scs8hd_inv_1 chany_top_in[8] mux_right_track_0.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_1_226 vgnd vgnd scs8hd_fill_2
XFILLER_32_119 vgnd vgnd scs8hd_decap_4
XFILLER_25_193 vgnd vgnd scs8hd_fill_2
XFILLER_17_127 vgnd vgnd scs8hd_fill_1
XFILLER_31_60 vgnd vgnd scs8hd_fill_1
XFILLER_15_83 vgnd vgnd scs8hd_decap_4
Xmem_right_track_8.LATCH_6_.latch vgnd mem_right_track_8.LATCH_6_.latch/Q _088_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_top_track_16.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mux_top_track_16.INVTX1_1_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_22_196 vgnd vgnd scs8hd_decap_4
XFILLER_22_141 vgnd vgnd scs8hd_fill_1
Xmem_left_track_17.LATCH_2_.latch vgnd vgnd _157_/Y vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mem_left_track_9.LATCH_7_.latch_SLEEPB _124_/Y vgnd vgnd scs8hd_diode_2
XFILLER_26_71 vgnd vgnd scs8hd_fill_2
XFILLER_26_60 vgnd vgnd scs8hd_fill_2
XFILLER_9_134 vgnd vgnd scs8hd_fill_2
XFILLER_27_222 vgnd vgnd scs8hd_fill_2
XFILLER_10_100 vgnd vgnd scs8hd_fill_2
X_082_ vgnd vgnd _082_/Y vgnd vgnd scs8hd_nor2_4
X_151_ vgnd _152_/B _151_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_148 vgnd vgnd scs8hd_fill_2
XFILLER_10_177 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.mux_l1_in_2_.TGATE_2_.scs8hd_ebufn_2_A _170_/HI vgnd vgnd
+ scs8hd_diode_2
Xmux_top_track_0.INVTX1_6_.scs8hd_inv_1 vgnd mux_top_track_0.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XANTENNA_mem_top_track_8.LATCH_4_.latch_D vgnd vgnd vgnd scs8hd_diode_2
Xmux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_bottom_track_17.INVTX1_3_.scs8hd_inv_1/Y
+ mem_bottom_track_17.LATCH_0_.latch/Q mux_bottom_track_17.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_3_107 vgnd vgnd scs8hd_fill_2
XFILLER_3_118 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_bottom_track_9.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
X_203_ _203_/A chany_top_out[4] vgnd vgnd scs8hd_buf_2
XANTENNA_mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_2_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
X_065_ address[2] address[1] address[0] vgnd vgnd vgnd scs8hd_or3_4
X_134_ vgnd vgnd _134_/Y vgnd vgnd scs8hd_nor2_4
Xmux_right_track_8.INVTX1_7_.scs8hd_inv_1 chanx_left_in[1] mux_right_track_8.INVTX1_7_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_24_7 vgnd vgnd scs8hd_fill_2
Xmem_bottom_track_1.LATCH_1_.latch vgnd mem_bottom_track_1.LATCH_1_.latch/Q _102_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_21_217 vgnd vgnd scs8hd_fill_1
XFILLER_9_52 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_8.LATCH_0_.latch_SLEEPB _094_/Y vgnd vgnd scs8hd_diode_2
XFILLER_12_228 vgnd vgnd scs8hd_fill_2
XFILLER_18_50 vgnd vgnd scs8hd_fill_2
XFILLER_18_72 vgnd vgnd scs8hd_decap_3
X_117_ _056_/B _114_/X _117_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA_mux_left_track_17.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_left_track_17.LATCH_0_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_7_210 vgnd vgnd scs8hd_decap_4
XFILLER_7_221 vgnd vgnd scs8hd_fill_2
X_048_ enable vgnd vgnd vgnd scs8hd_inv_8
Xmem_left_track_1.LATCH_0_.latch vgnd mem_left_track_1.LATCH_0_.latch/Q _122_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
Xmux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ mem_right_track_8.LATCH_0_.latch/Q mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_29_136 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_left_track_1.LATCH_3_.latch_SLEEPB _119_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_top_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_right_track_0.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_right_track_8.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_8.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_left_track_1.INVTX1_8_.scs8hd_inv_1_A left_top_grid_pin_10_ vgnd vgnd
+ scs8hd_diode_2
XANTENNA_mux_right_track_0.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_2_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_4_224 vgnd vgnd scs8hd_fill_2
XFILLER_4_213 vgnd vgnd scs8hd_fill_1
XFILLER_29_71 vgnd vgnd scs8hd_fill_2
XFILLER_28_180 vgnd vgnd scs8hd_decap_4
Xmem_right_track_16.LATCH_1_.latch vgnd mem_right_track_16.LATCH_1_.latch/Q _144_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_1.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_8_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_34_150 vgnd vgnd scs8hd_fill_1
XFILLER_26_106 vgnd vgnd scs8hd_fill_2
XFILLER_25_29 vgnd vgnd scs8hd_fill_2
XPHY_18 vgnd vgnd scs8hd_decap_3
XPHY_29 vgnd vgnd scs8hd_decap_3
XANTENNA_mux_left_track_17.mux_l1_in_2_.TGATE_0_.scs8hd_ebufn_2_A mux_left_track_17.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_15_51 vgnd vgnd scs8hd_fill_2
XFILLER_31_83 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_right_track_16.LATCH_3_.latch_SLEEPB _142_/Y vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_8.mux_l2_in_0_.TGATE_2_.scs8hd_ebufn_2_TEB mem_top_track_8.LATCH_6_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA__102__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_31_197 vgnd vgnd scs8hd_fill_2
XFILLER_31_153 vgnd vgnd scs8hd_fill_2
XFILLER_22_186 vgnd vgnd scs8hd_fill_1
Xmux_left_track_17.INVTX1_4_.scs8hd_inv_1 chanx_right_in[6] mux_left_track_17.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
Xmux_right_track_16.INVTX1_3_.scs8hd_inv_1 vgnd mux_right_track_16.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_inv_1
XFILLER_13_197 vgnd vgnd scs8hd_fill_2
XFILLER_9_179 vgnd vgnd scs8hd_fill_2
X_150_ vgnd _152_/B _150_/Y vgnd vgnd scs8hd_nor2_4
X_081_ chanx_right_in[2] vgnd _081_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_127 vgnd vgnd scs8hd_fill_2
XFILLER_12_30 vgnd vgnd scs8hd_fill_1
XANTENNA_mux_right_track_8.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2_A mux_right_track_8.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_33_226 vgnd vgnd scs8hd_decap_6
XFILLER_33_204 vgnd vgnd scs8hd_fill_2
XFILLER_18_212 vgnd vgnd scs8hd_fill_2
XFILLER_5_160 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_16.INVTX1_1_.scs8hd_inv_1_A chanx_right_in[3] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_17.LATCH_1_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA__200__A chany_bottom_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_15_204 vgnd vgnd scs8hd_fill_2
XFILLER_15_226 vgnd vgnd scs8hd_fill_2
XFILLER_23_95 vgnd vgnd scs8hd_decap_3
X_133_ _056_/B vgnd vgnd vgnd vgnd scs8hd_nor2_4
X_202_ chany_bottom_in[4] chany_top_out[5] vgnd vgnd scs8hd_buf_2
X_064_ _056_/B vgnd vgnd vgnd vgnd scs8hd_nor2_4
XFILLER_2_163 vgnd vgnd scs8hd_fill_2
Xmux_right_track_16.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_16.INVTX1_0_.scs8hd_inv_1/Y
+ vgnd mux_right_track_16.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2/Z vgnd vgnd scs8hd_ebufn_2
XANTENNA__110__A vgnd vgnd vgnd scs8hd_diode_2
Xmux_top_track_0.mux_l1_in_0_.TGATE_0_.scs8hd_ebufn_2 mux_top_track_0.INVTX1_0_.scs8hd_inv_1/Y
+ mem_top_track_0.LATCH_0_.latch/Q mux_top_track_0.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_bottom_track_1.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_bottom_track_1.LATCH_4_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_34_50 vgnd vgnd scs8hd_fill_2
XFILLER_18_84 vgnd vgnd scs8hd_fill_2
X_116_ _053_/X _114_/X _116_/Y vgnd vgnd scs8hd_nor2_4
XANTENNA__105__A vgnd vgnd vgnd scs8hd_diode_2
X_047_ vgnd vgnd vgnd vgnd scs8hd_inv_8
XANTENNA_mem_right_track_8.LATCH_5_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_1.LATCH_7_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_35_107 vgnd vgnd scs8hd_decap_3
XFILLER_6_32 vgnd vgnd scs8hd_fill_1
XPHY_19 vgnd vgnd scs8hd_decap_3
Xmem_right_track_0.LATCH_0_.latch vgnd mem_right_track_0.LATCH_0_.latch/Q _084_/Y
+ vgnd vgnd scs8hd_lpflow_inputisolatch_1
Xmem_top_track_8.LATCH_0_.latch vgnd mem_top_track_8.LATCH_0_.latch/Q _056_/B vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2_TEB mem_right_track_0.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_17_118 vgnd vgnd scs8hd_fill_2
XFILLER_25_173 vgnd vgnd scs8hd_fill_2
XFILLER_15_30 vgnd vgnd scs8hd_decap_4
XFILLER_31_40 vgnd vgnd scs8hd_fill_2
XANTENNA__102__B vgnd vgnd vgnd scs8hd_diode_2
Xmux_left_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2 _124_/Y mem_left_track_9.LATCH_1_.latch/Q
+ mux_left_track_9.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2/A vgnd vgnd scs8hd_ebufn_2
XPHY_190 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_31_132 vgnd vgnd scs8hd_fill_2
XFILLER_22_154 vgnd vgnd scs8hd_fill_2
XANTENNA__203__A _203_/A vgnd vgnd scs8hd_diode_2
XFILLER_26_84 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2_TEB mem_top_track_0.LATCH_5_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XANTENNA_mux_top_track_16.mux_l2_in_0_.TGATE_0_.scs8hd_ebufn_2_TEB mem_top_track_16.LATCH_3_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_9_114 vgnd vgnd scs8hd_fill_2
XFILLER_13_121 vgnd vgnd scs8hd_fill_1
XFILLER_13_132 vgnd vgnd scs8hd_fill_1
XFILLER_13_176 vgnd vgnd scs8hd_decap_4
XFILLER_3_22 vgnd vgnd scs8hd_fill_1
XANTENNA__113__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mux_bottom_track_1.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2_A mux_bottom_track_1.INVTX1_4_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
Xmux_top_track_8.mux_l1_in_0_.TGATE_2_.scs8hd_ebufn_2 mux_top_track_8.INVTX1_2_.scs8hd_inv_1/Y
+ mem_top_track_8.LATCH_2_.latch/Q mux_top_track_8.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
X_080_ vgnd vgnd _080_/Y vgnd vgnd scs8hd_nor2_4
XFILLER_6_106 vgnd vgnd scs8hd_fill_2
Xmux_bottom_track_17.INVTX1_7_.scs8hd_inv_1 chany_bottom_in[1] vgnd vgnd vgnd scs8hd_inv_1
XFILLER_12_97 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.tap_buf4_0_.scs8hd_inv_1 mux_right_track_0.tap_buf4_0_.scs8hd_inv_1/A
+ _189_/A vgnd vgnd scs8hd_inv_1
XANTENNA_mux_left_track_1.mux_l1_in_1_.TGATE_2_.scs8hd_ebufn_2_A mux_left_track_1.INVTX1_6_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_18_224 vgnd vgnd scs8hd_fill_2
XANTENNA__108__A vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_9.LATCH_2_.latch_SLEEPB vgnd vgnd vgnd scs8hd_diode_2
XANTENNA_mem_left_track_9.LATCH_1_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_24_205 vgnd vgnd scs8hd_fill_2
X_063_ address[2] address[1] _063_/C vgnd vgnd vgnd scs8hd_or3_4
X_201_ vgnd chany_top_out[6] vgnd vgnd scs8hd_buf_2
X_132_ chany_top_in[1] vgnd vgnd _067_/D vgnd vgnd vgnd scs8hd_or4_4
Xmem_top_track_0.LATCH_5_.latch vgnd mem_top_track_0.LATCH_5_.latch/Q vgnd vgnd vgnd
+ scs8hd_lpflow_inputisolatch_1
XFILLER_2_186 vgnd vgnd scs8hd_fill_2
XFILLER_2_142 vgnd vgnd scs8hd_fill_2
Xmem_bottom_track_9.LATCH_2_.latch vgnd mem_bottom_track_9.LATCH_2_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA__110__B _110_/B vgnd vgnd scs8hd_diode_2
Xmux_right_track_16.tap_buf4_0_.scs8hd_inv_1 vgnd _181_/A vgnd vgnd scs8hd_inv_1
XANTENNA_mux_left_track_1.INVTX1_3_.scs8hd_inv_1_A chanx_right_in[0] vgnd vgnd scs8hd_diode_2
XANTENNA_mem_bottom_track_1.LATCH_3_.latch_D vgnd vgnd vgnd scs8hd_diode_2
XFILLER_18_30 vgnd vgnd scs8hd_fill_1
XFILLER_18_41 vgnd vgnd scs8hd_decap_3
XFILLER_34_84 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_0.INVTX1_5_.scs8hd_inv_1_A chany_bottom_in[4] vgnd vgnd scs8hd_diode_2
X_115_ vgnd _114_/X _115_/Y vgnd vgnd scs8hd_nor2_4
X_046_ vgnd chany_top_in[1] vgnd vgnd scs8hd_inv_8
XANTENNA__105__B _110_/B vgnd vgnd scs8hd_diode_2
XANTENNA__121__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_22_6 vgnd vgnd scs8hd_fill_2
Xmem_left_track_9.LATCH_1_.latch vgnd mem_left_track_9.LATCH_1_.latch/Q _130_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XANTENNA_mux_left_track_9.INVTX1_5_.scs8hd_inv_1_A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_29_149 vgnd vgnd scs8hd_fill_2
XFILLER_29_116 vgnd vgnd scs8hd_decap_4
XANTENNA_mem_right_track_0.LATCH_4_.latch_SLEEPB _080_/Y vgnd vgnd scs8hd_diode_2
XANTENNA__206__A vgnd vgnd vgnd scs8hd_diode_2
XFILLER_20_20 vgnd vgnd scs8hd_fill_2
XFILLER_20_42 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_top_track_8.INVTX1_7_.scs8hd_inv_1_A chanx_left_in[6] vgnd vgnd scs8hd_diode_2
XFILLER_35_119 vgnd vgnd scs8hd_decap_3
XANTENNA__116__A _053_/X vgnd vgnd scs8hd_diode_2
XFILLER_6_77 vgnd vgnd scs8hd_fill_2
XFILLER_6_88 vgnd vgnd scs8hd_fill_2
XANTENNA_mux_bottom_track_9.mux_l1_in_0_.TGATE_1_.scs8hd_ebufn_2_A mem_bottom_track_9.LATCH_1_.latch/Q
+ vgnd vgnd scs8hd_diode_2
XFILLER_26_119 vgnd vgnd scs8hd_decap_4
Xmem_top_track_16.LATCH_2_.latch vgnd mem_top_track_16.LATCH_2_.latch/Q _136_/Y vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
XFILLER_20_3 vgnd vgnd scs8hd_fill_2
XFILLER_34_163 vgnd vgnd scs8hd_decap_8
XFILLER_19_193 vgnd vgnd scs8hd_fill_2
Xmux_right_track_8.mux_l2_in_0_.TGATE_1_.scs8hd_ebufn_2 mux_right_track_8.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2/Z
+ mem_right_track_8.LATCH_5_.latch/Q mux_right_track_8.tap_buf4_0_.scs8hd_inv_1/A
+ vgnd vgnd scs8hd_ebufn_2
XANTENNA_mux_left_track_9.mux_l1_in_0_.TGATE_3_.scs8hd_ebufn_2_A mux_left_track_9.INVTX1_3_.scs8hd_inv_1/Y
+ vgnd vgnd scs8hd_diode_2
XFILLER_15_75 vgnd vgnd scs8hd_fill_2
XFILLER_31_52 vgnd vgnd scs8hd_fill_2
Xmux_right_track_0.mux_l1_in_1_.TGATE_0_.scs8hd_ebufn_2 mux_right_track_0.INVTX1_4_.scs8hd_inv_1/Y
+ mem_right_track_0.LATCH_0_.latch/Q mux_right_track_0.mux_l1_in_1_.TGATE_1_.scs8hd_ebufn_2/Z
+ vgnd vgnd scs8hd_ebufn_2
XFILLER_31_100 vgnd vgnd scs8hd_fill_2
XANTENNA_mem_top_track_8.LATCH_6_.latch_SLEEPB _069_/Y vgnd vgnd scs8hd_diode_2
XFILLER_16_152 vgnd vgnd scs8hd_fill_1
XFILLER_16_174 vgnd vgnd scs8hd_fill_2
XPHY_191 vgnd vgnd scs8hd_tapvpwrvgnd_1
XFILLER_31_177 vgnd vgnd scs8hd_decap_4
XFILLER_31_166 vgnd vgnd scs8hd_decap_4
XPHY_180 vgnd vgnd scs8hd_tapvpwrvgnd_1
Xmem_bottom_track_1.LATCH_7_.latch vgnd mem_bottom_track_1.LATCH_7_.latch/Q vgnd vgnd
+ vgnd scs8hd_lpflow_inputisolatch_1
.ends

