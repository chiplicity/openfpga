magic
tech sky130A
magscale 1 2
timestamp 1604667756
<< locali >>
rect 7849 14807 7883 14909
rect 3249 12223 3283 12325
rect 26617 11543 26651 11713
<< viali >>
rect 12357 21097 12391 21131
rect 17509 21097 17543 21131
rect 12173 20961 12207 20995
rect 17325 20961 17359 20995
rect 18245 20961 18279 20995
rect 18705 20961 18739 20995
rect 18797 20893 18831 20927
rect 18889 20893 18923 20927
rect 4997 20757 5031 20791
rect 12725 20757 12759 20791
rect 18337 20757 18371 20791
rect 20177 20757 20211 20791
rect 1593 20553 1627 20587
rect 2605 20553 2639 20587
rect 7297 20553 7331 20587
rect 9505 20553 9539 20587
rect 14657 20553 14691 20587
rect 16957 20553 16991 20587
rect 18613 20553 18647 20587
rect 24317 20553 24351 20587
rect 26617 20553 26651 20587
rect 11345 20485 11379 20519
rect 12449 20485 12483 20519
rect 17509 20485 17543 20519
rect 19625 20485 19659 20519
rect 25421 20485 25455 20519
rect 5365 20417 5399 20451
rect 5457 20417 5491 20451
rect 12909 20417 12943 20451
rect 13001 20417 13035 20451
rect 17877 20417 17911 20451
rect 19165 20417 19199 20451
rect 20637 20417 20671 20451
rect 20729 20417 20763 20451
rect 1409 20349 1443 20383
rect 2421 20349 2455 20383
rect 2881 20349 2915 20383
rect 4813 20349 4847 20383
rect 7113 20349 7147 20383
rect 9321 20349 9355 20383
rect 12265 20349 12299 20383
rect 14473 20349 14507 20383
rect 14933 20349 14967 20383
rect 16773 20349 16807 20383
rect 24133 20349 24167 20383
rect 25237 20349 25271 20383
rect 26433 20349 26467 20383
rect 26893 20349 26927 20383
rect 5273 20281 5307 20315
rect 12817 20281 12851 20315
rect 13461 20281 13495 20315
rect 19073 20281 19107 20315
rect 19993 20281 20027 20315
rect 20545 20281 20579 20315
rect 1961 20213 1995 20247
rect 4353 20213 4387 20247
rect 4905 20213 4939 20247
rect 7573 20213 7607 20247
rect 9781 20213 9815 20247
rect 11713 20213 11747 20247
rect 16589 20213 16623 20247
rect 18521 20213 18555 20247
rect 18981 20213 19015 20247
rect 20177 20213 20211 20247
rect 24685 20213 24719 20247
rect 25789 20213 25823 20247
rect 4445 20009 4479 20043
rect 5273 20009 5307 20043
rect 5641 20009 5675 20043
rect 11621 20009 11655 20043
rect 16773 20009 16807 20043
rect 17325 20009 17359 20043
rect 17693 20009 17727 20043
rect 18889 20009 18923 20043
rect 21097 20009 21131 20043
rect 22109 20009 22143 20043
rect 11989 19941 12023 19975
rect 4261 19873 4295 19907
rect 11529 19873 11563 19907
rect 12081 19873 12115 19907
rect 15669 19873 15703 19907
rect 15761 19873 15795 19907
rect 17785 19873 17819 19907
rect 19257 19873 19291 19907
rect 20545 19873 20579 19907
rect 20913 19873 20947 19907
rect 21925 19873 21959 19907
rect 5733 19805 5767 19839
rect 5825 19805 5859 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 15853 19805 15887 19839
rect 17877 19805 17911 19839
rect 19349 19805 19383 19839
rect 19533 19805 19567 19839
rect 26525 19805 26559 19839
rect 27077 19805 27111 19839
rect 3525 19669 3559 19703
rect 5089 19669 5123 19703
rect 10885 19669 10919 19703
rect 14933 19669 14967 19703
rect 15301 19669 15335 19703
rect 18613 19669 18647 19703
rect 20177 19669 20211 19703
rect 6009 19465 6043 19499
rect 13829 19465 13863 19499
rect 16681 19465 16715 19499
rect 3341 19329 3375 19363
rect 3985 19329 4019 19363
rect 5549 19329 5583 19363
rect 6377 19329 6411 19363
rect 11345 19329 11379 19363
rect 11805 19329 11839 19363
rect 15485 19329 15519 19363
rect 27629 19329 27663 19363
rect 2973 19261 3007 19295
rect 3801 19261 3835 19295
rect 4537 19261 4571 19295
rect 10701 19261 10735 19295
rect 11253 19261 11287 19295
rect 12449 19261 12483 19295
rect 12705 19261 12739 19295
rect 14841 19261 14875 19295
rect 15301 19261 15335 19295
rect 17049 19261 17083 19295
rect 18889 19261 18923 19295
rect 19349 19261 19383 19295
rect 19605 19261 19639 19295
rect 21833 19261 21867 19295
rect 24593 19261 24627 19295
rect 27445 19261 27479 19295
rect 4905 19193 4939 19227
rect 5365 19193 5399 19227
rect 10333 19193 10367 19227
rect 11161 19193 11195 19227
rect 14473 19193 14507 19227
rect 17417 19193 17451 19227
rect 21281 19193 21315 19227
rect 24838 19193 24872 19227
rect 27537 19193 27571 19227
rect 1685 19125 1719 19159
rect 1961 19125 1995 19159
rect 3433 19125 3467 19159
rect 3893 19125 3927 19159
rect 4997 19125 5031 19159
rect 5457 19125 5491 19159
rect 6837 19125 6871 19159
rect 10793 19125 10827 19159
rect 12173 19125 12207 19159
rect 14933 19125 14967 19159
rect 15393 19125 15427 19159
rect 15945 19125 15979 19159
rect 17785 19125 17819 19159
rect 18337 19125 18371 19159
rect 19165 19125 19199 19159
rect 20729 19125 20763 19159
rect 22293 19125 22327 19159
rect 24409 19125 24443 19159
rect 25973 19125 26007 19159
rect 26525 19125 26559 19159
rect 26893 19125 26927 19159
rect 27077 19125 27111 19159
rect 2697 18921 2731 18955
rect 3893 18921 3927 18955
rect 4721 18921 4755 18955
rect 6193 18921 6227 18955
rect 7297 18921 7331 18955
rect 7757 18921 7791 18955
rect 9873 18921 9907 18955
rect 13645 18921 13679 18955
rect 14657 18921 14691 18955
rect 15117 18921 15151 18955
rect 15577 18921 15611 18955
rect 18889 18921 18923 18955
rect 18981 18921 19015 18955
rect 20361 18921 20395 18955
rect 24777 18921 24811 18955
rect 5058 18853 5092 18887
rect 18521 18853 18555 18887
rect 1409 18785 1443 18819
rect 2053 18785 2087 18819
rect 2513 18785 2547 18819
rect 2973 18785 3007 18819
rect 7665 18785 7699 18819
rect 9689 18785 9723 18819
rect 11428 18785 11462 18819
rect 14013 18785 14047 18819
rect 16764 18785 16798 18819
rect 19349 18785 19383 18819
rect 19441 18785 19475 18819
rect 21916 18785 21950 18819
rect 25145 18785 25179 18819
rect 26157 18785 26191 18819
rect 26893 18785 26927 18819
rect 26985 18785 27019 18819
rect 4813 18717 4847 18751
rect 7849 18717 7883 18751
rect 11161 18717 11195 18751
rect 14105 18717 14139 18751
rect 14197 18717 14231 18751
rect 16497 18717 16531 18751
rect 19533 18717 19567 18751
rect 21649 18717 21683 18751
rect 25237 18717 25271 18751
rect 25421 18717 25455 18751
rect 27077 18717 27111 18751
rect 1593 18649 1627 18683
rect 8677 18649 8711 18683
rect 12541 18649 12575 18683
rect 13553 18649 13587 18683
rect 19993 18649 20027 18683
rect 24225 18649 24259 18683
rect 26525 18649 26559 18683
rect 2329 18581 2363 18615
rect 3433 18581 3467 18615
rect 4353 18581 4387 18615
rect 6929 18581 6963 18615
rect 8953 18581 8987 18615
rect 10793 18581 10827 18615
rect 17877 18581 17911 18615
rect 23029 18581 23063 18615
rect 24685 18581 24719 18615
rect 25789 18581 25823 18615
rect 3341 18377 3375 18411
rect 4905 18377 4939 18411
rect 10609 18377 10643 18411
rect 10793 18377 10827 18411
rect 12449 18377 12483 18411
rect 18061 18377 18095 18411
rect 19441 18377 19475 18411
rect 19625 18377 19659 18411
rect 23121 18377 23155 18411
rect 25145 18377 25179 18411
rect 27077 18377 27111 18411
rect 27629 18377 27663 18411
rect 6837 18309 6871 18343
rect 8585 18309 8619 18343
rect 16957 18309 16991 18343
rect 17877 18309 17911 18343
rect 21189 18309 21223 18343
rect 24133 18309 24167 18343
rect 2053 18241 2087 18275
rect 2237 18241 2271 18275
rect 3893 18241 3927 18275
rect 5549 18241 5583 18275
rect 5917 18241 5951 18275
rect 7389 18241 7423 18275
rect 9137 18241 9171 18275
rect 10333 18241 10367 18275
rect 11437 18241 11471 18275
rect 13093 18241 13127 18275
rect 17509 18241 17543 18275
rect 18521 18241 18555 18275
rect 18613 18241 18647 18275
rect 20177 18241 20211 18275
rect 22201 18241 22235 18275
rect 22385 18241 22419 18275
rect 24041 18241 24075 18275
rect 24777 18241 24811 18275
rect 1961 18173 1995 18207
rect 3709 18173 3743 18207
rect 5365 18173 5399 18207
rect 7205 18173 7239 18207
rect 9689 18173 9723 18207
rect 11161 18173 11195 18207
rect 14013 18173 14047 18207
rect 14280 18173 14314 18207
rect 18429 18173 18463 18207
rect 19993 18173 20027 18207
rect 20637 18173 20671 18207
rect 22109 18173 22143 18207
rect 22753 18173 22787 18207
rect 25697 18173 25731 18207
rect 25964 18173 25998 18207
rect 4445 18105 4479 18139
rect 7849 18105 7883 18139
rect 8953 18105 8987 18139
rect 11897 18105 11931 18139
rect 12909 18105 12943 18139
rect 16497 18105 16531 18139
rect 19073 18105 19107 18139
rect 21649 18105 21683 18139
rect 27997 18105 28031 18139
rect 1593 18037 1627 18071
rect 2697 18037 2731 18071
rect 3249 18037 3283 18071
rect 3801 18037 3835 18071
rect 4813 18037 4847 18071
rect 5273 18037 5307 18071
rect 6561 18037 6595 18071
rect 7297 18037 7331 18071
rect 8493 18037 8527 18071
rect 9045 18037 9079 18071
rect 11253 18037 11287 18071
rect 12173 18037 12207 18071
rect 12817 18037 12851 18071
rect 13645 18037 13679 18071
rect 15393 18037 15427 18071
rect 20085 18037 20119 18071
rect 21741 18037 21775 18071
rect 24501 18037 24535 18071
rect 24593 18037 24627 18071
rect 25513 18037 25547 18071
rect 1685 17833 1719 17867
rect 2697 17833 2731 17867
rect 3433 17833 3467 17867
rect 4353 17833 4387 17867
rect 4813 17833 4847 17867
rect 6377 17833 6411 17867
rect 7665 17833 7699 17867
rect 10885 17833 10919 17867
rect 12909 17833 12943 17867
rect 13645 17833 13679 17867
rect 14013 17833 14047 17867
rect 15301 17833 15335 17867
rect 18061 17833 18095 17867
rect 19165 17833 19199 17867
rect 20177 17833 20211 17867
rect 21005 17833 21039 17867
rect 22385 17833 22419 17867
rect 25237 17833 25271 17867
rect 25697 17833 25731 17867
rect 26341 17833 26375 17867
rect 26525 17833 26559 17867
rect 5242 17765 5276 17799
rect 6929 17765 6963 17799
rect 7389 17765 7423 17799
rect 10425 17765 10459 17799
rect 13553 17765 13587 17799
rect 14657 17765 14691 17799
rect 21465 17765 21499 17799
rect 2053 17697 2087 17731
rect 4997 17697 5031 17731
rect 8401 17697 8435 17731
rect 11805 17697 11839 17731
rect 14105 17697 14139 17731
rect 16681 17697 16715 17731
rect 16948 17697 16982 17731
rect 19533 17697 19567 17731
rect 20729 17697 20763 17731
rect 21373 17697 21407 17731
rect 22569 17697 22603 17731
rect 22836 17697 22870 17731
rect 26893 17697 26927 17731
rect 2145 17629 2179 17663
rect 2329 17629 2363 17663
rect 8493 17629 8527 17663
rect 8677 17629 8711 17663
rect 11897 17629 11931 17663
rect 11989 17629 12023 17663
rect 14197 17629 14231 17663
rect 19625 17629 19659 17663
rect 19717 17629 19751 17663
rect 21649 17629 21683 17663
rect 26985 17629 27019 17663
rect 27169 17629 27203 17663
rect 11345 17561 11379 17595
rect 24593 17561 24627 17595
rect 3801 17493 3835 17527
rect 8033 17493 8067 17527
rect 9965 17493 9999 17527
rect 11437 17493 11471 17527
rect 12541 17493 12575 17527
rect 18797 17493 18831 17527
rect 22109 17493 22143 17527
rect 23949 17493 23983 17527
rect 24869 17493 24903 17527
rect 3709 17289 3743 17323
rect 5641 17289 5675 17323
rect 6193 17289 6227 17323
rect 7665 17289 7699 17323
rect 10609 17289 10643 17323
rect 12173 17289 12207 17323
rect 12449 17289 12483 17323
rect 13461 17289 13495 17323
rect 13921 17289 13955 17323
rect 16497 17289 16531 17323
rect 17417 17289 17451 17323
rect 17785 17289 17819 17323
rect 18245 17289 18279 17323
rect 20177 17289 20211 17323
rect 21097 17289 21131 17323
rect 23029 17289 23063 17323
rect 23397 17289 23431 17323
rect 23949 17289 23983 17323
rect 24133 17289 24167 17323
rect 27997 17289 28031 17323
rect 3157 17221 3191 17255
rect 7573 17221 7607 17255
rect 14933 17221 14967 17255
rect 25513 17221 25547 17255
rect 27629 17221 27663 17255
rect 8217 17153 8251 17187
rect 13093 17153 13127 17187
rect 15117 17153 15151 17187
rect 17049 17153 17083 17187
rect 21557 17153 21591 17187
rect 22661 17153 22695 17187
rect 24777 17153 24811 17187
rect 25697 17153 25731 17187
rect 1777 17085 1811 17119
rect 2044 17085 2078 17119
rect 4261 17085 4295 17119
rect 4517 17085 4551 17119
rect 6653 17085 6687 17119
rect 8033 17085 8067 17119
rect 8125 17085 8159 17119
rect 9229 17085 9263 17119
rect 9485 17085 9519 17119
rect 18797 17085 18831 17119
rect 19053 17085 19087 17119
rect 24501 17085 24535 17119
rect 4169 17017 4203 17051
rect 7205 17017 7239 17051
rect 12909 17017 12943 17051
rect 14197 17017 14231 17051
rect 15362 17017 15396 17051
rect 22477 17017 22511 17051
rect 25942 17017 25976 17051
rect 1685 16949 1719 16983
rect 8677 16949 8711 16983
rect 9045 16949 9079 16983
rect 11529 16949 11563 16983
rect 11897 16949 11931 16983
rect 12817 16949 12851 16983
rect 14565 16949 14599 16983
rect 18613 16949 18647 16983
rect 21833 16949 21867 16983
rect 22017 16949 22051 16983
rect 22385 16949 22419 16983
rect 24593 16949 24627 16983
rect 25145 16949 25179 16983
rect 27077 16949 27111 16983
rect 2881 16745 2915 16779
rect 4997 16745 5031 16779
rect 7941 16745 7975 16779
rect 8033 16745 8067 16779
rect 9229 16745 9263 16779
rect 9689 16745 9723 16779
rect 10149 16745 10183 16779
rect 12817 16745 12851 16779
rect 13553 16745 13587 16779
rect 14289 16745 14323 16779
rect 16681 16745 16715 16779
rect 18521 16745 18555 16779
rect 20729 16745 20763 16779
rect 22569 16745 22603 16779
rect 25329 16745 25363 16779
rect 25881 16745 25915 16779
rect 26985 16745 27019 16779
rect 1768 16677 1802 16711
rect 3801 16677 3835 16711
rect 5426 16677 5460 16711
rect 7205 16677 7239 16711
rect 10057 16677 10091 16711
rect 15117 16677 15151 16711
rect 15568 16677 15602 16711
rect 18981 16677 19015 16711
rect 1501 16609 1535 16643
rect 5181 16609 5215 16643
rect 7573 16609 7607 16643
rect 8401 16609 8435 16643
rect 8493 16609 8527 16643
rect 10793 16609 10827 16643
rect 11437 16609 11471 16643
rect 11704 16609 11738 16643
rect 13829 16609 13863 16643
rect 18889 16609 18923 16643
rect 19533 16609 19567 16643
rect 21189 16609 21223 16643
rect 21445 16609 21479 16643
rect 24216 16609 24250 16643
rect 26893 16609 26927 16643
rect 4077 16541 4111 16575
rect 8677 16541 8711 16575
rect 10333 16541 10367 16575
rect 15301 16541 15335 16575
rect 19073 16541 19107 16575
rect 23949 16541 23983 16575
rect 27169 16541 27203 16575
rect 26525 16473 26559 16507
rect 3525 16405 3559 16439
rect 4629 16405 4663 16439
rect 6561 16405 6595 16439
rect 11253 16405 11287 16439
rect 18153 16405 18187 16439
rect 26341 16405 26375 16439
rect 3065 16201 3099 16235
rect 3985 16201 4019 16235
rect 4169 16201 4203 16235
rect 5181 16201 5215 16235
rect 5549 16201 5583 16235
rect 8125 16201 8159 16235
rect 9689 16201 9723 16235
rect 10793 16201 10827 16235
rect 12173 16201 12207 16235
rect 15025 16201 15059 16235
rect 17509 16201 17543 16235
rect 19993 16201 20027 16235
rect 21189 16201 21223 16235
rect 21465 16201 21499 16235
rect 23121 16201 23155 16235
rect 23397 16201 23431 16235
rect 24409 16201 24443 16235
rect 24593 16201 24627 16235
rect 25973 16201 26007 16235
rect 28089 16201 28123 16235
rect 3617 16133 3651 16167
rect 13461 16133 13495 16167
rect 16037 16133 16071 16167
rect 20913 16133 20947 16167
rect 4721 16065 4755 16099
rect 7297 16065 7331 16099
rect 11437 16065 11471 16099
rect 13001 16065 13035 16099
rect 14105 16065 14139 16099
rect 14565 16065 14599 16099
rect 15669 16065 15703 16099
rect 18061 16065 18095 16099
rect 22017 16065 22051 16099
rect 22569 16065 22603 16099
rect 25053 16065 25087 16099
rect 25237 16065 25271 16099
rect 26157 16065 26191 16099
rect 1685 15997 1719 16031
rect 8309 15997 8343 16031
rect 11161 15997 11195 16031
rect 13829 15997 13863 16031
rect 18317 15997 18351 16031
rect 20545 15997 20579 16031
rect 21833 15997 21867 16031
rect 24133 15997 24167 16031
rect 24961 15997 24995 16031
rect 1952 15929 1986 15963
rect 4537 15929 4571 15963
rect 5917 15929 5951 15963
rect 8576 15929 8610 15963
rect 26424 15929 26458 15963
rect 4629 15861 4663 15895
rect 7205 15861 7239 15895
rect 10333 15861 10367 15895
rect 10609 15861 10643 15895
rect 11253 15861 11287 15895
rect 11897 15861 11931 15895
rect 13369 15861 13403 15895
rect 13921 15861 13955 15895
rect 14933 15861 14967 15895
rect 15393 15861 15427 15895
rect 15485 15861 15519 15895
rect 17785 15861 17819 15895
rect 19441 15861 19475 15895
rect 21925 15861 21959 15895
rect 25605 15861 25639 15895
rect 27537 15861 27571 15895
rect 2053 15657 2087 15691
rect 2421 15657 2455 15691
rect 3525 15657 3559 15691
rect 3801 15657 3835 15691
rect 6745 15657 6779 15691
rect 8033 15657 8067 15691
rect 8401 15657 8435 15691
rect 10333 15657 10367 15691
rect 10701 15657 10735 15691
rect 13277 15657 13311 15691
rect 14749 15657 14783 15691
rect 16681 15657 16715 15691
rect 18061 15657 18095 15691
rect 21189 15657 21223 15691
rect 22201 15657 22235 15691
rect 22753 15657 22787 15691
rect 23213 15657 23247 15691
rect 24225 15657 24259 15691
rect 24869 15657 24903 15691
rect 27629 15657 27663 15691
rect 5610 15589 5644 15623
rect 9505 15589 9539 15623
rect 15546 15589 15580 15623
rect 20729 15589 20763 15623
rect 21649 15589 21683 15623
rect 24777 15589 24811 15623
rect 25237 15589 25271 15623
rect 4077 15521 4111 15555
rect 5365 15521 5399 15555
rect 12153 15521 12187 15555
rect 15301 15521 15335 15555
rect 18337 15521 18371 15555
rect 18604 15521 18638 15555
rect 21557 15521 21591 15555
rect 23121 15521 23155 15555
rect 25329 15521 25363 15555
rect 26893 15521 26927 15555
rect 2513 15453 2547 15487
rect 2697 15453 2731 15487
rect 3157 15453 3191 15487
rect 8493 15453 8527 15487
rect 8677 15453 8711 15487
rect 10793 15453 10827 15487
rect 10885 15453 10919 15487
rect 11897 15453 11931 15487
rect 21741 15453 21775 15487
rect 23305 15453 23339 15487
rect 25421 15453 25455 15487
rect 26985 15453 27019 15487
rect 27169 15453 27203 15487
rect 7941 15385 7975 15419
rect 10241 15385 10275 15419
rect 23949 15385 23983 15419
rect 26249 15385 26283 15419
rect 1685 15317 1719 15351
rect 4261 15317 4295 15351
rect 4629 15317 4663 15351
rect 5273 15317 5307 15351
rect 9045 15317 9079 15351
rect 11437 15317 11471 15351
rect 11805 15317 11839 15351
rect 13829 15317 13863 15351
rect 15117 15317 15151 15351
rect 19717 15317 19751 15351
rect 26525 15317 26559 15351
rect 2053 15113 2087 15147
rect 3617 15113 3651 15147
rect 7941 15113 7975 15147
rect 9505 15113 9539 15147
rect 12633 15113 12667 15147
rect 13093 15113 13127 15147
rect 18429 15113 18463 15147
rect 19533 15113 19567 15147
rect 21005 15113 21039 15147
rect 22477 15113 22511 15147
rect 23489 15113 23523 15147
rect 24133 15113 24167 15147
rect 28089 15113 28123 15147
rect 14657 15045 14691 15079
rect 16037 15045 16071 15079
rect 27721 15045 27755 15079
rect 2697 14977 2731 15011
rect 4169 14977 4203 15011
rect 5825 14977 5859 15011
rect 6561 14977 6595 15011
rect 10425 14977 10459 15011
rect 11345 14977 11379 15011
rect 13737 14977 13771 15011
rect 15117 14977 15151 15011
rect 15209 14977 15243 15011
rect 16773 14977 16807 15011
rect 19441 14977 19475 15011
rect 20085 14977 20119 15011
rect 21104 14977 21138 15011
rect 24225 14977 24259 15011
rect 27261 14977 27295 15011
rect 3065 14909 3099 14943
rect 4077 14909 4111 14943
rect 5089 14909 5123 14943
rect 5641 14909 5675 14943
rect 7849 14909 7883 14943
rect 8125 14909 8159 14943
rect 8392 14909 8426 14943
rect 11161 14909 11195 14943
rect 13461 14909 13495 14943
rect 16681 14909 16715 14943
rect 26249 14909 26283 14943
rect 27169 14909 27203 14943
rect 28457 14909 28491 14943
rect 3525 14841 3559 14875
rect 3985 14841 4019 14875
rect 5549 14841 5583 14875
rect 7665 14841 7699 14875
rect 11897 14841 11931 14875
rect 14105 14841 14139 14875
rect 16589 14841 16623 14875
rect 18705 14841 18739 14875
rect 21342 14841 21376 14875
rect 24492 14841 24526 14875
rect 26617 14841 26651 14875
rect 1961 14773 1995 14807
rect 2421 14773 2455 14807
rect 2513 14773 2547 14807
rect 4721 14773 4755 14807
rect 5181 14773 5215 14807
rect 6193 14773 6227 14807
rect 7205 14773 7239 14807
rect 7849 14773 7883 14807
rect 10793 14773 10827 14807
rect 11253 14773 11287 14807
rect 13553 14773 13587 14807
rect 14473 14773 14507 14807
rect 15025 14773 15059 14807
rect 15669 14773 15703 14807
rect 16221 14773 16255 14807
rect 19901 14773 19935 14807
rect 19993 14773 20027 14807
rect 20545 14773 20579 14807
rect 23121 14773 23155 14807
rect 25605 14773 25639 14807
rect 26709 14773 26743 14807
rect 27077 14773 27111 14807
rect 1869 14569 1903 14603
rect 3249 14569 3283 14603
rect 3617 14569 3651 14603
rect 5273 14569 5307 14603
rect 7573 14569 7607 14603
rect 7941 14569 7975 14603
rect 8493 14569 8527 14603
rect 9137 14569 9171 14603
rect 10149 14569 10183 14603
rect 12725 14569 12759 14603
rect 13737 14569 13771 14603
rect 15301 14569 15335 14603
rect 15761 14569 15795 14603
rect 20361 14569 20395 14603
rect 21281 14569 21315 14603
rect 26525 14569 26559 14603
rect 11590 14501 11624 14535
rect 14289 14501 14323 14535
rect 14749 14501 14783 14535
rect 15669 14501 15703 14535
rect 17408 14501 17442 14535
rect 20729 14501 20763 14535
rect 24216 14501 24250 14535
rect 2237 14433 2271 14467
rect 4077 14433 4111 14467
rect 5549 14433 5583 14467
rect 5816 14433 5850 14467
rect 8401 14433 8435 14467
rect 10885 14433 10919 14467
rect 11345 14433 11379 14467
rect 15117 14433 15151 14467
rect 16313 14433 16347 14467
rect 21649 14433 21683 14467
rect 22293 14433 22327 14467
rect 23949 14433 23983 14467
rect 26893 14433 26927 14467
rect 2329 14365 2363 14399
rect 2513 14365 2547 14399
rect 2973 14365 3007 14399
rect 8677 14365 8711 14399
rect 10241 14365 10275 14399
rect 10425 14365 10459 14399
rect 13829 14365 13863 14399
rect 15853 14365 15887 14399
rect 17141 14365 17175 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 22753 14365 22787 14399
rect 22937 14365 22971 14399
rect 26985 14365 27019 14399
rect 27169 14365 27203 14399
rect 9781 14297 9815 14331
rect 19901 14297 19935 14331
rect 1777 14229 1811 14263
rect 4261 14229 4295 14263
rect 4813 14229 4847 14263
rect 6929 14229 6963 14263
rect 8033 14229 8067 14263
rect 9505 14229 9539 14263
rect 11253 14229 11287 14263
rect 13277 14229 13311 14263
rect 18521 14229 18555 14263
rect 19165 14229 19199 14263
rect 19625 14229 19659 14263
rect 21189 14229 21223 14263
rect 23489 14229 23523 14263
rect 23857 14229 23891 14263
rect 25329 14229 25363 14263
rect 27537 14229 27571 14263
rect 3617 14025 3651 14059
rect 4169 14025 4203 14059
rect 4721 14025 4755 14059
rect 5733 14025 5767 14059
rect 6561 14025 6595 14059
rect 8125 14025 8159 14059
rect 8953 14025 8987 14059
rect 11253 14025 11287 14059
rect 13829 14025 13863 14059
rect 14473 14025 14507 14059
rect 14749 14025 14783 14059
rect 15945 14025 15979 14059
rect 16313 14025 16347 14059
rect 17509 14025 17543 14059
rect 23857 14025 23891 14059
rect 24041 14025 24075 14059
rect 25145 14025 25179 14059
rect 27537 14025 27571 14059
rect 14933 13957 14967 13991
rect 19533 13957 19567 13991
rect 20637 13957 20671 13991
rect 20913 13957 20947 13991
rect 22477 13957 22511 13991
rect 23121 13957 23155 13991
rect 23489 13957 23523 13991
rect 28273 13957 28307 13991
rect 5273 13889 5307 13923
rect 7389 13889 7423 13923
rect 15393 13889 15427 13923
rect 15485 13889 15519 13923
rect 19441 13889 19475 13923
rect 20177 13889 20211 13923
rect 24501 13889 24535 13923
rect 24593 13889 24627 13923
rect 25605 13889 25639 13923
rect 27905 13889 27939 13923
rect 2237 13821 2271 13855
rect 4629 13821 4663 13855
rect 5181 13821 5215 13855
rect 7297 13821 7331 13855
rect 9229 13821 9263 13855
rect 9873 13821 9907 13855
rect 10140 13821 10174 13855
rect 12449 13821 12483 13855
rect 19073 13821 19107 13855
rect 19993 13821 20027 13855
rect 21097 13821 21131 13855
rect 24409 13821 24443 13855
rect 25861 13821 25895 13855
rect 2504 13753 2538 13787
rect 5089 13753 5123 13787
rect 11805 13753 11839 13787
rect 12173 13753 12207 13787
rect 12716 13753 12750 13787
rect 21364 13753 21398 13787
rect 25421 13753 25455 13787
rect 1961 13685 1995 13719
rect 6193 13685 6227 13719
rect 6837 13685 6871 13719
rect 7205 13685 7239 13719
rect 8401 13685 8435 13719
rect 9689 13685 9723 13719
rect 15301 13685 15335 13719
rect 17141 13685 17175 13719
rect 18245 13685 18279 13719
rect 19901 13685 19935 13719
rect 26985 13685 27019 13719
rect 4813 13481 4847 13515
rect 5641 13481 5675 13515
rect 5733 13481 5767 13515
rect 9137 13481 9171 13515
rect 9965 13481 9999 13515
rect 11345 13481 11379 13515
rect 11805 13481 11839 13515
rect 12265 13481 12299 13515
rect 12909 13481 12943 13515
rect 15853 13481 15887 13515
rect 19257 13481 19291 13515
rect 21465 13481 21499 13515
rect 24225 13481 24259 13515
rect 25881 13481 25915 13515
rect 3801 13413 3835 13447
rect 5181 13413 5215 13447
rect 7358 13413 7392 13447
rect 9505 13413 9539 13447
rect 13277 13413 13311 13447
rect 14013 13413 14047 13447
rect 1501 13345 1535 13379
rect 1768 13345 1802 13379
rect 4077 13345 4111 13379
rect 6377 13345 6411 13379
rect 10333 13345 10367 13379
rect 12173 13345 12207 13379
rect 14105 13345 14139 13379
rect 16589 13345 16623 13379
rect 16856 13345 16890 13379
rect 19625 13345 19659 13379
rect 20729 13345 20763 13379
rect 21833 13345 21867 13379
rect 24133 13345 24167 13379
rect 25329 13345 25363 13379
rect 26893 13345 26927 13379
rect 3525 13277 3559 13311
rect 5825 13277 5859 13311
rect 7113 13277 7147 13311
rect 10425 13277 10459 13311
rect 10609 13277 10643 13311
rect 12357 13277 12391 13311
rect 14289 13277 14323 13311
rect 19717 13277 19751 13311
rect 19809 13277 19843 13311
rect 20361 13277 20395 13311
rect 21925 13277 21959 13311
rect 22017 13277 22051 13311
rect 24317 13277 24351 13311
rect 26985 13277 27019 13311
rect 27077 13277 27111 13311
rect 2881 13209 2915 13243
rect 13645 13209 13679 13243
rect 15485 13209 15519 13243
rect 4261 13141 4295 13175
rect 5273 13141 5307 13175
rect 6929 13141 6963 13175
rect 8493 13141 8527 13175
rect 15025 13141 15059 13175
rect 16497 13141 16531 13175
rect 17969 13141 18003 13175
rect 21097 13141 21131 13175
rect 23305 13141 23339 13175
rect 23581 13141 23615 13175
rect 23765 13141 23799 13175
rect 24869 13141 24903 13175
rect 25145 13141 25179 13175
rect 25513 13141 25547 13175
rect 26341 13141 26375 13175
rect 26525 13141 26559 13175
rect 3065 12937 3099 12971
rect 4169 12937 4203 12971
rect 4997 12937 5031 12971
rect 6193 12937 6227 12971
rect 7849 12937 7883 12971
rect 8217 12937 8251 12971
rect 10701 12937 10735 12971
rect 11529 12937 11563 12971
rect 12449 12937 12483 12971
rect 13645 12937 13679 12971
rect 14105 12937 14139 12971
rect 16405 12937 16439 12971
rect 18613 12937 18647 12971
rect 22385 12937 22419 12971
rect 23029 12937 23063 12971
rect 23949 12937 23983 12971
rect 24961 12937 24995 12971
rect 25329 12937 25363 12971
rect 25973 12937 26007 12971
rect 6561 12869 6595 12903
rect 11069 12869 11103 12903
rect 11897 12869 11931 12903
rect 19441 12869 19475 12903
rect 20821 12869 20855 12903
rect 23489 12869 23523 12903
rect 28181 12869 28215 12903
rect 4629 12801 4663 12835
rect 5549 12801 5583 12835
rect 5733 12801 5767 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 8401 12801 8435 12835
rect 10425 12801 10459 12835
rect 13093 12801 13127 12835
rect 15301 12801 15335 12835
rect 15485 12801 15519 12835
rect 16865 12801 16899 12835
rect 17049 12801 17083 12835
rect 19993 12801 20027 12835
rect 24409 12801 24443 12835
rect 24593 12801 24627 12835
rect 26157 12801 26191 12835
rect 1685 12733 1719 12767
rect 5457 12733 5491 12767
rect 7205 12733 7239 12767
rect 8657 12733 8691 12767
rect 12817 12733 12851 12767
rect 16313 12733 16347 12767
rect 21005 12733 21039 12767
rect 24317 12733 24351 12767
rect 1952 12665 1986 12699
rect 12173 12665 12207 12699
rect 12909 12665 12943 12699
rect 16773 12665 16807 12699
rect 17785 12665 17819 12699
rect 19809 12665 19843 12699
rect 21272 12665 21306 12699
rect 26402 12665 26436 12699
rect 3709 12597 3743 12631
rect 5089 12597 5123 12631
rect 6837 12597 6871 12631
rect 9781 12597 9815 12631
rect 14473 12597 14507 12631
rect 14841 12597 14875 12631
rect 15209 12597 15243 12631
rect 15853 12597 15887 12631
rect 17417 12597 17451 12631
rect 18981 12597 19015 12631
rect 19349 12597 19383 12631
rect 19901 12597 19935 12631
rect 20453 12597 20487 12631
rect 27537 12597 27571 12631
rect 1685 12393 1719 12427
rect 1961 12393 1995 12427
rect 4537 12393 4571 12427
rect 5365 12393 5399 12427
rect 7021 12393 7055 12427
rect 8033 12393 8067 12427
rect 12909 12393 12943 12427
rect 15577 12393 15611 12427
rect 16681 12393 16715 12427
rect 19533 12393 19567 12427
rect 26157 12393 26191 12427
rect 26985 12393 27019 12427
rect 27537 12393 27571 12427
rect 3249 12325 3283 12359
rect 3525 12325 3559 12359
rect 5886 12325 5920 12359
rect 10302 12325 10336 12359
rect 2789 12257 2823 12291
rect 4445 12257 4479 12291
rect 13001 12257 13035 12291
rect 15945 12257 15979 12291
rect 17408 12257 17442 12291
rect 21169 12257 21203 12291
rect 23305 12257 23339 12291
rect 23664 12257 23698 12291
rect 25881 12257 25915 12291
rect 26893 12257 26927 12291
rect 2881 12189 2915 12223
rect 3065 12189 3099 12223
rect 3249 12189 3283 12223
rect 4721 12189 4755 12223
rect 5641 12189 5675 12223
rect 10057 12189 10091 12223
rect 13093 12189 13127 12223
rect 16037 12189 16071 12223
rect 16221 12189 16255 12223
rect 17141 12189 17175 12223
rect 19809 12189 19843 12223
rect 20913 12189 20947 12223
rect 23397 12189 23431 12223
rect 27169 12189 27203 12223
rect 7665 12121 7699 12155
rect 13645 12121 13679 12155
rect 14933 12121 14967 12155
rect 2421 12053 2455 12087
rect 3893 12053 3927 12087
rect 4077 12053 4111 12087
rect 8401 12053 8435 12087
rect 8769 12053 8803 12087
rect 11437 12053 11471 12087
rect 11989 12053 12023 12087
rect 12541 12053 12575 12087
rect 14565 12053 14599 12087
rect 17049 12053 17083 12087
rect 18521 12053 18555 12087
rect 20269 12053 20303 12087
rect 20637 12053 20671 12087
rect 22293 12053 22327 12087
rect 24777 12053 24811 12087
rect 25421 12053 25455 12087
rect 26525 12053 26559 12087
rect 2145 11849 2179 11883
rect 6653 11849 6687 11883
rect 7481 11849 7515 11883
rect 9781 11849 9815 11883
rect 10241 11849 10275 11883
rect 14841 11849 14875 11883
rect 21465 11849 21499 11883
rect 23029 11849 23063 11883
rect 25421 11849 25455 11883
rect 26801 11849 26835 11883
rect 4353 11781 4387 11815
rect 11897 11781 11931 11815
rect 12725 11781 12759 11815
rect 20637 11781 20671 11815
rect 23489 11781 23523 11815
rect 27997 11781 28031 11815
rect 1685 11713 1719 11747
rect 2329 11713 2363 11747
rect 5825 11713 5859 11747
rect 8585 11713 8619 11747
rect 8953 11713 8987 11747
rect 9413 11713 9447 11747
rect 10793 11713 10827 11747
rect 12265 11713 12299 11747
rect 13737 11713 13771 11747
rect 13921 11713 13955 11747
rect 15485 11713 15519 11747
rect 17049 11713 17083 11747
rect 17509 11713 17543 11747
rect 22109 11713 22143 11747
rect 22477 11713 22511 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 24961 11713 24995 11747
rect 25237 11713 25271 11747
rect 25881 11713 25915 11747
rect 25973 11713 26007 11747
rect 26617 11713 26651 11747
rect 27445 11713 27479 11747
rect 27537 11713 27571 11747
rect 6837 11645 6871 11679
rect 8309 11645 8343 11679
rect 10149 11645 10183 11679
rect 10609 11645 10643 11679
rect 13185 11645 13219 11679
rect 13645 11645 13679 11679
rect 14749 11645 14783 11679
rect 15209 11645 15243 11679
rect 15853 11645 15887 11679
rect 16773 11645 16807 11679
rect 17877 11645 17911 11679
rect 18153 11645 18187 11679
rect 18420 11645 18454 11679
rect 21005 11645 21039 11679
rect 21833 11645 21867 11679
rect 24225 11645 24259 11679
rect 2596 11577 2630 11611
rect 5089 11577 5123 11611
rect 7849 11577 7883 11611
rect 14381 11577 14415 11611
rect 16865 11577 16899 11611
rect 25789 11577 25823 11611
rect 27353 11577 27387 11611
rect 3709 11509 3743 11543
rect 4721 11509 4755 11543
rect 5181 11509 5215 11543
rect 5549 11509 5583 11543
rect 5641 11509 5675 11543
rect 6285 11509 6319 11543
rect 7021 11509 7055 11543
rect 7941 11509 7975 11543
rect 8401 11509 8435 11543
rect 10701 11509 10735 11543
rect 11253 11509 11287 11543
rect 13277 11509 13311 11543
rect 15301 11509 15335 11543
rect 16221 11509 16255 11543
rect 16405 11509 16439 11543
rect 19533 11509 19567 11543
rect 20177 11509 20211 11543
rect 21281 11509 21315 11543
rect 21925 11509 21959 11543
rect 23857 11509 23891 11543
rect 26433 11509 26467 11543
rect 26617 11509 26651 11543
rect 26985 11509 27019 11543
rect 2145 11305 2179 11339
rect 2789 11305 2823 11339
rect 3525 11305 3559 11339
rect 4629 11305 4663 11339
rect 6377 11305 6411 11339
rect 6929 11305 6963 11339
rect 7297 11305 7331 11339
rect 7941 11305 7975 11339
rect 8493 11305 8527 11339
rect 8861 11305 8895 11339
rect 11805 11305 11839 11339
rect 12173 11305 12207 11339
rect 13277 11305 13311 11339
rect 16129 11305 16163 11339
rect 16589 11305 16623 11339
rect 17233 11305 17267 11339
rect 18153 11305 18187 11339
rect 18705 11305 18739 11339
rect 19257 11305 19291 11339
rect 20913 11305 20947 11339
rect 23673 11305 23707 11339
rect 24869 11305 24903 11339
rect 25237 11305 25271 11339
rect 26525 11305 26559 11339
rect 26893 11305 26927 11339
rect 26985 11305 27019 11339
rect 27537 11305 27571 11339
rect 4353 11237 4387 11271
rect 10149 11237 10183 11271
rect 14933 11237 14967 11271
rect 15669 11237 15703 11271
rect 18061 11237 18095 11271
rect 24041 11237 24075 11271
rect 2881 11169 2915 11203
rect 5264 11169 5298 11203
rect 7849 11169 7883 11203
rect 10609 11169 10643 11203
rect 16497 11169 16531 11203
rect 19625 11169 19659 11203
rect 20729 11169 20763 11203
rect 21281 11169 21315 11203
rect 21373 11169 21407 11203
rect 22569 11169 22603 11203
rect 25329 11169 25363 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 4997 11101 5031 11135
rect 8125 11101 8159 11135
rect 10701 11101 10735 11135
rect 10885 11101 10919 11135
rect 12265 11101 12299 11135
rect 12357 11101 12391 11135
rect 16681 11101 16715 11135
rect 18337 11101 18371 11135
rect 19717 11101 19751 11135
rect 19809 11101 19843 11135
rect 21465 11101 21499 11135
rect 24133 11101 24167 11135
rect 24317 11101 24351 11135
rect 27077 11101 27111 11135
rect 2421 11033 2455 11067
rect 10241 11033 10275 11067
rect 16037 11033 16071 11067
rect 17693 11033 17727 11067
rect 19073 11033 19107 11067
rect 22753 11033 22787 11067
rect 25513 11033 25547 11067
rect 3893 10965 3927 10999
rect 7481 10965 7515 10999
rect 21925 10965 21959 10999
rect 23489 10965 23523 10999
rect 26249 10965 26283 10999
rect 3157 10761 3191 10795
rect 3617 10761 3651 10795
rect 5181 10761 5215 10795
rect 7297 10761 7331 10795
rect 8677 10761 8711 10795
rect 10149 10761 10183 10795
rect 10333 10761 10367 10795
rect 11437 10761 11471 10795
rect 11897 10761 11931 10795
rect 12173 10761 12207 10795
rect 12633 10761 12667 10795
rect 16405 10761 16439 10795
rect 17785 10761 17819 10795
rect 18981 10761 19015 10795
rect 19349 10761 19383 10795
rect 21465 10761 21499 10795
rect 22937 10761 22971 10795
rect 26157 10761 26191 10795
rect 27261 10761 27295 10795
rect 27629 10761 27663 10795
rect 4997 10693 5031 10727
rect 8309 10693 8343 10727
rect 15209 10693 15243 10727
rect 15577 10693 15611 10727
rect 25053 10693 25087 10727
rect 2513 10625 2547 10659
rect 2697 10625 2731 10659
rect 3525 10625 3559 10659
rect 4261 10625 4295 10659
rect 5641 10625 5675 10659
rect 5825 10625 5859 10659
rect 7205 10625 7239 10659
rect 7849 10625 7883 10659
rect 10977 10625 11011 10659
rect 17049 10625 17083 10659
rect 19441 10625 19475 10659
rect 22477 10625 22511 10659
rect 25973 10625 26007 10659
rect 26709 10625 26743 10659
rect 1961 10557 1995 10591
rect 2421 10557 2455 10591
rect 3985 10557 4019 10591
rect 7757 10557 7791 10591
rect 8861 10557 8895 10591
rect 9413 10557 9447 10591
rect 9781 10557 9815 10591
rect 10701 10557 10735 10591
rect 16313 10557 16347 10591
rect 16865 10557 16899 10591
rect 21833 10557 21867 10591
rect 22293 10557 22327 10591
rect 22385 10557 22419 10591
rect 23673 10557 23707 10591
rect 23940 10557 23974 10591
rect 25605 10557 25639 10591
rect 26525 10557 26559 10591
rect 4721 10489 4755 10523
rect 15945 10489 15979 10523
rect 16773 10489 16807 10523
rect 19708 10489 19742 10523
rect 23489 10489 23523 10523
rect 2053 10421 2087 10455
rect 4077 10421 4111 10455
rect 5549 10421 5583 10455
rect 6285 10421 6319 10455
rect 6561 10421 6595 10455
rect 7665 10421 7699 10455
rect 9045 10421 9079 10455
rect 10793 10421 10827 10455
rect 18337 10421 18371 10455
rect 20821 10421 20855 10455
rect 21925 10421 21959 10455
rect 26617 10421 26651 10455
rect 2421 10217 2455 10251
rect 2513 10217 2547 10251
rect 3065 10217 3099 10251
rect 5457 10217 5491 10251
rect 7021 10217 7055 10251
rect 8033 10217 8067 10251
rect 10333 10217 10367 10251
rect 11161 10217 11195 10251
rect 15761 10217 15795 10251
rect 16221 10217 16255 10251
rect 17693 10217 17727 10251
rect 18797 10217 18831 10251
rect 19257 10217 19291 10251
rect 19717 10217 19751 10251
rect 20361 10217 20395 10251
rect 20913 10217 20947 10251
rect 21373 10217 21407 10251
rect 23489 10217 23523 10251
rect 23581 10217 23615 10251
rect 24409 10217 24443 10251
rect 24593 10217 24627 10251
rect 25053 10217 25087 10251
rect 9045 10149 9079 10183
rect 20729 10149 20763 10183
rect 23121 10149 23155 10183
rect 24041 10149 24075 10183
rect 4344 10081 4378 10115
rect 6929 10081 6963 10115
rect 8125 10081 8159 10115
rect 10793 10081 10827 10115
rect 16865 10081 16899 10115
rect 19625 10081 19659 10115
rect 21281 10081 21315 10115
rect 24961 10081 24995 10115
rect 26525 10081 26559 10115
rect 2605 10013 2639 10047
rect 4077 10013 4111 10047
rect 7113 10013 7147 10047
rect 8677 10013 8711 10047
rect 16957 10013 16991 10047
rect 17141 10013 17175 10047
rect 19165 10013 19199 10047
rect 19901 10013 19935 10047
rect 21557 10013 21591 10047
rect 25237 10013 25271 10047
rect 27077 10013 27111 10047
rect 1961 9945 1995 9979
rect 6101 9945 6135 9979
rect 6469 9945 6503 9979
rect 26249 9945 26283 9979
rect 2053 9877 2087 9911
rect 3709 9877 3743 9911
rect 6561 9877 6595 9911
rect 7573 9877 7607 9911
rect 8309 9877 8343 9911
rect 16497 9877 16531 9911
rect 21925 9877 21959 9911
rect 26709 9877 26743 9911
rect 2421 9673 2455 9707
rect 6653 9673 6687 9707
rect 8125 9673 8159 9707
rect 21097 9673 21131 9707
rect 21741 9673 21775 9707
rect 25237 9673 25271 9707
rect 26985 9673 27019 9707
rect 2145 9605 2179 9639
rect 4169 9605 4203 9639
rect 5641 9605 5675 9639
rect 6837 9605 6871 9639
rect 15945 9605 15979 9639
rect 18613 9605 18647 9639
rect 24409 9605 24443 9639
rect 25513 9605 25547 9639
rect 3157 9537 3191 9571
rect 3709 9537 3743 9571
rect 4721 9537 4755 9571
rect 6193 9537 6227 9571
rect 7389 9537 7423 9571
rect 15577 9537 15611 9571
rect 17049 9537 17083 9571
rect 21373 9537 21407 9571
rect 1409 9469 1443 9503
rect 4537 9469 4571 9503
rect 16313 9469 16347 9503
rect 19073 9469 19107 9503
rect 24041 9469 24075 9503
rect 24225 9469 24259 9503
rect 25329 9469 25363 9503
rect 25881 9469 25915 9503
rect 26341 9469 26375 9503
rect 26433 9469 26467 9503
rect 27537 9469 27571 9503
rect 28089 9469 28123 9503
rect 3065 9401 3099 9435
rect 4077 9401 4111 9435
rect 5733 9401 5767 9435
rect 7205 9401 7239 9435
rect 16773 9401 16807 9435
rect 17417 9401 17451 9435
rect 17877 9401 17911 9435
rect 19340 9401 19374 9435
rect 1593 9333 1627 9367
rect 2605 9333 2639 9367
rect 2973 9333 3007 9367
rect 4629 9333 4663 9367
rect 5181 9333 5215 9367
rect 7297 9333 7331 9367
rect 16405 9333 16439 9367
rect 16865 9333 16899 9367
rect 18889 9333 18923 9367
rect 20453 9333 20487 9367
rect 24869 9333 24903 9367
rect 26617 9333 26651 9367
rect 27721 9333 27755 9367
rect 1593 9129 1627 9163
rect 2329 9129 2363 9163
rect 2881 9129 2915 9163
rect 3617 9129 3651 9163
rect 7205 9129 7239 9163
rect 15301 9129 15335 9163
rect 19165 9129 19199 9163
rect 19717 9129 19751 9163
rect 24685 9129 24719 9163
rect 2237 9061 2271 9095
rect 5172 9061 5206 9095
rect 16221 9061 16255 9095
rect 16580 9061 16614 9095
rect 19625 9061 19659 9095
rect 7757 8993 7791 9027
rect 16313 8993 16347 9027
rect 25329 8993 25363 9027
rect 26525 8993 26559 9027
rect 2513 8925 2547 8959
rect 3249 8925 3283 8959
rect 4905 8925 4939 8959
rect 7849 8925 7883 8959
rect 7941 8925 7975 8959
rect 19901 8925 19935 8959
rect 4353 8857 4387 8891
rect 18797 8857 18831 8891
rect 1869 8789 1903 8823
rect 4813 8789 4847 8823
rect 6285 8789 6319 8823
rect 6929 8789 6963 8823
rect 7389 8789 7423 8823
rect 17693 8789 17727 8823
rect 19257 8789 19291 8823
rect 25513 8789 25547 8823
rect 26709 8789 26743 8823
rect 1777 8585 1811 8619
rect 1961 8585 1995 8619
rect 3341 8585 3375 8619
rect 3709 8585 3743 8619
rect 4813 8585 4847 8619
rect 9137 8585 9171 8619
rect 16221 8585 16255 8619
rect 18613 8585 18647 8619
rect 19717 8585 19751 8619
rect 20177 8585 20211 8619
rect 25145 8585 25179 8619
rect 25881 8585 25915 8619
rect 27353 8585 27387 8619
rect 27721 8585 27755 8619
rect 28089 8585 28123 8619
rect 8217 8517 8251 8551
rect 8769 8517 8803 8551
rect 15853 8517 15887 8551
rect 25513 8517 25547 8551
rect 26617 8517 26651 8551
rect 2513 8449 2547 8483
rect 3065 8449 3099 8483
rect 4169 8449 4203 8483
rect 5273 8449 5307 8483
rect 5457 8449 5491 8483
rect 15485 8449 15519 8483
rect 16773 8449 16807 8483
rect 16865 8449 16899 8483
rect 17877 8449 17911 8483
rect 19165 8449 19199 8483
rect 19349 8449 19383 8483
rect 2329 8381 2363 8415
rect 3525 8381 3559 8415
rect 4721 8381 4755 8415
rect 6561 8381 6595 8415
rect 6837 8381 6871 8415
rect 16681 8381 16715 8415
rect 17325 8381 17359 8415
rect 25329 8381 25363 8415
rect 26433 8381 26467 8415
rect 26985 8381 27019 8415
rect 27537 8381 27571 8415
rect 5181 8313 5215 8347
rect 6285 8313 6319 8347
rect 7104 8313 7138 8347
rect 19073 8313 19107 8347
rect 20453 8313 20487 8347
rect 2421 8245 2455 8279
rect 5825 8245 5859 8279
rect 16313 8245 16347 8279
rect 18705 8245 18739 8279
rect 2329 8041 2363 8075
rect 2697 8041 2731 8075
rect 3433 8041 3467 8075
rect 4629 8041 4663 8075
rect 4997 8041 5031 8075
rect 5641 8041 5675 8075
rect 6653 8041 6687 8075
rect 8217 8041 8251 8075
rect 16405 8041 16439 8075
rect 20177 8041 20211 8075
rect 20913 8041 20947 8075
rect 21281 8041 21315 8075
rect 25513 8041 25547 8075
rect 3065 7973 3099 8007
rect 4537 7973 4571 8007
rect 8125 7973 8159 8007
rect 16926 7973 16960 8007
rect 1409 7905 1443 7939
rect 2053 7905 2087 7939
rect 2513 7905 2547 7939
rect 6561 7905 6595 7939
rect 16681 7905 16715 7939
rect 19533 7905 19567 7939
rect 25329 7905 25363 7939
rect 26525 7905 26559 7939
rect 5089 7837 5123 7871
rect 5273 7837 5307 7871
rect 6101 7837 6135 7871
rect 6837 7837 6871 7871
rect 7481 7837 7515 7871
rect 8309 7837 8343 7871
rect 19625 7837 19659 7871
rect 19717 7837 19751 7871
rect 21373 7837 21407 7871
rect 21465 7837 21499 7871
rect 6193 7769 6227 7803
rect 18797 7769 18831 7803
rect 1593 7701 1627 7735
rect 7757 7701 7791 7735
rect 18061 7701 18095 7735
rect 19165 7701 19199 7735
rect 26709 7701 26743 7735
rect 1961 7497 1995 7531
rect 2421 7497 2455 7531
rect 4261 7497 4295 7531
rect 4721 7497 4755 7531
rect 5181 7497 5215 7531
rect 6285 7497 6319 7531
rect 6837 7497 6871 7531
rect 7849 7497 7883 7531
rect 8217 7497 8251 7531
rect 16313 7497 16347 7531
rect 19165 7497 19199 7531
rect 21005 7497 21039 7531
rect 21649 7497 21683 7531
rect 25329 7497 25363 7531
rect 27077 7497 27111 7531
rect 2697 7429 2731 7463
rect 5089 7429 5123 7463
rect 18061 7429 18095 7463
rect 21281 7429 21315 7463
rect 27353 7429 27387 7463
rect 3157 7361 3191 7395
rect 5733 7361 5767 7395
rect 7481 7361 7515 7395
rect 15945 7361 15979 7395
rect 16865 7361 16899 7395
rect 17049 7361 17083 7395
rect 18613 7361 18647 7395
rect 20177 7361 20211 7395
rect 1409 7293 1443 7327
rect 2519 7293 2553 7327
rect 3617 7293 3651 7327
rect 5641 7293 5675 7327
rect 6653 7293 6687 7327
rect 15577 7293 15611 7327
rect 16773 7293 16807 7327
rect 18429 7293 18463 7327
rect 19993 7293 20027 7327
rect 26433 7293 26467 7327
rect 27537 7293 27571 7327
rect 28089 7293 28123 7327
rect 5549 7225 5583 7259
rect 17785 7225 17819 7259
rect 20085 7225 20119 7259
rect 1593 7157 1627 7191
rect 3801 7157 3835 7191
rect 7205 7157 7239 7191
rect 7297 7157 7331 7191
rect 8585 7157 8619 7191
rect 16405 7157 16439 7191
rect 17417 7157 17451 7191
rect 18521 7157 18555 7191
rect 19625 7157 19659 7191
rect 26617 7157 26651 7191
rect 27721 7157 27755 7191
rect 2053 6953 2087 6987
rect 4721 6953 4755 6987
rect 5181 6953 5215 6987
rect 5641 6953 5675 6987
rect 6285 6953 6319 6987
rect 7297 6953 7331 6987
rect 16773 6953 16807 6987
rect 18521 6953 18555 6987
rect 19257 6953 19291 6987
rect 19717 6953 19751 6987
rect 19993 6953 20027 6987
rect 18153 6885 18187 6919
rect 1409 6817 1443 6851
rect 2329 6817 2363 6851
rect 2513 6817 2547 6851
rect 15301 6817 15335 6851
rect 18889 6817 18923 6851
rect 26525 6817 26559 6851
rect 2697 6681 2731 6715
rect 1593 6613 1627 6647
rect 6929 6613 6963 6647
rect 15485 6613 15519 6647
rect 26709 6613 26743 6647
rect 1593 6409 1627 6443
rect 2421 6409 2455 6443
rect 3157 6409 3191 6443
rect 5273 6409 5307 6443
rect 15393 6409 15427 6443
rect 26525 6409 26559 6443
rect 2053 6341 2087 6375
rect 1409 6205 1443 6239
rect 2513 6205 2547 6239
rect 2697 6069 2731 6103
rect 2513 5865 2547 5899
rect 1409 5729 1443 5763
rect 1593 5525 1627 5559
rect 1593 5321 1627 5355
rect 26433 5117 26467 5151
rect 26985 5117 27019 5151
rect 26617 4981 26651 5015
rect 2053 3145 2087 3179
rect 1409 2941 1443 2975
rect 26433 2941 26467 2975
rect 26985 2941 27019 2975
rect 1593 2805 1627 2839
rect 26617 2805 26651 2839
rect 6377 2601 6411 2635
rect 8309 2601 8343 2635
rect 6745 2465 6779 2499
rect 7196 2465 7230 2499
rect 6929 2397 6963 2431
<< metal1 >>
rect 3326 22788 3332 22840
rect 3384 22828 3390 22840
rect 10594 22828 10600 22840
rect 3384 22800 10600 22828
rect 3384 22788 3390 22800
rect 10594 22788 10600 22800
rect 10652 22788 10658 22840
rect 3510 22516 3516 22568
rect 3568 22556 3574 22568
rect 7374 22556 7380 22568
rect 3568 22528 7380 22556
rect 3568 22516 3574 22528
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 12345 21131 12403 21137
rect 12345 21097 12357 21131
rect 12391 21128 12403 21131
rect 13998 21128 14004 21140
rect 12391 21100 14004 21128
rect 12391 21097 12403 21100
rect 12345 21091 12403 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 17497 21131 17555 21137
rect 17497 21097 17509 21131
rect 17543 21128 17555 21131
rect 19610 21128 19616 21140
rect 17543 21100 19616 21128
rect 17543 21097 17555 21100
rect 17497 21091 17555 21097
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 17954 21020 17960 21072
rect 18012 21060 18018 21072
rect 18012 21032 19104 21060
rect 18012 21020 18018 21032
rect 12158 20992 12164 21004
rect 12119 20964 12164 20992
rect 12158 20952 12164 20964
rect 12216 20952 12222 21004
rect 16574 20952 16580 21004
rect 16632 20992 16638 21004
rect 17313 20995 17371 21001
rect 17313 20992 17325 20995
rect 16632 20964 17325 20992
rect 16632 20952 16638 20964
rect 17313 20961 17325 20964
rect 17359 20961 17371 20995
rect 17313 20955 17371 20961
rect 18233 20995 18291 21001
rect 18233 20961 18245 20995
rect 18279 20992 18291 20995
rect 18693 20995 18751 21001
rect 18693 20992 18705 20995
rect 18279 20964 18705 20992
rect 18279 20961 18291 20964
rect 18233 20955 18291 20961
rect 18693 20961 18705 20964
rect 18739 20992 18751 20995
rect 18966 20992 18972 21004
rect 18739 20964 18972 20992
rect 18739 20961 18751 20964
rect 18693 20955 18751 20961
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 18506 20884 18512 20936
rect 18564 20924 18570 20936
rect 18785 20927 18843 20933
rect 18785 20924 18797 20927
rect 18564 20896 18797 20924
rect 18564 20884 18570 20896
rect 18785 20893 18797 20896
rect 18831 20893 18843 20927
rect 18785 20887 18843 20893
rect 4062 20816 4068 20868
rect 4120 20856 4126 20868
rect 5626 20856 5632 20868
rect 4120 20828 5632 20856
rect 4120 20816 4126 20828
rect 5626 20816 5632 20828
rect 5684 20816 5690 20868
rect 18800 20856 18828 20887
rect 18874 20884 18880 20936
rect 18932 20924 18938 20936
rect 19076 20924 19104 21032
rect 18932 20896 19104 20924
rect 18932 20884 18938 20896
rect 19242 20856 19248 20868
rect 18800 20828 19248 20856
rect 19242 20816 19248 20828
rect 19300 20816 19306 20868
rect 21726 20816 21732 20868
rect 21784 20856 21790 20868
rect 25038 20856 25044 20868
rect 21784 20828 25044 20856
rect 21784 20816 21790 20828
rect 25038 20816 25044 20828
rect 25096 20816 25102 20868
rect 4982 20788 4988 20800
rect 4943 20760 4988 20788
rect 4982 20748 4988 20760
rect 5040 20748 5046 20800
rect 12710 20788 12716 20800
rect 12671 20760 12716 20788
rect 12710 20748 12716 20760
rect 12768 20748 12774 20800
rect 18322 20788 18328 20800
rect 18283 20760 18328 20788
rect 18322 20748 18328 20760
rect 18380 20748 18386 20800
rect 20162 20788 20168 20800
rect 20123 20760 20168 20788
rect 20162 20748 20168 20760
rect 20220 20748 20226 20800
rect 22186 20748 22192 20800
rect 22244 20788 22250 20800
rect 24854 20788 24860 20800
rect 22244 20760 24860 20788
rect 22244 20748 22250 20760
rect 24854 20748 24860 20760
rect 24912 20748 24918 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 992 20556 1593 20584
rect 992 20544 998 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 1581 20547 1639 20553
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2682 20584 2688 20596
rect 2639 20556 2688 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2682 20544 2688 20556
rect 2740 20544 2746 20596
rect 7285 20587 7343 20593
rect 7285 20553 7297 20587
rect 7331 20584 7343 20587
rect 8202 20584 8208 20596
rect 7331 20556 8208 20584
rect 7331 20553 7343 20556
rect 7285 20547 7343 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9493 20587 9551 20593
rect 9493 20553 9505 20587
rect 9539 20584 9551 20587
rect 10226 20584 10232 20596
rect 9539 20556 10232 20584
rect 9539 20553 9551 20556
rect 9493 20547 9551 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 14645 20587 14703 20593
rect 14645 20553 14657 20587
rect 14691 20584 14703 20587
rect 15838 20584 15844 20596
rect 14691 20556 15844 20584
rect 14691 20553 14703 20556
rect 14645 20547 14703 20553
rect 15838 20544 15844 20556
rect 15896 20544 15902 20596
rect 16945 20587 17003 20593
rect 16945 20553 16957 20587
rect 16991 20584 17003 20587
rect 17770 20584 17776 20596
rect 16991 20556 17776 20584
rect 16991 20553 17003 20556
rect 16945 20547 17003 20553
rect 17770 20544 17776 20556
rect 17828 20544 17834 20596
rect 18601 20587 18659 20593
rect 18601 20553 18613 20587
rect 18647 20584 18659 20587
rect 20162 20584 20168 20596
rect 18647 20556 20168 20584
rect 18647 20553 18659 20556
rect 18601 20547 18659 20553
rect 20162 20544 20168 20556
rect 20220 20584 20226 20596
rect 24305 20587 24363 20593
rect 20220 20556 20668 20584
rect 20220 20544 20226 20556
rect 11333 20519 11391 20525
rect 11333 20485 11345 20519
rect 11379 20516 11391 20519
rect 12158 20516 12164 20528
rect 11379 20488 12164 20516
rect 11379 20485 11391 20488
rect 11333 20479 11391 20485
rect 12158 20476 12164 20488
rect 12216 20516 12222 20528
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 12216 20488 12449 20516
rect 12216 20476 12222 20488
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12437 20479 12495 20485
rect 17497 20519 17555 20525
rect 17497 20485 17509 20519
rect 17543 20516 17555 20519
rect 17954 20516 17960 20528
rect 17543 20488 17960 20516
rect 17543 20485 17555 20488
rect 17497 20479 17555 20485
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 19334 20476 19340 20528
rect 19392 20516 19398 20528
rect 19613 20519 19671 20525
rect 19613 20516 19625 20519
rect 19392 20488 19625 20516
rect 19392 20476 19398 20488
rect 19613 20485 19625 20488
rect 19659 20485 19671 20519
rect 19613 20479 19671 20485
rect 4982 20408 4988 20460
rect 5040 20448 5046 20460
rect 5353 20451 5411 20457
rect 5353 20448 5365 20451
rect 5040 20420 5365 20448
rect 5040 20408 5046 20420
rect 5353 20417 5365 20420
rect 5399 20417 5411 20451
rect 5353 20411 5411 20417
rect 5445 20451 5503 20457
rect 5445 20417 5457 20451
rect 5491 20417 5503 20451
rect 5445 20411 5503 20417
rect 1397 20383 1455 20389
rect 1397 20349 1409 20383
rect 1443 20380 1455 20383
rect 1443 20352 1992 20380
rect 1443 20349 1455 20352
rect 1397 20343 1455 20349
rect 1964 20256 1992 20352
rect 2130 20340 2136 20392
rect 2188 20380 2194 20392
rect 2409 20383 2467 20389
rect 2409 20380 2421 20383
rect 2188 20352 2421 20380
rect 2188 20340 2194 20352
rect 2409 20349 2421 20352
rect 2455 20380 2467 20383
rect 2869 20383 2927 20389
rect 2869 20380 2881 20383
rect 2455 20352 2881 20380
rect 2455 20349 2467 20352
rect 2409 20343 2467 20349
rect 2869 20349 2881 20352
rect 2915 20349 2927 20383
rect 2869 20343 2927 20349
rect 4706 20340 4712 20392
rect 4764 20380 4770 20392
rect 4801 20383 4859 20389
rect 4801 20380 4813 20383
rect 4764 20352 4813 20380
rect 4764 20340 4770 20352
rect 4801 20349 4813 20352
rect 4847 20380 4859 20383
rect 5460 20380 5488 20411
rect 12710 20408 12716 20460
rect 12768 20448 12774 20460
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12768 20420 12909 20448
rect 12768 20408 12774 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20417 13047 20451
rect 12989 20411 13047 20417
rect 4847 20352 5488 20380
rect 7101 20383 7159 20389
rect 4847 20349 4859 20352
rect 4801 20343 4859 20349
rect 7101 20349 7113 20383
rect 7147 20380 7159 20383
rect 9309 20383 9367 20389
rect 7147 20352 7512 20380
rect 7147 20349 7159 20352
rect 7101 20343 7159 20349
rect 5261 20315 5319 20321
rect 5261 20312 5273 20315
rect 4356 20284 5273 20312
rect 1946 20244 1952 20256
rect 1907 20216 1952 20244
rect 1946 20204 1952 20216
rect 2004 20204 2010 20256
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4356 20253 4384 20284
rect 5261 20281 5273 20284
rect 5307 20281 5319 20315
rect 5261 20275 5319 20281
rect 7484 20256 7512 20352
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 12253 20383 12311 20389
rect 9355 20352 9812 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 9784 20256 9812 20352
rect 12253 20349 12265 20383
rect 12299 20380 12311 20383
rect 13004 20380 13032 20411
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 20640 20457 20668 20556
rect 24305 20553 24317 20587
rect 24351 20584 24363 20587
rect 25222 20584 25228 20596
rect 24351 20556 25228 20584
rect 24351 20553 24363 20556
rect 24305 20547 24363 20553
rect 25222 20544 25228 20556
rect 25280 20544 25286 20596
rect 26602 20584 26608 20596
rect 26563 20556 26608 20584
rect 26602 20544 26608 20556
rect 26660 20544 26666 20596
rect 25406 20516 25412 20528
rect 25367 20488 25412 20516
rect 25406 20476 25412 20488
rect 25464 20476 25470 20528
rect 17865 20451 17923 20457
rect 17865 20448 17877 20451
rect 17644 20420 17877 20448
rect 17644 20408 17650 20420
rect 17865 20417 17877 20420
rect 17911 20448 17923 20451
rect 19153 20451 19211 20457
rect 19153 20448 19165 20451
rect 17911 20420 19165 20448
rect 17911 20417 17923 20420
rect 17865 20411 17923 20417
rect 19153 20417 19165 20420
rect 19199 20417 19211 20451
rect 19153 20411 19211 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 13630 20380 13636 20392
rect 12299 20352 13636 20380
rect 12299 20349 12311 20352
rect 12253 20343 12311 20349
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13814 20340 13820 20392
rect 13872 20380 13878 20392
rect 14461 20383 14519 20389
rect 14461 20380 14473 20383
rect 13872 20352 14473 20380
rect 13872 20340 13878 20352
rect 14461 20349 14473 20352
rect 14507 20380 14519 20383
rect 14921 20383 14979 20389
rect 14921 20380 14933 20383
rect 14507 20352 14933 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 14921 20349 14933 20352
rect 14967 20349 14979 20383
rect 16758 20380 16764 20392
rect 16719 20352 16764 20380
rect 14921 20343 14979 20349
rect 16758 20340 16764 20352
rect 16816 20340 16822 20392
rect 20162 20340 20168 20392
rect 20220 20380 20226 20392
rect 20732 20380 20760 20411
rect 20220 20352 20760 20380
rect 24121 20383 24179 20389
rect 20220 20340 20226 20352
rect 24121 20349 24133 20383
rect 24167 20380 24179 20383
rect 25225 20383 25283 20389
rect 24167 20352 24716 20380
rect 24167 20349 24179 20352
rect 24121 20343 24179 20349
rect 12802 20312 12808 20324
rect 12715 20284 12808 20312
rect 12802 20272 12808 20284
rect 12860 20312 12866 20324
rect 13449 20315 13507 20321
rect 13449 20312 13461 20315
rect 12860 20284 13461 20312
rect 12860 20272 12866 20284
rect 13449 20281 13461 20284
rect 13495 20281 13507 20315
rect 19061 20315 19119 20321
rect 19061 20312 19073 20315
rect 13449 20275 13507 20281
rect 18616 20284 19073 20312
rect 18616 20256 18644 20284
rect 19061 20281 19073 20284
rect 19107 20281 19119 20315
rect 19978 20312 19984 20324
rect 19939 20284 19984 20312
rect 19061 20275 19119 20281
rect 19978 20272 19984 20284
rect 20036 20312 20042 20324
rect 20533 20315 20591 20321
rect 20533 20312 20545 20315
rect 20036 20284 20545 20312
rect 20036 20272 20042 20284
rect 20533 20281 20545 20284
rect 20579 20281 20591 20315
rect 20533 20275 20591 20281
rect 4341 20247 4399 20253
rect 4341 20244 4353 20247
rect 4212 20216 4353 20244
rect 4212 20204 4218 20216
rect 4341 20213 4353 20216
rect 4387 20213 4399 20247
rect 4890 20244 4896 20256
rect 4851 20216 4896 20244
rect 4341 20207 4399 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 7466 20204 7472 20256
rect 7524 20244 7530 20256
rect 7561 20247 7619 20253
rect 7561 20244 7573 20247
rect 7524 20216 7573 20244
rect 7524 20204 7530 20216
rect 7561 20213 7573 20216
rect 7607 20213 7619 20247
rect 9766 20244 9772 20256
rect 9727 20216 9772 20244
rect 7561 20207 7619 20213
rect 9766 20204 9772 20216
rect 9824 20204 9830 20256
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 12250 20244 12256 20256
rect 11747 20216 12256 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 16574 20244 16580 20256
rect 16535 20216 16580 20244
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 18509 20247 18567 20253
rect 18509 20213 18521 20247
rect 18555 20244 18567 20247
rect 18598 20244 18604 20256
rect 18555 20216 18604 20244
rect 18555 20213 18567 20216
rect 18509 20207 18567 20213
rect 18598 20204 18604 20216
rect 18656 20204 18662 20256
rect 18690 20204 18696 20256
rect 18748 20244 18754 20256
rect 18969 20247 19027 20253
rect 18969 20244 18981 20247
rect 18748 20216 18981 20244
rect 18748 20204 18754 20216
rect 18969 20213 18981 20216
rect 19015 20213 19027 20247
rect 18969 20207 19027 20213
rect 19334 20204 19340 20256
rect 19392 20244 19398 20256
rect 24688 20253 24716 20352
rect 25225 20349 25237 20383
rect 25271 20380 25283 20383
rect 26421 20383 26479 20389
rect 25271 20352 25820 20380
rect 25271 20349 25283 20352
rect 25225 20343 25283 20349
rect 20165 20247 20223 20253
rect 20165 20244 20177 20247
rect 19392 20216 20177 20244
rect 19392 20204 19398 20216
rect 20165 20213 20177 20216
rect 20211 20213 20223 20247
rect 20165 20207 20223 20213
rect 24673 20247 24731 20253
rect 24673 20213 24685 20247
rect 24719 20244 24731 20247
rect 24762 20244 24768 20256
rect 24719 20216 24768 20244
rect 24719 20213 24731 20216
rect 24673 20207 24731 20213
rect 24762 20204 24768 20216
rect 24820 20204 24826 20256
rect 25792 20253 25820 20352
rect 26421 20349 26433 20383
rect 26467 20380 26479 20383
rect 26602 20380 26608 20392
rect 26467 20352 26608 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 26602 20340 26608 20352
rect 26660 20380 26666 20392
rect 26881 20383 26939 20389
rect 26881 20380 26893 20383
rect 26660 20352 26893 20380
rect 26660 20340 26666 20352
rect 26881 20349 26893 20352
rect 26927 20349 26939 20383
rect 26881 20343 26939 20349
rect 25777 20247 25835 20253
rect 25777 20213 25789 20247
rect 25823 20244 25835 20247
rect 25866 20244 25872 20256
rect 25823 20216 25872 20244
rect 25823 20213 25835 20216
rect 25777 20207 25835 20213
rect 25866 20204 25872 20216
rect 25924 20204 25930 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 4430 20040 4436 20052
rect 4391 20012 4436 20040
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 4982 20000 4988 20052
rect 5040 20040 5046 20052
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 5040 20012 5273 20040
rect 5040 20000 5046 20012
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5626 20040 5632 20052
rect 5587 20012 5632 20040
rect 5261 20003 5319 20009
rect 5626 20000 5632 20012
rect 5684 20000 5690 20052
rect 11609 20043 11667 20049
rect 11609 20009 11621 20043
rect 11655 20040 11667 20043
rect 12710 20040 12716 20052
rect 11655 20012 12716 20040
rect 11655 20009 11667 20012
rect 11609 20003 11667 20009
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 16758 20040 16764 20052
rect 16719 20012 16764 20040
rect 16758 20000 16764 20012
rect 16816 20040 16822 20052
rect 17313 20043 17371 20049
rect 17313 20040 17325 20043
rect 16816 20012 17325 20040
rect 16816 20000 16822 20012
rect 17313 20009 17325 20012
rect 17359 20009 17371 20043
rect 17678 20040 17684 20052
rect 17591 20012 17684 20040
rect 17313 20003 17371 20009
rect 17678 20000 17684 20012
rect 17736 20040 17742 20052
rect 18877 20043 18935 20049
rect 18877 20040 18889 20043
rect 17736 20012 18889 20040
rect 17736 20000 17742 20012
rect 18877 20009 18889 20012
rect 18923 20009 18935 20043
rect 18877 20003 18935 20009
rect 21085 20043 21143 20049
rect 21085 20009 21097 20043
rect 21131 20040 21143 20043
rect 21542 20040 21548 20052
rect 21131 20012 21548 20040
rect 21131 20009 21143 20012
rect 21085 20003 21143 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 22097 20043 22155 20049
rect 22097 20009 22109 20043
rect 22143 20040 22155 20043
rect 23382 20040 23388 20052
rect 22143 20012 23388 20040
rect 22143 20009 22155 20012
rect 22097 20003 22155 20009
rect 23382 20000 23388 20012
rect 23440 20000 23446 20052
rect 11977 19975 12035 19981
rect 11977 19941 11989 19975
rect 12023 19972 12035 19975
rect 12250 19972 12256 19984
rect 12023 19944 12256 19972
rect 12023 19941 12035 19944
rect 11977 19935 12035 19941
rect 12250 19932 12256 19944
rect 12308 19932 12314 19984
rect 4062 19864 4068 19916
rect 4120 19904 4126 19916
rect 4249 19907 4307 19913
rect 4249 19904 4261 19907
rect 4120 19876 4261 19904
rect 4120 19864 4126 19876
rect 4249 19873 4261 19876
rect 4295 19873 4307 19907
rect 4249 19867 4307 19873
rect 11517 19907 11575 19913
rect 11517 19873 11529 19907
rect 11563 19904 11575 19907
rect 12069 19907 12127 19913
rect 12069 19904 12081 19907
rect 11563 19876 12081 19904
rect 11563 19873 11575 19876
rect 11517 19867 11575 19873
rect 12069 19873 12081 19876
rect 12115 19904 12127 19907
rect 12342 19904 12348 19916
rect 12115 19876 12348 19904
rect 12115 19873 12127 19876
rect 12069 19867 12127 19873
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 15194 19864 15200 19916
rect 15252 19904 15258 19916
rect 15657 19907 15715 19913
rect 15657 19904 15669 19907
rect 15252 19876 15669 19904
rect 15252 19864 15258 19876
rect 15657 19873 15669 19876
rect 15703 19873 15715 19907
rect 15657 19867 15715 19873
rect 15746 19864 15752 19916
rect 15804 19904 15810 19916
rect 17770 19904 17776 19916
rect 15804 19876 15849 19904
rect 17731 19876 17776 19904
rect 15804 19864 15810 19876
rect 17770 19864 17776 19876
rect 17828 19864 17834 19916
rect 19245 19907 19303 19913
rect 19245 19873 19257 19907
rect 19291 19904 19303 19907
rect 19610 19904 19616 19916
rect 19291 19876 19616 19904
rect 19291 19873 19303 19876
rect 19245 19867 19303 19873
rect 19610 19864 19616 19876
rect 19668 19904 19674 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 19668 19876 20545 19904
rect 19668 19864 19674 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20898 19904 20904 19916
rect 20859 19876 20904 19904
rect 20533 19867 20591 19873
rect 20898 19864 20904 19876
rect 20956 19864 20962 19916
rect 21910 19904 21916 19916
rect 21871 19876 21916 19904
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 5718 19836 5724 19848
rect 5679 19808 5724 19836
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 5813 19839 5871 19845
rect 5813 19805 5825 19839
rect 5859 19805 5871 19839
rect 12158 19836 12164 19848
rect 12119 19808 12164 19836
rect 5813 19799 5871 19805
rect 5828 19768 5856 19799
rect 12158 19796 12164 19808
rect 12216 19836 12222 19848
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 12216 19808 12633 19836
rect 12216 19796 12222 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 15838 19836 15844 19848
rect 15799 19808 15844 19836
rect 12621 19799 12679 19805
rect 15838 19796 15844 19808
rect 15896 19796 15902 19848
rect 17862 19836 17868 19848
rect 17823 19808 17868 19836
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 19150 19796 19156 19848
rect 19208 19836 19214 19848
rect 19337 19839 19395 19845
rect 19337 19836 19349 19839
rect 19208 19808 19349 19836
rect 19208 19796 19214 19808
rect 19337 19805 19349 19808
rect 19383 19805 19395 19839
rect 19337 19799 19395 19805
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 20714 19836 20720 19848
rect 19567 19808 20720 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 5276 19740 5856 19768
rect 5276 19712 5304 19740
rect 18782 19728 18788 19780
rect 18840 19768 18846 19780
rect 19536 19768 19564 19799
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 26513 19839 26571 19845
rect 26513 19805 26525 19839
rect 26559 19836 26571 19839
rect 27065 19839 27123 19845
rect 27065 19836 27077 19839
rect 26559 19808 27077 19836
rect 26559 19805 26571 19808
rect 26513 19799 26571 19805
rect 27065 19805 27077 19808
rect 27111 19836 27123 19839
rect 27430 19836 27436 19848
rect 27111 19808 27436 19836
rect 27111 19805 27123 19808
rect 27065 19799 27123 19805
rect 27430 19796 27436 19808
rect 27488 19796 27494 19848
rect 18840 19740 19564 19768
rect 18840 19728 18846 19740
rect 3513 19703 3571 19709
rect 3513 19669 3525 19703
rect 3559 19700 3571 19703
rect 3878 19700 3884 19712
rect 3559 19672 3884 19700
rect 3559 19669 3571 19672
rect 3513 19663 3571 19669
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 5077 19703 5135 19709
rect 5077 19669 5089 19703
rect 5123 19700 5135 19703
rect 5258 19700 5264 19712
rect 5123 19672 5264 19700
rect 5123 19669 5135 19672
rect 5077 19663 5135 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 10870 19700 10876 19712
rect 10831 19672 10876 19700
rect 10870 19660 10876 19672
rect 10928 19660 10934 19712
rect 14918 19700 14924 19712
rect 14879 19672 14924 19700
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15286 19700 15292 19712
rect 15247 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 18230 19660 18236 19712
rect 18288 19700 18294 19712
rect 18601 19703 18659 19709
rect 18601 19700 18613 19703
rect 18288 19672 18613 19700
rect 18288 19660 18294 19672
rect 18601 19669 18613 19672
rect 18647 19700 18659 19703
rect 18690 19700 18696 19712
rect 18647 19672 18696 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 18690 19660 18696 19672
rect 18748 19660 18754 19712
rect 20162 19700 20168 19712
rect 20123 19672 20168 19700
rect 20162 19660 20168 19672
rect 20220 19660 20226 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 5626 19456 5632 19508
rect 5684 19496 5690 19508
rect 5997 19499 6055 19505
rect 5997 19496 6009 19499
rect 5684 19468 6009 19496
rect 5684 19456 5690 19468
rect 5997 19465 6009 19468
rect 6043 19496 6055 19499
rect 6362 19496 6368 19508
rect 6043 19468 6368 19496
rect 6043 19465 6055 19468
rect 5997 19459 6055 19465
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 13630 19456 13636 19508
rect 13688 19496 13694 19508
rect 13814 19496 13820 19508
rect 13688 19468 13820 19496
rect 13688 19456 13694 19468
rect 13814 19456 13820 19468
rect 13872 19456 13878 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 17678 19496 17684 19508
rect 16715 19468 17684 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 17678 19456 17684 19468
rect 17736 19456 17742 19508
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 14918 19428 14924 19440
rect 14608 19400 14924 19428
rect 14608 19388 14614 19400
rect 14918 19388 14924 19400
rect 14976 19428 14982 19440
rect 14976 19400 15516 19428
rect 14976 19388 14982 19400
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19360 3387 19363
rect 3694 19360 3700 19372
rect 3375 19332 3700 19360
rect 3375 19329 3387 19332
rect 3329 19323 3387 19329
rect 3694 19320 3700 19332
rect 3752 19360 3758 19372
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 3752 19332 3985 19360
rect 3752 19320 3758 19332
rect 3973 19329 3985 19332
rect 4019 19329 4031 19363
rect 4890 19360 4896 19372
rect 3973 19323 4031 19329
rect 4080 19332 4896 19360
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 3789 19295 3847 19301
rect 3789 19292 3801 19295
rect 3007 19264 3801 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 3789 19261 3801 19264
rect 3835 19292 3847 19295
rect 4080 19292 4108 19332
rect 4890 19320 4896 19332
rect 4948 19320 4954 19372
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5316 19332 5549 19360
rect 5316 19320 5322 19332
rect 5537 19329 5549 19332
rect 5583 19360 5595 19363
rect 6365 19363 6423 19369
rect 6365 19360 6377 19363
rect 5583 19332 6377 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 6365 19329 6377 19332
rect 6411 19329 6423 19363
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 6365 19323 6423 19329
rect 10796 19332 11345 19360
rect 3835 19264 4108 19292
rect 4525 19295 4583 19301
rect 3835 19261 3847 19264
rect 3789 19255 3847 19261
rect 4525 19261 4537 19295
rect 4571 19292 4583 19295
rect 5718 19292 5724 19304
rect 4571 19264 5724 19292
rect 4571 19261 4583 19264
rect 4525 19255 4583 19261
rect 5718 19252 5724 19264
rect 5776 19252 5782 19304
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10796 19292 10824 19332
rect 11333 19329 11345 19332
rect 11379 19360 11391 19363
rect 11793 19363 11851 19369
rect 11793 19360 11805 19363
rect 11379 19332 11805 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11793 19329 11805 19332
rect 11839 19360 11851 19363
rect 12158 19360 12164 19372
rect 11839 19332 12164 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 12158 19320 12164 19332
rect 12216 19360 12222 19372
rect 15194 19360 15200 19372
rect 12216 19332 12572 19360
rect 12216 19320 12222 19332
rect 12544 19304 12572 19332
rect 15120 19332 15200 19360
rect 10735 19264 10824 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 10870 19252 10876 19304
rect 10928 19292 10934 19304
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 10928 19264 11253 19292
rect 10928 19252 10934 19264
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11241 19255 11299 19261
rect 12176 19264 12449 19292
rect 4062 19224 4068 19236
rect 3436 19196 4068 19224
rect 1670 19156 1676 19168
rect 1631 19128 1676 19156
rect 1670 19116 1676 19128
rect 1728 19116 1734 19168
rect 1946 19156 1952 19168
rect 1907 19128 1952 19156
rect 1946 19116 1952 19128
rect 2004 19116 2010 19168
rect 3436 19165 3464 19196
rect 4062 19184 4068 19196
rect 4120 19184 4126 19236
rect 4890 19224 4896 19236
rect 4851 19196 4896 19224
rect 4890 19184 4896 19196
rect 4948 19224 4954 19236
rect 5353 19227 5411 19233
rect 5353 19224 5365 19227
rect 4948 19196 5365 19224
rect 4948 19184 4954 19196
rect 5353 19193 5365 19196
rect 5399 19193 5411 19227
rect 5353 19187 5411 19193
rect 10321 19227 10379 19233
rect 10321 19193 10333 19227
rect 10367 19224 10379 19227
rect 11149 19227 11207 19233
rect 11149 19224 11161 19227
rect 10367 19196 11161 19224
rect 10367 19193 10379 19196
rect 10321 19187 10379 19193
rect 11149 19193 11161 19196
rect 11195 19224 11207 19227
rect 11330 19224 11336 19236
rect 11195 19196 11336 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 11330 19184 11336 19196
rect 11388 19184 11394 19236
rect 3421 19159 3479 19165
rect 3421 19125 3433 19159
rect 3467 19125 3479 19159
rect 3878 19156 3884 19168
rect 3839 19128 3884 19156
rect 3421 19119 3479 19125
rect 3878 19116 3884 19128
rect 3936 19116 3942 19168
rect 4982 19156 4988 19168
rect 4943 19128 4988 19156
rect 4982 19116 4988 19128
rect 5040 19116 5046 19168
rect 5442 19156 5448 19168
rect 5403 19128 5448 19156
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 6822 19156 6828 19168
rect 6783 19128 6828 19156
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 10778 19156 10784 19168
rect 10739 19128 10784 19156
rect 10778 19116 10784 19128
rect 10836 19116 10842 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12176 19165 12204 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 12693 19295 12751 19301
rect 12693 19292 12705 19295
rect 12584 19264 12705 19292
rect 12584 19252 12590 19264
rect 12693 19261 12705 19264
rect 12739 19261 12751 19295
rect 12693 19255 12751 19261
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19292 14887 19295
rect 15120 19292 15148 19332
rect 15194 19320 15200 19332
rect 15252 19320 15258 19372
rect 15488 19369 15516 19400
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 19260 19332 19472 19360
rect 15286 19292 15292 19304
rect 14875 19264 15148 19292
rect 15247 19264 15292 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 17037 19295 17095 19301
rect 17037 19261 17049 19295
rect 17083 19292 17095 19295
rect 17770 19292 17776 19304
rect 17083 19264 17776 19292
rect 17083 19261 17095 19264
rect 17037 19255 17095 19261
rect 17770 19252 17776 19264
rect 17828 19252 17834 19304
rect 18874 19292 18880 19304
rect 18835 19264 18880 19292
rect 18874 19252 18880 19264
rect 18932 19292 18938 19304
rect 19260 19292 19288 19332
rect 18932 19264 19288 19292
rect 19337 19295 19395 19301
rect 18932 19252 18938 19264
rect 19337 19261 19349 19295
rect 19383 19261 19395 19295
rect 19444 19292 19472 19332
rect 26510 19320 26516 19372
rect 26568 19360 26574 19372
rect 27617 19363 27675 19369
rect 27617 19360 27629 19363
rect 26568 19332 27629 19360
rect 26568 19320 26574 19332
rect 27617 19329 27629 19332
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 19593 19295 19651 19301
rect 19593 19292 19605 19295
rect 19444 19264 19605 19292
rect 19337 19255 19395 19261
rect 19593 19261 19605 19264
rect 19639 19292 19651 19295
rect 20162 19292 20168 19304
rect 19639 19264 20168 19292
rect 19639 19261 19651 19264
rect 19593 19255 19651 19261
rect 14461 19227 14519 19233
rect 14461 19193 14473 19227
rect 14507 19224 14519 19227
rect 17405 19227 17463 19233
rect 14507 19196 15056 19224
rect 14507 19193 14519 19196
rect 14461 19187 14519 19193
rect 15028 19168 15056 19196
rect 17405 19193 17417 19227
rect 17451 19224 17463 19227
rect 17862 19224 17868 19236
rect 17451 19196 17868 19224
rect 17451 19193 17463 19196
rect 17405 19187 17463 19193
rect 17862 19184 17868 19196
rect 17920 19184 17926 19236
rect 18414 19224 18420 19236
rect 18248 19196 18420 19224
rect 12161 19159 12219 19165
rect 12161 19156 12173 19159
rect 11940 19128 12173 19156
rect 11940 19116 11946 19128
rect 12161 19125 12173 19128
rect 12207 19125 12219 19159
rect 14918 19156 14924 19168
rect 14879 19128 14924 19156
rect 12161 19119 12219 19125
rect 14918 19116 14924 19128
rect 14976 19116 14982 19168
rect 15010 19116 15016 19168
rect 15068 19156 15074 19168
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 15068 19128 15393 19156
rect 15068 19116 15074 19128
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15381 19119 15439 19125
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 15933 19159 15991 19165
rect 15933 19156 15945 19159
rect 15804 19128 15945 19156
rect 15804 19116 15810 19128
rect 15933 19125 15945 19128
rect 15979 19125 15991 19159
rect 15933 19119 15991 19125
rect 17773 19159 17831 19165
rect 17773 19125 17785 19159
rect 17819 19156 17831 19159
rect 18248 19156 18276 19196
rect 18414 19184 18420 19196
rect 18472 19224 18478 19236
rect 19242 19224 19248 19236
rect 18472 19196 19248 19224
rect 18472 19184 18478 19196
rect 19242 19184 19248 19196
rect 19300 19184 19306 19236
rect 19352 19168 19380 19255
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 21821 19295 21879 19301
rect 21821 19261 21833 19295
rect 21867 19292 21879 19295
rect 22278 19292 22284 19304
rect 21867 19264 22284 19292
rect 21867 19261 21879 19264
rect 21821 19255 21879 19261
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 24581 19295 24639 19301
rect 24581 19292 24593 19295
rect 24412 19264 24593 19292
rect 20346 19184 20352 19236
rect 20404 19224 20410 19236
rect 20898 19224 20904 19236
rect 20404 19196 20904 19224
rect 20404 19184 20410 19196
rect 20898 19184 20904 19196
rect 20956 19224 20962 19236
rect 21269 19227 21327 19233
rect 21269 19224 21281 19227
rect 20956 19196 21281 19224
rect 20956 19184 20962 19196
rect 21269 19193 21281 19196
rect 21315 19193 21327 19227
rect 21269 19187 21327 19193
rect 17819 19128 18276 19156
rect 18325 19159 18383 19165
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 18325 19125 18337 19159
rect 18371 19156 18383 19159
rect 18690 19156 18696 19168
rect 18371 19128 18696 19156
rect 18371 19125 18383 19128
rect 18325 19119 18383 19125
rect 18690 19116 18696 19128
rect 18748 19116 18754 19168
rect 19153 19159 19211 19165
rect 19153 19125 19165 19159
rect 19199 19156 19211 19159
rect 19334 19156 19340 19168
rect 19199 19128 19340 19156
rect 19199 19125 19211 19128
rect 19153 19119 19211 19125
rect 19334 19116 19340 19128
rect 19392 19156 19398 19168
rect 20714 19156 20720 19168
rect 19392 19128 19485 19156
rect 20675 19128 20720 19156
rect 19392 19116 19398 19128
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 22094 19116 22100 19168
rect 22152 19156 22158 19168
rect 22281 19159 22339 19165
rect 22281 19156 22293 19159
rect 22152 19128 22293 19156
rect 22152 19116 22158 19128
rect 22281 19125 22293 19128
rect 22327 19125 22339 19159
rect 22281 19119 22339 19125
rect 22554 19116 22560 19168
rect 22612 19156 22618 19168
rect 24412 19165 24440 19264
rect 24581 19261 24593 19264
rect 24627 19261 24639 19295
rect 27430 19292 27436 19304
rect 27391 19264 27436 19292
rect 24581 19255 24639 19261
rect 27430 19252 27436 19264
rect 27488 19252 27494 19304
rect 24670 19184 24676 19236
rect 24728 19224 24734 19236
rect 24826 19227 24884 19233
rect 24826 19224 24838 19227
rect 24728 19196 24838 19224
rect 24728 19184 24734 19196
rect 24826 19193 24838 19196
rect 24872 19193 24884 19227
rect 27525 19227 27583 19233
rect 27525 19224 27537 19227
rect 24826 19187 24884 19193
rect 26896 19196 27537 19224
rect 26896 19168 26924 19196
rect 27525 19193 27537 19196
rect 27571 19193 27583 19227
rect 27525 19187 27583 19193
rect 24397 19159 24455 19165
rect 24397 19156 24409 19159
rect 22612 19128 24409 19156
rect 22612 19116 22618 19128
rect 24397 19125 24409 19128
rect 24443 19125 24455 19159
rect 25958 19156 25964 19168
rect 25919 19128 25964 19156
rect 24397 19119 24455 19125
rect 25958 19116 25964 19128
rect 26016 19116 26022 19168
rect 26510 19156 26516 19168
rect 26471 19128 26516 19156
rect 26510 19116 26516 19128
rect 26568 19116 26574 19168
rect 26878 19156 26884 19168
rect 26839 19128 26884 19156
rect 26878 19116 26884 19128
rect 26936 19116 26942 19168
rect 27062 19156 27068 19168
rect 27023 19128 27068 19156
rect 27062 19116 27068 19128
rect 27120 19116 27126 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 2682 18952 2688 18964
rect 2643 18924 2688 18952
rect 2682 18912 2688 18924
rect 2740 18912 2746 18964
rect 3881 18955 3939 18961
rect 3881 18921 3893 18955
rect 3927 18952 3939 18955
rect 4062 18952 4068 18964
rect 3927 18924 4068 18952
rect 3927 18921 3939 18924
rect 3881 18915 3939 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4706 18952 4712 18964
rect 4667 18924 4712 18952
rect 4706 18912 4712 18924
rect 4764 18912 4770 18964
rect 6178 18952 6184 18964
rect 6139 18924 6184 18952
rect 6178 18912 6184 18924
rect 6236 18912 6242 18964
rect 7282 18952 7288 18964
rect 7243 18924 7288 18952
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 7742 18952 7748 18964
rect 7703 18924 7748 18952
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 9858 18952 9864 18964
rect 9819 18924 9864 18952
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 11330 18912 11336 18964
rect 11388 18952 11394 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 11388 18924 13645 18952
rect 11388 18912 11394 18924
rect 13633 18921 13645 18924
rect 13679 18921 13691 18955
rect 13633 18915 13691 18921
rect 13814 18912 13820 18964
rect 13872 18952 13878 18964
rect 14274 18952 14280 18964
rect 13872 18924 14280 18952
rect 13872 18912 13878 18924
rect 14274 18912 14280 18924
rect 14332 18952 14338 18964
rect 14645 18955 14703 18961
rect 14645 18952 14657 18955
rect 14332 18924 14657 18952
rect 14332 18912 14338 18924
rect 14645 18921 14657 18924
rect 14691 18921 14703 18955
rect 14645 18915 14703 18921
rect 15105 18955 15163 18961
rect 15105 18921 15117 18955
rect 15151 18952 15163 18955
rect 15286 18952 15292 18964
rect 15151 18924 15292 18952
rect 15151 18921 15163 18924
rect 15105 18915 15163 18921
rect 15286 18912 15292 18924
rect 15344 18912 15350 18964
rect 15565 18955 15623 18961
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 15838 18952 15844 18964
rect 15611 18924 15844 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15838 18912 15844 18924
rect 15896 18912 15902 18964
rect 18874 18952 18880 18964
rect 18835 18924 18880 18952
rect 18874 18912 18880 18924
rect 18932 18912 18938 18964
rect 18969 18955 19027 18961
rect 18969 18921 18981 18955
rect 19015 18952 19027 18955
rect 19150 18952 19156 18964
rect 19015 18924 19156 18952
rect 19015 18921 19027 18924
rect 18969 18915 19027 18921
rect 19150 18912 19156 18924
rect 19208 18952 19214 18964
rect 20349 18955 20407 18961
rect 20349 18952 20361 18955
rect 19208 18924 20361 18952
rect 19208 18912 19214 18924
rect 20349 18921 20361 18924
rect 20395 18921 20407 18955
rect 24762 18952 24768 18964
rect 24723 18924 24768 18952
rect 20349 18915 20407 18921
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 2866 18844 2872 18896
rect 2924 18884 2930 18896
rect 4724 18884 4752 18912
rect 5046 18887 5104 18893
rect 5046 18884 5058 18887
rect 2924 18856 3096 18884
rect 4724 18856 5058 18884
rect 2924 18844 2930 18856
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 2038 18816 2044 18828
rect 1443 18788 2044 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 2038 18776 2044 18788
rect 2096 18776 2102 18828
rect 2498 18816 2504 18828
rect 2459 18788 2504 18816
rect 2498 18776 2504 18788
rect 2556 18816 2562 18828
rect 2961 18819 3019 18825
rect 2961 18816 2973 18819
rect 2556 18788 2973 18816
rect 2556 18776 2562 18788
rect 2961 18785 2973 18788
rect 3007 18785 3019 18819
rect 3068 18816 3096 18856
rect 5046 18853 5058 18856
rect 5092 18884 5104 18887
rect 5534 18884 5540 18896
rect 5092 18856 5540 18884
rect 5092 18853 5104 18856
rect 5046 18847 5104 18853
rect 5534 18844 5540 18856
rect 5592 18844 5598 18896
rect 18509 18887 18567 18893
rect 18509 18853 18521 18887
rect 18555 18884 18567 18887
rect 18782 18884 18788 18896
rect 18555 18856 18788 18884
rect 18555 18853 18567 18856
rect 18509 18847 18567 18853
rect 18782 18844 18788 18856
rect 18840 18844 18846 18896
rect 27062 18884 27068 18896
rect 26896 18856 27068 18884
rect 6454 18816 6460 18828
rect 3068 18788 6460 18816
rect 2961 18779 3019 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 7650 18816 7656 18828
rect 7611 18788 7656 18816
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 9674 18816 9680 18828
rect 9635 18788 9680 18816
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 11422 18825 11428 18828
rect 11416 18816 11428 18825
rect 11383 18788 11428 18816
rect 11416 18779 11428 18788
rect 11422 18776 11428 18779
rect 11480 18776 11486 18828
rect 13906 18776 13912 18828
rect 13964 18816 13970 18828
rect 16758 18825 16764 18828
rect 14001 18819 14059 18825
rect 14001 18816 14013 18819
rect 13964 18788 14013 18816
rect 13964 18776 13970 18788
rect 14001 18785 14013 18788
rect 14047 18785 14059 18819
rect 16752 18816 16764 18825
rect 16719 18788 16764 18816
rect 14001 18779 14059 18785
rect 16752 18779 16764 18788
rect 16758 18776 16764 18779
rect 16816 18776 16822 18828
rect 19058 18776 19064 18828
rect 19116 18816 19122 18828
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 19116 18788 19349 18816
rect 19116 18776 19122 18788
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 19426 18776 19432 18828
rect 19484 18816 19490 18828
rect 21904 18819 21962 18825
rect 19484 18788 19529 18816
rect 19484 18776 19490 18788
rect 21904 18785 21916 18819
rect 21950 18816 21962 18819
rect 23106 18816 23112 18828
rect 21950 18788 23112 18816
rect 21950 18785 21962 18788
rect 21904 18779 21962 18785
rect 23106 18776 23112 18788
rect 23164 18776 23170 18828
rect 25133 18819 25191 18825
rect 25133 18785 25145 18819
rect 25179 18816 25191 18819
rect 26145 18819 26203 18825
rect 26145 18816 26157 18819
rect 25179 18788 26157 18816
rect 25179 18785 25191 18788
rect 25133 18779 25191 18785
rect 26145 18785 26157 18788
rect 26191 18785 26203 18819
rect 26145 18779 26203 18785
rect 4798 18748 4804 18760
rect 4759 18720 4804 18748
rect 4798 18708 4804 18720
rect 4856 18708 4862 18760
rect 7834 18748 7840 18760
rect 7795 18720 7840 18748
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18717 11207 18751
rect 11149 18711 11207 18717
rect 1581 18683 1639 18689
rect 1581 18649 1593 18683
rect 1627 18680 1639 18683
rect 3234 18680 3240 18692
rect 1627 18652 3240 18680
rect 1627 18649 1639 18652
rect 1581 18643 1639 18649
rect 3234 18640 3240 18652
rect 3292 18640 3298 18692
rect 8665 18683 8723 18689
rect 8665 18649 8677 18683
rect 8711 18680 8723 18683
rect 9030 18680 9036 18692
rect 8711 18652 9036 18680
rect 8711 18649 8723 18652
rect 8665 18643 8723 18649
rect 9030 18640 9036 18652
rect 9088 18640 9094 18692
rect 2222 18572 2228 18624
rect 2280 18612 2286 18624
rect 2317 18615 2375 18621
rect 2317 18612 2329 18615
rect 2280 18584 2329 18612
rect 2280 18572 2286 18584
rect 2317 18581 2329 18584
rect 2363 18581 2375 18615
rect 2317 18575 2375 18581
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 3878 18612 3884 18624
rect 3467 18584 3884 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 3878 18572 3884 18584
rect 3936 18572 3942 18624
rect 4341 18615 4399 18621
rect 4341 18581 4353 18615
rect 4387 18612 4399 18615
rect 5442 18612 5448 18624
rect 4387 18584 5448 18612
rect 4387 18581 4399 18584
rect 4341 18575 4399 18581
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 6917 18615 6975 18621
rect 6917 18581 6929 18615
rect 6963 18612 6975 18615
rect 7006 18612 7012 18624
rect 6963 18584 7012 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 8938 18612 8944 18624
rect 8899 18584 8944 18612
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 10778 18612 10784 18624
rect 10739 18584 10784 18612
rect 10778 18572 10784 18584
rect 10836 18572 10842 18624
rect 11164 18612 11192 18711
rect 13630 18708 13636 18760
rect 13688 18748 13694 18760
rect 14090 18748 14096 18760
rect 13688 18720 14096 18748
rect 13688 18708 13694 18720
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14185 18751 14243 18757
rect 14185 18717 14197 18751
rect 14231 18717 14243 18751
rect 16482 18748 16488 18760
rect 16443 18720 16488 18748
rect 14185 18711 14243 18717
rect 12526 18680 12532 18692
rect 12487 18652 12532 18680
rect 12526 18640 12532 18652
rect 12584 18640 12590 18692
rect 13078 18640 13084 18692
rect 13136 18680 13142 18692
rect 13541 18683 13599 18689
rect 13541 18680 13553 18683
rect 13136 18652 13553 18680
rect 13136 18640 13142 18652
rect 13541 18649 13553 18652
rect 13587 18680 13599 18683
rect 14200 18680 14228 18711
rect 16482 18708 16488 18720
rect 16540 18708 16546 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 18932 18720 19533 18748
rect 18932 18708 18938 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 21634 18748 21640 18760
rect 21595 18720 21640 18748
rect 19521 18711 19579 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 25222 18748 25228 18760
rect 25183 18720 25228 18748
rect 25222 18708 25228 18720
rect 25280 18708 25286 18760
rect 25406 18748 25412 18760
rect 25319 18720 25412 18748
rect 25406 18708 25412 18720
rect 25464 18748 25470 18760
rect 25958 18748 25964 18760
rect 25464 18720 25964 18748
rect 25464 18708 25470 18720
rect 25958 18708 25964 18720
rect 26016 18708 26022 18760
rect 19978 18680 19984 18692
rect 13587 18652 14228 18680
rect 19939 18652 19984 18680
rect 13587 18649 13599 18652
rect 13541 18643 13599 18649
rect 19978 18640 19984 18652
rect 20036 18640 20042 18692
rect 24213 18683 24271 18689
rect 24213 18649 24225 18683
rect 24259 18680 24271 18683
rect 24578 18680 24584 18692
rect 24259 18652 24584 18680
rect 24259 18649 24271 18652
rect 24213 18643 24271 18649
rect 24578 18640 24584 18652
rect 24636 18640 24642 18692
rect 26160 18680 26188 18779
rect 26326 18776 26332 18828
rect 26384 18816 26390 18828
rect 26896 18825 26924 18856
rect 27062 18844 27068 18856
rect 27120 18844 27126 18896
rect 26881 18819 26939 18825
rect 26881 18816 26893 18819
rect 26384 18788 26893 18816
rect 26384 18776 26390 18788
rect 26881 18785 26893 18788
rect 26927 18785 26939 18819
rect 26881 18779 26939 18785
rect 26970 18776 26976 18828
rect 27028 18816 27034 18828
rect 27028 18788 27073 18816
rect 27028 18776 27034 18788
rect 27062 18748 27068 18760
rect 27023 18720 27068 18748
rect 27062 18708 27068 18720
rect 27120 18708 27126 18760
rect 26513 18683 26571 18689
rect 26513 18680 26525 18683
rect 26160 18652 26525 18680
rect 26513 18649 26525 18652
rect 26559 18649 26571 18683
rect 26513 18643 26571 18649
rect 11882 18612 11888 18624
rect 11164 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 17862 18612 17868 18624
rect 17823 18584 17868 18612
rect 17862 18572 17868 18584
rect 17920 18572 17926 18624
rect 23017 18615 23075 18621
rect 23017 18581 23029 18615
rect 23063 18612 23075 18615
rect 23382 18612 23388 18624
rect 23063 18584 23388 18612
rect 23063 18581 23075 18584
rect 23017 18575 23075 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 24670 18612 24676 18624
rect 24631 18584 24676 18612
rect 24670 18572 24676 18584
rect 24728 18572 24734 18624
rect 25774 18612 25780 18624
rect 25735 18584 25780 18612
rect 25774 18572 25780 18584
rect 25832 18572 25838 18624
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 3329 18411 3387 18417
rect 3329 18377 3341 18411
rect 3375 18408 3387 18411
rect 3970 18408 3976 18420
rect 3375 18380 3976 18408
rect 3375 18377 3387 18380
rect 3329 18371 3387 18377
rect 3970 18368 3976 18380
rect 4028 18368 4034 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 5442 18408 5448 18420
rect 4939 18380 5448 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 10594 18408 10600 18420
rect 10555 18380 10600 18408
rect 10594 18368 10600 18380
rect 10652 18368 10658 18420
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 10870 18408 10876 18420
rect 10827 18380 10876 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 12250 18368 12256 18420
rect 12308 18408 12314 18420
rect 12437 18411 12495 18417
rect 12437 18408 12449 18411
rect 12308 18380 12449 18408
rect 12308 18368 12314 18380
rect 12437 18377 12449 18380
rect 12483 18377 12495 18411
rect 12437 18371 12495 18377
rect 17770 18368 17776 18420
rect 17828 18408 17834 18420
rect 18049 18411 18107 18417
rect 18049 18408 18061 18411
rect 17828 18380 18061 18408
rect 17828 18368 17834 18380
rect 18049 18377 18061 18380
rect 18095 18377 18107 18411
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 18049 18371 18107 18377
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19610 18408 19616 18420
rect 19571 18380 19616 18408
rect 19610 18368 19616 18380
rect 19668 18368 19674 18420
rect 23106 18408 23112 18420
rect 23067 18380 23112 18408
rect 23106 18368 23112 18380
rect 23164 18368 23170 18420
rect 25133 18411 25191 18417
rect 25133 18377 25145 18411
rect 25179 18408 25191 18411
rect 25406 18408 25412 18420
rect 25179 18380 25412 18408
rect 25179 18377 25191 18380
rect 25133 18371 25191 18377
rect 25406 18368 25412 18380
rect 25464 18368 25470 18420
rect 27062 18408 27068 18420
rect 25700 18380 27068 18408
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 7650 18340 7656 18352
rect 6871 18312 7656 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 7650 18300 7656 18312
rect 7708 18300 7714 18352
rect 8110 18300 8116 18352
rect 8168 18340 8174 18352
rect 8573 18343 8631 18349
rect 8573 18340 8585 18343
rect 8168 18312 8585 18340
rect 8168 18300 8174 18312
rect 8573 18309 8585 18312
rect 8619 18309 8631 18343
rect 8573 18303 8631 18309
rect 16758 18300 16764 18352
rect 16816 18340 16822 18352
rect 16945 18343 17003 18349
rect 16945 18340 16957 18343
rect 16816 18312 16957 18340
rect 16816 18300 16822 18312
rect 16945 18309 16957 18312
rect 16991 18340 17003 18343
rect 17865 18343 17923 18349
rect 17865 18340 17877 18343
rect 16991 18312 17877 18340
rect 16991 18309 17003 18312
rect 16945 18303 17003 18309
rect 17865 18309 17877 18312
rect 17911 18340 17923 18343
rect 17911 18312 18644 18340
rect 17911 18309 17923 18312
rect 17865 18303 17923 18309
rect 1670 18232 1676 18284
rect 1728 18272 1734 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1728 18244 2053 18272
rect 1728 18232 1734 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2222 18272 2228 18284
rect 2183 18244 2228 18272
rect 2041 18235 2099 18241
rect 1946 18204 1952 18216
rect 1907 18176 1952 18204
rect 1946 18164 1952 18176
rect 2004 18164 2010 18216
rect 2056 18204 2084 18235
rect 2222 18232 2228 18244
rect 2280 18232 2286 18284
rect 3878 18272 3884 18284
rect 3839 18244 3884 18272
rect 3878 18232 3884 18244
rect 3936 18272 3942 18284
rect 4154 18272 4160 18284
rect 3936 18244 4160 18272
rect 3936 18232 3942 18244
rect 4154 18232 4160 18244
rect 4212 18232 4218 18284
rect 4338 18232 4344 18284
rect 4396 18272 4402 18284
rect 5537 18275 5595 18281
rect 5537 18272 5549 18275
rect 4396 18244 5549 18272
rect 4396 18232 4402 18244
rect 5537 18241 5549 18244
rect 5583 18272 5595 18275
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 5583 18244 5917 18272
rect 5583 18241 5595 18244
rect 5537 18235 5595 18241
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 7282 18232 7288 18284
rect 7340 18272 7346 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7340 18244 7389 18272
rect 7340 18232 7346 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 8662 18232 8668 18284
rect 8720 18272 8726 18284
rect 9125 18275 9183 18281
rect 9125 18272 9137 18275
rect 8720 18244 9137 18272
rect 8720 18232 8726 18244
rect 9125 18241 9137 18244
rect 9171 18241 9183 18275
rect 9125 18235 9183 18241
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10870 18272 10876 18284
rect 10367 18244 10876 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10870 18232 10876 18244
rect 10928 18272 10934 18284
rect 11422 18272 11428 18284
rect 10928 18244 11428 18272
rect 10928 18232 10934 18244
rect 11422 18232 11428 18244
rect 11480 18272 11486 18284
rect 13078 18272 13084 18284
rect 11480 18244 13084 18272
rect 11480 18232 11486 18244
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 17497 18275 17555 18281
rect 17497 18241 17509 18275
rect 17543 18272 17555 18275
rect 18322 18272 18328 18284
rect 17543 18244 18328 18272
rect 17543 18241 17555 18244
rect 17497 18235 17555 18241
rect 18322 18232 18328 18244
rect 18380 18272 18386 18284
rect 18616 18281 18644 18312
rect 18874 18300 18880 18352
rect 18932 18340 18938 18352
rect 19242 18340 19248 18352
rect 18932 18312 19248 18340
rect 18932 18300 18938 18312
rect 19242 18300 19248 18312
rect 19300 18340 19306 18352
rect 21177 18343 21235 18349
rect 21177 18340 21189 18343
rect 19300 18312 21189 18340
rect 19300 18300 19306 18312
rect 21177 18309 21189 18312
rect 21223 18340 21235 18343
rect 21266 18340 21272 18352
rect 21223 18312 21272 18340
rect 21223 18309 21235 18312
rect 21177 18303 21235 18309
rect 21266 18300 21272 18312
rect 21324 18340 21330 18352
rect 21634 18340 21640 18352
rect 21324 18312 21640 18340
rect 21324 18300 21330 18312
rect 21634 18300 21640 18312
rect 21692 18340 21698 18352
rect 22554 18340 22560 18352
rect 21692 18312 22560 18340
rect 21692 18300 21698 18312
rect 22554 18300 22560 18312
rect 22612 18300 22618 18352
rect 24121 18343 24179 18349
rect 24121 18309 24133 18343
rect 24167 18340 24179 18343
rect 25222 18340 25228 18352
rect 24167 18312 25228 18340
rect 24167 18309 24179 18312
rect 24121 18303 24179 18309
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 18509 18275 18567 18281
rect 18509 18272 18521 18275
rect 18380 18244 18521 18272
rect 18380 18232 18386 18244
rect 18509 18241 18521 18244
rect 18555 18241 18567 18275
rect 18509 18235 18567 18241
rect 18601 18275 18659 18281
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 18782 18272 18788 18284
rect 18647 18244 18788 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 20162 18272 20168 18284
rect 20123 18244 20168 18272
rect 20162 18232 20168 18244
rect 20220 18232 20226 18284
rect 22186 18272 22192 18284
rect 21468 18244 22192 18272
rect 2406 18204 2412 18216
rect 2056 18176 2412 18204
rect 2406 18164 2412 18176
rect 2464 18164 2470 18216
rect 3694 18204 3700 18216
rect 3655 18176 3700 18204
rect 3694 18164 3700 18176
rect 3752 18164 3758 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 4948 18176 5365 18204
rect 4948 18164 4954 18176
rect 5353 18173 5365 18176
rect 5399 18173 5411 18207
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 5353 18167 5411 18173
rect 6564 18176 7205 18204
rect 2130 18136 2136 18148
rect 1596 18108 2136 18136
rect 1596 18077 1624 18108
rect 2130 18096 2136 18108
rect 2188 18096 2194 18148
rect 4433 18139 4491 18145
rect 4433 18105 4445 18139
rect 4479 18136 4491 18139
rect 4479 18108 5120 18136
rect 4479 18105 4491 18108
rect 4433 18099 4491 18105
rect 5092 18080 5120 18108
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18037 1639 18071
rect 2682 18068 2688 18080
rect 2643 18040 2688 18068
rect 1581 18031 1639 18037
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 3237 18071 3295 18077
rect 3237 18037 3249 18071
rect 3283 18068 3295 18071
rect 3789 18071 3847 18077
rect 3789 18068 3801 18071
rect 3283 18040 3801 18068
rect 3283 18037 3295 18040
rect 3237 18031 3295 18037
rect 3789 18037 3801 18040
rect 3835 18068 3847 18071
rect 3970 18068 3976 18080
rect 3835 18040 3976 18068
rect 3835 18037 3847 18040
rect 3789 18031 3847 18037
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 4801 18071 4859 18077
rect 4801 18037 4813 18071
rect 4847 18068 4859 18071
rect 4890 18068 4896 18080
rect 4847 18040 4896 18068
rect 4847 18037 4859 18040
rect 4801 18031 4859 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 5074 18028 5080 18080
rect 5132 18068 5138 18080
rect 5261 18071 5319 18077
rect 5261 18068 5273 18071
rect 5132 18040 5273 18068
rect 5132 18028 5138 18040
rect 5261 18037 5273 18040
rect 5307 18037 5319 18071
rect 5261 18031 5319 18037
rect 5718 18028 5724 18080
rect 5776 18068 5782 18080
rect 6564 18077 6592 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 9306 18204 9312 18216
rect 7193 18167 7251 18173
rect 7944 18176 9312 18204
rect 6914 18096 6920 18148
rect 6972 18136 6978 18148
rect 7834 18136 7840 18148
rect 6972 18108 7840 18136
rect 6972 18096 6978 18108
rect 7834 18096 7840 18108
rect 7892 18096 7898 18148
rect 6549 18071 6607 18077
rect 6549 18068 6561 18071
rect 5776 18040 6561 18068
rect 5776 18028 5782 18040
rect 6549 18037 6561 18040
rect 6595 18037 6607 18071
rect 6549 18031 6607 18037
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 7285 18071 7343 18077
rect 7285 18068 7297 18071
rect 7064 18040 7297 18068
rect 7064 18028 7070 18040
rect 7285 18037 7297 18040
rect 7331 18068 7343 18071
rect 7944 18068 7972 18176
rect 9306 18164 9312 18176
rect 9364 18164 9370 18216
rect 9674 18204 9680 18216
rect 9635 18176 9680 18204
rect 9674 18164 9680 18176
rect 9732 18164 9738 18216
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 11146 18204 11152 18216
rect 10652 18176 11152 18204
rect 10652 18164 10658 18176
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 14274 18213 14280 18216
rect 14001 18207 14059 18213
rect 14001 18204 14013 18207
rect 11900 18176 14013 18204
rect 11900 18148 11928 18176
rect 14001 18173 14013 18176
rect 14047 18173 14059 18207
rect 14268 18204 14280 18213
rect 14235 18176 14280 18204
rect 14001 18167 14059 18173
rect 14268 18167 14280 18176
rect 8294 18096 8300 18148
rect 8352 18136 8358 18148
rect 8938 18136 8944 18148
rect 8352 18108 8944 18136
rect 8352 18096 8358 18108
rect 8938 18096 8944 18108
rect 8996 18096 9002 18148
rect 11882 18136 11888 18148
rect 11843 18108 11888 18136
rect 11882 18096 11888 18108
rect 11940 18096 11946 18148
rect 12526 18096 12532 18148
rect 12584 18136 12590 18148
rect 12897 18139 12955 18145
rect 12897 18136 12909 18139
rect 12584 18108 12909 18136
rect 12584 18096 12590 18108
rect 12897 18105 12909 18108
rect 12943 18105 12955 18139
rect 14016 18136 14044 18167
rect 14274 18164 14280 18167
rect 14332 18164 14338 18216
rect 18414 18204 18420 18216
rect 18375 18176 18420 18204
rect 18414 18164 18420 18176
rect 18472 18164 18478 18216
rect 18690 18164 18696 18216
rect 18748 18204 18754 18216
rect 19981 18207 20039 18213
rect 19981 18204 19993 18207
rect 18748 18176 19993 18204
rect 18748 18164 18754 18176
rect 19981 18173 19993 18176
rect 20027 18204 20039 18207
rect 20625 18207 20683 18213
rect 20625 18204 20637 18207
rect 20027 18176 20637 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20625 18173 20637 18176
rect 20671 18173 20683 18207
rect 20625 18167 20683 18173
rect 14642 18136 14648 18148
rect 14016 18108 14648 18136
rect 12897 18099 12955 18105
rect 14642 18096 14648 18108
rect 14700 18136 14706 18148
rect 16482 18136 16488 18148
rect 14700 18108 16488 18136
rect 14700 18096 14706 18108
rect 16482 18096 16488 18108
rect 16540 18096 16546 18148
rect 19058 18136 19064 18148
rect 19019 18108 19064 18136
rect 19058 18096 19064 18108
rect 19116 18136 19122 18148
rect 19610 18136 19616 18148
rect 19116 18108 19616 18136
rect 19116 18096 19122 18108
rect 19610 18096 19616 18108
rect 19668 18096 19674 18148
rect 21468 18136 21496 18244
rect 22186 18232 22192 18244
rect 22244 18232 22250 18284
rect 22370 18272 22376 18284
rect 22331 18244 22376 18272
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 24029 18275 24087 18281
rect 24029 18241 24041 18275
rect 24075 18272 24087 18275
rect 24670 18272 24676 18284
rect 24075 18244 24676 18272
rect 24075 18241 24087 18244
rect 24029 18235 24087 18241
rect 24670 18232 24676 18244
rect 24728 18272 24734 18284
rect 24765 18275 24823 18281
rect 24765 18272 24777 18275
rect 24728 18244 24777 18272
rect 24728 18232 24734 18244
rect 24765 18241 24777 18244
rect 24811 18272 24823 18275
rect 25700 18272 25728 18380
rect 27062 18368 27068 18380
rect 27120 18408 27126 18420
rect 27617 18411 27675 18417
rect 27617 18408 27629 18411
rect 27120 18380 27629 18408
rect 27120 18368 27126 18380
rect 27617 18377 27629 18380
rect 27663 18377 27675 18411
rect 27617 18371 27675 18377
rect 24811 18244 25728 18272
rect 24811 18241 24823 18244
rect 24765 18235 24823 18241
rect 22097 18207 22155 18213
rect 22097 18173 22109 18207
rect 22143 18204 22155 18207
rect 22278 18204 22284 18216
rect 22143 18176 22284 18204
rect 22143 18173 22155 18176
rect 22097 18167 22155 18173
rect 22278 18164 22284 18176
rect 22336 18204 22342 18216
rect 22741 18207 22799 18213
rect 22741 18204 22753 18207
rect 22336 18176 22753 18204
rect 22336 18164 22342 18176
rect 22741 18173 22753 18176
rect 22787 18173 22799 18207
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 22741 18167 22799 18173
rect 25516 18176 25697 18204
rect 21634 18136 21640 18148
rect 21468 18108 21640 18136
rect 21634 18096 21640 18108
rect 21692 18096 21698 18148
rect 25516 18080 25544 18176
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 25685 18167 25743 18173
rect 25774 18164 25780 18216
rect 25832 18204 25838 18216
rect 25952 18207 26010 18213
rect 25952 18204 25964 18207
rect 25832 18176 25964 18204
rect 25832 18164 25838 18176
rect 25952 18173 25964 18176
rect 25998 18204 26010 18207
rect 26510 18204 26516 18216
rect 25998 18176 26516 18204
rect 25998 18173 26010 18176
rect 25952 18167 26010 18173
rect 26510 18164 26516 18176
rect 26568 18204 26574 18216
rect 27154 18204 27160 18216
rect 26568 18176 27160 18204
rect 26568 18164 26574 18176
rect 27154 18164 27160 18176
rect 27212 18164 27218 18216
rect 26970 18096 26976 18148
rect 27028 18136 27034 18148
rect 27985 18139 28043 18145
rect 27985 18136 27997 18139
rect 27028 18108 27997 18136
rect 27028 18096 27034 18108
rect 27985 18105 27997 18108
rect 28031 18105 28043 18139
rect 27985 18099 28043 18105
rect 7331 18040 7972 18068
rect 8481 18071 8539 18077
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 8481 18037 8493 18071
rect 8527 18068 8539 18071
rect 8662 18068 8668 18080
rect 8527 18040 8668 18068
rect 8527 18037 8539 18040
rect 8481 18031 8539 18037
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9030 18028 9036 18080
rect 9088 18068 9094 18080
rect 9582 18068 9588 18080
rect 9088 18040 9588 18068
rect 9088 18028 9094 18040
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10042 18028 10048 18080
rect 10100 18068 10106 18080
rect 10778 18068 10784 18080
rect 10100 18040 10784 18068
rect 10100 18028 10106 18040
rect 10778 18028 10784 18040
rect 10836 18068 10842 18080
rect 11241 18071 11299 18077
rect 11241 18068 11253 18071
rect 10836 18040 11253 18068
rect 10836 18028 10842 18040
rect 11241 18037 11253 18040
rect 11287 18037 11299 18071
rect 11241 18031 11299 18037
rect 11330 18028 11336 18080
rect 11388 18068 11394 18080
rect 12161 18071 12219 18077
rect 12161 18068 12173 18071
rect 11388 18040 12173 18068
rect 11388 18028 11394 18040
rect 12161 18037 12173 18040
rect 12207 18068 12219 18071
rect 12805 18071 12863 18077
rect 12805 18068 12817 18071
rect 12207 18040 12817 18068
rect 12207 18037 12219 18040
rect 12161 18031 12219 18037
rect 12805 18037 12817 18040
rect 12851 18068 12863 18071
rect 12986 18068 12992 18080
rect 12851 18040 12992 18068
rect 12851 18037 12863 18040
rect 12805 18031 12863 18037
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13630 18068 13636 18080
rect 13591 18040 13636 18068
rect 13630 18028 13636 18040
rect 13688 18028 13694 18080
rect 15381 18071 15439 18077
rect 15381 18037 15393 18071
rect 15427 18068 15439 18071
rect 15470 18068 15476 18080
rect 15427 18040 15476 18068
rect 15427 18037 15439 18040
rect 15381 18031 15439 18037
rect 15470 18028 15476 18040
rect 15528 18028 15534 18080
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20073 18071 20131 18077
rect 20073 18068 20085 18071
rect 20036 18040 20085 18068
rect 20036 18028 20042 18040
rect 20073 18037 20085 18040
rect 20119 18037 20131 18071
rect 20073 18031 20131 18037
rect 21542 18028 21548 18080
rect 21600 18068 21606 18080
rect 21729 18071 21787 18077
rect 21729 18068 21741 18071
rect 21600 18040 21741 18068
rect 21600 18028 21606 18040
rect 21729 18037 21741 18040
rect 21775 18037 21787 18071
rect 24486 18068 24492 18080
rect 24447 18040 24492 18068
rect 21729 18031 21787 18037
rect 24486 18028 24492 18040
rect 24544 18028 24550 18080
rect 24578 18028 24584 18080
rect 24636 18068 24642 18080
rect 25498 18068 25504 18080
rect 24636 18040 24681 18068
rect 25459 18040 25504 18068
rect 24636 18028 24642 18040
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 1673 17867 1731 17873
rect 1673 17833 1685 17867
rect 1719 17864 1731 17867
rect 2498 17864 2504 17876
rect 1719 17836 2504 17864
rect 1719 17833 1731 17836
rect 1673 17827 1731 17833
rect 2498 17824 2504 17836
rect 2556 17824 2562 17876
rect 2682 17864 2688 17876
rect 2643 17836 2688 17864
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 3421 17867 3479 17873
rect 3421 17833 3433 17867
rect 3467 17864 3479 17867
rect 3694 17864 3700 17876
rect 3467 17836 3700 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 3694 17824 3700 17836
rect 3752 17824 3758 17876
rect 4338 17864 4344 17876
rect 4299 17836 4344 17864
rect 4338 17824 4344 17836
rect 4396 17824 4402 17876
rect 4798 17864 4804 17876
rect 4759 17836 4804 17864
rect 4798 17824 4804 17836
rect 4856 17824 4862 17876
rect 5534 17824 5540 17876
rect 5592 17864 5598 17876
rect 6365 17867 6423 17873
rect 6365 17864 6377 17867
rect 5592 17836 6377 17864
rect 5592 17824 5598 17836
rect 6365 17833 6377 17836
rect 6411 17864 6423 17867
rect 6822 17864 6828 17876
rect 6411 17836 6828 17864
rect 6411 17833 6423 17836
rect 6365 17827 6423 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 7650 17864 7656 17876
rect 7611 17836 7656 17864
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 10870 17864 10876 17876
rect 10831 17836 10876 17864
rect 10870 17824 10876 17836
rect 10928 17824 10934 17876
rect 12897 17867 12955 17873
rect 12897 17833 12909 17867
rect 12943 17864 12955 17867
rect 13078 17864 13084 17876
rect 12943 17836 13084 17864
rect 12943 17833 12955 17836
rect 12897 17827 12955 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13722 17864 13728 17876
rect 13679 17836 13728 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13722 17824 13728 17836
rect 13780 17824 13786 17876
rect 14001 17867 14059 17873
rect 14001 17833 14013 17867
rect 14047 17864 14059 17867
rect 14274 17864 14280 17876
rect 14047 17836 14280 17864
rect 14047 17833 14059 17836
rect 14001 17827 14059 17833
rect 14274 17824 14280 17836
rect 14332 17864 14338 17876
rect 14918 17864 14924 17876
rect 14332 17836 14924 17864
rect 14332 17824 14338 17836
rect 14918 17824 14924 17836
rect 14976 17824 14982 17876
rect 15194 17824 15200 17876
rect 15252 17864 15258 17876
rect 15289 17867 15347 17873
rect 15289 17864 15301 17867
rect 15252 17836 15301 17864
rect 15252 17824 15258 17836
rect 15289 17833 15301 17836
rect 15335 17833 15347 17867
rect 15289 17827 15347 17833
rect 17586 17824 17592 17876
rect 17644 17864 17650 17876
rect 18049 17867 18107 17873
rect 18049 17864 18061 17867
rect 17644 17836 18061 17864
rect 17644 17824 17650 17836
rect 18049 17833 18061 17836
rect 18095 17833 18107 17867
rect 18049 17827 18107 17833
rect 18966 17824 18972 17876
rect 19024 17864 19030 17876
rect 19153 17867 19211 17873
rect 19153 17864 19165 17867
rect 19024 17836 19165 17864
rect 19024 17824 19030 17836
rect 19153 17833 19165 17836
rect 19199 17833 19211 17867
rect 20162 17864 20168 17876
rect 20123 17836 20168 17864
rect 19153 17827 19211 17833
rect 20162 17824 20168 17836
rect 20220 17824 20226 17876
rect 20993 17867 21051 17873
rect 20993 17833 21005 17867
rect 21039 17864 21051 17867
rect 21910 17864 21916 17876
rect 21039 17836 21916 17864
rect 21039 17833 21051 17836
rect 20993 17827 21051 17833
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 22370 17864 22376 17876
rect 22331 17836 22376 17864
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 25222 17864 25228 17876
rect 25183 17836 25228 17864
rect 25222 17824 25228 17836
rect 25280 17824 25286 17876
rect 25406 17824 25412 17876
rect 25464 17864 25470 17876
rect 25685 17867 25743 17873
rect 25685 17864 25697 17867
rect 25464 17836 25697 17864
rect 25464 17824 25470 17836
rect 25685 17833 25697 17836
rect 25731 17833 25743 17867
rect 26326 17864 26332 17876
rect 26287 17836 26332 17864
rect 25685 17827 25743 17833
rect 26326 17824 26332 17836
rect 26384 17824 26390 17876
rect 26513 17867 26571 17873
rect 26513 17833 26525 17867
rect 26559 17864 26571 17867
rect 26970 17864 26976 17876
rect 26559 17836 26976 17864
rect 26559 17833 26571 17836
rect 26513 17827 26571 17833
rect 26970 17824 26976 17836
rect 27028 17824 27034 17876
rect 4154 17756 4160 17808
rect 4212 17796 4218 17808
rect 5258 17805 5264 17808
rect 5230 17799 5264 17805
rect 5230 17796 5242 17799
rect 4212 17768 5242 17796
rect 4212 17756 4218 17768
rect 5230 17765 5242 17768
rect 5316 17796 5322 17808
rect 6917 17799 6975 17805
rect 6917 17796 6929 17799
rect 5316 17768 6929 17796
rect 5230 17759 5264 17765
rect 5258 17756 5264 17759
rect 5316 17756 5322 17768
rect 6917 17765 6929 17768
rect 6963 17796 6975 17799
rect 7282 17796 7288 17808
rect 6963 17768 7288 17796
rect 6963 17765 6975 17768
rect 6917 17759 6975 17765
rect 7282 17756 7288 17768
rect 7340 17756 7346 17808
rect 7377 17799 7435 17805
rect 7377 17765 7389 17799
rect 7423 17796 7435 17799
rect 7742 17796 7748 17808
rect 7423 17768 7748 17796
rect 7423 17765 7435 17768
rect 7377 17759 7435 17765
rect 7742 17756 7748 17768
rect 7800 17756 7806 17808
rect 10413 17799 10471 17805
rect 10413 17765 10425 17799
rect 10459 17796 10471 17799
rect 13541 17799 13599 17805
rect 13541 17796 13553 17799
rect 10459 17768 13553 17796
rect 10459 17765 10471 17768
rect 10413 17759 10471 17765
rect 13541 17765 13553 17768
rect 13587 17796 13599 17799
rect 13906 17796 13912 17808
rect 13587 17768 13912 17796
rect 13587 17765 13599 17768
rect 13541 17759 13599 17765
rect 13906 17756 13912 17768
rect 13964 17756 13970 17808
rect 14642 17796 14648 17808
rect 14603 17768 14648 17796
rect 14642 17756 14648 17768
rect 14700 17756 14706 17808
rect 21450 17796 21456 17808
rect 21411 17768 21456 17796
rect 21450 17756 21456 17768
rect 21508 17756 21514 17808
rect 21652 17768 22784 17796
rect 2041 17731 2099 17737
rect 2041 17697 2053 17731
rect 2087 17728 2099 17731
rect 2087 17700 3832 17728
rect 2087 17697 2099 17700
rect 2041 17691 2099 17697
rect 2130 17660 2136 17672
rect 2091 17632 2136 17660
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2314 17660 2320 17672
rect 2227 17632 2320 17660
rect 2314 17620 2320 17632
rect 2372 17660 2378 17672
rect 2682 17660 2688 17672
rect 2372 17632 2688 17660
rect 2372 17620 2378 17632
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 3804 17533 3832 17700
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 4856 17700 4997 17728
rect 4856 17688 4862 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 4985 17691 5043 17697
rect 8294 17688 8300 17740
rect 8352 17728 8358 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 8352 17700 8401 17728
rect 8352 17688 8358 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 12066 17728 12072 17740
rect 11839 17700 12072 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 12066 17688 12072 17700
rect 12124 17688 12130 17740
rect 13814 17688 13820 17740
rect 13872 17728 13878 17740
rect 14093 17731 14151 17737
rect 14093 17728 14105 17731
rect 13872 17700 14105 17728
rect 13872 17688 13878 17700
rect 14093 17697 14105 17700
rect 14139 17697 14151 17731
rect 14093 17691 14151 17697
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 16942 17737 16948 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16540 17700 16681 17728
rect 16540 17688 16546 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16936 17728 16948 17737
rect 16903 17700 16948 17728
rect 16669 17691 16727 17697
rect 16936 17691 16948 17700
rect 16942 17688 16948 17691
rect 17000 17688 17006 17740
rect 19518 17728 19524 17740
rect 19479 17700 19524 17728
rect 19518 17688 19524 17700
rect 19576 17688 19582 17740
rect 20717 17731 20775 17737
rect 20717 17697 20729 17731
rect 20763 17728 20775 17731
rect 21358 17728 21364 17740
rect 20763 17700 21364 17728
rect 20763 17697 20775 17700
rect 20717 17691 20775 17697
rect 21358 17688 21364 17700
rect 21416 17688 21422 17740
rect 8478 17660 8484 17672
rect 8439 17632 8484 17660
rect 8478 17620 8484 17632
rect 8536 17620 8542 17672
rect 8662 17660 8668 17672
rect 8623 17632 8668 17660
rect 8662 17620 8668 17632
rect 8720 17620 8726 17672
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11885 17663 11943 17669
rect 11885 17660 11897 17663
rect 11664 17632 11897 17660
rect 11664 17620 11670 17632
rect 11885 17629 11897 17632
rect 11931 17629 11943 17663
rect 11885 17623 11943 17629
rect 11977 17663 12035 17669
rect 11977 17629 11989 17663
rect 12023 17660 12035 17663
rect 12158 17660 12164 17672
rect 12023 17632 12164 17660
rect 12023 17629 12035 17632
rect 11977 17623 12035 17629
rect 10594 17552 10600 17604
rect 10652 17592 10658 17604
rect 11333 17595 11391 17601
rect 11333 17592 11345 17595
rect 10652 17564 11345 17592
rect 10652 17552 10658 17564
rect 11333 17561 11345 17564
rect 11379 17592 11391 17595
rect 11992 17592 12020 17623
rect 12158 17620 12164 17632
rect 12216 17620 12222 17672
rect 14182 17660 14188 17672
rect 14143 17632 14188 17660
rect 14182 17620 14188 17632
rect 14240 17620 14246 17672
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 19613 17663 19671 17669
rect 19613 17660 19625 17663
rect 18656 17632 19625 17660
rect 18656 17620 18662 17632
rect 19613 17629 19625 17632
rect 19659 17629 19671 17663
rect 19613 17623 19671 17629
rect 19705 17663 19763 17669
rect 19705 17629 19717 17663
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 11379 17564 12020 17592
rect 11379 17561 11391 17564
rect 11333 17555 11391 17561
rect 19058 17552 19064 17604
rect 19116 17592 19122 17604
rect 19720 17592 19748 17623
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 21652 17669 21680 17768
rect 22554 17728 22560 17740
rect 22515 17700 22560 17728
rect 22554 17688 22560 17700
rect 22612 17688 22618 17740
rect 22756 17728 22784 17768
rect 22824 17731 22882 17737
rect 22824 17728 22836 17731
rect 22756 17700 22836 17728
rect 22824 17697 22836 17700
rect 22870 17728 22882 17731
rect 23382 17728 23388 17740
rect 22870 17700 23388 17728
rect 22870 17697 22882 17700
rect 22824 17691 22882 17697
rect 23382 17688 23388 17700
rect 23440 17688 23446 17740
rect 26878 17728 26884 17740
rect 26839 17700 26884 17728
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 21637 17663 21695 17669
rect 21637 17660 21649 17663
rect 21140 17632 21649 17660
rect 21140 17620 21146 17632
rect 21637 17629 21649 17632
rect 21683 17629 21695 17663
rect 21637 17623 21695 17629
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 26973 17663 27031 17669
rect 26973 17660 26985 17663
rect 26844 17632 26985 17660
rect 26844 17620 26850 17632
rect 26973 17629 26985 17632
rect 27019 17629 27031 17663
rect 27154 17660 27160 17672
rect 27115 17632 27160 17660
rect 26973 17623 27031 17629
rect 27154 17620 27160 17632
rect 27212 17620 27218 17672
rect 19116 17564 19748 17592
rect 24581 17595 24639 17601
rect 19116 17552 19122 17564
rect 24581 17561 24593 17595
rect 24627 17592 24639 17595
rect 24762 17592 24768 17604
rect 24627 17564 24768 17592
rect 24627 17561 24639 17564
rect 24581 17555 24639 17561
rect 24762 17552 24768 17564
rect 24820 17552 24826 17604
rect 3789 17527 3847 17533
rect 3789 17493 3801 17527
rect 3835 17524 3847 17527
rect 4062 17524 4068 17536
rect 3835 17496 4068 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 4062 17484 4068 17496
rect 4120 17484 4126 17536
rect 7834 17484 7840 17536
rect 7892 17524 7898 17536
rect 8021 17527 8079 17533
rect 8021 17524 8033 17527
rect 7892 17496 8033 17524
rect 7892 17484 7898 17496
rect 8021 17493 8033 17496
rect 8067 17493 8079 17527
rect 9950 17524 9956 17536
rect 9911 17496 9956 17524
rect 8021 17487 8079 17493
rect 9950 17484 9956 17496
rect 10008 17484 10014 17536
rect 11422 17524 11428 17536
rect 11383 17496 11428 17524
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 12526 17524 12532 17536
rect 12487 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 18782 17524 18788 17536
rect 18743 17496 18788 17524
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22278 17524 22284 17536
rect 22143 17496 22284 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 23842 17484 23848 17536
rect 23900 17524 23906 17536
rect 23937 17527 23995 17533
rect 23937 17524 23949 17527
rect 23900 17496 23949 17524
rect 23900 17484 23906 17496
rect 23937 17493 23949 17496
rect 23983 17493 23995 17527
rect 24854 17524 24860 17536
rect 24815 17496 24860 17524
rect 23937 17487 23995 17493
rect 24854 17484 24860 17496
rect 24912 17484 24918 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2130 17280 2136 17332
rect 2188 17320 2194 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 2188 17292 3709 17320
rect 2188 17280 2194 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 5258 17280 5264 17332
rect 5316 17320 5322 17332
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 5316 17292 5641 17320
rect 5316 17280 5322 17292
rect 5629 17289 5641 17292
rect 5675 17320 5687 17323
rect 6181 17323 6239 17329
rect 6181 17320 6193 17323
rect 5675 17292 6193 17320
rect 5675 17289 5687 17292
rect 5629 17283 5687 17289
rect 6181 17289 6193 17292
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 7653 17323 7711 17329
rect 7653 17289 7665 17323
rect 7699 17320 7711 17323
rect 7926 17320 7932 17332
rect 7699 17292 7932 17320
rect 7699 17289 7711 17292
rect 7653 17283 7711 17289
rect 7926 17280 7932 17292
rect 7984 17280 7990 17332
rect 10594 17320 10600 17332
rect 8036 17292 8248 17320
rect 10555 17292 10600 17320
rect 3145 17255 3203 17261
rect 3145 17221 3157 17255
rect 3191 17221 3203 17255
rect 3145 17215 3203 17221
rect 7561 17255 7619 17261
rect 7561 17221 7573 17255
rect 7607 17252 7619 17255
rect 8036 17252 8064 17292
rect 7607 17224 8064 17252
rect 7607 17221 7619 17224
rect 7561 17215 7619 17221
rect 3160 17184 3188 17215
rect 8110 17212 8116 17264
rect 8168 17212 8174 17264
rect 3160 17156 4384 17184
rect 4356 17128 4384 17156
rect 1765 17119 1823 17125
rect 1765 17116 1777 17119
rect 1688 17088 1777 17116
rect 1688 16992 1716 17088
rect 1765 17085 1777 17088
rect 1811 17085 1823 17119
rect 1765 17079 1823 17085
rect 2032 17119 2090 17125
rect 2032 17085 2044 17119
rect 2078 17116 2090 17119
rect 2314 17116 2320 17128
rect 2078 17088 2320 17116
rect 2078 17085 2090 17088
rect 2032 17079 2090 17085
rect 2314 17076 2320 17088
rect 2372 17076 2378 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 4157 17051 4215 17057
rect 4157 17017 4169 17051
rect 4203 17048 4215 17051
rect 4264 17048 4292 17079
rect 4338 17076 4344 17128
rect 4396 17116 4402 17128
rect 4505 17119 4563 17125
rect 4505 17116 4517 17119
rect 4396 17088 4517 17116
rect 4396 17076 4402 17088
rect 4505 17085 4517 17088
rect 4551 17085 4563 17119
rect 4505 17079 4563 17085
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17116 6699 17119
rect 7834 17116 7840 17128
rect 6687 17088 7840 17116
rect 6687 17085 6699 17088
rect 6641 17079 6699 17085
rect 7834 17076 7840 17088
rect 7892 17116 7898 17128
rect 8128 17125 8156 17212
rect 8220 17193 8248 17292
rect 10594 17280 10600 17292
rect 10652 17280 10658 17332
rect 11974 17280 11980 17332
rect 12032 17320 12038 17332
rect 12161 17323 12219 17329
rect 12161 17320 12173 17323
rect 12032 17292 12173 17320
rect 12032 17280 12038 17292
rect 12161 17289 12173 17292
rect 12207 17289 12219 17323
rect 12161 17283 12219 17289
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12492 17292 12537 17320
rect 12492 17280 12498 17292
rect 13078 17280 13084 17332
rect 13136 17320 13142 17332
rect 13449 17323 13507 17329
rect 13449 17320 13461 17323
rect 13136 17292 13461 17320
rect 13136 17280 13142 17292
rect 13449 17289 13461 17292
rect 13495 17289 13507 17323
rect 13449 17283 13507 17289
rect 13909 17323 13967 17329
rect 13909 17289 13921 17323
rect 13955 17320 13967 17323
rect 14182 17320 14188 17332
rect 13955 17292 14188 17320
rect 13955 17289 13967 17292
rect 13909 17283 13967 17289
rect 14182 17280 14188 17292
rect 14240 17320 14246 17332
rect 16485 17323 16543 17329
rect 16485 17320 16497 17323
rect 14240 17292 16497 17320
rect 14240 17280 14246 17292
rect 16485 17289 16497 17292
rect 16531 17320 16543 17323
rect 16942 17320 16948 17332
rect 16531 17292 16948 17320
rect 16531 17289 16543 17292
rect 16485 17283 16543 17289
rect 16942 17280 16948 17292
rect 17000 17320 17006 17332
rect 17405 17323 17463 17329
rect 17405 17320 17417 17323
rect 17000 17292 17417 17320
rect 17000 17280 17006 17292
rect 17405 17289 17417 17292
rect 17451 17289 17463 17323
rect 17405 17283 17463 17289
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 17773 17323 17831 17329
rect 17773 17320 17785 17323
rect 17644 17292 17785 17320
rect 17644 17280 17650 17292
rect 17773 17289 17785 17292
rect 17819 17320 17831 17323
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 17819 17292 18245 17320
rect 17819 17289 17831 17292
rect 17773 17283 17831 17289
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 18233 17283 18291 17289
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 9122 17184 9128 17196
rect 8251 17156 9128 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 9122 17144 9128 17156
rect 9180 17184 9186 17196
rect 9180 17156 9352 17184
rect 9180 17144 9186 17156
rect 8021 17119 8079 17125
rect 8021 17116 8033 17119
rect 7892 17088 8033 17116
rect 7892 17076 7898 17088
rect 8021 17085 8033 17088
rect 8067 17085 8079 17119
rect 8021 17079 8079 17085
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8113 17079 8171 17085
rect 9048 17088 9229 17116
rect 4798 17048 4804 17060
rect 4203 17020 4804 17048
rect 4203 17017 4215 17020
rect 4157 17011 4215 17017
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 7193 17051 7251 17057
rect 7193 17017 7205 17051
rect 7239 17048 7251 17051
rect 8478 17048 8484 17060
rect 7239 17020 8484 17048
rect 7239 17017 7251 17020
rect 7193 17011 7251 17017
rect 8478 17008 8484 17020
rect 8536 17008 8542 17060
rect 9048 16992 9076 17088
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 9324 17116 9352 17156
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 13096 17193 13124 17280
rect 14642 17212 14648 17264
rect 14700 17252 14706 17264
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 14700 17224 14933 17252
rect 14700 17212 14706 17224
rect 14921 17221 14933 17224
rect 14967 17252 14979 17255
rect 14967 17224 15148 17252
rect 14967 17221 14979 17224
rect 14921 17215 14979 17221
rect 15120 17196 15148 17224
rect 13081 17187 13139 17193
rect 11480 17156 12940 17184
rect 11480 17144 11486 17156
rect 9473 17119 9531 17125
rect 9473 17116 9485 17119
rect 9324 17088 9485 17116
rect 9217 17079 9275 17085
rect 9473 17085 9485 17088
rect 9519 17085 9531 17119
rect 9473 17079 9531 17085
rect 11974 17008 11980 17060
rect 12032 17048 12038 17060
rect 12912 17057 12940 17156
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 15102 17184 15108 17196
rect 15015 17156 15108 17184
rect 13081 17147 13139 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 17037 17187 17095 17193
rect 17037 17184 17049 17187
rect 16540 17156 17049 17184
rect 16540 17144 16546 17156
rect 17037 17153 17049 17156
rect 17083 17153 17095 17187
rect 18248 17184 18276 17283
rect 20162 17280 20168 17292
rect 20220 17280 20226 17332
rect 21082 17320 21088 17332
rect 21043 17292 21088 17320
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 22554 17280 22560 17332
rect 22612 17320 22618 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22612 17292 23029 17320
rect 22612 17280 22618 17292
rect 23017 17289 23029 17292
rect 23063 17320 23075 17323
rect 23198 17320 23204 17332
rect 23063 17292 23204 17320
rect 23063 17289 23075 17292
rect 23017 17283 23075 17289
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 23382 17320 23388 17332
rect 23343 17292 23388 17320
rect 23382 17280 23388 17292
rect 23440 17280 23446 17332
rect 23934 17320 23940 17332
rect 23895 17292 23940 17320
rect 23934 17280 23940 17292
rect 23992 17280 23998 17332
rect 24121 17323 24179 17329
rect 24121 17289 24133 17323
rect 24167 17320 24179 17323
rect 24486 17320 24492 17332
rect 24167 17292 24492 17320
rect 24167 17289 24179 17292
rect 24121 17283 24179 17289
rect 24486 17280 24492 17292
rect 24544 17320 24550 17332
rect 24854 17320 24860 17332
rect 24544 17292 24860 17320
rect 24544 17280 24550 17292
rect 24854 17280 24860 17292
rect 24912 17280 24918 17332
rect 26786 17280 26792 17332
rect 26844 17320 26850 17332
rect 27985 17323 28043 17329
rect 27985 17320 27997 17323
rect 26844 17292 27997 17320
rect 26844 17280 26850 17292
rect 27985 17289 27997 17292
rect 28031 17289 28043 17323
rect 27985 17283 28043 17289
rect 23216 17252 23244 17280
rect 25498 17252 25504 17264
rect 23216 17224 25504 17252
rect 25498 17212 25504 17224
rect 25556 17252 25562 17264
rect 25556 17224 25728 17252
rect 25556 17212 25562 17224
rect 25700 17196 25728 17224
rect 26878 17212 26884 17264
rect 26936 17252 26942 17264
rect 27617 17255 27675 17261
rect 27617 17252 27629 17255
rect 26936 17224 27629 17252
rect 26936 17212 26942 17224
rect 27617 17221 27629 17224
rect 27663 17252 27675 17255
rect 27663 17224 28028 17252
rect 27663 17221 27675 17224
rect 27617 17215 27675 17221
rect 28000 17196 28028 17224
rect 21545 17187 21603 17193
rect 18248 17156 18920 17184
rect 17037 17147 17095 17153
rect 17052 17116 17080 17147
rect 18782 17116 18788 17128
rect 17052 17088 18788 17116
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 18892 17116 18920 17156
rect 21545 17153 21557 17187
rect 21591 17184 21603 17187
rect 22649 17187 22707 17193
rect 22649 17184 22661 17187
rect 21591 17156 22661 17184
rect 21591 17153 21603 17156
rect 21545 17147 21603 17153
rect 22649 17153 22661 17156
rect 22695 17184 22707 17187
rect 23014 17184 23020 17196
rect 22695 17156 23020 17184
rect 22695 17153 22707 17156
rect 22649 17147 22707 17153
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 24762 17184 24768 17196
rect 24723 17156 24768 17184
rect 24762 17144 24768 17156
rect 24820 17144 24826 17196
rect 25682 17184 25688 17196
rect 25595 17156 25688 17184
rect 25682 17144 25688 17156
rect 25740 17144 25746 17196
rect 27982 17144 27988 17196
rect 28040 17144 28046 17196
rect 19058 17125 19064 17128
rect 19041 17119 19064 17125
rect 19041 17116 19053 17119
rect 18892 17088 19053 17116
rect 19041 17085 19053 17088
rect 19116 17116 19122 17128
rect 19116 17088 19189 17116
rect 19041 17079 19064 17085
rect 19058 17076 19064 17079
rect 19116 17076 19122 17088
rect 23934 17076 23940 17128
rect 23992 17116 23998 17128
rect 24489 17119 24547 17125
rect 24489 17116 24501 17119
rect 23992 17088 24501 17116
rect 23992 17076 23998 17088
rect 24489 17085 24501 17088
rect 24535 17085 24547 17119
rect 24489 17079 24547 17085
rect 12897 17051 12955 17057
rect 12032 17020 12756 17048
rect 12032 17008 12038 17020
rect 12728 16992 12756 17020
rect 12897 17017 12909 17051
rect 12943 17048 12955 17051
rect 14185 17051 14243 17057
rect 14185 17048 14197 17051
rect 12943 17020 14197 17048
rect 12943 17017 12955 17020
rect 12897 17011 12955 17017
rect 14185 17017 14197 17020
rect 14231 17017 14243 17051
rect 15350 17051 15408 17057
rect 15350 17048 15362 17051
rect 14185 17011 14243 17017
rect 14568 17020 15362 17048
rect 14568 16992 14596 17020
rect 15350 17017 15362 17020
rect 15396 17048 15408 17051
rect 16666 17048 16672 17060
rect 15396 17020 16672 17048
rect 15396 17017 15408 17020
rect 15350 17011 15408 17017
rect 16666 17008 16672 17020
rect 16724 17008 16730 17060
rect 22462 17048 22468 17060
rect 21836 17020 22468 17048
rect 1670 16980 1676 16992
rect 1631 16952 1676 16980
rect 1670 16940 1676 16952
rect 1728 16940 1734 16992
rect 7926 16940 7932 16992
rect 7984 16980 7990 16992
rect 8662 16980 8668 16992
rect 7984 16952 8668 16980
rect 7984 16940 7990 16952
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 11517 16983 11575 16989
rect 11517 16949 11529 16983
rect 11563 16980 11575 16983
rect 11606 16980 11612 16992
rect 11563 16952 11612 16980
rect 11563 16949 11575 16952
rect 11517 16943 11575 16949
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 12066 16980 12072 16992
rect 11931 16952 12072 16980
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12710 16940 12716 16992
rect 12768 16980 12774 16992
rect 12805 16983 12863 16989
rect 12805 16980 12817 16983
rect 12768 16952 12817 16980
rect 12768 16940 12774 16952
rect 12805 16949 12817 16952
rect 12851 16949 12863 16983
rect 14550 16980 14556 16992
rect 14511 16952 14556 16980
rect 12805 16943 12863 16949
rect 14550 16940 14556 16952
rect 14608 16940 14614 16992
rect 18598 16980 18604 16992
rect 18559 16952 18604 16980
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 20806 16940 20812 16992
rect 20864 16980 20870 16992
rect 21836 16989 21864 17020
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 25406 17008 25412 17060
rect 25464 17048 25470 17060
rect 25930 17051 25988 17057
rect 25930 17048 25942 17051
rect 25464 17020 25942 17048
rect 25464 17008 25470 17020
rect 25930 17017 25942 17020
rect 25976 17017 25988 17051
rect 25930 17011 25988 17017
rect 21821 16983 21879 16989
rect 21821 16980 21833 16983
rect 20864 16952 21833 16980
rect 20864 16940 20870 16952
rect 21821 16949 21833 16952
rect 21867 16949 21879 16983
rect 22002 16980 22008 16992
rect 21963 16952 22008 16980
rect 21821 16943 21879 16949
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 22278 16940 22284 16992
rect 22336 16980 22342 16992
rect 22373 16983 22431 16989
rect 22373 16980 22385 16983
rect 22336 16952 22385 16980
rect 22336 16940 22342 16952
rect 22373 16949 22385 16952
rect 22419 16949 22431 16983
rect 22373 16943 22431 16949
rect 24578 16940 24584 16992
rect 24636 16980 24642 16992
rect 25133 16983 25191 16989
rect 25133 16980 25145 16983
rect 24636 16952 25145 16980
rect 24636 16940 24642 16952
rect 25133 16949 25145 16952
rect 25179 16949 25191 16983
rect 25133 16943 25191 16949
rect 26418 16940 26424 16992
rect 26476 16980 26482 16992
rect 27065 16983 27123 16989
rect 27065 16980 27077 16983
rect 26476 16952 27077 16980
rect 26476 16940 26482 16952
rect 27065 16949 27077 16952
rect 27111 16949 27123 16983
rect 27065 16943 27123 16949
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16736 1676 16788
rect 1728 16736 1734 16788
rect 2314 16736 2320 16788
rect 2372 16776 2378 16788
rect 2869 16779 2927 16785
rect 2869 16776 2881 16779
rect 2372 16748 2881 16776
rect 2372 16736 2378 16748
rect 2869 16745 2881 16748
rect 2915 16745 2927 16779
rect 2869 16739 2927 16745
rect 4798 16736 4804 16788
rect 4856 16776 4862 16788
rect 4985 16779 5043 16785
rect 4985 16776 4997 16779
rect 4856 16748 4997 16776
rect 4856 16736 4862 16748
rect 4985 16745 4997 16748
rect 5031 16745 5043 16779
rect 7926 16776 7932 16788
rect 7887 16748 7932 16776
rect 4985 16739 5043 16745
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16640 1547 16643
rect 1688 16640 1716 16736
rect 1756 16711 1814 16717
rect 1756 16677 1768 16711
rect 1802 16708 1814 16711
rect 2222 16708 2228 16720
rect 1802 16680 2228 16708
rect 1802 16677 1814 16680
rect 1756 16671 1814 16677
rect 2222 16668 2228 16680
rect 2280 16708 2286 16720
rect 3050 16708 3056 16720
rect 2280 16680 3056 16708
rect 2280 16668 2286 16680
rect 3050 16668 3056 16680
rect 3108 16708 3114 16720
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 3108 16680 3801 16708
rect 3108 16668 3114 16680
rect 3789 16677 3801 16680
rect 3835 16677 3847 16711
rect 3789 16671 3847 16677
rect 1535 16612 1716 16640
rect 5000 16640 5028 16739
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8021 16779 8079 16785
rect 8021 16745 8033 16779
rect 8067 16776 8079 16779
rect 8478 16776 8484 16788
rect 8067 16748 8484 16776
rect 8067 16745 8079 16748
rect 8021 16739 8079 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 9122 16736 9128 16788
rect 9180 16776 9186 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 9180 16748 9229 16776
rect 9180 16736 9186 16748
rect 9217 16745 9229 16748
rect 9263 16745 9275 16779
rect 9674 16776 9680 16788
rect 9635 16748 9680 16776
rect 9217 16739 9275 16745
rect 5350 16668 5356 16720
rect 5408 16717 5414 16720
rect 5408 16711 5472 16717
rect 5408 16677 5426 16711
rect 5460 16677 5472 16711
rect 5408 16671 5472 16677
rect 7193 16711 7251 16717
rect 7193 16677 7205 16711
rect 7239 16708 7251 16711
rect 8110 16708 8116 16720
rect 7239 16680 8116 16708
rect 7239 16677 7251 16680
rect 7193 16671 7251 16677
rect 5408 16668 5414 16671
rect 8110 16668 8116 16680
rect 8168 16668 8174 16720
rect 8294 16708 8300 16720
rect 8207 16680 8300 16708
rect 8294 16668 8300 16680
rect 8352 16708 8358 16720
rect 9232 16708 9260 16739
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 10137 16779 10195 16785
rect 10137 16776 10149 16779
rect 10008 16748 10149 16776
rect 10008 16736 10014 16748
rect 10137 16745 10149 16748
rect 10183 16745 10195 16779
rect 10137 16739 10195 16745
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 13078 16776 13084 16788
rect 12851 16748 13084 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 13538 16776 13544 16788
rect 13499 16748 13544 16776
rect 13538 16736 13544 16748
rect 13596 16776 13602 16788
rect 13906 16776 13912 16788
rect 13596 16748 13912 16776
rect 13596 16736 13602 16748
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 14274 16776 14280 16788
rect 14235 16748 14280 16776
rect 14274 16736 14280 16748
rect 14332 16736 14338 16788
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 18506 16776 18512 16788
rect 18467 16748 18512 16776
rect 18506 16736 18512 16748
rect 18564 16736 18570 16788
rect 20717 16779 20775 16785
rect 20717 16745 20729 16779
rect 20763 16776 20775 16779
rect 21450 16776 21456 16788
rect 20763 16748 21456 16776
rect 20763 16745 20775 16748
rect 20717 16739 20775 16745
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 22554 16776 22560 16788
rect 22467 16748 22560 16776
rect 22554 16736 22560 16748
rect 22612 16776 22618 16788
rect 23106 16776 23112 16788
rect 22612 16748 23112 16776
rect 22612 16736 22618 16748
rect 23106 16736 23112 16748
rect 23164 16736 23170 16788
rect 24762 16736 24768 16788
rect 24820 16776 24826 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 24820 16748 25329 16776
rect 24820 16736 24826 16748
rect 25317 16745 25329 16748
rect 25363 16745 25375 16779
rect 25866 16776 25872 16788
rect 25827 16748 25872 16776
rect 25317 16739 25375 16745
rect 9582 16708 9588 16720
rect 8352 16680 8892 16708
rect 9232 16680 9588 16708
rect 8352 16668 8358 16680
rect 5166 16640 5172 16652
rect 5000 16612 5172 16640
rect 1535 16609 1547 16612
rect 1489 16603 1547 16609
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 7561 16643 7619 16649
rect 7561 16609 7573 16643
rect 7607 16640 7619 16643
rect 8312 16640 8340 16668
rect 7607 16612 8340 16640
rect 8389 16643 8447 16649
rect 7607 16609 7619 16612
rect 7561 16603 7619 16609
rect 8389 16609 8401 16643
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 8481 16643 8539 16649
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 8864 16640 8892 16680
rect 9582 16668 9588 16680
rect 9640 16668 9646 16720
rect 10045 16711 10103 16717
rect 10045 16677 10057 16711
rect 10091 16708 10103 16711
rect 10318 16708 10324 16720
rect 10091 16680 10324 16708
rect 10091 16677 10103 16680
rect 10045 16671 10103 16677
rect 10318 16668 10324 16680
rect 10376 16668 10382 16720
rect 11882 16708 11888 16720
rect 11440 16680 11888 16708
rect 10778 16640 10784 16652
rect 8527 16612 8800 16640
rect 8864 16612 9628 16640
rect 10739 16612 10784 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 3510 16532 3516 16584
rect 3568 16572 3574 16584
rect 4065 16575 4123 16581
rect 4065 16572 4077 16575
rect 3568 16544 4077 16572
rect 3568 16532 3574 16544
rect 4065 16541 4077 16544
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 8110 16532 8116 16584
rect 8168 16572 8174 16584
rect 8404 16572 8432 16603
rect 8168 16544 8432 16572
rect 8665 16575 8723 16581
rect 8168 16532 8174 16544
rect 8665 16541 8677 16575
rect 8711 16541 8723 16575
rect 8772 16572 8800 16612
rect 8846 16572 8852 16584
rect 8772 16544 8852 16572
rect 8665 16535 8723 16541
rect 8680 16504 8708 16535
rect 8846 16532 8852 16544
rect 8904 16532 8910 16584
rect 9600 16572 9628 16612
rect 10778 16600 10784 16612
rect 10836 16600 10842 16652
rect 11440 16649 11468 16680
rect 11882 16668 11888 16680
rect 11940 16668 11946 16720
rect 15105 16711 15163 16717
rect 15105 16677 15117 16711
rect 15151 16708 15163 16711
rect 15556 16711 15614 16717
rect 15556 16708 15568 16711
rect 15151 16680 15568 16708
rect 15151 16677 15163 16680
rect 15105 16671 15163 16677
rect 15556 16677 15568 16680
rect 15602 16708 15614 16711
rect 15838 16708 15844 16720
rect 15602 16680 15844 16708
rect 15602 16677 15614 16680
rect 15556 16671 15614 16677
rect 15838 16668 15844 16680
rect 15896 16668 15902 16720
rect 18966 16708 18972 16720
rect 18708 16680 18972 16708
rect 11425 16643 11483 16649
rect 11425 16609 11437 16643
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 11692 16643 11750 16649
rect 11692 16609 11704 16643
rect 11738 16640 11750 16643
rect 12158 16640 12164 16652
rect 11738 16612 12164 16640
rect 11738 16609 11750 16612
rect 11692 16603 11750 16609
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 13814 16640 13820 16652
rect 13775 16612 13820 16640
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 18708 16640 18736 16680
rect 18966 16668 18972 16680
rect 19024 16668 19030 16720
rect 25332 16708 25360 16739
rect 25866 16736 25872 16748
rect 25924 16776 25930 16788
rect 26973 16779 27031 16785
rect 26973 16776 26985 16779
rect 25924 16748 26985 16776
rect 25924 16736 25930 16748
rect 26973 16745 26985 16748
rect 27019 16745 27031 16779
rect 26973 16739 27031 16745
rect 25332 16680 26372 16708
rect 18874 16640 18880 16652
rect 17880 16612 18736 16640
rect 18835 16612 18880 16640
rect 9858 16572 9864 16584
rect 9600 16544 9864 16572
rect 9858 16532 9864 16544
rect 9916 16532 9922 16584
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 10367 16544 11284 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10336 16504 10364 16535
rect 8680 16476 10364 16504
rect 3513 16439 3571 16445
rect 3513 16405 3525 16439
rect 3559 16436 3571 16439
rect 3602 16436 3608 16448
rect 3559 16408 3608 16436
rect 3559 16405 3571 16408
rect 3513 16399 3571 16405
rect 3602 16396 3608 16408
rect 3660 16396 3666 16448
rect 4614 16436 4620 16448
rect 4575 16408 4620 16436
rect 4614 16396 4620 16408
rect 4672 16396 4678 16448
rect 6270 16396 6276 16448
rect 6328 16436 6334 16448
rect 11256 16445 11284 16544
rect 15102 16532 15108 16584
rect 15160 16572 15166 16584
rect 15289 16575 15347 16581
rect 15289 16572 15301 16575
rect 15160 16544 15301 16572
rect 15160 16532 15166 16544
rect 15289 16541 15301 16544
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 17770 16532 17776 16584
rect 17828 16572 17834 16584
rect 17880 16572 17908 16612
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 19518 16640 19524 16652
rect 19479 16612 19524 16640
rect 19518 16600 19524 16612
rect 19576 16600 19582 16652
rect 21174 16640 21180 16652
rect 21135 16612 21180 16640
rect 21174 16600 21180 16612
rect 21232 16600 21238 16652
rect 21266 16600 21272 16652
rect 21324 16640 21330 16652
rect 21433 16643 21491 16649
rect 21433 16640 21445 16643
rect 21324 16612 21445 16640
rect 21324 16600 21330 16612
rect 21433 16609 21445 16612
rect 21479 16640 21491 16643
rect 22370 16640 22376 16652
rect 21479 16612 22376 16640
rect 21479 16609 21491 16612
rect 21433 16603 21491 16609
rect 22370 16600 22376 16612
rect 22428 16600 22434 16652
rect 23106 16600 23112 16652
rect 23164 16640 23170 16652
rect 23842 16640 23848 16652
rect 23164 16612 23848 16640
rect 23164 16600 23170 16612
rect 23842 16600 23848 16612
rect 23900 16640 23906 16652
rect 24204 16643 24262 16649
rect 24204 16640 24216 16643
rect 23900 16612 24216 16640
rect 23900 16600 23906 16612
rect 24204 16609 24216 16612
rect 24250 16640 24262 16643
rect 24250 16612 24992 16640
rect 24250 16609 24262 16612
rect 24204 16603 24262 16609
rect 17828 16544 17908 16572
rect 17828 16532 17834 16544
rect 19058 16532 19064 16584
rect 19116 16572 19122 16584
rect 19116 16544 19161 16572
rect 19116 16532 19122 16544
rect 23198 16532 23204 16584
rect 23256 16572 23262 16584
rect 23750 16572 23756 16584
rect 23256 16544 23756 16572
rect 23256 16532 23262 16544
rect 23750 16532 23756 16544
rect 23808 16572 23814 16584
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 23808 16544 23949 16572
rect 23808 16532 23814 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 24964 16572 24992 16612
rect 25406 16572 25412 16584
rect 24964 16544 25412 16572
rect 23937 16535 23995 16541
rect 25406 16532 25412 16544
rect 25464 16532 25470 16584
rect 6549 16439 6607 16445
rect 6549 16436 6561 16439
rect 6328 16408 6561 16436
rect 6328 16396 6334 16408
rect 6549 16405 6561 16408
rect 6595 16405 6607 16439
rect 6549 16399 6607 16405
rect 11241 16439 11299 16445
rect 11241 16405 11253 16439
rect 11287 16436 11299 16439
rect 11422 16436 11428 16448
rect 11287 16408 11428 16436
rect 11287 16405 11299 16408
rect 11241 16399 11299 16405
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 18138 16436 18144 16448
rect 18099 16408 18144 16436
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 26344 16445 26372 16680
rect 26510 16600 26516 16652
rect 26568 16600 26574 16652
rect 26878 16640 26884 16652
rect 26839 16612 26884 16640
rect 26878 16600 26884 16612
rect 26936 16600 26942 16652
rect 26528 16513 26556 16600
rect 27154 16572 27160 16584
rect 27115 16544 27160 16572
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 26513 16507 26571 16513
rect 26513 16473 26525 16507
rect 26559 16473 26571 16507
rect 26513 16467 26571 16473
rect 26329 16439 26387 16445
rect 26329 16405 26341 16439
rect 26375 16436 26387 16439
rect 27154 16436 27160 16448
rect 26375 16408 27160 16436
rect 26375 16405 26387 16408
rect 26329 16399 26387 16405
rect 27154 16396 27160 16408
rect 27212 16396 27218 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 3050 16232 3056 16244
rect 3011 16204 3056 16232
rect 3050 16192 3056 16204
rect 3108 16232 3114 16244
rect 3973 16235 4031 16241
rect 3973 16232 3985 16235
rect 3108 16204 3985 16232
rect 3108 16192 3114 16204
rect 3973 16201 3985 16204
rect 4019 16201 4031 16235
rect 4154 16232 4160 16244
rect 4115 16204 4160 16232
rect 3973 16195 4031 16201
rect 3602 16164 3608 16176
rect 3563 16136 3608 16164
rect 3602 16124 3608 16136
rect 3660 16124 3666 16176
rect 3988 16096 4016 16195
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 5166 16232 5172 16244
rect 5127 16204 5172 16232
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 5534 16232 5540 16244
rect 5495 16204 5540 16232
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 8110 16232 8116 16244
rect 7432 16204 8116 16232
rect 7432 16192 7438 16204
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 10781 16235 10839 16241
rect 10781 16232 10793 16235
rect 9916 16204 10793 16232
rect 9916 16192 9922 16204
rect 10781 16201 10793 16204
rect 10827 16201 10839 16235
rect 12158 16232 12164 16244
rect 12119 16204 12164 16232
rect 10781 16195 10839 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 15010 16232 15016 16244
rect 14971 16204 15016 16232
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16232 17555 16235
rect 17586 16232 17592 16244
rect 17543 16204 17592 16232
rect 17543 16201 17555 16204
rect 17497 16195 17555 16201
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 19978 16232 19984 16244
rect 19939 16204 19984 16232
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 21174 16232 21180 16244
rect 21135 16204 21180 16232
rect 21174 16192 21180 16204
rect 21232 16192 21238 16244
rect 21358 16192 21364 16244
rect 21416 16232 21422 16244
rect 21453 16235 21511 16241
rect 21453 16232 21465 16235
rect 21416 16204 21465 16232
rect 21416 16192 21422 16204
rect 21453 16201 21465 16204
rect 21499 16201 21511 16235
rect 23106 16232 23112 16244
rect 23067 16204 23112 16232
rect 21453 16195 21511 16201
rect 23106 16192 23112 16204
rect 23164 16192 23170 16244
rect 23198 16192 23204 16244
rect 23256 16232 23262 16244
rect 23385 16235 23443 16241
rect 23385 16232 23397 16235
rect 23256 16204 23397 16232
rect 23256 16192 23262 16204
rect 23385 16201 23397 16204
rect 23431 16201 23443 16235
rect 24394 16232 24400 16244
rect 24355 16204 24400 16232
rect 23385 16195 23443 16201
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 24578 16232 24584 16244
rect 24539 16204 24584 16232
rect 24578 16192 24584 16204
rect 24636 16192 24642 16244
rect 25682 16192 25688 16244
rect 25740 16232 25746 16244
rect 25961 16235 26019 16241
rect 25961 16232 25973 16235
rect 25740 16204 25973 16232
rect 25740 16192 25746 16204
rect 25961 16201 25973 16204
rect 26007 16201 26019 16235
rect 25961 16195 26019 16201
rect 13449 16167 13507 16173
rect 13449 16133 13461 16167
rect 13495 16164 13507 16167
rect 13906 16164 13912 16176
rect 13495 16136 13912 16164
rect 13495 16133 13507 16136
rect 13449 16127 13507 16133
rect 13906 16124 13912 16136
rect 13964 16124 13970 16176
rect 15102 16124 15108 16176
rect 15160 16164 15166 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15160 16136 16037 16164
rect 15160 16124 15166 16136
rect 16025 16133 16037 16136
rect 16071 16164 16083 16167
rect 20901 16167 20959 16173
rect 16071 16136 18092 16164
rect 16071 16133 16083 16136
rect 16025 16127 16083 16133
rect 18064 16108 18092 16136
rect 20901 16133 20913 16167
rect 20947 16164 20959 16167
rect 21266 16164 21272 16176
rect 20947 16136 21272 16164
rect 20947 16133 20959 16136
rect 20901 16127 20959 16133
rect 21266 16124 21272 16136
rect 21324 16124 21330 16176
rect 4709 16099 4767 16105
rect 4709 16096 4721 16099
rect 3988 16068 4721 16096
rect 4709 16065 4721 16068
rect 4755 16065 4767 16099
rect 7282 16096 7288 16108
rect 7243 16068 7288 16096
rect 4709 16059 4767 16065
rect 7282 16056 7288 16068
rect 7340 16056 7346 16108
rect 11422 16096 11428 16108
rect 11383 16068 11428 16096
rect 11422 16056 11428 16068
rect 11480 16056 11486 16108
rect 12989 16099 13047 16105
rect 12989 16065 13001 16099
rect 13035 16096 13047 16099
rect 14093 16099 14151 16105
rect 14093 16096 14105 16099
rect 13035 16068 14105 16096
rect 13035 16065 13047 16068
rect 12989 16059 13047 16065
rect 14093 16065 14105 16068
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 14734 16096 14740 16108
rect 14599 16068 14740 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 1670 16028 1676 16040
rect 1631 16000 1676 16028
rect 1670 15988 1676 16000
rect 1728 15988 1734 16040
rect 8294 16028 8300 16040
rect 8255 16000 8300 16028
rect 8294 15988 8300 16000
rect 8352 15988 8358 16040
rect 11146 16028 11152 16040
rect 11107 16000 11152 16028
rect 11146 15988 11152 16000
rect 11204 15988 11210 16040
rect 13814 16028 13820 16040
rect 13775 16000 13820 16028
rect 13814 15988 13820 16000
rect 13872 15988 13878 16040
rect 14108 16028 14136 16059
rect 14734 16056 14740 16068
rect 14792 16096 14798 16108
rect 15657 16099 15715 16105
rect 15657 16096 15669 16099
rect 14792 16068 15669 16096
rect 14792 16056 14798 16068
rect 15657 16065 15669 16068
rect 15703 16096 15715 16099
rect 15838 16096 15844 16108
rect 15703 16068 15844 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 15838 16056 15844 16068
rect 15896 16056 15902 16108
rect 18046 16096 18052 16108
rect 17959 16068 18052 16096
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 22002 16096 22008 16108
rect 21963 16068 22008 16096
rect 22002 16056 22008 16068
rect 22060 16096 22066 16108
rect 22554 16096 22560 16108
rect 22060 16068 22560 16096
rect 22060 16056 22066 16068
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 24412 16096 24440 16192
rect 25041 16099 25099 16105
rect 25041 16096 25053 16099
rect 24412 16068 25053 16096
rect 25041 16065 25053 16068
rect 25087 16065 25099 16099
rect 25041 16059 25099 16065
rect 25225 16099 25283 16105
rect 25225 16065 25237 16099
rect 25271 16096 25283 16099
rect 25406 16096 25412 16108
rect 25271 16068 25412 16096
rect 25271 16065 25283 16068
rect 25225 16059 25283 16065
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 25976 16096 26004 16195
rect 27154 16192 27160 16244
rect 27212 16232 27218 16244
rect 28077 16235 28135 16241
rect 28077 16232 28089 16235
rect 27212 16204 28089 16232
rect 27212 16192 27218 16204
rect 28077 16201 28089 16204
rect 28123 16201 28135 16235
rect 28077 16195 28135 16201
rect 26145 16099 26203 16105
rect 26145 16096 26157 16099
rect 25976 16068 26157 16096
rect 26145 16065 26157 16068
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 15470 16028 15476 16040
rect 14108 16000 15476 16028
rect 15470 15988 15476 16000
rect 15528 15988 15534 16040
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18305 16031 18363 16037
rect 18305 16028 18317 16031
rect 18196 16000 18317 16028
rect 18196 15988 18202 16000
rect 18305 15997 18317 16000
rect 18351 15997 18363 16031
rect 18305 15991 18363 15997
rect 20533 16031 20591 16037
rect 20533 15997 20545 16031
rect 20579 16028 20591 16031
rect 21542 16028 21548 16040
rect 20579 16000 21548 16028
rect 20579 15997 20591 16000
rect 20533 15991 20591 15997
rect 21542 15988 21548 16000
rect 21600 16028 21606 16040
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 21600 16000 21833 16028
rect 21600 15988 21606 16000
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 23566 15988 23572 16040
rect 23624 16028 23630 16040
rect 24121 16031 24179 16037
rect 24121 16028 24133 16031
rect 23624 16000 24133 16028
rect 23624 15988 23630 16000
rect 24121 15997 24133 16000
rect 24167 16028 24179 16031
rect 24946 16028 24952 16040
rect 24167 16000 24952 16028
rect 24167 15997 24179 16000
rect 24121 15991 24179 15997
rect 24946 15988 24952 16000
rect 25004 15988 25010 16040
rect 1940 15963 1998 15969
rect 1940 15929 1952 15963
rect 1986 15960 1998 15963
rect 2682 15960 2688 15972
rect 1986 15932 2688 15960
rect 1986 15929 1998 15932
rect 1940 15923 1998 15929
rect 2682 15920 2688 15932
rect 2740 15920 2746 15972
rect 4522 15960 4528 15972
rect 4483 15932 4528 15960
rect 4522 15920 4528 15932
rect 4580 15960 4586 15972
rect 5905 15963 5963 15969
rect 5905 15960 5917 15963
rect 4580 15932 5917 15960
rect 4580 15920 4586 15932
rect 5905 15929 5917 15932
rect 5951 15929 5963 15963
rect 5905 15923 5963 15929
rect 8564 15963 8622 15969
rect 8564 15929 8576 15963
rect 8610 15960 8622 15963
rect 8662 15960 8668 15972
rect 8610 15932 8668 15960
rect 8610 15929 8622 15932
rect 8564 15923 8622 15929
rect 8662 15920 8668 15932
rect 8720 15960 8726 15972
rect 9490 15960 9496 15972
rect 8720 15932 9496 15960
rect 8720 15920 8726 15932
rect 9490 15920 9496 15932
rect 9548 15920 9554 15972
rect 26418 15969 26424 15972
rect 26412 15960 26424 15969
rect 26379 15932 26424 15960
rect 26412 15923 26424 15932
rect 26418 15920 26424 15923
rect 26476 15920 26482 15972
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 7193 15895 7251 15901
rect 7193 15861 7205 15895
rect 7239 15892 7251 15895
rect 8846 15892 8852 15904
rect 7239 15864 8852 15892
rect 7239 15861 7251 15864
rect 7193 15855 7251 15861
rect 8846 15852 8852 15864
rect 8904 15852 8910 15904
rect 10318 15892 10324 15904
rect 10279 15864 10324 15892
rect 10318 15852 10324 15864
rect 10376 15852 10382 15904
rect 10594 15892 10600 15904
rect 10555 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15892 10658 15904
rect 11241 15895 11299 15901
rect 11241 15892 11253 15895
rect 10652 15864 11253 15892
rect 10652 15852 10658 15864
rect 11241 15861 11253 15864
rect 11287 15892 11299 15895
rect 11514 15892 11520 15904
rect 11287 15864 11520 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11514 15852 11520 15864
rect 11572 15852 11578 15904
rect 11882 15892 11888 15904
rect 11843 15864 11888 15892
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 13354 15892 13360 15904
rect 13267 15864 13360 15892
rect 13354 15852 13360 15864
rect 13412 15892 13418 15904
rect 13909 15895 13967 15901
rect 13909 15892 13921 15895
rect 13412 15864 13921 15892
rect 13412 15852 13418 15864
rect 13909 15861 13921 15864
rect 13955 15861 13967 15895
rect 13909 15855 13967 15861
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15378 15892 15384 15904
rect 14967 15864 15384 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15473 15895 15531 15901
rect 15473 15861 15485 15895
rect 15519 15892 15531 15895
rect 15562 15892 15568 15904
rect 15519 15864 15568 15892
rect 15519 15861 15531 15864
rect 15473 15855 15531 15861
rect 15562 15852 15568 15864
rect 15620 15852 15626 15904
rect 17770 15892 17776 15904
rect 17731 15864 17776 15892
rect 17770 15852 17776 15864
rect 17828 15852 17834 15904
rect 18598 15852 18604 15904
rect 18656 15892 18662 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 18656 15864 19441 15892
rect 18656 15852 18662 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19429 15855 19487 15861
rect 21913 15895 21971 15901
rect 21913 15861 21925 15895
rect 21959 15892 21971 15895
rect 22186 15892 22192 15904
rect 21959 15864 22192 15892
rect 21959 15861 21971 15864
rect 21913 15855 21971 15861
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 25406 15852 25412 15904
rect 25464 15892 25470 15904
rect 25593 15895 25651 15901
rect 25593 15892 25605 15895
rect 25464 15864 25605 15892
rect 25464 15852 25470 15864
rect 25593 15861 25605 15864
rect 25639 15861 25651 15895
rect 25593 15855 25651 15861
rect 27246 15852 27252 15904
rect 27304 15892 27310 15904
rect 27525 15895 27583 15901
rect 27525 15892 27537 15895
rect 27304 15864 27537 15892
rect 27304 15852 27310 15864
rect 27525 15861 27537 15864
rect 27571 15861 27583 15895
rect 27525 15855 27583 15861
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 2038 15688 2044 15700
rect 1999 15660 2044 15688
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2409 15691 2467 15697
rect 2409 15657 2421 15691
rect 2455 15688 2467 15691
rect 3510 15688 3516 15700
rect 2455 15660 3516 15688
rect 2455 15657 2467 15660
rect 2409 15651 2467 15657
rect 3510 15648 3516 15660
rect 3568 15648 3574 15700
rect 3602 15648 3608 15700
rect 3660 15688 3666 15700
rect 3789 15691 3847 15697
rect 3789 15688 3801 15691
rect 3660 15660 3801 15688
rect 3660 15648 3666 15660
rect 3789 15657 3801 15660
rect 3835 15657 3847 15691
rect 3789 15651 3847 15657
rect 5810 15648 5816 15700
rect 5868 15688 5874 15700
rect 6733 15691 6791 15697
rect 6733 15688 6745 15691
rect 5868 15660 6745 15688
rect 5868 15648 5874 15660
rect 6733 15657 6745 15660
rect 6779 15657 6791 15691
rect 6733 15651 6791 15657
rect 8021 15691 8079 15697
rect 8021 15657 8033 15691
rect 8067 15688 8079 15691
rect 8202 15688 8208 15700
rect 8067 15660 8208 15688
rect 8067 15657 8079 15660
rect 8021 15651 8079 15657
rect 8202 15648 8208 15660
rect 8260 15648 8266 15700
rect 8386 15688 8392 15700
rect 8347 15660 8392 15688
rect 8386 15648 8392 15660
rect 8444 15648 8450 15700
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10321 15691 10379 15697
rect 10321 15688 10333 15691
rect 10008 15660 10333 15688
rect 10008 15648 10014 15660
rect 10321 15657 10333 15660
rect 10367 15657 10379 15691
rect 10321 15651 10379 15657
rect 10689 15691 10747 15697
rect 10689 15657 10701 15691
rect 10735 15688 10747 15691
rect 10870 15688 10876 15700
rect 10735 15660 10876 15688
rect 10735 15657 10747 15660
rect 10689 15651 10747 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 11422 15648 11428 15700
rect 11480 15688 11486 15700
rect 13265 15691 13323 15697
rect 13265 15688 13277 15691
rect 11480 15660 13277 15688
rect 11480 15648 11486 15660
rect 13265 15657 13277 15660
rect 13311 15657 13323 15691
rect 14734 15688 14740 15700
rect 14695 15660 14740 15688
rect 13265 15651 13323 15657
rect 14734 15648 14740 15660
rect 14792 15648 14798 15700
rect 15838 15648 15844 15700
rect 15896 15688 15902 15700
rect 16669 15691 16727 15697
rect 16669 15688 16681 15691
rect 15896 15660 16681 15688
rect 15896 15648 15902 15660
rect 16669 15657 16681 15660
rect 16715 15657 16727 15691
rect 18046 15688 18052 15700
rect 18007 15660 18052 15688
rect 16669 15651 16727 15657
rect 18046 15648 18052 15660
rect 18104 15648 18110 15700
rect 21177 15691 21235 15697
rect 21177 15657 21189 15691
rect 21223 15688 21235 15691
rect 21450 15688 21456 15700
rect 21223 15660 21456 15688
rect 21223 15657 21235 15660
rect 21177 15651 21235 15657
rect 21450 15648 21456 15660
rect 21508 15648 21514 15700
rect 22186 15688 22192 15700
rect 22147 15660 22192 15688
rect 22186 15648 22192 15660
rect 22244 15688 22250 15700
rect 22741 15691 22799 15697
rect 22741 15688 22753 15691
rect 22244 15660 22753 15688
rect 22244 15648 22250 15660
rect 22741 15657 22753 15660
rect 22787 15657 22799 15691
rect 23198 15688 23204 15700
rect 23159 15660 23204 15688
rect 22741 15651 22799 15657
rect 23198 15648 23204 15660
rect 23256 15688 23262 15700
rect 23474 15688 23480 15700
rect 23256 15660 23480 15688
rect 23256 15648 23262 15660
rect 23474 15648 23480 15660
rect 23532 15648 23538 15700
rect 23750 15648 23756 15700
rect 23808 15688 23814 15700
rect 24213 15691 24271 15697
rect 24213 15688 24225 15691
rect 23808 15660 24225 15688
rect 23808 15648 23814 15660
rect 24213 15657 24225 15660
rect 24259 15657 24271 15691
rect 24213 15651 24271 15657
rect 24857 15691 24915 15697
rect 24857 15657 24869 15691
rect 24903 15688 24915 15691
rect 26878 15688 26884 15700
rect 24903 15660 26884 15688
rect 24903 15657 24915 15660
rect 24857 15651 24915 15657
rect 26878 15648 26884 15660
rect 26936 15688 26942 15700
rect 27617 15691 27675 15697
rect 27617 15688 27629 15691
rect 26936 15660 27629 15688
rect 26936 15648 26942 15660
rect 27617 15657 27629 15660
rect 27663 15657 27675 15691
rect 27617 15651 27675 15657
rect 5258 15580 5264 15632
rect 5316 15620 5322 15632
rect 5598 15623 5656 15629
rect 5598 15620 5610 15623
rect 5316 15592 5610 15620
rect 5316 15580 5322 15592
rect 5598 15589 5610 15592
rect 5644 15589 5656 15623
rect 5598 15583 5656 15589
rect 9493 15623 9551 15629
rect 9493 15589 9505 15623
rect 9539 15620 9551 15623
rect 11440 15620 11468 15648
rect 9539 15592 11468 15620
rect 9539 15589 9551 15592
rect 9493 15583 9551 15589
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4706 15552 4712 15564
rect 4111 15524 4712 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4706 15512 4712 15524
rect 4764 15512 4770 15564
rect 5166 15512 5172 15564
rect 5224 15552 5230 15564
rect 5353 15555 5411 15561
rect 5353 15552 5365 15555
rect 5224 15524 5365 15552
rect 5224 15512 5230 15524
rect 5353 15521 5365 15524
rect 5399 15552 5411 15555
rect 5442 15552 5448 15564
rect 5399 15524 5448 15552
rect 5399 15521 5411 15524
rect 5353 15515 5411 15521
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 2498 15484 2504 15496
rect 2459 15456 2504 15484
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2682 15484 2688 15496
rect 2643 15456 2688 15484
rect 2682 15444 2688 15456
rect 2740 15444 2746 15496
rect 3145 15487 3203 15493
rect 3145 15453 3157 15487
rect 3191 15484 3203 15487
rect 5184 15484 5212 15512
rect 3191 15456 5212 15484
rect 8481 15487 8539 15493
rect 3191 15453 3203 15456
rect 3145 15447 3203 15453
rect 8481 15453 8493 15487
rect 8527 15484 8539 15487
rect 8570 15484 8576 15496
rect 8527 15456 8576 15484
rect 8527 15453 8539 15456
rect 8481 15447 8539 15453
rect 1670 15348 1676 15360
rect 1583 15320 1676 15348
rect 1670 15308 1676 15320
rect 1728 15348 1734 15360
rect 3050 15348 3056 15360
rect 1728 15320 3056 15348
rect 1728 15308 1734 15320
rect 3050 15308 3056 15320
rect 3108 15348 3114 15360
rect 3160 15348 3188 15447
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 9508 15484 9536 15583
rect 15470 15580 15476 15632
rect 15528 15629 15534 15632
rect 15528 15623 15592 15629
rect 15528 15589 15546 15623
rect 15580 15589 15592 15623
rect 15528 15583 15592 15589
rect 15528 15580 15534 15583
rect 12141 15555 12199 15561
rect 12141 15552 12153 15555
rect 10888 15524 12153 15552
rect 8711 15456 9536 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 7929 15419 7987 15425
rect 7929 15385 7941 15419
rect 7975 15416 7987 15419
rect 8386 15416 8392 15428
rect 7975 15388 8392 15416
rect 7975 15385 7987 15388
rect 7929 15379 7987 15385
rect 8386 15376 8392 15388
rect 8444 15416 8450 15428
rect 8680 15416 8708 15447
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10888 15493 10916 15524
rect 12141 15521 12153 15524
rect 12187 15552 12199 15555
rect 12526 15552 12532 15564
rect 12187 15524 12532 15552
rect 12187 15521 12199 15524
rect 12141 15515 12199 15521
rect 12526 15512 12532 15524
rect 12584 15512 12590 15564
rect 15102 15512 15108 15564
rect 15160 15552 15166 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 15160 15524 15301 15552
rect 15160 15512 15166 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 18064 15552 18092 15648
rect 20714 15620 20720 15632
rect 20627 15592 20720 15620
rect 20714 15580 20720 15592
rect 20772 15620 20778 15632
rect 21637 15623 21695 15629
rect 21637 15620 21649 15623
rect 20772 15592 21649 15620
rect 20772 15580 20778 15592
rect 21637 15589 21649 15592
rect 21683 15589 21695 15623
rect 24762 15620 24768 15632
rect 24675 15592 24768 15620
rect 21637 15583 21695 15589
rect 24762 15580 24768 15592
rect 24820 15620 24826 15632
rect 25225 15623 25283 15629
rect 25225 15620 25237 15623
rect 24820 15592 25237 15620
rect 24820 15580 24826 15592
rect 25225 15589 25237 15592
rect 25271 15620 25283 15623
rect 25866 15620 25872 15632
rect 25271 15592 25872 15620
rect 25271 15589 25283 15592
rect 25225 15583 25283 15589
rect 25866 15580 25872 15592
rect 25924 15580 25930 15632
rect 18325 15555 18383 15561
rect 18325 15552 18337 15555
rect 18064 15524 18337 15552
rect 15289 15515 15347 15521
rect 18325 15521 18337 15524
rect 18371 15552 18383 15555
rect 18414 15552 18420 15564
rect 18371 15524 18420 15552
rect 18371 15521 18383 15524
rect 18325 15515 18383 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 18598 15561 18604 15564
rect 18592 15552 18604 15561
rect 18559 15524 18604 15552
rect 18592 15515 18604 15524
rect 18598 15512 18604 15515
rect 18656 15512 18662 15564
rect 21542 15552 21548 15564
rect 21503 15524 21548 15552
rect 21542 15512 21548 15524
rect 21600 15512 21606 15564
rect 23106 15552 23112 15564
rect 23067 15524 23112 15552
rect 23106 15512 23112 15524
rect 23164 15512 23170 15564
rect 25317 15555 25375 15561
rect 25317 15521 25329 15555
rect 25363 15552 25375 15555
rect 26602 15552 26608 15564
rect 25363 15524 26608 15552
rect 25363 15521 25375 15524
rect 25317 15515 25375 15521
rect 10781 15487 10839 15493
rect 10781 15484 10793 15487
rect 10468 15456 10793 15484
rect 10468 15444 10474 15456
rect 10781 15453 10793 15456
rect 10827 15453 10839 15487
rect 10781 15447 10839 15453
rect 10873 15487 10931 15493
rect 10873 15453 10885 15487
rect 10919 15453 10931 15487
rect 11882 15484 11888 15496
rect 11843 15456 11888 15484
rect 10873 15447 10931 15453
rect 8444 15388 8708 15416
rect 10229 15419 10287 15425
rect 8444 15376 8450 15388
rect 10229 15385 10241 15419
rect 10275 15416 10287 15419
rect 10888 15416 10916 15447
rect 11882 15444 11888 15456
rect 11940 15444 11946 15496
rect 21726 15484 21732 15496
rect 21687 15456 21732 15484
rect 21726 15444 21732 15456
rect 21784 15484 21790 15496
rect 22002 15484 22008 15496
rect 21784 15456 22008 15484
rect 21784 15444 21790 15456
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15453 23351 15487
rect 23293 15447 23351 15453
rect 10275 15388 10916 15416
rect 10275 15385 10287 15388
rect 10229 15379 10287 15385
rect 22370 15376 22376 15428
rect 22428 15416 22434 15428
rect 23308 15416 23336 15447
rect 24578 15444 24584 15496
rect 24636 15484 24642 15496
rect 25332 15484 25360 15515
rect 26602 15512 26608 15524
rect 26660 15512 26666 15564
rect 26878 15552 26884 15564
rect 26839 15524 26884 15552
rect 26878 15512 26884 15524
rect 26936 15512 26942 15564
rect 24636 15456 25360 15484
rect 24636 15444 24642 15456
rect 25406 15444 25412 15496
rect 25464 15484 25470 15496
rect 26970 15484 26976 15496
rect 25464 15456 25509 15484
rect 26931 15456 26976 15484
rect 25464 15444 25470 15456
rect 26970 15444 26976 15456
rect 27028 15444 27034 15496
rect 27157 15487 27215 15493
rect 27157 15453 27169 15487
rect 27203 15484 27215 15487
rect 27522 15484 27528 15496
rect 27203 15456 27528 15484
rect 27203 15453 27215 15456
rect 27157 15447 27215 15453
rect 22428 15388 23336 15416
rect 23937 15419 23995 15425
rect 22428 15376 22434 15388
rect 23937 15385 23949 15419
rect 23983 15416 23995 15419
rect 24486 15416 24492 15428
rect 23983 15388 24492 15416
rect 23983 15385 23995 15388
rect 23937 15379 23995 15385
rect 24486 15376 24492 15388
rect 24544 15376 24550 15428
rect 26237 15419 26295 15425
rect 26237 15385 26249 15419
rect 26283 15416 26295 15419
rect 26418 15416 26424 15428
rect 26283 15388 26424 15416
rect 26283 15385 26295 15388
rect 26237 15379 26295 15385
rect 26418 15376 26424 15388
rect 26476 15416 26482 15428
rect 27172 15416 27200 15447
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 26476 15388 27200 15416
rect 26476 15376 26482 15388
rect 3108 15320 3188 15348
rect 4249 15351 4307 15357
rect 3108 15308 3114 15320
rect 4249 15317 4261 15351
rect 4295 15348 4307 15351
rect 4338 15348 4344 15360
rect 4295 15320 4344 15348
rect 4295 15317 4307 15320
rect 4249 15311 4307 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 4614 15348 4620 15360
rect 4575 15320 4620 15348
rect 4614 15308 4620 15320
rect 4672 15308 4678 15360
rect 5258 15348 5264 15360
rect 5219 15320 5264 15348
rect 5258 15308 5264 15320
rect 5316 15308 5322 15360
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9030 15348 9036 15360
rect 8352 15320 9036 15348
rect 8352 15308 8358 15320
rect 9030 15308 9036 15320
rect 9088 15308 9094 15360
rect 11422 15348 11428 15360
rect 11383 15320 11428 15348
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 11793 15351 11851 15357
rect 11793 15317 11805 15351
rect 11839 15348 11851 15351
rect 12250 15348 12256 15360
rect 11839 15320 12256 15348
rect 11839 15317 11851 15320
rect 11793 15311 11851 15317
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 13814 15348 13820 15360
rect 13775 15320 13820 15348
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14366 15308 14372 15360
rect 14424 15348 14430 15360
rect 15105 15351 15163 15357
rect 15105 15348 15117 15351
rect 14424 15320 15117 15348
rect 14424 15308 14430 15320
rect 15105 15317 15117 15320
rect 15151 15348 15163 15351
rect 15562 15348 15568 15360
rect 15151 15320 15568 15348
rect 15151 15317 15163 15320
rect 15105 15311 15163 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 19702 15348 19708 15360
rect 19663 15320 19708 15348
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 26513 15351 26571 15357
rect 26513 15317 26525 15351
rect 26559 15348 26571 15351
rect 27154 15348 27160 15360
rect 26559 15320 27160 15348
rect 26559 15317 26571 15320
rect 26513 15311 26571 15317
rect 27154 15308 27160 15320
rect 27212 15308 27218 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 2038 15144 2044 15156
rect 1999 15116 2044 15144
rect 2038 15104 2044 15116
rect 2096 15104 2102 15156
rect 2406 15104 2412 15156
rect 2464 15144 2470 15156
rect 3605 15147 3663 15153
rect 3605 15144 3617 15147
rect 2464 15116 3617 15144
rect 2464 15104 2470 15116
rect 3605 15113 3617 15116
rect 3651 15113 3663 15147
rect 7926 15144 7932 15156
rect 7887 15116 7932 15144
rect 3605 15107 3663 15113
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 12621 15147 12679 15153
rect 12621 15144 12633 15147
rect 12584 15116 12633 15144
rect 12584 15104 12590 15116
rect 12621 15113 12633 15116
rect 12667 15113 12679 15147
rect 12621 15107 12679 15113
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 13722 15144 13728 15156
rect 13127 15116 13728 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 18414 15104 18420 15156
rect 18472 15144 18478 15156
rect 19521 15147 19579 15153
rect 18472 15116 18517 15144
rect 18472 15104 18478 15116
rect 19521 15113 19533 15147
rect 19567 15144 19579 15147
rect 20622 15144 20628 15156
rect 19567 15116 20628 15144
rect 19567 15113 19579 15116
rect 19521 15107 19579 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21266 15144 21272 15156
rect 21039 15116 21272 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 14645 15079 14703 15085
rect 14645 15076 14657 15079
rect 13872 15048 14657 15076
rect 13872 15036 13878 15048
rect 14645 15045 14657 15048
rect 14691 15045 14703 15079
rect 14645 15039 14703 15045
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 16022 15076 16028 15088
rect 14792 15048 15240 15076
rect 15983 15048 16028 15076
rect 14792 15036 14798 15048
rect 15212 15020 15240 15048
rect 16022 15036 16028 15048
rect 16080 15036 16086 15088
rect 18432 15076 18460 15104
rect 21008 15076 21036 15107
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 22370 15104 22376 15156
rect 22428 15144 22434 15156
rect 22465 15147 22523 15153
rect 22465 15144 22477 15147
rect 22428 15116 22477 15144
rect 22428 15104 22434 15116
rect 22465 15113 22477 15116
rect 22511 15113 22523 15147
rect 23474 15144 23480 15156
rect 23435 15116 23480 15144
rect 22465 15107 22523 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 24121 15147 24179 15153
rect 24121 15113 24133 15147
rect 24167 15144 24179 15147
rect 24578 15144 24584 15156
rect 24167 15116 24584 15144
rect 24167 15113 24179 15116
rect 24121 15107 24179 15113
rect 24578 15104 24584 15116
rect 24636 15104 24642 15156
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 28077 15147 28135 15153
rect 28077 15144 28089 15147
rect 27672 15116 28089 15144
rect 27672 15104 27678 15116
rect 28077 15113 28089 15116
rect 28123 15113 28135 15147
rect 28077 15107 28135 15113
rect 18432 15048 21036 15076
rect 2682 15008 2688 15020
rect 2595 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 15008 2746 15020
rect 3602 15008 3608 15020
rect 2740 14980 3608 15008
rect 2740 14968 2746 14980
rect 3602 14968 3608 14980
rect 3660 15008 3666 15020
rect 4157 15011 4215 15017
rect 4157 15008 4169 15011
rect 3660 14980 4169 15008
rect 3660 14968 3666 14980
rect 4157 14977 4169 14980
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 5258 14968 5264 15020
rect 5316 15008 5322 15020
rect 5813 15011 5871 15017
rect 5813 15008 5825 15011
rect 5316 14980 5825 15008
rect 5316 14968 5322 14980
rect 5813 14977 5825 14980
rect 5859 15008 5871 15011
rect 6270 15008 6276 15020
rect 5859 14980 6276 15008
rect 5859 14977 5871 14980
rect 5813 14971 5871 14977
rect 6270 14968 6276 14980
rect 6328 15008 6334 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 6328 14980 6561 15008
rect 6328 14968 6334 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 10410 15008 10416 15020
rect 10371 14980 10416 15008
rect 6549 14971 6607 14977
rect 10410 14968 10416 14980
rect 10468 14968 10474 15020
rect 11330 15008 11336 15020
rect 11291 14980 11336 15008
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 13722 15008 13728 15020
rect 13683 14980 13728 15008
rect 13722 14968 13728 14980
rect 13780 14968 13786 15020
rect 13906 14968 13912 15020
rect 13964 15008 13970 15020
rect 15105 15011 15163 15017
rect 15105 15008 15117 15011
rect 13964 14980 15117 15008
rect 13964 14968 13970 14980
rect 15105 14977 15117 14980
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 15194 14968 15200 15020
rect 15252 15008 15258 15020
rect 15252 14980 15345 15008
rect 15252 14968 15258 14980
rect 15470 14968 15476 15020
rect 15528 15008 15534 15020
rect 16761 15011 16819 15017
rect 16761 15008 16773 15011
rect 15528 14980 16773 15008
rect 15528 14968 15534 14980
rect 16761 14977 16773 14980
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 19429 15011 19487 15017
rect 19429 14977 19441 15011
rect 19475 15008 19487 15011
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19475 14980 20085 15008
rect 19475 14977 19487 14980
rect 19429 14971 19487 14977
rect 20073 14977 20085 14980
rect 20119 15008 20131 15011
rect 20622 15008 20628 15020
rect 20119 14980 20628 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 21008 15008 21036 15048
rect 26878 15036 26884 15088
rect 26936 15076 26942 15088
rect 27706 15076 27712 15088
rect 26936 15048 27712 15076
rect 26936 15036 26942 15048
rect 27706 15036 27712 15048
rect 27764 15036 27770 15088
rect 21092 15011 21150 15017
rect 21092 15008 21104 15011
rect 21008 14980 21104 15008
rect 21092 14977 21104 14980
rect 21138 14977 21150 15011
rect 21092 14971 21150 14977
rect 23750 14968 23756 15020
rect 23808 15008 23814 15020
rect 24213 15011 24271 15017
rect 24213 15008 24225 15011
rect 23808 14980 24225 15008
rect 23808 14968 23814 14980
rect 24213 14977 24225 14980
rect 24259 14977 24271 15011
rect 27246 15008 27252 15020
rect 27207 14980 27252 15008
rect 24213 14971 24271 14977
rect 27246 14968 27252 14980
rect 27304 14968 27310 15020
rect 2498 14900 2504 14952
rect 2556 14940 2562 14952
rect 3053 14943 3111 14949
rect 3053 14940 3065 14943
rect 2556 14912 3065 14940
rect 2556 14900 2562 14912
rect 3053 14909 3065 14912
rect 3099 14909 3111 14943
rect 3053 14903 3111 14909
rect 4065 14943 4123 14949
rect 4065 14909 4077 14943
rect 4111 14940 4123 14943
rect 4614 14940 4620 14952
rect 4111 14912 4620 14940
rect 4111 14909 4123 14912
rect 4065 14903 4123 14909
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14940 5135 14943
rect 5626 14940 5632 14952
rect 5123 14912 5632 14940
rect 5123 14909 5135 14912
rect 5077 14903 5135 14909
rect 3510 14872 3516 14884
rect 3423 14844 3516 14872
rect 3510 14832 3516 14844
rect 3568 14872 3574 14884
rect 3973 14875 4031 14881
rect 3973 14872 3985 14875
rect 3568 14844 3985 14872
rect 3568 14832 3574 14844
rect 3973 14841 3985 14844
rect 4019 14872 4031 14875
rect 5092 14872 5120 14903
rect 5626 14900 5632 14912
rect 5684 14900 5690 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 7883 14912 8125 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 8113 14909 8125 14912
rect 8159 14940 8171 14943
rect 8202 14940 8208 14952
rect 8159 14912 8208 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8386 14949 8392 14952
rect 8380 14940 8392 14949
rect 8347 14912 8392 14940
rect 8380 14903 8392 14912
rect 8386 14900 8392 14903
rect 8444 14900 8450 14952
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 12250 14940 12256 14952
rect 11195 14912 12256 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13814 14940 13820 14952
rect 13495 14912 13820 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 16022 14900 16028 14952
rect 16080 14940 16086 14952
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16080 14912 16681 14940
rect 16080 14900 16086 14912
rect 16669 14909 16681 14912
rect 16715 14940 16727 14943
rect 16942 14940 16948 14952
rect 16715 14912 16948 14940
rect 16715 14909 16727 14912
rect 16669 14903 16727 14909
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 26237 14943 26295 14949
rect 26237 14909 26249 14943
rect 26283 14940 26295 14943
rect 26786 14940 26792 14952
rect 26283 14912 26792 14940
rect 26283 14909 26295 14912
rect 26237 14903 26295 14909
rect 26786 14900 26792 14912
rect 26844 14900 26850 14952
rect 27154 14940 27160 14952
rect 27115 14912 27160 14940
rect 27154 14900 27160 14912
rect 27212 14940 27218 14952
rect 28445 14943 28503 14949
rect 28445 14940 28457 14943
rect 27212 14912 28457 14940
rect 27212 14900 27218 14912
rect 28445 14909 28457 14912
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 4019 14844 5120 14872
rect 4019 14841 4031 14844
rect 3973 14835 4031 14841
rect 5258 14832 5264 14884
rect 5316 14872 5322 14884
rect 5537 14875 5595 14881
rect 5537 14872 5549 14875
rect 5316 14844 5549 14872
rect 5316 14832 5322 14844
rect 5537 14841 5549 14844
rect 5583 14872 5595 14875
rect 7653 14875 7711 14881
rect 7653 14872 7665 14875
rect 5583 14844 7665 14872
rect 5583 14841 5595 14844
rect 5537 14835 5595 14841
rect 7653 14841 7665 14844
rect 7699 14872 7711 14875
rect 8478 14872 8484 14884
rect 7699 14844 8484 14872
rect 7699 14841 7711 14844
rect 7653 14835 7711 14841
rect 8478 14832 8484 14844
rect 8536 14832 8542 14884
rect 11514 14832 11520 14884
rect 11572 14872 11578 14884
rect 11882 14872 11888 14884
rect 11572 14844 11888 14872
rect 11572 14832 11578 14844
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 13722 14832 13728 14884
rect 13780 14872 13786 14884
rect 14093 14875 14151 14881
rect 14093 14872 14105 14875
rect 13780 14844 14105 14872
rect 13780 14832 13786 14844
rect 14093 14841 14105 14844
rect 14139 14872 14151 14875
rect 14550 14872 14556 14884
rect 14139 14844 14556 14872
rect 14139 14841 14151 14844
rect 14093 14835 14151 14841
rect 14550 14832 14556 14844
rect 14608 14832 14614 14884
rect 16574 14872 16580 14884
rect 15672 14844 16580 14872
rect 15672 14816 15700 14844
rect 16574 14832 16580 14844
rect 16632 14832 16638 14884
rect 18138 14832 18144 14884
rect 18196 14872 18202 14884
rect 18598 14872 18604 14884
rect 18196 14844 18604 14872
rect 18196 14832 18202 14844
rect 18598 14832 18604 14844
rect 18656 14872 18662 14884
rect 24486 14881 24492 14884
rect 18693 14875 18751 14881
rect 18693 14872 18705 14875
rect 18656 14844 18705 14872
rect 18656 14832 18662 14844
rect 18693 14841 18705 14844
rect 18739 14841 18751 14875
rect 21330 14875 21388 14881
rect 21330 14872 21342 14875
rect 18693 14835 18751 14841
rect 20548 14844 21342 14872
rect 1949 14807 2007 14813
rect 1949 14773 1961 14807
rect 1995 14804 2007 14807
rect 2406 14804 2412 14816
rect 1995 14776 2412 14804
rect 1995 14773 2007 14776
rect 1949 14767 2007 14773
rect 2406 14764 2412 14776
rect 2464 14764 2470 14816
rect 2501 14807 2559 14813
rect 2501 14773 2513 14807
rect 2547 14804 2559 14807
rect 2958 14804 2964 14816
rect 2547 14776 2964 14804
rect 2547 14773 2559 14776
rect 2501 14767 2559 14773
rect 2958 14764 2964 14776
rect 3016 14764 3022 14816
rect 4706 14804 4712 14816
rect 4667 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 5166 14804 5172 14816
rect 5127 14776 5172 14804
rect 5166 14764 5172 14776
rect 5224 14764 5230 14816
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 6181 14807 6239 14813
rect 6181 14804 6193 14807
rect 5684 14776 6193 14804
rect 5684 14764 5690 14776
rect 6181 14773 6193 14776
rect 6227 14804 6239 14807
rect 6730 14804 6736 14816
rect 6227 14776 6736 14804
rect 6227 14773 6239 14776
rect 6181 14767 6239 14773
rect 6730 14764 6736 14776
rect 6788 14804 6794 14816
rect 7193 14807 7251 14813
rect 7193 14804 7205 14807
rect 6788 14776 7205 14804
rect 6788 14764 6794 14776
rect 7193 14773 7205 14776
rect 7239 14804 7251 14807
rect 7837 14807 7895 14813
rect 7837 14804 7849 14807
rect 7239 14776 7849 14804
rect 7239 14773 7251 14776
rect 7193 14767 7251 14773
rect 7837 14773 7849 14776
rect 7883 14773 7895 14807
rect 10778 14804 10784 14816
rect 10739 14776 10784 14804
rect 7837 14767 7895 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11241 14807 11299 14813
rect 11241 14773 11253 14807
rect 11287 14804 11299 14807
rect 11422 14804 11428 14816
rect 11287 14776 11428 14804
rect 11287 14773 11299 14776
rect 11241 14767 11299 14773
rect 11422 14764 11428 14776
rect 11480 14804 11486 14816
rect 11790 14804 11796 14816
rect 11480 14776 11796 14804
rect 11480 14764 11486 14776
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 13538 14804 13544 14816
rect 13499 14776 13544 14804
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 14458 14804 14464 14816
rect 14419 14776 14464 14804
rect 14458 14764 14464 14776
rect 14516 14804 14522 14816
rect 15010 14804 15016 14816
rect 14516 14776 15016 14804
rect 14516 14764 14522 14776
rect 15010 14764 15016 14776
rect 15068 14764 15074 14816
rect 15654 14804 15660 14816
rect 15615 14776 15660 14804
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 16206 14804 16212 14816
rect 16167 14776 16212 14804
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 19886 14804 19892 14816
rect 19847 14776 19892 14804
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 19981 14807 20039 14813
rect 19981 14773 19993 14807
rect 20027 14804 20039 14807
rect 20070 14804 20076 14816
rect 20027 14776 20076 14804
rect 20027 14773 20039 14776
rect 19981 14767 20039 14773
rect 20070 14764 20076 14776
rect 20128 14764 20134 14816
rect 20438 14764 20444 14816
rect 20496 14804 20502 14816
rect 20548 14813 20576 14844
rect 21330 14841 21342 14844
rect 21376 14841 21388 14875
rect 24480 14872 24492 14881
rect 24447 14844 24492 14872
rect 21330 14835 21388 14841
rect 24480 14835 24492 14844
rect 24486 14832 24492 14835
rect 24544 14832 24550 14884
rect 26605 14875 26663 14881
rect 26605 14841 26617 14875
rect 26651 14872 26663 14875
rect 26970 14872 26976 14884
rect 26651 14844 26976 14872
rect 26651 14841 26663 14844
rect 26605 14835 26663 14841
rect 26970 14832 26976 14844
rect 27028 14832 27034 14884
rect 20533 14807 20591 14813
rect 20533 14804 20545 14807
rect 20496 14776 20545 14804
rect 20496 14764 20502 14776
rect 20533 14773 20545 14776
rect 20579 14773 20591 14807
rect 23106 14804 23112 14816
rect 23067 14776 23112 14804
rect 20533 14767 20591 14773
rect 23106 14764 23112 14776
rect 23164 14764 23170 14816
rect 25590 14804 25596 14816
rect 25551 14776 25596 14804
rect 25590 14764 25596 14776
rect 25648 14764 25654 14816
rect 26694 14804 26700 14816
rect 26655 14776 26700 14804
rect 26694 14764 26700 14776
rect 26752 14764 26758 14816
rect 26786 14764 26792 14816
rect 26844 14804 26850 14816
rect 27065 14807 27123 14813
rect 27065 14804 27077 14807
rect 26844 14776 27077 14804
rect 26844 14764 26850 14776
rect 27065 14773 27077 14776
rect 27111 14773 27123 14807
rect 27065 14767 27123 14773
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 1854 14600 1860 14612
rect 1815 14572 1860 14600
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 3050 14560 3056 14612
rect 3108 14600 3114 14612
rect 3237 14603 3295 14609
rect 3237 14600 3249 14603
rect 3108 14572 3249 14600
rect 3108 14560 3114 14572
rect 3237 14569 3249 14572
rect 3283 14569 3295 14603
rect 3602 14600 3608 14612
rect 3563 14572 3608 14600
rect 3237 14563 3295 14569
rect 3602 14560 3608 14572
rect 3660 14560 3666 14612
rect 5258 14600 5264 14612
rect 5219 14572 5264 14600
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 7561 14603 7619 14609
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7607 14572 7941 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7929 14569 7941 14572
rect 7975 14600 7987 14603
rect 8386 14600 8392 14612
rect 7975 14572 8392 14600
rect 7975 14569 7987 14572
rect 7929 14563 7987 14569
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 8481 14603 8539 14609
rect 8481 14569 8493 14603
rect 8527 14600 8539 14603
rect 8938 14600 8944 14612
rect 8527 14572 8944 14600
rect 8527 14569 8539 14572
rect 8481 14563 8539 14569
rect 8938 14560 8944 14572
rect 8996 14560 9002 14612
rect 9125 14603 9183 14609
rect 9125 14569 9137 14603
rect 9171 14600 9183 14603
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9171 14572 10149 14600
rect 9171 14569 9183 14572
rect 9125 14563 9183 14569
rect 10137 14569 10149 14572
rect 10183 14600 10195 14603
rect 10778 14600 10784 14612
rect 10183 14572 10784 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12584 14572 12725 14600
rect 12584 14560 12590 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 13538 14560 13544 14612
rect 13596 14600 13602 14612
rect 13725 14603 13783 14609
rect 13725 14600 13737 14603
rect 13596 14572 13737 14600
rect 13596 14560 13602 14572
rect 13725 14569 13737 14572
rect 13771 14600 13783 14603
rect 15289 14603 15347 14609
rect 15289 14600 15301 14603
rect 13771 14572 15301 14600
rect 13771 14569 13783 14572
rect 13725 14563 13783 14569
rect 15289 14569 15301 14572
rect 15335 14569 15347 14603
rect 15289 14563 15347 14569
rect 15749 14603 15807 14609
rect 15749 14569 15761 14603
rect 15795 14600 15807 14603
rect 16206 14600 16212 14612
rect 15795 14572 16212 14600
rect 15795 14569 15807 14572
rect 15749 14563 15807 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 20349 14603 20407 14609
rect 20349 14569 20361 14603
rect 20395 14600 20407 14603
rect 21269 14603 21327 14609
rect 21269 14600 21281 14603
rect 20395 14572 21281 14600
rect 20395 14569 20407 14572
rect 20349 14563 20407 14569
rect 21269 14569 21281 14572
rect 21315 14600 21327 14603
rect 21542 14600 21548 14612
rect 21315 14572 21548 14600
rect 21315 14569 21327 14572
rect 21269 14563 21327 14569
rect 21542 14560 21548 14572
rect 21600 14560 21606 14612
rect 26326 14560 26332 14612
rect 26384 14600 26390 14612
rect 26513 14603 26571 14609
rect 26513 14600 26525 14603
rect 26384 14572 26525 14600
rect 26384 14560 26390 14572
rect 26513 14569 26525 14572
rect 26559 14569 26571 14603
rect 26513 14563 26571 14569
rect 11146 14492 11152 14544
rect 11204 14532 11210 14544
rect 11578 14535 11636 14541
rect 11578 14532 11590 14535
rect 11204 14504 11590 14532
rect 11204 14492 11210 14504
rect 11578 14501 11590 14504
rect 11624 14501 11636 14535
rect 11578 14495 11636 14501
rect 13906 14492 13912 14544
rect 13964 14532 13970 14544
rect 14277 14535 14335 14541
rect 14277 14532 14289 14535
rect 13964 14504 14289 14532
rect 13964 14492 13970 14504
rect 14277 14501 14289 14504
rect 14323 14501 14335 14535
rect 14277 14495 14335 14501
rect 14458 14492 14464 14544
rect 14516 14532 14522 14544
rect 14737 14535 14795 14541
rect 14737 14532 14749 14535
rect 14516 14504 14749 14532
rect 14516 14492 14522 14504
rect 14737 14501 14749 14504
rect 14783 14532 14795 14535
rect 15470 14532 15476 14544
rect 14783 14504 15476 14532
rect 14783 14501 14795 14504
rect 14737 14495 14795 14501
rect 15470 14492 15476 14504
rect 15528 14492 15534 14544
rect 15657 14535 15715 14541
rect 15657 14501 15669 14535
rect 15703 14532 15715 14535
rect 15838 14532 15844 14544
rect 15703 14504 15844 14532
rect 15703 14501 15715 14504
rect 15657 14495 15715 14501
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 17402 14541 17408 14544
rect 17396 14532 17408 14541
rect 17363 14504 17408 14532
rect 17396 14495 17408 14504
rect 17402 14492 17408 14495
rect 17460 14492 17466 14544
rect 20717 14535 20775 14541
rect 20717 14501 20729 14535
rect 20763 14532 20775 14535
rect 21726 14532 21732 14544
rect 20763 14504 21732 14532
rect 20763 14501 20775 14504
rect 20717 14495 20775 14501
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 24204 14535 24262 14541
rect 24204 14501 24216 14535
rect 24250 14532 24262 14535
rect 24578 14532 24584 14544
rect 24250 14504 24584 14532
rect 24250 14501 24262 14504
rect 24204 14495 24262 14501
rect 24578 14492 24584 14504
rect 24636 14532 24642 14544
rect 25590 14532 25596 14544
rect 24636 14504 25596 14532
rect 24636 14492 24642 14504
rect 25590 14492 25596 14504
rect 25648 14492 25654 14544
rect 750 14424 756 14476
rect 808 14464 814 14476
rect 2038 14464 2044 14476
rect 808 14436 2044 14464
rect 808 14424 814 14436
rect 2038 14424 2044 14436
rect 2096 14464 2102 14476
rect 2225 14467 2283 14473
rect 2225 14464 2237 14467
rect 2096 14436 2237 14464
rect 2096 14424 2102 14436
rect 2225 14433 2237 14436
rect 2271 14433 2283 14467
rect 4062 14464 4068 14476
rect 4023 14436 4068 14464
rect 2225 14427 2283 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 5442 14424 5448 14476
rect 5500 14464 5506 14476
rect 5537 14467 5595 14473
rect 5537 14464 5549 14467
rect 5500 14436 5549 14464
rect 5500 14424 5506 14436
rect 5537 14433 5549 14436
rect 5583 14464 5595 14467
rect 5626 14464 5632 14476
rect 5583 14436 5632 14464
rect 5583 14433 5595 14436
rect 5537 14427 5595 14433
rect 5626 14424 5632 14436
rect 5684 14424 5690 14476
rect 5810 14473 5816 14476
rect 5804 14464 5816 14473
rect 5771 14436 5816 14464
rect 5804 14427 5816 14436
rect 5810 14424 5816 14427
rect 5868 14424 5874 14476
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 8389 14467 8447 14473
rect 8389 14464 8401 14467
rect 8352 14436 8401 14464
rect 8352 14424 8358 14436
rect 8389 14433 8401 14436
rect 8435 14433 8447 14467
rect 10870 14464 10876 14476
rect 10831 14436 10876 14464
rect 8389 14427 8447 14433
rect 10870 14424 10876 14436
rect 10928 14424 10934 14476
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14464 11391 14467
rect 11422 14464 11428 14476
rect 11379 14436 11428 14464
rect 11379 14433 11391 14436
rect 11333 14427 11391 14433
rect 11422 14424 11428 14436
rect 11480 14424 11486 14476
rect 15102 14464 15108 14476
rect 15063 14436 15108 14464
rect 15102 14424 15108 14436
rect 15160 14424 15166 14476
rect 15488 14464 15516 14492
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15488 14436 16313 14464
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 20898 14424 20904 14476
rect 20956 14464 20962 14476
rect 21637 14467 21695 14473
rect 21637 14464 21649 14467
rect 20956 14436 21649 14464
rect 20956 14424 20962 14436
rect 21637 14433 21649 14436
rect 21683 14433 21695 14467
rect 22281 14467 22339 14473
rect 22281 14464 22293 14467
rect 21637 14427 21695 14433
rect 21744 14436 22293 14464
rect 21744 14408 21772 14436
rect 22281 14433 22293 14436
rect 22327 14433 22339 14467
rect 22281 14427 22339 14433
rect 23750 14424 23756 14476
rect 23808 14464 23814 14476
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 23808 14436 23949 14464
rect 23808 14424 23814 14436
rect 23937 14433 23949 14436
rect 23983 14433 23995 14467
rect 26878 14464 26884 14476
rect 26839 14436 26884 14464
rect 23937 14427 23995 14433
rect 26878 14424 26884 14436
rect 26936 14424 26942 14476
rect 2317 14399 2375 14405
rect 2317 14396 2329 14399
rect 1780 14368 2329 14396
rect 1486 14220 1492 14272
rect 1544 14260 1550 14272
rect 1780 14269 1808 14368
rect 2317 14365 2329 14368
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 2682 14396 2688 14408
rect 2547 14368 2688 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 2332 14328 2360 14359
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 2958 14396 2964 14408
rect 2871 14368 2964 14396
rect 2958 14356 2964 14368
rect 3016 14396 3022 14408
rect 4706 14396 4712 14408
rect 3016 14368 4712 14396
rect 3016 14356 3022 14368
rect 4706 14356 4712 14368
rect 4764 14356 4770 14408
rect 8662 14396 8668 14408
rect 8623 14368 8668 14396
rect 8662 14356 8668 14368
rect 8720 14356 8726 14408
rect 9674 14356 9680 14408
rect 9732 14396 9738 14408
rect 10226 14396 10232 14408
rect 9732 14368 10088 14396
rect 10187 14368 10232 14396
rect 9732 14356 9738 14368
rect 5258 14328 5264 14340
rect 2332 14300 5264 14328
rect 5258 14288 5264 14300
rect 5316 14288 5322 14340
rect 9766 14328 9772 14340
rect 9727 14300 9772 14328
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 10060 14328 10088 14368
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10413 14399 10471 14405
rect 10413 14365 10425 14399
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10428 14328 10456 14359
rect 13722 14356 13728 14408
rect 13780 14396 13786 14408
rect 13817 14399 13875 14405
rect 13817 14396 13829 14399
rect 13780 14368 13829 14396
rect 13780 14356 13786 14368
rect 13817 14365 13829 14368
rect 13863 14365 13875 14399
rect 13817 14359 13875 14365
rect 15194 14356 15200 14408
rect 15252 14396 15258 14408
rect 15746 14396 15752 14408
rect 15252 14368 15752 14396
rect 15252 14356 15258 14368
rect 15746 14356 15752 14368
rect 15804 14396 15810 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15804 14368 15853 14396
rect 15804 14356 15810 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 17126 14396 17132 14408
rect 17087 14368 17132 14396
rect 15841 14359 15899 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 21726 14396 21732 14408
rect 21687 14368 21732 14396
rect 21726 14356 21732 14368
rect 21784 14356 21790 14408
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22370 14396 22376 14408
rect 21867 14368 22376 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 11146 14328 11152 14340
rect 10060 14300 11152 14328
rect 11146 14288 11152 14300
rect 11204 14288 11210 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19886 14328 19892 14340
rect 19392 14300 19892 14328
rect 19392 14288 19398 14300
rect 19886 14288 19892 14300
rect 19944 14288 19950 14340
rect 20622 14288 20628 14340
rect 20680 14328 20686 14340
rect 21836 14328 21864 14359
rect 22370 14356 22376 14368
rect 22428 14396 22434 14408
rect 22741 14399 22799 14405
rect 22741 14396 22753 14399
rect 22428 14368 22753 14396
rect 22428 14356 22434 14368
rect 22741 14365 22753 14368
rect 22787 14365 22799 14399
rect 22922 14396 22928 14408
rect 22883 14368 22928 14396
rect 22741 14359 22799 14365
rect 22922 14356 22928 14368
rect 22980 14356 22986 14408
rect 26694 14356 26700 14408
rect 26752 14396 26758 14408
rect 26973 14399 27031 14405
rect 26973 14396 26985 14399
rect 26752 14368 26985 14396
rect 26752 14356 26758 14368
rect 26973 14365 26985 14368
rect 27019 14365 27031 14399
rect 26973 14359 27031 14365
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14365 27215 14399
rect 27157 14359 27215 14365
rect 20680 14300 21864 14328
rect 20680 14288 20686 14300
rect 27172 14272 27200 14359
rect 1765 14263 1823 14269
rect 1765 14260 1777 14263
rect 1544 14232 1777 14260
rect 1544 14220 1550 14232
rect 1765 14229 1777 14232
rect 1811 14229 1823 14263
rect 1765 14223 1823 14229
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 3050 14260 3056 14272
rect 2372 14232 3056 14260
rect 2372 14220 2378 14232
rect 3050 14220 3056 14232
rect 3108 14220 3114 14272
rect 4154 14220 4160 14272
rect 4212 14260 4218 14272
rect 4249 14263 4307 14269
rect 4249 14260 4261 14263
rect 4212 14232 4261 14260
rect 4212 14220 4218 14232
rect 4249 14229 4261 14232
rect 4295 14229 4307 14263
rect 4798 14260 4804 14272
rect 4759 14232 4804 14260
rect 4249 14223 4307 14229
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 6914 14260 6920 14272
rect 6875 14232 6920 14260
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 8018 14260 8024 14272
rect 7979 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 9493 14263 9551 14269
rect 9493 14229 9505 14263
rect 9539 14260 9551 14263
rect 9950 14260 9956 14272
rect 9539 14232 9956 14260
rect 9539 14229 9551 14232
rect 9493 14223 9551 14229
rect 9950 14220 9956 14232
rect 10008 14220 10014 14272
rect 11241 14263 11299 14269
rect 11241 14229 11253 14263
rect 11287 14260 11299 14263
rect 11330 14260 11336 14272
rect 11287 14232 11336 14260
rect 11287 14229 11299 14232
rect 11241 14223 11299 14229
rect 11330 14220 11336 14232
rect 11388 14220 11394 14272
rect 13262 14260 13268 14272
rect 13223 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18509 14263 18567 14269
rect 18509 14260 18521 14263
rect 18104 14232 18521 14260
rect 18104 14220 18110 14232
rect 18509 14229 18521 14232
rect 18555 14229 18567 14263
rect 19150 14260 19156 14272
rect 19111 14232 19156 14260
rect 18509 14223 18567 14229
rect 19150 14220 19156 14232
rect 19208 14220 19214 14272
rect 19613 14263 19671 14269
rect 19613 14229 19625 14263
rect 19659 14260 19671 14263
rect 20070 14260 20076 14272
rect 19659 14232 20076 14260
rect 19659 14229 19671 14232
rect 19613 14223 19671 14229
rect 20070 14220 20076 14232
rect 20128 14260 20134 14272
rect 20530 14260 20536 14272
rect 20128 14232 20536 14260
rect 20128 14220 20134 14232
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 21174 14260 21180 14272
rect 21135 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 23474 14260 23480 14272
rect 23435 14232 23480 14260
rect 23474 14220 23480 14232
rect 23532 14220 23538 14272
rect 23842 14260 23848 14272
rect 23803 14232 23848 14260
rect 23842 14220 23848 14232
rect 23900 14220 23906 14272
rect 25317 14263 25375 14269
rect 25317 14229 25329 14263
rect 25363 14260 25375 14263
rect 25682 14260 25688 14272
rect 25363 14232 25688 14260
rect 25363 14229 25375 14232
rect 25317 14223 25375 14229
rect 25682 14220 25688 14232
rect 25740 14260 25746 14272
rect 27154 14260 27160 14272
rect 25740 14232 27160 14260
rect 25740 14220 25746 14232
rect 27154 14220 27160 14232
rect 27212 14220 27218 14272
rect 27246 14220 27252 14272
rect 27304 14260 27310 14272
rect 27525 14263 27583 14269
rect 27525 14260 27537 14263
rect 27304 14232 27537 14260
rect 27304 14220 27310 14232
rect 27525 14229 27537 14232
rect 27571 14229 27583 14263
rect 27525 14223 27583 14229
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 3602 14056 3608 14068
rect 3563 14028 3608 14056
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 4062 14016 4068 14068
rect 4120 14056 4126 14068
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 4120 14028 4169 14056
rect 4120 14016 4126 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4157 14019 4215 14025
rect 4614 14016 4620 14068
rect 4672 14056 4678 14068
rect 4709 14059 4767 14065
rect 4709 14056 4721 14059
rect 4672 14028 4721 14056
rect 4672 14016 4678 14028
rect 4709 14025 4721 14028
rect 4755 14025 4767 14059
rect 4709 14019 4767 14025
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5684 14028 5733 14056
rect 5684 14016 5690 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 5721 14019 5779 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8294 14056 8300 14068
rect 8159 14028 8300 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8938 14056 8944 14068
rect 8899 14028 8944 14056
rect 8938 14016 8944 14028
rect 8996 14016 9002 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11204 14028 11253 14056
rect 11204 14016 11210 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 11241 14019 11299 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14458 14056 14464 14068
rect 14419 14028 14464 14056
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 14734 14056 14740 14068
rect 14695 14028 14740 14056
rect 14734 14016 14740 14028
rect 14792 14016 14798 14068
rect 15746 14016 15752 14068
rect 15804 14056 15810 14068
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15804 14028 15945 14056
rect 15804 14016 15810 14028
rect 15933 14025 15945 14028
rect 15979 14025 15991 14059
rect 16298 14056 16304 14068
rect 16259 14028 16304 14056
rect 15933 14019 15991 14025
rect 16298 14016 16304 14028
rect 16356 14016 16362 14068
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 17402 14056 17408 14068
rect 16632 14028 17408 14056
rect 16632 14016 16638 14028
rect 17402 14016 17408 14028
rect 17460 14056 17466 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 17460 14028 17509 14056
rect 17460 14016 17466 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 20456 14028 23152 14056
rect 4798 13880 4804 13932
rect 4856 13920 4862 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 4856 13892 5273 13920
rect 4856 13880 4862 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 6328 13892 7389 13920
rect 6328 13880 6334 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 11330 13880 11336 13932
rect 11388 13880 11394 13932
rect 14752 13920 14780 14016
rect 14921 13991 14979 13997
rect 14921 13957 14933 13991
rect 14967 13988 14979 13991
rect 15838 13988 15844 14000
rect 14967 13960 15844 13988
rect 14967 13957 14979 13960
rect 14921 13951 14979 13957
rect 15838 13948 15844 13960
rect 15896 13948 15902 14000
rect 19518 13988 19524 14000
rect 19479 13960 19524 13988
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 15378 13920 15384 13932
rect 14752 13892 15384 13920
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 19429 13923 19487 13929
rect 15528 13892 15573 13920
rect 15528 13880 15534 13892
rect 19429 13889 19441 13923
rect 19475 13920 19487 13923
rect 20165 13923 20223 13929
rect 20165 13920 20177 13923
rect 19475 13892 20177 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 20165 13889 20177 13892
rect 20211 13920 20223 13923
rect 20456 13920 20484 14028
rect 20622 13988 20628 14000
rect 20583 13960 20628 13988
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 20898 13988 20904 14000
rect 20859 13960 20904 13988
rect 20898 13948 20904 13960
rect 20956 13948 20962 14000
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 23124 13997 23152 14028
rect 23750 14016 23756 14068
rect 23808 14056 23814 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23808 14028 23857 14056
rect 23808 14016 23814 14028
rect 23845 14025 23857 14028
rect 23891 14025 23903 14059
rect 24026 14056 24032 14068
rect 23987 14028 24032 14056
rect 23845 14019 23903 14025
rect 24026 14016 24032 14028
rect 24084 14016 24090 14068
rect 25133 14059 25191 14065
rect 25133 14025 25145 14059
rect 25179 14056 25191 14059
rect 25406 14056 25412 14068
rect 25179 14028 25412 14056
rect 25179 14025 25191 14028
rect 25133 14019 25191 14025
rect 25406 14016 25412 14028
rect 25464 14016 25470 14068
rect 27154 14016 27160 14068
rect 27212 14056 27218 14068
rect 27525 14059 27583 14065
rect 27525 14056 27537 14059
rect 27212 14028 27537 14056
rect 27212 14016 27218 14028
rect 27525 14025 27537 14028
rect 27571 14025 27583 14059
rect 27525 14019 27583 14025
rect 22465 13991 22523 13997
rect 22465 13988 22477 13991
rect 22152 13960 22477 13988
rect 22152 13948 22158 13960
rect 22465 13957 22477 13960
rect 22511 13957 22523 13991
rect 22465 13951 22523 13957
rect 23109 13991 23167 13997
rect 23109 13957 23121 13991
rect 23155 13988 23167 13991
rect 23477 13991 23535 13997
rect 23477 13988 23489 13991
rect 23155 13960 23489 13988
rect 23155 13957 23167 13960
rect 23109 13951 23167 13957
rect 23477 13957 23489 13960
rect 23523 13988 23535 13991
rect 23523 13960 24624 13988
rect 23523 13957 23535 13960
rect 23477 13951 23535 13957
rect 24596 13932 24624 13960
rect 26878 13948 26884 14000
rect 26936 13988 26942 14000
rect 28261 13991 28319 13997
rect 28261 13988 28273 13991
rect 26936 13960 28273 13988
rect 26936 13948 26942 13960
rect 28261 13957 28273 13960
rect 28307 13957 28319 13991
rect 28261 13951 28319 13957
rect 20211 13892 20484 13920
rect 21008 13892 21200 13920
rect 20211 13889 20223 13892
rect 20165 13883 20223 13889
rect 2225 13855 2283 13861
rect 2225 13821 2237 13855
rect 2271 13852 2283 13855
rect 2314 13852 2320 13864
rect 2271 13824 2320 13852
rect 2271 13821 2283 13824
rect 2225 13815 2283 13821
rect 2314 13812 2320 13824
rect 2372 13812 2378 13864
rect 4614 13852 4620 13864
rect 4527 13824 4620 13852
rect 4614 13812 4620 13824
rect 4672 13852 4678 13864
rect 5169 13855 5227 13861
rect 5169 13852 5181 13855
rect 4672 13824 5181 13852
rect 4672 13812 4678 13824
rect 5169 13821 5181 13824
rect 5215 13852 5227 13855
rect 5215 13824 5764 13852
rect 5215 13821 5227 13824
rect 5169 13815 5227 13821
rect 2498 13793 2504 13796
rect 2492 13784 2504 13793
rect 2459 13756 2504 13784
rect 2492 13747 2504 13756
rect 2498 13744 2504 13747
rect 2556 13744 2562 13796
rect 5077 13787 5135 13793
rect 5077 13753 5089 13787
rect 5123 13784 5135 13787
rect 5626 13784 5632 13796
rect 5123 13756 5632 13784
rect 5123 13753 5135 13756
rect 5077 13747 5135 13753
rect 5626 13744 5632 13756
rect 5684 13744 5690 13796
rect 5736 13784 5764 13824
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6822 13852 6828 13864
rect 6604 13824 6828 13852
rect 6604 13812 6610 13824
rect 6822 13812 6828 13824
rect 6880 13852 6886 13864
rect 7285 13855 7343 13861
rect 7285 13852 7297 13855
rect 6880 13824 7297 13852
rect 6880 13812 6886 13824
rect 7285 13821 7297 13824
rect 7331 13821 7343 13855
rect 7285 13815 7343 13821
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9217 13855 9275 13861
rect 9217 13852 9229 13855
rect 8720 13824 9229 13852
rect 8720 13812 8726 13824
rect 9217 13821 9229 13824
rect 9263 13821 9275 13855
rect 9861 13855 9919 13861
rect 9861 13852 9873 13855
rect 9217 13815 9275 13821
rect 9600 13824 9873 13852
rect 5902 13784 5908 13796
rect 5736 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13744 5966 13796
rect 9030 13744 9036 13796
rect 9088 13784 9094 13796
rect 9600 13784 9628 13824
rect 9088 13756 9628 13784
rect 9692 13784 9720 13824
rect 9861 13821 9873 13824
rect 9907 13821 9919 13855
rect 9861 13815 9919 13821
rect 9950 13812 9956 13864
rect 10008 13852 10014 13864
rect 10128 13855 10186 13861
rect 10128 13852 10140 13855
rect 10008 13824 10140 13852
rect 10008 13812 10014 13824
rect 10128 13821 10140 13824
rect 10174 13852 10186 13855
rect 10594 13852 10600 13864
rect 10174 13824 10600 13852
rect 10174 13821 10186 13824
rect 10128 13815 10186 13821
rect 10594 13812 10600 13824
rect 10652 13852 10658 13864
rect 11348 13852 11376 13880
rect 10652 13824 11376 13852
rect 12437 13855 12495 13861
rect 10652 13812 10658 13824
rect 12437 13821 12449 13855
rect 12483 13821 12495 13855
rect 12437 13815 12495 13821
rect 19061 13855 19119 13861
rect 19061 13821 19073 13855
rect 19107 13852 19119 13855
rect 19978 13852 19984 13864
rect 19107 13824 19984 13852
rect 19107 13821 19119 13824
rect 19061 13815 19119 13821
rect 11422 13784 11428 13796
rect 9692 13756 11428 13784
rect 9088 13744 9094 13756
rect 9692 13728 9720 13756
rect 11422 13744 11428 13756
rect 11480 13784 11486 13796
rect 11793 13787 11851 13793
rect 11793 13784 11805 13787
rect 11480 13756 11805 13784
rect 11480 13744 11486 13756
rect 11793 13753 11805 13756
rect 11839 13784 11851 13787
rect 12161 13787 12219 13793
rect 12161 13784 12173 13787
rect 11839 13756 12173 13784
rect 11839 13753 11851 13756
rect 11793 13747 11851 13753
rect 12161 13753 12173 13756
rect 12207 13784 12219 13787
rect 12452 13784 12480 13815
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 20070 13812 20076 13864
rect 20128 13852 20134 13864
rect 21008 13852 21036 13892
rect 21172 13864 21200 13892
rect 23842 13880 23848 13932
rect 23900 13920 23906 13932
rect 24489 13923 24547 13929
rect 24489 13920 24501 13923
rect 23900 13892 24501 13920
rect 23900 13880 23906 13892
rect 24489 13889 24501 13892
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 20128 13824 21036 13852
rect 21085 13855 21143 13861
rect 20128 13812 20134 13824
rect 21085 13821 21097 13855
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 12207 13756 12480 13784
rect 12704 13787 12762 13793
rect 12207 13753 12219 13756
rect 12161 13747 12219 13753
rect 12704 13753 12716 13787
rect 12750 13784 12762 13787
rect 13262 13784 13268 13796
rect 12750 13756 13268 13784
rect 12750 13753 12762 13756
rect 12704 13747 12762 13753
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 1949 13719 2007 13725
rect 1949 13685 1961 13719
rect 1995 13716 2007 13719
rect 2038 13716 2044 13728
rect 1995 13688 2044 13716
rect 1995 13685 2007 13688
rect 1949 13679 2007 13685
rect 2038 13676 2044 13688
rect 2096 13676 2102 13728
rect 6178 13716 6184 13728
rect 6139 13688 6184 13716
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6825 13719 6883 13725
rect 6825 13685 6837 13719
rect 6871 13716 6883 13719
rect 7006 13716 7012 13728
rect 6871 13688 7012 13716
rect 6871 13685 6883 13688
rect 6825 13679 6883 13685
rect 7006 13676 7012 13688
rect 7064 13676 7070 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7193 13719 7251 13725
rect 7193 13716 7205 13719
rect 7156 13688 7205 13716
rect 7156 13676 7162 13688
rect 7193 13685 7205 13688
rect 7239 13685 7251 13719
rect 8386 13716 8392 13728
rect 8347 13688 8392 13716
rect 7193 13679 7251 13685
rect 8386 13676 8392 13688
rect 8444 13676 8450 13728
rect 9674 13676 9680 13728
rect 9732 13716 9738 13728
rect 9732 13688 9777 13716
rect 9732 13676 9738 13688
rect 15102 13676 15108 13728
rect 15160 13716 15166 13728
rect 15289 13719 15347 13725
rect 15289 13716 15301 13719
rect 15160 13688 15301 13716
rect 15160 13676 15166 13688
rect 15289 13685 15301 13688
rect 15335 13685 15347 13719
rect 17126 13716 17132 13728
rect 17087 13688 17132 13716
rect 15289 13679 15347 13685
rect 17126 13676 17132 13688
rect 17184 13676 17190 13728
rect 18230 13716 18236 13728
rect 18191 13688 18236 13716
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 19886 13716 19892 13728
rect 19208 13688 19892 13716
rect 19208 13676 19214 13688
rect 19886 13676 19892 13688
rect 19944 13676 19950 13728
rect 21100 13716 21128 13815
rect 21172 13812 21180 13864
rect 21232 13852 21238 13864
rect 21232 13824 21305 13852
rect 21232 13812 21238 13824
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 24394 13852 24400 13864
rect 23532 13824 24400 13852
rect 23532 13812 23538 13824
rect 24394 13812 24400 13824
rect 24452 13812 24458 13864
rect 24504 13852 24532 13883
rect 24578 13880 24584 13932
rect 24636 13920 24642 13932
rect 25590 13920 25596 13932
rect 24636 13892 24681 13920
rect 25424 13892 25596 13920
rect 24636 13880 24642 13892
rect 24762 13852 24768 13864
rect 24504 13824 24768 13852
rect 24762 13812 24768 13824
rect 24820 13812 24826 13864
rect 21172 13784 21200 13812
rect 21352 13787 21410 13793
rect 21352 13784 21364 13787
rect 21172 13756 21364 13784
rect 21352 13753 21364 13756
rect 21398 13753 21410 13787
rect 21352 13747 21410 13753
rect 23750 13744 23756 13796
rect 23808 13784 23814 13796
rect 25424 13793 25452 13892
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 26694 13880 26700 13932
rect 26752 13920 26758 13932
rect 27893 13923 27951 13929
rect 27893 13920 27905 13923
rect 26752 13892 27905 13920
rect 26752 13880 26758 13892
rect 27893 13889 27905 13892
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 25682 13812 25688 13864
rect 25740 13852 25746 13864
rect 25849 13855 25907 13861
rect 25849 13852 25861 13855
rect 25740 13824 25861 13852
rect 25740 13812 25746 13824
rect 25849 13821 25861 13824
rect 25895 13821 25907 13855
rect 25849 13815 25907 13821
rect 25409 13787 25467 13793
rect 25409 13784 25421 13787
rect 23808 13756 25421 13784
rect 23808 13744 23814 13756
rect 25409 13753 25421 13756
rect 25455 13753 25467 13787
rect 25409 13747 25467 13753
rect 21266 13716 21272 13728
rect 21100 13688 21272 13716
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 26973 13719 27031 13725
rect 26973 13685 26985 13719
rect 27019 13716 27031 13719
rect 27062 13716 27068 13728
rect 27019 13688 27068 13716
rect 27019 13685 27031 13688
rect 26973 13679 27031 13685
rect 27062 13676 27068 13688
rect 27120 13676 27126 13728
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 4801 13515 4859 13521
rect 4801 13481 4813 13515
rect 4847 13512 4859 13515
rect 4982 13512 4988 13524
rect 4847 13484 4988 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 4982 13472 4988 13484
rect 5040 13512 5046 13524
rect 5626 13512 5632 13524
rect 5040 13484 5632 13512
rect 5040 13472 5046 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 5902 13512 5908 13524
rect 5767 13484 5908 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 5902 13472 5908 13484
rect 5960 13512 5966 13524
rect 6638 13512 6644 13524
rect 5960 13484 6644 13512
rect 5960 13472 5966 13484
rect 6638 13472 6644 13484
rect 6696 13472 6702 13524
rect 9125 13515 9183 13521
rect 9125 13481 9137 13515
rect 9171 13512 9183 13515
rect 9953 13515 10011 13521
rect 9953 13512 9965 13515
rect 9171 13484 9965 13512
rect 9171 13481 9183 13484
rect 9125 13475 9183 13481
rect 9953 13481 9965 13484
rect 9999 13512 10011 13515
rect 10226 13512 10232 13524
rect 9999 13484 10232 13512
rect 9999 13481 10011 13484
rect 9953 13475 10011 13481
rect 10226 13472 10232 13484
rect 10284 13472 10290 13524
rect 11330 13512 11336 13524
rect 11291 13484 11336 13512
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11790 13512 11796 13524
rect 11751 13484 11796 13512
rect 11790 13472 11796 13484
rect 11848 13472 11854 13524
rect 12250 13512 12256 13524
rect 12211 13484 12256 13512
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12860 13484 12909 13512
rect 12860 13472 12866 13484
rect 12897 13481 12909 13484
rect 12943 13512 12955 13515
rect 13722 13512 13728 13524
rect 12943 13484 13728 13512
rect 12943 13481 12955 13484
rect 12897 13475 12955 13481
rect 13722 13472 13728 13484
rect 13780 13472 13786 13524
rect 15838 13512 15844 13524
rect 15799 13484 15844 13512
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 19242 13512 19248 13524
rect 19203 13484 19248 13512
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 21453 13515 21511 13521
rect 21453 13481 21465 13515
rect 21499 13512 21511 13515
rect 21726 13512 21732 13524
rect 21499 13484 21732 13512
rect 21499 13481 21511 13484
rect 21453 13475 21511 13481
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 24210 13512 24216 13524
rect 24171 13484 24216 13512
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 25869 13515 25927 13521
rect 25869 13512 25881 13515
rect 25740 13484 25881 13512
rect 25740 13472 25746 13484
rect 25869 13481 25881 13484
rect 25915 13481 25927 13515
rect 25869 13475 25927 13481
rect 3602 13404 3608 13456
rect 3660 13444 3666 13456
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 3660 13416 3801 13444
rect 3660 13404 3666 13416
rect 3789 13413 3801 13416
rect 3835 13413 3847 13447
rect 3789 13407 3847 13413
rect 5169 13447 5227 13453
rect 5169 13413 5181 13447
rect 5215 13444 5227 13447
rect 5810 13444 5816 13456
rect 5215 13416 5816 13444
rect 5215 13413 5227 13416
rect 5169 13407 5227 13413
rect 5810 13404 5816 13416
rect 5868 13444 5874 13456
rect 5868 13416 6408 13444
rect 5868 13404 5874 13416
rect 6380 13388 6408 13416
rect 6914 13404 6920 13456
rect 6972 13444 6978 13456
rect 7190 13444 7196 13456
rect 6972 13416 7196 13444
rect 6972 13404 6978 13416
rect 7190 13404 7196 13416
rect 7248 13444 7254 13456
rect 7346 13447 7404 13453
rect 7346 13444 7358 13447
rect 7248 13416 7358 13444
rect 7248 13404 7254 13416
rect 7346 13413 7358 13416
rect 7392 13413 7404 13447
rect 7346 13407 7404 13413
rect 9493 13447 9551 13453
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 9582 13444 9588 13456
rect 9539 13416 9588 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 13262 13444 13268 13456
rect 13223 13416 13268 13444
rect 13262 13404 13268 13416
rect 13320 13404 13326 13456
rect 13538 13404 13544 13456
rect 13596 13444 13602 13456
rect 14001 13447 14059 13453
rect 14001 13444 14013 13447
rect 13596 13416 14013 13444
rect 13596 13404 13602 13416
rect 14001 13413 14013 13416
rect 14047 13413 14059 13447
rect 17126 13444 17132 13456
rect 14001 13407 14059 13413
rect 16592 13416 17132 13444
rect 1489 13379 1547 13385
rect 1489 13345 1501 13379
rect 1535 13376 1547 13379
rect 1578 13376 1584 13388
rect 1535 13348 1584 13376
rect 1535 13345 1547 13348
rect 1489 13339 1547 13345
rect 1578 13336 1584 13348
rect 1636 13336 1642 13388
rect 1762 13385 1768 13388
rect 1756 13376 1768 13385
rect 1675 13348 1768 13376
rect 1756 13339 1768 13348
rect 1820 13376 1826 13388
rect 3050 13376 3056 13388
rect 1820 13348 3056 13376
rect 1762 13336 1768 13339
rect 1820 13336 1826 13348
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 4065 13379 4123 13385
rect 4065 13345 4077 13379
rect 4111 13376 4123 13379
rect 4246 13376 4252 13388
rect 4111 13348 4252 13376
rect 4111 13345 4123 13348
rect 4065 13339 4123 13345
rect 4246 13336 4252 13348
rect 4304 13336 4310 13388
rect 6362 13376 6368 13388
rect 6275 13348 6368 13376
rect 6362 13336 6368 13348
rect 6420 13376 6426 13388
rect 7650 13376 7656 13388
rect 6420 13348 7656 13376
rect 6420 13336 6426 13348
rect 7650 13336 7656 13348
rect 7708 13336 7714 13388
rect 10321 13379 10379 13385
rect 10321 13345 10333 13379
rect 10367 13376 10379 13379
rect 11054 13376 11060 13388
rect 10367 13348 11060 13376
rect 10367 13345 10379 13348
rect 10321 13339 10379 13345
rect 11054 13336 11060 13348
rect 11112 13336 11118 13388
rect 12158 13376 12164 13388
rect 12119 13348 12164 13376
rect 12158 13336 12164 13348
rect 12216 13336 12222 13388
rect 14090 13376 14096 13388
rect 14051 13348 14096 13376
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 16592 13385 16620 13416
rect 17126 13404 17132 13416
rect 17184 13404 17190 13456
rect 21652 13416 25360 13444
rect 16850 13385 16856 13388
rect 16577 13379 16635 13385
rect 16577 13345 16589 13379
rect 16623 13345 16635 13379
rect 16844 13376 16856 13385
rect 16763 13348 16856 13376
rect 16577 13339 16635 13345
rect 16844 13339 16856 13348
rect 16908 13376 16914 13388
rect 17862 13376 17868 13388
rect 16908 13348 17868 13376
rect 16850 13336 16856 13339
rect 16908 13336 16914 13348
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 18966 13336 18972 13388
rect 19024 13376 19030 13388
rect 19613 13379 19671 13385
rect 19613 13376 19625 13379
rect 19024 13348 19625 13376
rect 19024 13336 19030 13348
rect 19613 13345 19625 13348
rect 19659 13345 19671 13379
rect 20438 13376 20444 13388
rect 19613 13339 19671 13345
rect 19812 13348 20444 13376
rect 19812 13320 19840 13348
rect 20438 13336 20444 13348
rect 20496 13376 20502 13388
rect 20717 13379 20775 13385
rect 20717 13376 20729 13379
rect 20496 13348 20729 13376
rect 20496 13336 20502 13348
rect 20717 13345 20729 13348
rect 20763 13345 20775 13379
rect 20717 13339 20775 13345
rect 2498 13268 2504 13320
rect 2556 13308 2562 13320
rect 3513 13311 3571 13317
rect 3513 13308 3525 13311
rect 2556 13280 3525 13308
rect 2556 13268 2562 13280
rect 2884 13249 2912 13280
rect 3513 13277 3525 13280
rect 3559 13308 3571 13311
rect 4798 13308 4804 13320
rect 3559 13280 4804 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 5442 13268 5448 13320
rect 5500 13308 5506 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5500 13280 5825 13308
rect 5500 13268 5506 13280
rect 5813 13277 5825 13280
rect 5859 13308 5871 13311
rect 6178 13308 6184 13320
rect 5859 13280 6184 13308
rect 5859 13277 5871 13280
rect 5813 13271 5871 13277
rect 6178 13268 6184 13280
rect 6236 13268 6242 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 7101 13311 7159 13317
rect 7101 13308 7113 13311
rect 6788 13280 7113 13308
rect 6788 13268 6794 13280
rect 7101 13277 7113 13280
rect 7147 13277 7159 13311
rect 10410 13308 10416 13320
rect 10371 13280 10416 13308
rect 7101 13271 7159 13277
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 10594 13308 10600 13320
rect 10555 13280 10600 13308
rect 10594 13268 10600 13280
rect 10652 13268 10658 13320
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 14277 13311 14335 13317
rect 12391 13280 12425 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14458 13308 14464 13320
rect 14323 13280 14464 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 2869 13243 2927 13249
rect 2869 13209 2881 13243
rect 2915 13209 2927 13243
rect 2869 13203 2927 13209
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 12360 13240 12388 13271
rect 14458 13268 14464 13280
rect 14516 13268 14522 13320
rect 19702 13308 19708 13320
rect 19663 13280 19708 13308
rect 19702 13268 19708 13280
rect 19760 13268 19766 13320
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20349 13311 20407 13317
rect 19852 13280 19897 13308
rect 19852 13268 19858 13280
rect 20349 13277 20361 13311
rect 20395 13308 20407 13311
rect 20622 13308 20628 13320
rect 20395 13280 20628 13308
rect 20395 13277 20407 13280
rect 20349 13271 20407 13277
rect 20622 13268 20628 13280
rect 20680 13268 20686 13320
rect 13262 13240 13268 13252
rect 11940 13212 13268 13240
rect 11940 13200 11946 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13633 13243 13691 13249
rect 13633 13209 13645 13243
rect 13679 13240 13691 13243
rect 15286 13240 15292 13252
rect 13679 13212 15292 13240
rect 13679 13209 13691 13212
rect 13633 13203 13691 13209
rect 15286 13200 15292 13212
rect 15344 13240 15350 13252
rect 15473 13243 15531 13249
rect 15473 13240 15485 13243
rect 15344 13212 15485 13240
rect 15344 13200 15350 13212
rect 15473 13209 15485 13212
rect 15519 13209 15531 13243
rect 20732 13240 20760 13339
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21652 13308 21680 13416
rect 25332 13388 25360 13416
rect 21818 13376 21824 13388
rect 21779 13348 21824 13376
rect 21818 13336 21824 13348
rect 21876 13376 21882 13388
rect 23014 13376 23020 13388
rect 21876 13348 23020 13376
rect 21876 13336 21882 13348
rect 23014 13336 23020 13348
rect 23072 13336 23078 13388
rect 24118 13376 24124 13388
rect 24079 13348 24124 13376
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 25314 13376 25320 13388
rect 25227 13348 25320 13376
rect 25314 13336 25320 13348
rect 25372 13336 25378 13388
rect 25498 13336 25504 13388
rect 25556 13376 25562 13388
rect 26881 13379 26939 13385
rect 26881 13376 26893 13379
rect 25556 13348 26893 13376
rect 25556 13336 25562 13348
rect 26881 13345 26893 13348
rect 26927 13376 26939 13379
rect 28166 13376 28172 13388
rect 26927 13348 28172 13376
rect 26927 13345 26939 13348
rect 26881 13339 26939 13345
rect 28166 13336 28172 13348
rect 28224 13336 28230 13388
rect 21913 13311 21971 13317
rect 21913 13308 21925 13311
rect 21048 13280 21925 13308
rect 21048 13268 21054 13280
rect 21913 13277 21925 13280
rect 21959 13277 21971 13311
rect 21913 13271 21971 13277
rect 22005 13311 22063 13317
rect 22005 13277 22017 13311
rect 22051 13308 22063 13311
rect 22094 13308 22100 13320
rect 22051 13280 22100 13308
rect 22051 13277 22063 13280
rect 22005 13271 22063 13277
rect 22020 13240 22048 13271
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 24305 13311 24363 13317
rect 24305 13277 24317 13311
rect 24351 13277 24363 13311
rect 24305 13271 24363 13277
rect 24320 13240 24348 13271
rect 26418 13268 26424 13320
rect 26476 13308 26482 13320
rect 26973 13311 27031 13317
rect 26973 13308 26985 13311
rect 26476 13280 26985 13308
rect 26476 13268 26482 13280
rect 26973 13277 26985 13280
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27062 13268 27068 13320
rect 27120 13308 27126 13320
rect 27120 13280 27213 13308
rect 27120 13268 27126 13280
rect 27080 13240 27108 13268
rect 20732 13212 22048 13240
rect 23584 13212 24348 13240
rect 26344 13212 27108 13240
rect 15473 13203 15531 13209
rect 4154 13132 4160 13184
rect 4212 13172 4218 13184
rect 4249 13175 4307 13181
rect 4249 13172 4261 13175
rect 4212 13144 4261 13172
rect 4212 13132 4218 13144
rect 4249 13141 4261 13144
rect 4295 13141 4307 13175
rect 5258 13172 5264 13184
rect 5219 13144 5264 13172
rect 4249 13135 4307 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 6917 13175 6975 13181
rect 6917 13141 6929 13175
rect 6963 13172 6975 13175
rect 7098 13172 7104 13184
rect 6963 13144 7104 13172
rect 6963 13141 6975 13144
rect 6917 13135 6975 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 8478 13172 8484 13184
rect 8439 13144 8484 13172
rect 8478 13132 8484 13144
rect 8536 13132 8542 13184
rect 15013 13175 15071 13181
rect 15013 13141 15025 13175
rect 15059 13172 15071 13175
rect 15102 13172 15108 13184
rect 15059 13144 15108 13172
rect 15059 13141 15071 13144
rect 15013 13135 15071 13141
rect 15102 13132 15108 13144
rect 15160 13132 15166 13184
rect 16482 13172 16488 13184
rect 16443 13144 16488 13172
rect 16482 13132 16488 13144
rect 16540 13132 16546 13184
rect 17954 13172 17960 13184
rect 17915 13144 17960 13172
rect 17954 13132 17960 13144
rect 18012 13132 18018 13184
rect 21082 13172 21088 13184
rect 21043 13144 21088 13172
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 23290 13172 23296 13184
rect 23251 13144 23296 13172
rect 23290 13132 23296 13144
rect 23348 13132 23354 13184
rect 23474 13132 23480 13184
rect 23532 13172 23538 13184
rect 23584 13181 23612 13212
rect 26344 13184 26372 13212
rect 23569 13175 23627 13181
rect 23569 13172 23581 13175
rect 23532 13144 23581 13172
rect 23532 13132 23538 13144
rect 23569 13141 23581 13144
rect 23615 13141 23627 13175
rect 23750 13172 23756 13184
rect 23711 13144 23756 13172
rect 23569 13135 23627 13141
rect 23750 13132 23756 13144
rect 23808 13132 23814 13184
rect 24857 13175 24915 13181
rect 24857 13141 24869 13175
rect 24903 13172 24915 13175
rect 25038 13172 25044 13184
rect 24903 13144 25044 13172
rect 24903 13141 24915 13144
rect 24857 13135 24915 13141
rect 25038 13132 25044 13144
rect 25096 13132 25102 13184
rect 25130 13132 25136 13184
rect 25188 13172 25194 13184
rect 25188 13144 25233 13172
rect 25188 13132 25194 13144
rect 25406 13132 25412 13184
rect 25464 13172 25470 13184
rect 25501 13175 25559 13181
rect 25501 13172 25513 13175
rect 25464 13144 25513 13172
rect 25464 13132 25470 13144
rect 25501 13141 25513 13144
rect 25547 13141 25559 13175
rect 26326 13172 26332 13184
rect 26287 13144 26332 13172
rect 25501 13135 25559 13141
rect 26326 13132 26332 13144
rect 26384 13132 26390 13184
rect 26510 13172 26516 13184
rect 26471 13144 26516 13172
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 3050 12968 3056 12980
rect 3011 12940 3056 12968
rect 3050 12928 3056 12940
rect 3108 12928 3114 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4246 12968 4252 12980
rect 4203 12940 4252 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4982 12968 4988 12980
rect 4943 12940 4988 12968
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6454 12968 6460 12980
rect 6227 12940 6460 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6454 12928 6460 12940
rect 6512 12968 6518 12980
rect 6638 12968 6644 12980
rect 6512 12940 6644 12968
rect 6512 12928 6518 12940
rect 6638 12928 6644 12940
rect 6696 12928 6702 12980
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 6788 12940 7849 12968
rect 6788 12928 6794 12940
rect 7837 12937 7849 12940
rect 7883 12968 7895 12971
rect 8205 12971 8263 12977
rect 8205 12968 8217 12971
rect 7883 12940 8217 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 8205 12937 8217 12940
rect 8251 12937 8263 12971
rect 8205 12931 8263 12937
rect 6546 12900 6552 12912
rect 6507 12872 6552 12900
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 5258 12832 5264 12844
rect 4663 12804 5264 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 5258 12792 5264 12804
rect 5316 12832 5322 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5316 12804 5549 12832
rect 5316 12792 5322 12804
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 6362 12832 6368 12844
rect 5767 12804 6368 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 1670 12764 1676 12776
rect 1631 12736 1676 12764
rect 1670 12724 1676 12736
rect 1728 12724 1734 12776
rect 5166 12724 5172 12776
rect 5224 12764 5230 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5224 12736 5457 12764
rect 5224 12724 5230 12736
rect 5445 12733 5457 12736
rect 5491 12733 5503 12767
rect 6564 12764 6592 12860
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7285 12835 7343 12841
rect 7285 12832 7297 12835
rect 7064 12804 7297 12832
rect 7064 12792 7070 12804
rect 7285 12801 7297 12804
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12832 7527 12835
rect 7650 12832 7656 12844
rect 7515 12804 7656 12832
rect 7515 12801 7527 12804
rect 7469 12795 7527 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 8220 12832 8248 12931
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10689 12971 10747 12977
rect 10689 12968 10701 12971
rect 10468 12940 10701 12968
rect 10468 12928 10474 12940
rect 10689 12937 10701 12940
rect 10735 12968 10747 12971
rect 11330 12968 11336 12980
rect 10735 12940 11336 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 11330 12928 11336 12940
rect 11388 12928 11394 12980
rect 11514 12928 11520 12980
rect 11572 12968 11578 12980
rect 12250 12968 12256 12980
rect 11572 12940 12256 12968
rect 11572 12928 11578 12940
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 12492 12940 12537 12968
rect 12492 12928 12498 12940
rect 13538 12928 13544 12980
rect 13596 12968 13602 12980
rect 13633 12971 13691 12977
rect 13633 12968 13645 12971
rect 13596 12940 13645 12968
rect 13596 12928 13602 12940
rect 13633 12937 13645 12940
rect 13679 12968 13691 12971
rect 13814 12968 13820 12980
rect 13679 12940 13820 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 13814 12928 13820 12940
rect 13872 12928 13878 12980
rect 14090 12968 14096 12980
rect 14051 12940 14096 12968
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 16390 12968 16396 12980
rect 16351 12940 16396 12968
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 19794 12968 19800 12980
rect 18647 12940 19800 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 19794 12928 19800 12940
rect 19852 12928 19858 12980
rect 20070 12928 20076 12980
rect 20128 12968 20134 12980
rect 22373 12971 22431 12977
rect 22373 12968 22385 12971
rect 20128 12940 22385 12968
rect 20128 12928 20134 12940
rect 22373 12937 22385 12940
rect 22419 12937 22431 12971
rect 23014 12968 23020 12980
rect 22975 12940 23020 12968
rect 22373 12931 22431 12937
rect 23014 12928 23020 12940
rect 23072 12928 23078 12980
rect 23934 12968 23940 12980
rect 23895 12940 23940 12968
rect 23934 12928 23940 12940
rect 23992 12928 23998 12980
rect 24118 12928 24124 12980
rect 24176 12968 24182 12980
rect 24949 12971 25007 12977
rect 24949 12968 24961 12971
rect 24176 12940 24961 12968
rect 24176 12928 24182 12940
rect 24949 12937 24961 12940
rect 24995 12937 25007 12971
rect 25314 12968 25320 12980
rect 25275 12940 25320 12968
rect 24949 12931 25007 12937
rect 25314 12928 25320 12940
rect 25372 12928 25378 12980
rect 25774 12928 25780 12980
rect 25832 12968 25838 12980
rect 25961 12971 26019 12977
rect 25961 12968 25973 12971
rect 25832 12940 25973 12968
rect 25832 12928 25838 12940
rect 25961 12937 25973 12940
rect 26007 12968 26019 12971
rect 26418 12968 26424 12980
rect 26007 12940 26424 12968
rect 26007 12937 26019 12940
rect 25961 12931 26019 12937
rect 26418 12928 26424 12940
rect 26476 12928 26482 12980
rect 11054 12900 11060 12912
rect 11015 12872 11060 12900
rect 11054 12860 11060 12872
rect 11112 12860 11118 12912
rect 11885 12903 11943 12909
rect 11885 12869 11897 12903
rect 11931 12900 11943 12903
rect 11974 12900 11980 12912
rect 11931 12872 11980 12900
rect 11931 12869 11943 12872
rect 11885 12863 11943 12869
rect 11974 12860 11980 12872
rect 12032 12900 12038 12912
rect 12158 12900 12164 12912
rect 12032 12872 12164 12900
rect 12032 12860 12038 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 16758 12900 16764 12912
rect 15488 12872 16764 12900
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 8220 12804 8401 12832
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 10413 12835 10471 12841
rect 10413 12801 10425 12835
rect 10459 12832 10471 12835
rect 10594 12832 10600 12844
rect 10459 12804 10600 12832
rect 10459 12801 10471 12804
rect 10413 12795 10471 12801
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 13262 12832 13268 12844
rect 13127 12804 13268 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 13262 12792 13268 12804
rect 13320 12792 13326 12844
rect 15286 12832 15292 12844
rect 15247 12804 15292 12832
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15488 12841 15516 12872
rect 16758 12860 16764 12872
rect 16816 12860 16822 12912
rect 19429 12903 19487 12909
rect 19429 12869 19441 12903
rect 19475 12900 19487 12903
rect 20346 12900 20352 12912
rect 19475 12872 20352 12900
rect 19475 12869 19487 12872
rect 19429 12863 19487 12869
rect 20346 12860 20352 12872
rect 20404 12860 20410 12912
rect 20622 12860 20628 12912
rect 20680 12900 20686 12912
rect 20809 12903 20867 12909
rect 20809 12900 20821 12903
rect 20680 12872 20821 12900
rect 20680 12860 20686 12872
rect 20809 12869 20821 12872
rect 20855 12900 20867 12903
rect 20990 12900 20996 12912
rect 20855 12872 20996 12900
rect 20855 12869 20867 12872
rect 20809 12863 20867 12869
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 23477 12903 23535 12909
rect 23477 12869 23489 12903
rect 23523 12900 23535 12903
rect 24210 12900 24216 12912
rect 23523 12872 24216 12900
rect 23523 12869 23535 12872
rect 23477 12863 23535 12869
rect 24210 12860 24216 12872
rect 24268 12860 24274 12912
rect 24854 12900 24860 12912
rect 24412 12872 24860 12900
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12801 15531 12835
rect 15473 12795 15531 12801
rect 16482 12792 16488 12844
rect 16540 12832 16546 12844
rect 16853 12835 16911 12841
rect 16853 12832 16865 12835
rect 16540 12804 16865 12832
rect 16540 12792 16546 12804
rect 16853 12801 16865 12804
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17402 12832 17408 12844
rect 17083 12804 17408 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6564 12736 7205 12764
rect 5445 12727 5503 12733
rect 7193 12733 7205 12736
rect 7239 12764 7251 12767
rect 7374 12764 7380 12776
rect 7239 12736 7380 12764
rect 7239 12733 7251 12736
rect 7193 12727 7251 12733
rect 7374 12724 7380 12736
rect 7432 12724 7438 12776
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 8645 12767 8703 12773
rect 8645 12764 8657 12767
rect 8536 12736 8657 12764
rect 8536 12724 8542 12736
rect 8645 12733 8657 12736
rect 8691 12733 8703 12767
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 8645 12727 8703 12733
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 16301 12767 16359 12773
rect 16301 12733 16313 12767
rect 16347 12764 16359 12767
rect 17052 12764 17080 12795
rect 17402 12792 17408 12804
rect 17460 12832 17466 12844
rect 17954 12832 17960 12844
rect 17460 12804 17960 12832
rect 17460 12792 17466 12804
rect 17954 12792 17960 12804
rect 18012 12792 18018 12844
rect 19978 12832 19984 12844
rect 19939 12804 19984 12832
rect 19978 12792 19984 12804
rect 20036 12792 20042 12844
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 24412 12841 24440 12872
rect 24854 12860 24860 12872
rect 24912 12860 24918 12912
rect 28166 12900 28172 12912
rect 28127 12872 28172 12900
rect 28166 12860 28172 12872
rect 28224 12860 28230 12912
rect 24397 12835 24455 12841
rect 24397 12832 24409 12835
rect 23348 12804 24409 12832
rect 23348 12792 23354 12804
rect 24397 12801 24409 12804
rect 24443 12801 24455 12835
rect 24397 12795 24455 12801
rect 24581 12835 24639 12841
rect 24581 12801 24593 12835
rect 24627 12832 24639 12835
rect 25038 12832 25044 12844
rect 24627 12804 25044 12832
rect 24627 12801 24639 12804
rect 24581 12795 24639 12801
rect 25038 12792 25044 12804
rect 25096 12792 25102 12844
rect 25590 12792 25596 12844
rect 25648 12832 25654 12844
rect 26142 12832 26148 12844
rect 25648 12804 26148 12832
rect 25648 12792 25654 12804
rect 26142 12792 26148 12804
rect 26200 12792 26206 12844
rect 16347 12736 17080 12764
rect 20993 12767 21051 12773
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 20993 12733 21005 12767
rect 21039 12764 21051 12767
rect 21082 12764 21088 12776
rect 21039 12736 21088 12764
rect 21039 12733 21051 12736
rect 20993 12727 21051 12733
rect 1940 12699 1998 12705
rect 1940 12665 1952 12699
rect 1986 12665 1998 12699
rect 1940 12659 1998 12665
rect 1955 12628 1983 12659
rect 2866 12656 2872 12708
rect 2924 12696 2930 12708
rect 3326 12696 3332 12708
rect 2924 12668 3332 12696
rect 2924 12656 2930 12668
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8496 12696 8524 12724
rect 12158 12696 12164 12708
rect 8352 12668 8524 12696
rect 12119 12668 12164 12696
rect 8352 12656 8358 12668
rect 12158 12656 12164 12668
rect 12216 12696 12222 12708
rect 12897 12699 12955 12705
rect 12897 12696 12909 12699
rect 12216 12668 12909 12696
rect 12216 12656 12222 12668
rect 12897 12665 12909 12668
rect 12943 12665 12955 12699
rect 16761 12699 16819 12705
rect 16761 12696 16773 12699
rect 12897 12659 12955 12665
rect 14844 12668 16773 12696
rect 3694 12628 3700 12640
rect 1955 12600 3700 12628
rect 3694 12588 3700 12600
rect 3752 12588 3758 12640
rect 5077 12631 5135 12637
rect 5077 12597 5089 12631
rect 5123 12628 5135 12631
rect 5350 12628 5356 12640
rect 5123 12600 5356 12628
rect 5123 12597 5135 12600
rect 5077 12591 5135 12597
rect 5350 12588 5356 12600
rect 5408 12588 5414 12640
rect 6730 12588 6736 12640
rect 6788 12628 6794 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6788 12600 6837 12628
rect 6788 12588 6794 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 6825 12591 6883 12597
rect 9769 12631 9827 12637
rect 9769 12597 9781 12631
rect 9815 12628 9827 12631
rect 10226 12628 10232 12640
rect 9815 12600 10232 12628
rect 9815 12597 9827 12600
rect 9769 12591 9827 12597
rect 10226 12588 10232 12600
rect 10284 12588 10290 12640
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 14844 12637 14872 12668
rect 16761 12665 16773 12668
rect 16807 12696 16819 12699
rect 17773 12699 17831 12705
rect 17773 12696 17785 12699
rect 16807 12668 17785 12696
rect 16807 12665 16819 12668
rect 16761 12659 16819 12665
rect 17773 12665 17785 12668
rect 17819 12665 17831 12699
rect 17773 12659 17831 12665
rect 19797 12699 19855 12705
rect 19797 12665 19809 12699
rect 19843 12696 19855 12699
rect 20622 12696 20628 12708
rect 19843 12668 20628 12696
rect 19843 12665 19855 12668
rect 19797 12659 19855 12665
rect 20622 12656 20628 12668
rect 20680 12656 20686 12708
rect 14829 12631 14887 12637
rect 14829 12597 14841 12631
rect 14875 12597 14887 12631
rect 15194 12628 15200 12640
rect 15155 12600 15200 12628
rect 14829 12591 14887 12597
rect 15194 12588 15200 12600
rect 15252 12588 15258 12640
rect 15838 12628 15844 12640
rect 15799 12600 15844 12628
rect 15838 12588 15844 12600
rect 15896 12588 15902 12640
rect 17126 12588 17132 12640
rect 17184 12628 17190 12640
rect 17405 12631 17463 12637
rect 17405 12628 17417 12631
rect 17184 12600 17417 12628
rect 17184 12588 17190 12600
rect 17405 12597 17417 12600
rect 17451 12597 17463 12631
rect 18966 12628 18972 12640
rect 18927 12600 18972 12628
rect 17405 12591 17463 12597
rect 18966 12588 18972 12600
rect 19024 12588 19030 12640
rect 19337 12631 19395 12637
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 19702 12628 19708 12640
rect 19383 12600 19708 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12628 19947 12631
rect 20254 12628 20260 12640
rect 19935 12600 20260 12628
rect 19935 12597 19947 12600
rect 19889 12591 19947 12597
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20346 12588 20352 12640
rect 20404 12628 20410 12640
rect 20441 12631 20499 12637
rect 20441 12628 20453 12631
rect 20404 12600 20453 12628
rect 20404 12588 20410 12600
rect 20441 12597 20453 12600
rect 20487 12628 20499 12631
rect 21008 12628 21036 12727
rect 21082 12724 21088 12736
rect 21140 12724 21146 12776
rect 23658 12724 23664 12776
rect 23716 12764 23722 12776
rect 24305 12767 24363 12773
rect 24305 12764 24317 12767
rect 23716 12736 24317 12764
rect 23716 12724 23722 12736
rect 24305 12733 24317 12736
rect 24351 12764 24363 12767
rect 25130 12764 25136 12776
rect 24351 12736 25136 12764
rect 24351 12733 24363 12736
rect 24305 12727 24363 12733
rect 25130 12724 25136 12736
rect 25188 12724 25194 12776
rect 21266 12705 21272 12708
rect 21260 12659 21272 12705
rect 21324 12696 21330 12708
rect 21324 12668 21360 12696
rect 21266 12656 21272 12659
rect 21324 12656 21330 12668
rect 26234 12656 26240 12708
rect 26292 12696 26298 12708
rect 26390 12699 26448 12705
rect 26390 12696 26402 12699
rect 26292 12668 26402 12696
rect 26292 12656 26298 12668
rect 26390 12665 26402 12668
rect 26436 12665 26448 12699
rect 26390 12659 26448 12665
rect 27522 12628 27528 12640
rect 20487 12600 21036 12628
rect 27483 12600 27528 12628
rect 20487 12597 20499 12600
rect 20441 12591 20499 12597
rect 27522 12588 27528 12600
rect 27580 12588 27586 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 1670 12424 1676 12436
rect 1631 12396 1676 12424
rect 1670 12384 1676 12396
rect 1728 12424 1734 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1728 12396 1961 12424
rect 1728 12384 1734 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 4522 12424 4528 12436
rect 4435 12396 4528 12424
rect 1949 12387 2007 12393
rect 4522 12384 4528 12396
rect 4580 12424 4586 12436
rect 5258 12424 5264 12436
rect 4580 12396 5264 12424
rect 4580 12384 4586 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 5353 12427 5411 12433
rect 5353 12393 5365 12427
rect 5399 12424 5411 12427
rect 5442 12424 5448 12436
rect 5399 12396 5448 12424
rect 5399 12393 5411 12396
rect 5353 12387 5411 12393
rect 5442 12384 5448 12396
rect 5500 12384 5506 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 5552 12396 7021 12424
rect 3237 12359 3295 12365
rect 3237 12325 3249 12359
rect 3283 12356 3295 12359
rect 3510 12356 3516 12368
rect 3283 12328 3516 12356
rect 3283 12325 3295 12328
rect 3237 12319 3295 12325
rect 3510 12316 3516 12328
rect 3568 12356 3574 12368
rect 5552 12356 5580 12396
rect 7009 12393 7021 12396
rect 7055 12393 7067 12427
rect 7009 12387 7067 12393
rect 8021 12427 8079 12433
rect 8021 12393 8033 12427
rect 8067 12424 8079 12427
rect 8386 12424 8392 12436
rect 8067 12396 8392 12424
rect 8067 12393 8079 12396
rect 8021 12387 8079 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 12894 12424 12900 12436
rect 12855 12396 12900 12424
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 15565 12427 15623 12433
rect 15565 12393 15577 12427
rect 15611 12424 15623 12427
rect 16482 12424 16488 12436
rect 15611 12396 16488 12424
rect 15611 12393 15623 12396
rect 15565 12387 15623 12393
rect 16482 12384 16488 12396
rect 16540 12384 16546 12436
rect 16669 12427 16727 12433
rect 16669 12393 16681 12427
rect 16715 12424 16727 12427
rect 16758 12424 16764 12436
rect 16715 12396 16764 12424
rect 16715 12393 16727 12396
rect 16669 12387 16727 12393
rect 3568 12328 5580 12356
rect 3568 12316 3574 12328
rect 5810 12316 5816 12368
rect 5868 12365 5874 12368
rect 5868 12359 5932 12365
rect 5868 12325 5886 12359
rect 5920 12325 5932 12359
rect 5868 12319 5932 12325
rect 5868 12316 5874 12319
rect 10226 12316 10232 12368
rect 10284 12365 10290 12368
rect 10284 12359 10348 12365
rect 10284 12325 10302 12359
rect 10336 12325 10348 12359
rect 10284 12319 10348 12325
rect 10284 12316 10290 12319
rect 2777 12291 2835 12297
rect 2777 12257 2789 12291
rect 2823 12288 2835 12291
rect 4062 12288 4068 12300
rect 2823 12260 4068 12288
rect 2823 12257 2835 12260
rect 2777 12251 2835 12257
rect 4062 12248 4068 12260
rect 4120 12248 4126 12300
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 5828 12288 5856 12316
rect 4433 12251 4491 12257
rect 4724 12260 5856 12288
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 3053 12223 3111 12229
rect 3053 12189 3065 12223
rect 3099 12220 3111 12223
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3099 12192 3249 12220
rect 3099 12189 3111 12192
rect 3053 12183 3111 12189
rect 3237 12189 3249 12192
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 2884 12152 2912 12183
rect 4448 12152 4476 12251
rect 4724 12229 4752 12260
rect 12710 12248 12716 12300
rect 12768 12288 12774 12300
rect 12986 12288 12992 12300
rect 12768 12260 12992 12288
rect 12768 12248 12774 12260
rect 12986 12248 12992 12260
rect 13044 12248 13050 12300
rect 15378 12248 15384 12300
rect 15436 12288 15442 12300
rect 15933 12291 15991 12297
rect 15933 12288 15945 12291
rect 15436 12260 15945 12288
rect 15436 12248 15442 12260
rect 15933 12257 15945 12260
rect 15979 12257 15991 12291
rect 15933 12251 15991 12257
rect 4709 12223 4767 12229
rect 4709 12189 4721 12223
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5629 12223 5687 12229
rect 5629 12189 5641 12223
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 4798 12152 4804 12164
rect 2884 12124 3924 12152
rect 4448 12124 4804 12152
rect 3896 12096 3924 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 2409 12087 2467 12093
rect 2409 12053 2421 12087
rect 2455 12084 2467 12087
rect 2590 12084 2596 12096
rect 2455 12056 2596 12084
rect 2455 12053 2467 12056
rect 2409 12047 2467 12053
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 3878 12084 3884 12096
rect 3839 12056 3884 12084
rect 3878 12044 3884 12056
rect 3936 12044 3942 12096
rect 4062 12084 4068 12096
rect 4023 12056 4068 12084
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 5644 12084 5672 12183
rect 7190 12180 7196 12232
rect 7248 12220 7254 12232
rect 7248 12192 8800 12220
rect 7248 12180 7254 12192
rect 7650 12152 7656 12164
rect 7563 12124 7656 12152
rect 7650 12112 7656 12124
rect 7708 12152 7714 12164
rect 8662 12152 8668 12164
rect 7708 12124 8668 12152
rect 7708 12112 7714 12124
rect 8662 12112 8668 12124
rect 8720 12112 8726 12164
rect 8772 12096 8800 12192
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9824 12192 10057 12220
rect 9824 12180 9830 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 12158 12180 12164 12232
rect 12216 12220 12222 12232
rect 13081 12223 13139 12229
rect 13081 12220 13093 12223
rect 12216 12192 13093 12220
rect 12216 12180 12222 12192
rect 13081 12189 13093 12192
rect 13127 12189 13139 12223
rect 13081 12183 13139 12189
rect 14826 12180 14832 12232
rect 14884 12220 14890 12232
rect 15838 12220 15844 12232
rect 14884 12192 15844 12220
rect 14884 12180 14890 12192
rect 15838 12180 15844 12192
rect 15896 12220 15902 12232
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15896 12192 16037 12220
rect 15896 12180 15902 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12220 16267 12223
rect 16684 12220 16712 12387
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 19978 12424 19984 12436
rect 19567 12396 19984 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 26142 12424 26148 12436
rect 26103 12396 26148 12424
rect 26142 12384 26148 12396
rect 26200 12384 26206 12436
rect 26510 12384 26516 12436
rect 26568 12424 26574 12436
rect 26973 12427 27031 12433
rect 26973 12424 26985 12427
rect 26568 12396 26985 12424
rect 26568 12384 26574 12396
rect 26973 12393 26985 12396
rect 27019 12424 27031 12427
rect 27525 12427 27583 12433
rect 27525 12424 27537 12427
rect 27019 12396 27537 12424
rect 27019 12393 27031 12396
rect 26973 12387 27031 12393
rect 27525 12393 27537 12396
rect 27571 12393 27583 12427
rect 27525 12387 27583 12393
rect 17402 12297 17408 12300
rect 17396 12288 17408 12297
rect 17363 12260 17408 12288
rect 17396 12251 17408 12260
rect 17402 12248 17408 12251
rect 17460 12248 17466 12300
rect 20162 12248 20168 12300
rect 20220 12288 20226 12300
rect 21157 12291 21215 12297
rect 21157 12288 21169 12291
rect 20220 12260 21169 12288
rect 20220 12248 20226 12260
rect 21157 12257 21169 12260
rect 21203 12257 21215 12291
rect 21157 12251 21215 12257
rect 23293 12291 23351 12297
rect 23293 12257 23305 12291
rect 23339 12288 23351 12291
rect 23474 12288 23480 12300
rect 23339 12260 23480 12288
rect 23339 12257 23351 12260
rect 23293 12251 23351 12257
rect 23474 12248 23480 12260
rect 23532 12288 23538 12300
rect 23652 12291 23710 12297
rect 23652 12288 23664 12291
rect 23532 12260 23664 12288
rect 23532 12248 23538 12260
rect 23652 12257 23664 12260
rect 23698 12288 23710 12291
rect 24486 12288 24492 12300
rect 23698 12260 24492 12288
rect 23698 12257 23710 12260
rect 23652 12251 23710 12257
rect 24486 12248 24492 12260
rect 24544 12248 24550 12300
rect 25869 12291 25927 12297
rect 25869 12257 25881 12291
rect 25915 12288 25927 12291
rect 26142 12288 26148 12300
rect 25915 12260 26148 12288
rect 25915 12257 25927 12260
rect 25869 12251 25927 12257
rect 26142 12248 26148 12260
rect 26200 12248 26206 12300
rect 26602 12248 26608 12300
rect 26660 12288 26666 12300
rect 26881 12291 26939 12297
rect 26881 12288 26893 12291
rect 26660 12260 26893 12288
rect 26660 12248 26666 12260
rect 26881 12257 26893 12260
rect 26927 12257 26939 12291
rect 26881 12251 26939 12257
rect 17126 12220 17132 12232
rect 16255 12192 16712 12220
rect 17087 12192 17132 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 13633 12155 13691 12161
rect 13633 12121 13645 12155
rect 13679 12152 13691 12155
rect 14458 12152 14464 12164
rect 13679 12124 14464 12152
rect 13679 12121 13691 12124
rect 13633 12115 13691 12121
rect 14458 12112 14464 12124
rect 14516 12112 14522 12164
rect 14921 12155 14979 12161
rect 14921 12121 14933 12155
rect 14967 12152 14979 12155
rect 15654 12152 15660 12164
rect 14967 12124 15660 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 15654 12112 15660 12124
rect 15712 12152 15718 12164
rect 16224 12152 16252 12183
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 20622 12220 20628 12232
rect 19843 12192 20628 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 20898 12220 20904 12232
rect 20859 12192 20904 12220
rect 20898 12180 20904 12192
rect 20956 12180 20962 12232
rect 23385 12223 23443 12229
rect 23385 12189 23397 12223
rect 23431 12189 23443 12223
rect 23385 12183 23443 12189
rect 27157 12223 27215 12229
rect 27157 12189 27169 12223
rect 27203 12220 27215 12223
rect 27522 12220 27528 12232
rect 27203 12192 27528 12220
rect 27203 12189 27215 12192
rect 27157 12183 27215 12189
rect 15712 12124 16252 12152
rect 15712 12112 15718 12124
rect 23290 12112 23296 12164
rect 23348 12152 23354 12164
rect 23400 12152 23428 12183
rect 27522 12180 27528 12192
rect 27580 12180 27586 12232
rect 23348 12124 23428 12152
rect 23348 12112 23354 12124
rect 6362 12084 6368 12096
rect 5644 12056 6368 12084
rect 6362 12044 6368 12056
rect 6420 12084 6426 12096
rect 6546 12084 6552 12096
rect 6420 12056 6552 12084
rect 6420 12044 6426 12056
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8352 12056 8401 12084
rect 8352 12044 8358 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8754 12084 8760 12096
rect 8715 12056 8760 12084
rect 8389 12047 8447 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 11422 12084 11428 12096
rect 11383 12056 11428 12084
rect 11422 12044 11428 12056
rect 11480 12084 11486 12096
rect 11882 12084 11888 12096
rect 11480 12056 11888 12084
rect 11480 12044 11486 12056
rect 11882 12044 11888 12056
rect 11940 12084 11946 12096
rect 11977 12087 12035 12093
rect 11977 12084 11989 12087
rect 11940 12056 11989 12084
rect 11940 12044 11946 12056
rect 11977 12053 11989 12056
rect 12023 12053 12035 12087
rect 12526 12084 12532 12096
rect 12487 12056 12532 12084
rect 11977 12047 12035 12053
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 14550 12084 14556 12096
rect 14511 12056 14556 12084
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 17034 12084 17040 12096
rect 16995 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12084 17098 12096
rect 18414 12084 18420 12096
rect 17092 12056 18420 12084
rect 17092 12044 17098 12056
rect 18414 12044 18420 12056
rect 18472 12084 18478 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 18472 12056 18521 12084
rect 18472 12044 18478 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 20254 12084 20260 12096
rect 20215 12056 20260 12084
rect 18509 12047 18567 12053
rect 20254 12044 20260 12056
rect 20312 12044 20318 12096
rect 20438 12044 20444 12096
rect 20496 12084 20502 12096
rect 20625 12087 20683 12093
rect 20625 12084 20637 12087
rect 20496 12056 20637 12084
rect 20496 12044 20502 12056
rect 20625 12053 20637 12056
rect 20671 12084 20683 12087
rect 21266 12084 21272 12096
rect 20671 12056 21272 12084
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 21266 12044 21272 12056
rect 21324 12084 21330 12096
rect 22281 12087 22339 12093
rect 22281 12084 22293 12087
rect 21324 12056 22293 12084
rect 21324 12044 21330 12056
rect 22281 12053 22293 12056
rect 22327 12053 22339 12087
rect 22281 12047 22339 12053
rect 24302 12044 24308 12096
rect 24360 12084 24366 12096
rect 24765 12087 24823 12093
rect 24765 12084 24777 12087
rect 24360 12056 24777 12084
rect 24360 12044 24366 12056
rect 24765 12053 24777 12056
rect 24811 12084 24823 12087
rect 25409 12087 25467 12093
rect 25409 12084 25421 12087
rect 24811 12056 25421 12084
rect 24811 12053 24823 12056
rect 24765 12047 24823 12053
rect 25409 12053 25421 12056
rect 25455 12084 25467 12087
rect 25774 12084 25780 12096
rect 25455 12056 25780 12084
rect 25455 12053 25467 12056
rect 25409 12047 25467 12053
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 25866 12044 25872 12096
rect 25924 12084 25930 12096
rect 26513 12087 26571 12093
rect 26513 12084 26525 12087
rect 25924 12056 26525 12084
rect 25924 12044 25930 12056
rect 26513 12053 26525 12056
rect 26559 12053 26571 12087
rect 26513 12047 26571 12053
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1728 11852 2145 11880
rect 1728 11840 1734 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 6641 11883 6699 11889
rect 6641 11849 6653 11883
rect 6687 11880 6699 11883
rect 7190 11880 7196 11892
rect 6687 11852 7196 11880
rect 6687 11849 6699 11852
rect 6641 11843 6699 11849
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1762 11744 1768 11756
rect 1719 11716 1768 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 1762 11704 1768 11716
rect 1820 11704 1826 11756
rect 2148 11744 2176 11843
rect 4341 11815 4399 11821
rect 4341 11781 4353 11815
rect 4387 11812 4399 11815
rect 4522 11812 4528 11824
rect 4387 11784 4528 11812
rect 4387 11781 4399 11784
rect 4341 11775 4399 11781
rect 4522 11772 4528 11784
rect 4580 11772 4586 11824
rect 2314 11744 2320 11756
rect 2148 11716 2320 11744
rect 2314 11704 2320 11716
rect 2372 11704 2378 11756
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6656 11744 6684 11843
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7469 11883 7527 11889
rect 7469 11849 7481 11883
rect 7515 11880 7527 11883
rect 7558 11880 7564 11892
rect 7515 11852 7564 11880
rect 7515 11849 7527 11852
rect 7469 11843 7527 11849
rect 5859 11716 6684 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 2406 11636 2412 11688
rect 2464 11676 2470 11688
rect 6825 11679 6883 11685
rect 2464 11648 5948 11676
rect 2464 11636 2470 11648
rect 2584 11611 2642 11617
rect 2584 11577 2596 11611
rect 2630 11608 2642 11611
rect 3510 11608 3516 11620
rect 2630 11580 3516 11608
rect 2630 11577 2642 11580
rect 2584 11571 2642 11577
rect 3510 11568 3516 11580
rect 3568 11568 3574 11620
rect 5077 11611 5135 11617
rect 5077 11577 5089 11611
rect 5123 11608 5135 11611
rect 5810 11608 5816 11620
rect 5123 11580 5816 11608
rect 5123 11577 5135 11580
rect 5077 11571 5135 11577
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 5920 11608 5948 11648
rect 6825 11645 6837 11679
rect 6871 11676 6883 11679
rect 7484 11676 7512 11843
rect 7558 11840 7564 11852
rect 7616 11840 7622 11892
rect 9766 11880 9772 11892
rect 9727 11852 9772 11880
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10229 11883 10287 11889
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10870 11880 10876 11892
rect 10275 11852 10876 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 14826 11880 14832 11892
rect 14787 11852 14832 11880
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 20530 11840 20536 11892
rect 20588 11880 20594 11892
rect 21453 11883 21511 11889
rect 21453 11880 21465 11883
rect 20588 11852 21465 11880
rect 20588 11840 20594 11852
rect 21453 11849 21465 11852
rect 21499 11849 21511 11883
rect 21453 11843 21511 11849
rect 22830 11840 22836 11892
rect 22888 11880 22894 11892
rect 23017 11883 23075 11889
rect 23017 11880 23029 11883
rect 22888 11852 23029 11880
rect 22888 11840 22894 11852
rect 23017 11849 23029 11852
rect 23063 11880 23075 11883
rect 23063 11852 24348 11880
rect 23063 11849 23075 11852
rect 23017 11843 23075 11849
rect 11698 11772 11704 11824
rect 11756 11812 11762 11824
rect 11885 11815 11943 11821
rect 11885 11812 11897 11815
rect 11756 11784 11897 11812
rect 11756 11772 11762 11784
rect 11885 11781 11897 11784
rect 11931 11812 11943 11815
rect 12158 11812 12164 11824
rect 11931 11784 12164 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 12158 11772 12164 11784
rect 12216 11772 12222 11824
rect 12710 11812 12716 11824
rect 12671 11784 12716 11812
rect 12710 11772 12716 11784
rect 12768 11772 12774 11824
rect 20346 11772 20352 11824
rect 20404 11812 20410 11824
rect 20625 11815 20683 11821
rect 20625 11812 20637 11815
rect 20404 11784 20637 11812
rect 20404 11772 20410 11784
rect 20625 11781 20637 11784
rect 20671 11812 20683 11815
rect 20898 11812 20904 11824
rect 20671 11784 20904 11812
rect 20671 11781 20683 11784
rect 20625 11775 20683 11781
rect 20898 11772 20904 11784
rect 20956 11812 20962 11824
rect 23290 11812 23296 11824
rect 20956 11784 23296 11812
rect 20956 11772 20962 11784
rect 23290 11772 23296 11784
rect 23348 11772 23354 11824
rect 23474 11812 23480 11824
rect 23435 11784 23480 11812
rect 23474 11772 23480 11784
rect 23532 11772 23538 11824
rect 8573 11747 8631 11753
rect 8573 11713 8585 11747
rect 8619 11744 8631 11747
rect 8662 11744 8668 11756
rect 8619 11716 8668 11744
rect 8619 11713 8631 11716
rect 8573 11707 8631 11713
rect 8662 11704 8668 11716
rect 8720 11744 8726 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8720 11716 8953 11744
rect 8720 11704 8726 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 10781 11747 10839 11753
rect 10781 11744 10793 11747
rect 9447 11716 10793 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 10781 11713 10793 11716
rect 10827 11744 10839 11747
rect 11422 11744 11428 11756
rect 10827 11716 11428 11744
rect 10827 11713 10839 11716
rect 10781 11707 10839 11713
rect 11422 11704 11428 11716
rect 11480 11704 11486 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12894 11744 12900 11756
rect 12299 11716 12900 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12894 11704 12900 11716
rect 12952 11704 12958 11756
rect 12986 11704 12992 11756
rect 13044 11744 13050 11756
rect 13725 11747 13783 11753
rect 13725 11744 13737 11747
rect 13044 11716 13737 11744
rect 13044 11704 13050 11716
rect 13725 11713 13737 11716
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 13909 11747 13967 11753
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 14458 11744 14464 11756
rect 13955 11716 14464 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 14458 11704 14464 11716
rect 14516 11744 14522 11756
rect 14918 11744 14924 11756
rect 14516 11716 14924 11744
rect 14516 11704 14522 11716
rect 14918 11704 14924 11716
rect 14976 11744 14982 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14976 11716 15485 11744
rect 14976 11704 14982 11716
rect 15473 11713 15485 11716
rect 15519 11744 15531 11747
rect 15746 11744 15752 11756
rect 15519 11716 15752 11744
rect 15519 11713 15531 11716
rect 15473 11707 15531 11713
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 16482 11744 16488 11756
rect 15804 11716 16488 11744
rect 15804 11704 15810 11716
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 17034 11744 17040 11756
rect 16995 11716 17040 11744
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 17126 11704 17132 11756
rect 17184 11744 17190 11756
rect 17497 11747 17555 11753
rect 17497 11744 17509 11747
rect 17184 11716 17509 11744
rect 17184 11704 17190 11716
rect 17497 11713 17509 11716
rect 17543 11744 17555 11747
rect 17543 11716 17908 11744
rect 17543 11713 17555 11716
rect 17497 11707 17555 11713
rect 6871 11648 7512 11676
rect 8297 11679 8355 11685
rect 6871 11645 6883 11648
rect 6825 11639 6883 11645
rect 8297 11645 8309 11679
rect 8343 11676 8355 11679
rect 8386 11676 8392 11688
rect 8343 11648 8392 11676
rect 8343 11645 8355 11648
rect 8297 11639 8355 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10502 11676 10508 11688
rect 10183 11648 10508 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 10502 11636 10508 11648
rect 10560 11676 10566 11688
rect 10597 11679 10655 11685
rect 10597 11676 10609 11679
rect 10560 11648 10609 11676
rect 10560 11636 10566 11648
rect 10597 11645 10609 11648
rect 10643 11645 10655 11679
rect 10597 11639 10655 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11676 13231 11679
rect 13630 11676 13636 11688
rect 13219 11648 13636 11676
rect 13219 11645 13231 11648
rect 13173 11639 13231 11645
rect 13630 11636 13636 11648
rect 13688 11636 13694 11688
rect 14737 11679 14795 11685
rect 14737 11645 14749 11679
rect 14783 11676 14795 11679
rect 15197 11679 15255 11685
rect 15197 11676 15209 11679
rect 14783 11648 15209 11676
rect 14783 11645 14795 11648
rect 14737 11639 14795 11645
rect 15197 11645 15209 11648
rect 15243 11676 15255 11679
rect 15286 11676 15292 11688
rect 15243 11648 15292 11676
rect 15243 11645 15255 11648
rect 15197 11639 15255 11645
rect 15286 11636 15292 11648
rect 15344 11636 15350 11688
rect 15838 11676 15844 11688
rect 15799 11648 15844 11676
rect 15838 11636 15844 11648
rect 15896 11676 15902 11688
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 15896 11648 16773 11676
rect 15896 11636 15902 11648
rect 16761 11645 16773 11648
rect 16807 11676 16819 11679
rect 16942 11676 16948 11688
rect 16807 11648 16948 11676
rect 16807 11645 16819 11648
rect 16761 11639 16819 11645
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 17770 11636 17776 11688
rect 17828 11636 17834 11688
rect 17880 11685 17908 11716
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 22465 11747 22523 11753
rect 22465 11744 22477 11747
rect 22152 11716 22477 11744
rect 22152 11704 22158 11716
rect 22465 11713 22477 11716
rect 22511 11713 22523 11747
rect 22465 11707 22523 11713
rect 18414 11685 18420 11688
rect 17865 11679 17923 11685
rect 17865 11645 17877 11679
rect 17911 11676 17923 11679
rect 18141 11679 18199 11685
rect 18141 11676 18153 11679
rect 17911 11648 18153 11676
rect 17911 11645 17923 11648
rect 17865 11639 17923 11645
rect 18141 11645 18153 11648
rect 18187 11645 18199 11679
rect 18408 11676 18420 11685
rect 18375 11648 18420 11676
rect 18141 11639 18199 11645
rect 18408 11639 18420 11648
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 5920 11580 7849 11608
rect 7837 11577 7849 11580
rect 7883 11608 7895 11611
rect 14369 11611 14427 11617
rect 7883 11580 8432 11608
rect 7883 11577 7895 11580
rect 7837 11571 7895 11577
rect 8404 11552 8432 11580
rect 14369 11577 14381 11611
rect 14415 11608 14427 11611
rect 16853 11611 16911 11617
rect 16853 11608 16865 11611
rect 14415 11580 15332 11608
rect 14415 11577 14427 11580
rect 14369 11571 14427 11577
rect 15304 11552 15332 11580
rect 16224 11580 16865 11608
rect 16224 11552 16252 11580
rect 16853 11577 16865 11580
rect 16899 11608 16911 11611
rect 17788 11608 17816 11636
rect 16899 11580 17816 11608
rect 18156 11608 18184 11639
rect 18414 11636 18420 11639
rect 18472 11636 18478 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20530 11676 20536 11688
rect 20036 11648 20536 11676
rect 20036 11636 20042 11648
rect 20530 11636 20536 11648
rect 20588 11676 20594 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20588 11648 21005 11676
rect 20588 11636 20594 11648
rect 20993 11645 21005 11648
rect 21039 11676 21051 11679
rect 21818 11676 21824 11688
rect 21039 11648 21824 11676
rect 21039 11645 21051 11648
rect 20993 11639 21051 11645
rect 21818 11636 21824 11648
rect 21876 11636 21882 11688
rect 23492 11676 23520 11772
rect 24320 11753 24348 11852
rect 24854 11840 24860 11892
rect 24912 11880 24918 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 24912 11852 25421 11880
rect 24912 11840 24918 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 26786 11880 26792 11892
rect 26747 11852 26792 11880
rect 25409 11843 25467 11849
rect 26786 11840 26792 11852
rect 26844 11880 26850 11892
rect 27154 11880 27160 11892
rect 26844 11852 27160 11880
rect 26844 11840 26850 11852
rect 27154 11840 27160 11852
rect 27212 11840 27218 11892
rect 25774 11772 25780 11824
rect 25832 11812 25838 11824
rect 27985 11815 28043 11821
rect 27985 11812 27997 11815
rect 25832 11784 26004 11812
rect 25832 11772 25838 11784
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11713 24363 11747
rect 24486 11744 24492 11756
rect 24399 11716 24492 11744
rect 24305 11707 24363 11713
rect 24486 11704 24492 11716
rect 24544 11744 24550 11756
rect 24949 11747 25007 11753
rect 24949 11744 24961 11747
rect 24544 11716 24961 11744
rect 24544 11704 24550 11716
rect 24949 11713 24961 11716
rect 24995 11744 25007 11747
rect 25225 11747 25283 11753
rect 25225 11744 25237 11747
rect 24995 11716 25237 11744
rect 24995 11713 25007 11716
rect 24949 11707 25007 11713
rect 25225 11713 25237 11716
rect 25271 11744 25283 11747
rect 25866 11744 25872 11756
rect 25271 11716 25452 11744
rect 25827 11716 25872 11744
rect 25271 11713 25283 11716
rect 25225 11707 25283 11713
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 23492 11648 24225 11676
rect 24213 11645 24225 11648
rect 24259 11676 24271 11679
rect 25314 11676 25320 11688
rect 24259 11648 25320 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 25314 11636 25320 11648
rect 25372 11636 25378 11688
rect 25424 11676 25452 11716
rect 25866 11704 25872 11716
rect 25924 11704 25930 11756
rect 25976 11753 26004 11784
rect 27448 11784 27997 11812
rect 27448 11756 27476 11784
rect 27985 11781 27997 11784
rect 28031 11781 28043 11815
rect 27985 11775 28043 11781
rect 25961 11747 26019 11753
rect 25961 11713 25973 11747
rect 26007 11713 26019 11747
rect 26602 11744 26608 11756
rect 26563 11716 26608 11744
rect 25961 11707 26019 11713
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 27430 11744 27436 11756
rect 27391 11716 27436 11744
rect 27430 11704 27436 11716
rect 27488 11704 27494 11756
rect 27522 11704 27528 11756
rect 27580 11744 27586 11756
rect 27580 11716 27625 11744
rect 27580 11704 27586 11716
rect 27540 11676 27568 11704
rect 25424 11648 27568 11676
rect 20346 11608 20352 11620
rect 18156 11580 20352 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 20346 11568 20352 11580
rect 20404 11568 20410 11620
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 21634 11608 21640 11620
rect 20864 11580 21640 11608
rect 20864 11568 20870 11580
rect 21634 11568 21640 11580
rect 21692 11568 21698 11620
rect 24946 11568 24952 11620
rect 25004 11608 25010 11620
rect 25777 11611 25835 11617
rect 25777 11608 25789 11611
rect 25004 11580 25789 11608
rect 25004 11568 25010 11580
rect 25777 11577 25789 11580
rect 25823 11608 25835 11611
rect 25823 11580 27016 11608
rect 25823 11577 25835 11580
rect 25777 11571 25835 11577
rect 3694 11540 3700 11552
rect 3655 11512 3700 11540
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 4709 11543 4767 11549
rect 4709 11509 4721 11543
rect 4755 11540 4767 11543
rect 4798 11540 4804 11552
rect 4755 11512 4804 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 4798 11500 4804 11512
rect 4856 11500 4862 11552
rect 5166 11540 5172 11552
rect 5127 11512 5172 11540
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5534 11540 5540 11552
rect 5495 11512 5540 11540
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 6273 11543 6331 11549
rect 5684 11512 5729 11540
rect 5684 11500 5690 11512
rect 6273 11509 6285 11543
rect 6319 11540 6331 11543
rect 6362 11540 6368 11552
rect 6319 11512 6368 11540
rect 6319 11509 6331 11512
rect 6273 11503 6331 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 7009 11543 7067 11549
rect 7009 11509 7021 11543
rect 7055 11540 7067 11543
rect 7098 11540 7104 11552
rect 7055 11512 7104 11540
rect 7055 11509 7067 11512
rect 7009 11503 7067 11509
rect 7098 11500 7104 11512
rect 7156 11500 7162 11552
rect 7929 11543 7987 11549
rect 7929 11509 7941 11543
rect 7975 11540 7987 11543
rect 8202 11540 8208 11552
rect 7975 11512 8208 11540
rect 7975 11509 7987 11512
rect 7929 11503 7987 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8386 11540 8392 11552
rect 8347 11512 8392 11540
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 10318 11500 10324 11552
rect 10376 11540 10382 11552
rect 10689 11543 10747 11549
rect 10689 11540 10701 11543
rect 10376 11512 10701 11540
rect 10376 11500 10382 11512
rect 10689 11509 10701 11512
rect 10735 11540 10747 11543
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 10735 11512 11253 11540
rect 10735 11509 10747 11512
rect 10689 11503 10747 11509
rect 11241 11509 11253 11512
rect 11287 11509 11299 11543
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 11241 11503 11299 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 15286 11540 15292 11552
rect 15247 11512 15292 11540
rect 15286 11500 15292 11512
rect 15344 11500 15350 11552
rect 16206 11540 16212 11552
rect 16167 11512 16212 11540
rect 16206 11500 16212 11512
rect 16264 11500 16270 11552
rect 16390 11540 16396 11552
rect 16351 11512 16396 11540
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 19521 11543 19579 11549
rect 19521 11509 19533 11543
rect 19567 11540 19579 11543
rect 20162 11540 20168 11552
rect 19567 11512 20168 11540
rect 19567 11509 19579 11512
rect 19521 11503 19579 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 21266 11540 21272 11552
rect 21227 11512 21272 11540
rect 21266 11500 21272 11512
rect 21324 11540 21330 11552
rect 21913 11543 21971 11549
rect 21913 11540 21925 11543
rect 21324 11512 21925 11540
rect 21324 11500 21330 11512
rect 21913 11509 21925 11512
rect 21959 11509 21971 11543
rect 23842 11540 23848 11552
rect 23803 11512 23848 11540
rect 21913 11503 21971 11509
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 26418 11540 26424 11552
rect 26379 11512 26424 11540
rect 26418 11500 26424 11512
rect 26476 11540 26482 11552
rect 26988 11549 27016 11580
rect 27154 11568 27160 11620
rect 27212 11608 27218 11620
rect 27341 11611 27399 11617
rect 27341 11608 27353 11611
rect 27212 11580 27353 11608
rect 27212 11568 27218 11580
rect 27341 11577 27353 11580
rect 27387 11577 27399 11611
rect 27341 11571 27399 11577
rect 26605 11543 26663 11549
rect 26605 11540 26617 11543
rect 26476 11512 26617 11540
rect 26476 11500 26482 11512
rect 26605 11509 26617 11512
rect 26651 11509 26663 11543
rect 26605 11503 26663 11509
rect 26973 11543 27031 11549
rect 26973 11509 26985 11543
rect 27019 11509 27031 11543
rect 26973 11503 27031 11509
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 2130 11336 2136 11348
rect 2091 11308 2136 11336
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 2777 11339 2835 11345
rect 2777 11305 2789 11339
rect 2823 11336 2835 11339
rect 3142 11336 3148 11348
rect 2823 11308 3148 11336
rect 2823 11305 2835 11308
rect 2777 11299 2835 11305
rect 3142 11296 3148 11308
rect 3200 11296 3206 11348
rect 3510 11336 3516 11348
rect 3471 11308 3516 11336
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4617 11339 4675 11345
rect 4617 11336 4629 11339
rect 4120 11308 4629 11336
rect 4120 11296 4126 11308
rect 4617 11305 4629 11308
rect 4663 11305 4675 11339
rect 4617 11299 4675 11305
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6365 11339 6423 11345
rect 6365 11336 6377 11339
rect 5868 11308 6377 11336
rect 5868 11296 5874 11308
rect 6365 11305 6377 11308
rect 6411 11305 6423 11339
rect 6914 11336 6920 11348
rect 6875 11308 6920 11336
rect 6365 11299 6423 11305
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7006 11296 7012 11348
rect 7064 11336 7070 11348
rect 7285 11339 7343 11345
rect 7285 11336 7297 11339
rect 7064 11308 7297 11336
rect 7064 11296 7070 11308
rect 7285 11305 7297 11308
rect 7331 11305 7343 11339
rect 7285 11299 7343 11305
rect 7929 11339 7987 11345
rect 7929 11305 7941 11339
rect 7975 11336 7987 11339
rect 8018 11336 8024 11348
rect 7975 11308 8024 11336
rect 7975 11305 7987 11308
rect 7929 11299 7987 11305
rect 8018 11296 8024 11308
rect 8076 11296 8082 11348
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 11330 11296 11336 11348
rect 11388 11336 11394 11348
rect 11793 11339 11851 11345
rect 11793 11336 11805 11339
rect 11388 11308 11805 11336
rect 11388 11296 11394 11308
rect 11793 11305 11805 11308
rect 11839 11305 11851 11339
rect 11793 11299 11851 11305
rect 12161 11339 12219 11345
rect 12161 11305 12173 11339
rect 12207 11336 12219 11339
rect 12526 11336 12532 11348
rect 12207 11308 12532 11336
rect 12207 11305 12219 11308
rect 12161 11299 12219 11305
rect 12526 11296 12532 11308
rect 12584 11296 12590 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13265 11339 13323 11345
rect 13265 11336 13277 11339
rect 13044 11308 13277 11336
rect 13044 11296 13050 11308
rect 13265 11305 13277 11308
rect 13311 11305 13323 11339
rect 13265 11299 13323 11305
rect 14550 11296 14556 11348
rect 14608 11336 14614 11348
rect 15194 11336 15200 11348
rect 14608 11308 15200 11336
rect 14608 11296 14614 11308
rect 15194 11296 15200 11308
rect 15252 11336 15258 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 15252 11308 16129 11336
rect 15252 11296 15258 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16577 11339 16635 11345
rect 16577 11336 16589 11339
rect 16540 11308 16589 11336
rect 16540 11296 16546 11308
rect 16577 11305 16589 11308
rect 16623 11305 16635 11339
rect 16577 11299 16635 11305
rect 17221 11339 17279 11345
rect 17221 11305 17233 11339
rect 17267 11336 17279 11339
rect 17402 11336 17408 11348
rect 17267 11308 17408 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 17402 11296 17408 11308
rect 17460 11296 17466 11348
rect 18138 11336 18144 11348
rect 18099 11308 18144 11336
rect 18138 11296 18144 11308
rect 18196 11296 18202 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18472 11308 18705 11336
rect 18472 11296 18478 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 18693 11299 18751 11305
rect 19245 11339 19303 11345
rect 19245 11305 19257 11339
rect 19291 11336 19303 11339
rect 20254 11336 20260 11348
rect 19291 11308 20260 11336
rect 19291 11305 19303 11308
rect 19245 11299 19303 11305
rect 20254 11296 20260 11308
rect 20312 11296 20318 11348
rect 20714 11296 20720 11348
rect 20772 11336 20778 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20772 11308 20913 11336
rect 20772 11296 20778 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 23658 11336 23664 11348
rect 23619 11308 23664 11336
rect 20901 11299 20959 11305
rect 23658 11296 23664 11308
rect 23716 11296 23722 11348
rect 24857 11339 24915 11345
rect 24857 11305 24869 11339
rect 24903 11336 24915 11339
rect 24946 11336 24952 11348
rect 24903 11308 24952 11336
rect 24903 11305 24915 11308
rect 24857 11299 24915 11305
rect 24946 11296 24952 11308
rect 25004 11296 25010 11348
rect 25225 11339 25283 11345
rect 25225 11305 25237 11339
rect 25271 11336 25283 11339
rect 25866 11336 25872 11348
rect 25271 11308 25872 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 25866 11296 25872 11308
rect 25924 11296 25930 11348
rect 26510 11336 26516 11348
rect 26471 11308 26516 11336
rect 26510 11296 26516 11308
rect 26568 11296 26574 11348
rect 26878 11336 26884 11348
rect 26839 11308 26884 11336
rect 26878 11296 26884 11308
rect 26936 11296 26942 11348
rect 26973 11339 27031 11345
rect 26973 11305 26985 11339
rect 27019 11336 27031 11339
rect 27338 11336 27344 11348
rect 27019 11308 27344 11336
rect 27019 11305 27031 11308
rect 26973 11299 27031 11305
rect 27338 11296 27344 11308
rect 27396 11296 27402 11348
rect 27522 11336 27528 11348
rect 27483 11308 27528 11336
rect 27522 11296 27528 11308
rect 27580 11296 27586 11348
rect 4341 11271 4399 11277
rect 4341 11237 4353 11271
rect 4387 11268 4399 11271
rect 5828 11268 5856 11296
rect 4387 11240 5856 11268
rect 10137 11271 10195 11277
rect 4387 11237 4399 11240
rect 4341 11231 4399 11237
rect 10137 11237 10149 11271
rect 10183 11268 10195 11271
rect 10226 11268 10232 11280
rect 10183 11240 10232 11268
rect 10183 11237 10195 11240
rect 10137 11231 10195 11237
rect 10226 11228 10232 11240
rect 10284 11268 10290 11280
rect 14918 11268 14924 11280
rect 10284 11240 10916 11268
rect 14879 11240 14924 11268
rect 10284 11228 10290 11240
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 3050 11200 3056 11212
rect 2915 11172 3056 11200
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3050 11160 3056 11172
rect 3108 11200 3114 11212
rect 4062 11200 4068 11212
rect 3108 11172 4068 11200
rect 3108 11160 3114 11172
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 5258 11209 5264 11212
rect 5252 11200 5264 11209
rect 5219 11172 5264 11200
rect 5252 11163 5264 11172
rect 5258 11160 5264 11163
rect 5316 11160 5322 11212
rect 7837 11203 7895 11209
rect 7837 11169 7849 11203
rect 7883 11200 7895 11203
rect 8202 11200 8208 11212
rect 7883 11172 8208 11200
rect 7883 11169 7895 11172
rect 7837 11163 7895 11169
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 10594 11200 10600 11212
rect 10555 11172 10600 11200
rect 10594 11160 10600 11172
rect 10652 11160 10658 11212
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11092 1458 11144
rect 2314 11092 2320 11144
rect 2372 11132 2378 11144
rect 2958 11132 2964 11144
rect 2372 11104 2820 11132
rect 2871 11104 2964 11132
rect 2372 11092 2378 11104
rect 2409 11067 2467 11073
rect 2409 11033 2421 11067
rect 2455 11064 2467 11067
rect 2682 11064 2688 11076
rect 2455 11036 2688 11064
rect 2455 11033 2467 11036
rect 2409 11027 2467 11033
rect 2682 11024 2688 11036
rect 2740 11024 2746 11076
rect 2792 10996 2820 11104
rect 2958 11092 2964 11104
rect 3016 11132 3022 11144
rect 3510 11132 3516 11144
rect 3016 11104 3516 11132
rect 3016 11092 3022 11104
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4985 11135 5043 11141
rect 4985 11101 4997 11135
rect 5031 11101 5043 11135
rect 4985 11095 5043 11101
rect 8113 11135 8171 11141
rect 8113 11101 8125 11135
rect 8159 11132 8171 11135
rect 8294 11132 8300 11144
rect 8159 11104 8300 11132
rect 8159 11101 8171 11104
rect 8113 11095 8171 11101
rect 5000 11064 5028 11095
rect 8294 11092 8300 11104
rect 8352 11132 8358 11144
rect 8754 11132 8760 11144
rect 8352 11104 8760 11132
rect 8352 11092 8358 11104
rect 8754 11092 8760 11104
rect 8812 11092 8818 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10686 11132 10692 11144
rect 10192 11104 10692 11132
rect 10192 11092 10198 11104
rect 10686 11092 10692 11104
rect 10744 11092 10750 11144
rect 10888 11141 10916 11240
rect 14918 11228 14924 11240
rect 14976 11228 14982 11280
rect 15654 11268 15660 11280
rect 15615 11240 15660 11268
rect 15654 11228 15660 11240
rect 15712 11228 15718 11280
rect 17770 11228 17776 11280
rect 17828 11268 17834 11280
rect 18049 11271 18107 11277
rect 18049 11268 18061 11271
rect 17828 11240 18061 11268
rect 17828 11228 17834 11240
rect 18049 11237 18061 11240
rect 18095 11268 18107 11271
rect 18506 11268 18512 11280
rect 18095 11240 18512 11268
rect 18095 11237 18107 11240
rect 18049 11231 18107 11237
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 19886 11228 19892 11280
rect 19944 11268 19950 11280
rect 22094 11268 22100 11280
rect 19944 11240 22100 11268
rect 19944 11228 19950 11240
rect 22094 11228 22100 11240
rect 22152 11228 22158 11280
rect 23474 11228 23480 11280
rect 23532 11268 23538 11280
rect 23750 11268 23756 11280
rect 23532 11240 23756 11268
rect 23532 11228 23538 11240
rect 23750 11228 23756 11240
rect 23808 11268 23814 11280
rect 24029 11271 24087 11277
rect 24029 11268 24041 11271
rect 23808 11240 24041 11268
rect 23808 11228 23814 11240
rect 24029 11237 24041 11240
rect 24075 11237 24087 11271
rect 26896 11268 26924 11296
rect 27614 11268 27620 11280
rect 26896 11240 27620 11268
rect 24029 11231 24087 11237
rect 27614 11228 27620 11240
rect 27672 11228 27678 11280
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 11940 11172 12388 11200
rect 11940 11160 11946 11172
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11698 11132 11704 11144
rect 10919 11104 11704 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12360 11141 12388 11172
rect 15562 11160 15568 11212
rect 15620 11200 15626 11212
rect 16298 11200 16304 11212
rect 15620 11172 16304 11200
rect 15620 11160 15626 11172
rect 16298 11160 16304 11172
rect 16356 11200 16362 11212
rect 16485 11203 16543 11209
rect 16485 11200 16497 11203
rect 16356 11172 16497 11200
rect 16356 11160 16362 11172
rect 16485 11169 16497 11172
rect 16531 11169 16543 11203
rect 16485 11163 16543 11169
rect 19242 11160 19248 11212
rect 19300 11200 19306 11212
rect 19613 11203 19671 11209
rect 19613 11200 19625 11203
rect 19300 11172 19625 11200
rect 19300 11160 19306 11172
rect 19613 11169 19625 11172
rect 19659 11169 19671 11203
rect 19613 11163 19671 11169
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 20806 11200 20812 11212
rect 20763 11172 20812 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 20806 11160 20812 11172
rect 20864 11200 20870 11212
rect 21269 11203 21327 11209
rect 21269 11200 21281 11203
rect 20864 11172 21281 11200
rect 20864 11160 20870 11172
rect 21269 11169 21281 11172
rect 21315 11169 21327 11203
rect 21269 11163 21327 11169
rect 21361 11203 21419 11209
rect 21361 11169 21373 11203
rect 21407 11200 21419 11203
rect 21910 11200 21916 11212
rect 21407 11172 21916 11200
rect 21407 11169 21419 11172
rect 21361 11163 21419 11169
rect 21910 11160 21916 11172
rect 21968 11160 21974 11212
rect 22554 11200 22560 11212
rect 22515 11172 22560 11200
rect 22554 11160 22560 11172
rect 22612 11160 22618 11212
rect 25317 11203 25375 11209
rect 25317 11169 25329 11203
rect 25363 11200 25375 11203
rect 25590 11200 25596 11212
rect 25363 11172 25596 11200
rect 25363 11169 25375 11172
rect 25317 11163 25375 11169
rect 25590 11160 25596 11172
rect 25648 11160 25654 11212
rect 12253 11135 12311 11141
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 3712 11036 5028 11064
rect 10229 11067 10287 11073
rect 3712 10996 3740 11036
rect 3878 10996 3884 11008
rect 2792 10968 3740 10996
rect 3839 10968 3884 10996
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 3970 10956 3976 11008
rect 4028 10996 4034 11008
rect 4080 10996 4108 11036
rect 10229 11033 10241 11067
rect 10275 11064 10287 11067
rect 12158 11064 12164 11076
rect 10275 11036 12164 11064
rect 10275 11033 10287 11036
rect 10229 11027 10287 11033
rect 12158 11024 12164 11036
rect 12216 11064 12222 11076
rect 12268 11064 12296 11095
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 18322 11132 18328 11144
rect 16724 11104 16769 11132
rect 18283 11104 18328 11132
rect 16724 11092 16730 11104
rect 18322 11092 18328 11104
rect 18380 11092 18386 11144
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 19797 11135 19855 11141
rect 19797 11101 19809 11135
rect 19843 11132 19855 11135
rect 20438 11132 20444 11144
rect 19843 11104 20444 11132
rect 19843 11101 19855 11104
rect 19797 11095 19855 11101
rect 12216 11036 12296 11064
rect 16025 11067 16083 11073
rect 12216 11024 12222 11036
rect 16025 11033 16037 11067
rect 16071 11064 16083 11067
rect 16482 11064 16488 11076
rect 16071 11036 16488 11064
rect 16071 11033 16083 11036
rect 16025 11027 16083 11033
rect 16482 11024 16488 11036
rect 16540 11024 16546 11076
rect 17681 11067 17739 11073
rect 17681 11033 17693 11067
rect 17727 11064 17739 11067
rect 19061 11067 19119 11073
rect 19061 11064 19073 11067
rect 17727 11036 19073 11064
rect 17727 11033 17739 11036
rect 17681 11027 17739 11033
rect 19061 11033 19073 11036
rect 19107 11064 19119 11067
rect 19720 11064 19748 11095
rect 19107 11036 19748 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 4028 10968 4108 10996
rect 4028 10956 4034 10968
rect 4982 10956 4988 11008
rect 5040 10996 5046 11008
rect 7006 10996 7012 11008
rect 5040 10968 7012 10996
rect 5040 10956 5046 10968
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 7469 10999 7527 11005
rect 7469 10965 7481 10999
rect 7515 10996 7527 10999
rect 7650 10996 7656 11008
rect 7515 10968 7656 10996
rect 7515 10965 7527 10968
rect 7469 10959 7527 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 18966 10956 18972 11008
rect 19024 10996 19030 11008
rect 19812 10996 19840 11095
rect 20438 11092 20444 11104
rect 20496 11132 20502 11144
rect 21450 11132 21456 11144
rect 20496 11104 21456 11132
rect 20496 11092 20502 11104
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 23474 11092 23480 11144
rect 23532 11132 23538 11144
rect 23842 11132 23848 11144
rect 23532 11104 23848 11132
rect 23532 11092 23538 11104
rect 23842 11092 23848 11104
rect 23900 11132 23906 11144
rect 24121 11135 24179 11141
rect 24121 11132 24133 11135
rect 23900 11104 24133 11132
rect 23900 11092 23906 11104
rect 24121 11101 24133 11104
rect 24167 11101 24179 11135
rect 24302 11132 24308 11144
rect 24263 11104 24308 11132
rect 24121 11095 24179 11101
rect 24302 11092 24308 11104
rect 24360 11092 24366 11144
rect 27065 11135 27123 11141
rect 27065 11132 27077 11135
rect 26712 11104 27077 11132
rect 22738 11064 22744 11076
rect 22699 11036 22744 11064
rect 22738 11024 22744 11036
rect 22796 11024 22802 11076
rect 25501 11067 25559 11073
rect 25501 11033 25513 11067
rect 25547 11064 25559 11067
rect 25682 11064 25688 11076
rect 25547 11036 25688 11064
rect 25547 11033 25559 11036
rect 25501 11027 25559 11033
rect 25682 11024 25688 11036
rect 25740 11024 25746 11076
rect 26712 11008 26740 11104
rect 27065 11101 27077 11104
rect 27111 11132 27123 11135
rect 27246 11132 27252 11144
rect 27111 11104 27252 11132
rect 27111 11101 27123 11104
rect 27065 11095 27123 11101
rect 27246 11092 27252 11104
rect 27304 11092 27310 11144
rect 19024 10968 19840 10996
rect 19024 10956 19030 10968
rect 21726 10956 21732 11008
rect 21784 10996 21790 11008
rect 21913 10999 21971 11005
rect 21913 10996 21925 10999
rect 21784 10968 21925 10996
rect 21784 10956 21790 10968
rect 21913 10965 21925 10968
rect 21959 10965 21971 10999
rect 21913 10959 21971 10965
rect 23290 10956 23296 11008
rect 23348 10996 23354 11008
rect 23477 10999 23535 11005
rect 23477 10996 23489 10999
rect 23348 10968 23489 10996
rect 23348 10956 23354 10968
rect 23477 10965 23489 10968
rect 23523 10996 23535 10999
rect 23658 10996 23664 11008
rect 23523 10968 23664 10996
rect 23523 10965 23535 10968
rect 23477 10959 23535 10965
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 26237 10999 26295 11005
rect 26237 10965 26249 10999
rect 26283 10996 26295 10999
rect 26694 10996 26700 11008
rect 26283 10968 26700 10996
rect 26283 10965 26295 10968
rect 26237 10959 26295 10965
rect 26694 10956 26700 10968
rect 26752 10956 26758 11008
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 3142 10792 3148 10804
rect 3103 10764 3148 10792
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 3602 10792 3608 10804
rect 3563 10764 3608 10792
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4212 10764 5181 10792
rect 4212 10752 4218 10764
rect 5169 10761 5181 10764
rect 5215 10761 5227 10795
rect 5169 10755 5227 10761
rect 7285 10795 7343 10801
rect 7285 10761 7297 10795
rect 7331 10792 7343 10795
rect 7466 10792 7472 10804
rect 7331 10764 7472 10792
rect 7331 10761 7343 10764
rect 7285 10755 7343 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 8665 10795 8723 10801
rect 8665 10792 8677 10795
rect 8260 10764 8677 10792
rect 8260 10752 8266 10764
rect 8665 10761 8677 10764
rect 8711 10761 8723 10795
rect 10134 10792 10140 10804
rect 10095 10764 10140 10792
rect 8665 10755 8723 10761
rect 10134 10752 10140 10764
rect 10192 10752 10198 10804
rect 10318 10792 10324 10804
rect 10279 10764 10324 10792
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11425 10795 11483 10801
rect 11425 10761 11437 10795
rect 11471 10792 11483 10795
rect 11698 10792 11704 10804
rect 11471 10764 11704 10792
rect 11471 10761 11483 10764
rect 11425 10755 11483 10761
rect 3786 10684 3792 10736
rect 3844 10724 3850 10736
rect 4985 10727 5043 10733
rect 4985 10724 4997 10727
rect 3844 10696 4997 10724
rect 3844 10684 3850 10696
rect 4985 10693 4997 10696
rect 5031 10724 5043 10727
rect 8294 10724 8300 10736
rect 5031 10696 5672 10724
rect 8255 10696 8300 10724
rect 5031 10693 5043 10696
rect 4985 10687 5043 10693
rect 5644 10668 5672 10696
rect 8294 10684 8300 10696
rect 8352 10684 8358 10736
rect 1578 10616 1584 10668
rect 1636 10656 1642 10668
rect 2130 10656 2136 10668
rect 1636 10628 2136 10656
rect 1636 10616 1642 10628
rect 2130 10616 2136 10628
rect 2188 10656 2194 10668
rect 2501 10659 2559 10665
rect 2501 10656 2513 10659
rect 2188 10628 2513 10656
rect 2188 10616 2194 10628
rect 2501 10625 2513 10628
rect 2547 10625 2559 10659
rect 2501 10619 2559 10625
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2958 10656 2964 10668
rect 2731 10628 2964 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 3559 10628 4261 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 4249 10625 4261 10628
rect 4295 10656 4307 10659
rect 5258 10656 5264 10668
rect 4295 10628 5264 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5626 10656 5632 10668
rect 5539 10628 5632 10656
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5810 10616 5816 10628
rect 5868 10616 5874 10668
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 7837 10659 7895 10665
rect 7837 10656 7849 10659
rect 7239 10628 7849 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7837 10625 7849 10628
rect 7883 10656 7895 10659
rect 8110 10656 8116 10668
rect 7883 10628 8116 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 10965 10659 11023 10665
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11330 10656 11336 10668
rect 11011 10628 11336 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11330 10616 11336 10628
rect 11388 10656 11394 10668
rect 11440 10656 11468 10755
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 11882 10792 11888 10804
rect 11843 10764 11888 10792
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12158 10792 12164 10804
rect 12119 10764 12164 10792
rect 12158 10752 12164 10764
rect 12216 10752 12222 10804
rect 12526 10752 12532 10804
rect 12584 10792 12590 10804
rect 12621 10795 12679 10801
rect 12621 10792 12633 10795
rect 12584 10764 12633 10792
rect 12584 10752 12590 10764
rect 12621 10761 12633 10764
rect 12667 10761 12679 10795
rect 12621 10755 12679 10761
rect 15286 10752 15292 10804
rect 15344 10792 15350 10804
rect 16393 10795 16451 10801
rect 16393 10792 16405 10795
rect 15344 10764 16405 10792
rect 15344 10752 15350 10764
rect 16393 10761 16405 10764
rect 16439 10761 16451 10795
rect 17770 10792 17776 10804
rect 17731 10764 17776 10792
rect 16393 10755 16451 10761
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 18966 10792 18972 10804
rect 18927 10764 18972 10792
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 19337 10795 19395 10801
rect 19337 10761 19349 10795
rect 19383 10792 19395 10795
rect 20346 10792 20352 10804
rect 19383 10764 20352 10792
rect 19383 10761 19395 10764
rect 19337 10755 19395 10761
rect 15197 10727 15255 10733
rect 15197 10693 15209 10727
rect 15243 10724 15255 10727
rect 15378 10724 15384 10736
rect 15243 10696 15384 10724
rect 15243 10693 15255 10696
rect 15197 10687 15255 10693
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 15562 10724 15568 10736
rect 15523 10696 15568 10724
rect 15562 10684 15568 10696
rect 15620 10684 15626 10736
rect 11388 10628 11468 10656
rect 11388 10616 11394 10628
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16632 10628 17049 10656
rect 16632 10616 16638 10628
rect 17037 10625 17049 10628
rect 17083 10656 17095 10659
rect 17862 10656 17868 10668
rect 17083 10628 17868 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 19334 10616 19340 10668
rect 19392 10656 19398 10668
rect 19444 10665 19472 10764
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 21450 10792 21456 10804
rect 21411 10764 21456 10792
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 22554 10752 22560 10804
rect 22612 10792 22618 10804
rect 22925 10795 22983 10801
rect 22925 10792 22937 10795
rect 22612 10764 22937 10792
rect 22612 10752 22618 10764
rect 22925 10761 22937 10764
rect 22971 10792 22983 10795
rect 22971 10764 24624 10792
rect 22971 10761 22983 10764
rect 22925 10755 22983 10761
rect 24596 10724 24624 10764
rect 24762 10752 24768 10804
rect 24820 10792 24826 10804
rect 26145 10795 26203 10801
rect 26145 10792 26157 10795
rect 24820 10764 26157 10792
rect 24820 10752 24826 10764
rect 26145 10761 26157 10764
rect 26191 10761 26203 10795
rect 26145 10755 26203 10761
rect 27249 10795 27307 10801
rect 27249 10761 27261 10795
rect 27295 10792 27307 10795
rect 27338 10792 27344 10804
rect 27295 10764 27344 10792
rect 27295 10761 27307 10764
rect 27249 10755 27307 10761
rect 27338 10752 27344 10764
rect 27396 10752 27402 10804
rect 27614 10792 27620 10804
rect 27575 10764 27620 10792
rect 27614 10752 27620 10764
rect 27672 10752 27678 10804
rect 24596 10696 24900 10724
rect 19429 10659 19487 10665
rect 19429 10656 19441 10659
rect 19392 10628 19441 10656
rect 19392 10616 19398 10628
rect 19429 10625 19441 10628
rect 19475 10625 19487 10659
rect 19429 10619 19487 10625
rect 21726 10616 21732 10668
rect 21784 10656 21790 10668
rect 22465 10659 22523 10665
rect 22465 10656 22477 10659
rect 21784 10628 22477 10656
rect 21784 10616 21790 10628
rect 22465 10625 22477 10628
rect 22511 10625 22523 10659
rect 24872 10656 24900 10696
rect 24946 10684 24952 10736
rect 25004 10724 25010 10736
rect 25041 10727 25099 10733
rect 25041 10724 25053 10727
rect 25004 10696 25053 10724
rect 25004 10684 25010 10696
rect 25041 10693 25053 10696
rect 25087 10724 25099 10727
rect 25222 10724 25228 10736
rect 25087 10696 25228 10724
rect 25087 10693 25099 10696
rect 25041 10687 25099 10693
rect 25222 10684 25228 10696
rect 25280 10684 25286 10736
rect 25961 10659 26019 10665
rect 25961 10656 25973 10659
rect 24872 10628 25973 10656
rect 22465 10619 22523 10625
rect 25961 10625 25973 10628
rect 26007 10656 26019 10659
rect 26694 10656 26700 10668
rect 26007 10628 26556 10656
rect 26655 10628 26700 10656
rect 26007 10625 26019 10628
rect 25961 10619 26019 10625
rect 1949 10591 2007 10597
rect 1949 10557 1961 10591
rect 1995 10588 2007 10591
rect 2409 10591 2467 10597
rect 2409 10588 2421 10591
rect 1995 10560 2421 10588
rect 1995 10557 2007 10560
rect 1949 10551 2007 10557
rect 2409 10557 2421 10560
rect 2455 10588 2467 10591
rect 2774 10588 2780 10600
rect 2455 10560 2780 10588
rect 2455 10557 2467 10560
rect 2409 10551 2467 10557
rect 2774 10548 2780 10560
rect 2832 10548 2838 10600
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 3973 10591 4031 10597
rect 3973 10588 3985 10591
rect 3936 10560 3985 10588
rect 3936 10548 3942 10560
rect 3973 10557 3985 10560
rect 4019 10557 4031 10591
rect 7742 10588 7748 10600
rect 7703 10560 7748 10588
rect 3973 10551 4031 10557
rect 7742 10548 7748 10560
rect 7800 10548 7806 10600
rect 8849 10591 8907 10597
rect 8849 10557 8861 10591
rect 8895 10588 8907 10591
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 8895 10560 9413 10588
rect 8895 10557 8907 10560
rect 8849 10551 8907 10557
rect 9401 10557 9413 10560
rect 9447 10588 9459 10591
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9447 10560 9781 10588
rect 9447 10557 9459 10560
rect 9401 10551 9459 10557
rect 9769 10557 9781 10560
rect 9815 10588 9827 10591
rect 10594 10588 10600 10600
rect 9815 10560 10600 10588
rect 9815 10557 9827 10560
rect 9769 10551 9827 10557
rect 4246 10480 4252 10532
rect 4304 10520 4310 10532
rect 4709 10523 4767 10529
rect 4709 10520 4721 10523
rect 4304 10492 4721 10520
rect 4304 10480 4310 10492
rect 4709 10489 4721 10492
rect 4755 10520 4767 10523
rect 4755 10492 5580 10520
rect 4755 10489 4767 10492
rect 4709 10483 4767 10489
rect 5552 10464 5580 10492
rect 6914 10480 6920 10532
rect 6972 10520 6978 10532
rect 8864 10520 8892 10551
rect 10594 10548 10600 10560
rect 10652 10548 10658 10600
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10588 10747 10591
rect 10778 10588 10784 10600
rect 10735 10560 10784 10588
rect 10735 10557 10747 10560
rect 10689 10551 10747 10557
rect 10778 10548 10784 10560
rect 10836 10548 10842 10600
rect 16301 10591 16359 10597
rect 16301 10557 16313 10591
rect 16347 10588 16359 10591
rect 16850 10588 16856 10600
rect 16347 10560 16856 10588
rect 16347 10557 16359 10560
rect 16301 10551 16359 10557
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 21818 10588 21824 10600
rect 21731 10560 21824 10588
rect 21818 10548 21824 10560
rect 21876 10588 21882 10600
rect 22281 10591 22339 10597
rect 22281 10588 22293 10591
rect 21876 10560 22293 10588
rect 21876 10548 21882 10560
rect 22281 10557 22293 10560
rect 22327 10557 22339 10591
rect 22281 10551 22339 10557
rect 22370 10548 22376 10600
rect 22428 10588 22434 10600
rect 23566 10588 23572 10600
rect 22428 10560 23572 10588
rect 22428 10548 22434 10560
rect 23566 10548 23572 10560
rect 23624 10548 23630 10600
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 23928 10591 23986 10597
rect 23716 10560 23809 10588
rect 23716 10548 23722 10560
rect 23928 10557 23940 10591
rect 23974 10588 23986 10591
rect 24302 10588 24308 10600
rect 23974 10560 24308 10588
rect 23974 10557 23986 10560
rect 23928 10551 23986 10557
rect 24302 10548 24308 10560
rect 24360 10548 24366 10600
rect 25590 10588 25596 10600
rect 25551 10560 25596 10588
rect 25590 10548 25596 10560
rect 25648 10548 25654 10600
rect 26528 10597 26556 10628
rect 26694 10616 26700 10628
rect 26752 10616 26758 10668
rect 26513 10591 26571 10597
rect 26513 10557 26525 10591
rect 26559 10557 26571 10591
rect 26513 10551 26571 10557
rect 6972 10492 8892 10520
rect 15933 10523 15991 10529
rect 6972 10480 6978 10492
rect 15933 10489 15945 10523
rect 15979 10520 15991 10523
rect 16758 10520 16764 10532
rect 15979 10492 16764 10520
rect 15979 10489 15991 10492
rect 15933 10483 15991 10489
rect 16758 10480 16764 10492
rect 16816 10480 16822 10532
rect 19696 10523 19754 10529
rect 19696 10489 19708 10523
rect 19742 10520 19754 10523
rect 20346 10520 20352 10532
rect 19742 10492 20352 10520
rect 19742 10489 19754 10492
rect 19696 10483 19754 10489
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 23477 10523 23535 10529
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23676 10520 23704 10548
rect 25774 10520 25780 10532
rect 23523 10492 25780 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 25774 10480 25780 10492
rect 25832 10480 25838 10532
rect 2038 10452 2044 10464
rect 1999 10424 2044 10452
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 4062 10452 4068 10464
rect 4023 10424 4068 10452
rect 4062 10412 4068 10424
rect 4120 10412 4126 10464
rect 5534 10452 5540 10464
rect 5495 10424 5540 10452
rect 5534 10412 5540 10424
rect 5592 10412 5598 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6362 10452 6368 10464
rect 6319 10424 6368 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6362 10412 6368 10424
rect 6420 10412 6426 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 7650 10452 7656 10464
rect 7611 10424 7656 10452
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 9030 10452 9036 10464
rect 8991 10424 9036 10452
rect 9030 10412 9036 10424
rect 9088 10412 9094 10464
rect 10318 10412 10324 10464
rect 10376 10452 10382 10464
rect 10781 10455 10839 10461
rect 10781 10452 10793 10455
rect 10376 10424 10793 10452
rect 10376 10412 10382 10424
rect 10781 10421 10793 10424
rect 10827 10421 10839 10455
rect 18322 10452 18328 10464
rect 18283 10424 18328 10452
rect 10781 10415 10839 10421
rect 18322 10412 18328 10424
rect 18380 10412 18386 10464
rect 20622 10412 20628 10464
rect 20680 10452 20686 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20680 10424 20821 10452
rect 20680 10412 20686 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 21910 10452 21916 10464
rect 21871 10424 21916 10452
rect 20809 10415 20867 10421
rect 21910 10412 21916 10424
rect 21968 10412 21974 10464
rect 26510 10412 26516 10464
rect 26568 10452 26574 10464
rect 26605 10455 26663 10461
rect 26605 10452 26617 10455
rect 26568 10424 26617 10452
rect 26568 10412 26574 10424
rect 26605 10421 26617 10424
rect 26651 10421 26663 10455
rect 26605 10415 26663 10421
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 2406 10248 2412 10260
rect 1452 10220 2412 10248
rect 1452 10208 1458 10220
rect 2406 10208 2412 10220
rect 2464 10208 2470 10260
rect 2498 10208 2504 10260
rect 2556 10248 2562 10260
rect 2556 10220 2601 10248
rect 2556 10208 2562 10220
rect 2958 10208 2964 10260
rect 3016 10248 3022 10260
rect 3053 10251 3111 10257
rect 3053 10248 3065 10251
rect 3016 10220 3065 10248
rect 3016 10208 3022 10220
rect 3053 10217 3065 10220
rect 3099 10217 3111 10251
rect 3053 10211 3111 10217
rect 5258 10208 5264 10260
rect 5316 10248 5322 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5316 10220 5457 10248
rect 5316 10208 5322 10220
rect 5445 10217 5457 10220
rect 5491 10248 5503 10251
rect 6546 10248 6552 10260
rect 5491 10220 6552 10248
rect 5491 10217 5503 10220
rect 5445 10211 5503 10217
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 7006 10248 7012 10260
rect 6967 10220 7012 10248
rect 7006 10208 7012 10220
rect 7064 10208 7070 10260
rect 8018 10248 8024 10260
rect 7979 10220 8024 10248
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 10318 10248 10324 10260
rect 10279 10220 10324 10248
rect 10318 10208 10324 10220
rect 10376 10208 10382 10260
rect 11149 10251 11207 10257
rect 11149 10217 11161 10251
rect 11195 10248 11207 10251
rect 11330 10248 11336 10260
rect 11195 10220 11336 10248
rect 11195 10217 11207 10220
rect 11149 10211 11207 10217
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 16209 10251 16267 10257
rect 16209 10217 16221 10251
rect 16255 10248 16267 10251
rect 16390 10248 16396 10260
rect 16255 10220 16396 10248
rect 16255 10217 16267 10220
rect 16209 10211 16267 10217
rect 16390 10208 16396 10220
rect 16448 10208 16454 10260
rect 17678 10248 17684 10260
rect 17639 10220 17684 10248
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 18785 10251 18843 10257
rect 18785 10217 18797 10251
rect 18831 10248 18843 10251
rect 19242 10248 19248 10260
rect 18831 10220 19248 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 19518 10208 19524 10260
rect 19576 10248 19582 10260
rect 19705 10251 19763 10257
rect 19705 10248 19717 10251
rect 19576 10220 19717 10248
rect 19576 10208 19582 10220
rect 19705 10217 19717 10220
rect 19751 10217 19763 10251
rect 20346 10248 20352 10260
rect 20307 10220 20352 10248
rect 19705 10211 19763 10217
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20864 10220 20913 10248
rect 20864 10208 20870 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 21358 10248 21364 10260
rect 21319 10220 21364 10248
rect 20901 10211 20959 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 23474 10248 23480 10260
rect 23435 10220 23480 10248
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 23569 10251 23627 10257
rect 23569 10217 23581 10251
rect 23615 10248 23627 10251
rect 24118 10248 24124 10260
rect 23615 10220 24124 10248
rect 23615 10217 23627 10220
rect 23569 10211 23627 10217
rect 24118 10208 24124 10220
rect 24176 10208 24182 10260
rect 24302 10208 24308 10260
rect 24360 10248 24366 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 24360 10220 24409 10248
rect 24360 10208 24366 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 24578 10248 24584 10260
rect 24539 10220 24584 10248
rect 24397 10211 24455 10217
rect 24578 10208 24584 10220
rect 24636 10208 24642 10260
rect 25041 10251 25099 10257
rect 25041 10217 25053 10251
rect 25087 10248 25099 10251
rect 25222 10248 25228 10260
rect 25087 10220 25228 10248
rect 25087 10217 25099 10220
rect 25041 10211 25099 10217
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 4856 10152 7052 10180
rect 4856 10140 4862 10152
rect 4332 10115 4390 10121
rect 4332 10081 4344 10115
rect 4378 10112 4390 10115
rect 4706 10112 4712 10124
rect 4378 10084 4712 10112
rect 4378 10081 4390 10084
rect 4332 10075 4390 10081
rect 4706 10072 4712 10084
rect 4764 10072 4770 10124
rect 6914 10112 6920 10124
rect 6875 10084 6920 10112
rect 6914 10072 6920 10084
rect 6972 10072 6978 10124
rect 7024 10112 7052 10152
rect 7650 10140 7656 10192
rect 7708 10180 7714 10192
rect 9033 10183 9091 10189
rect 9033 10180 9045 10183
rect 7708 10152 9045 10180
rect 7708 10140 7714 10152
rect 9033 10149 9045 10152
rect 9079 10149 9091 10183
rect 9033 10143 9091 10149
rect 20717 10183 20775 10189
rect 20717 10149 20729 10183
rect 20763 10180 20775 10183
rect 21910 10180 21916 10192
rect 20763 10152 21916 10180
rect 20763 10149 20775 10152
rect 20717 10143 20775 10149
rect 21910 10140 21916 10152
rect 21968 10140 21974 10192
rect 23109 10183 23167 10189
rect 23109 10149 23121 10183
rect 23155 10180 23167 10183
rect 23382 10180 23388 10192
rect 23155 10152 23388 10180
rect 23155 10149 23167 10152
rect 23109 10143 23167 10149
rect 23382 10140 23388 10152
rect 23440 10140 23446 10192
rect 24029 10183 24087 10189
rect 24029 10149 24041 10183
rect 24075 10180 24087 10183
rect 24320 10180 24348 10208
rect 25056 10180 25084 10211
rect 25222 10208 25228 10220
rect 25280 10248 25286 10260
rect 25866 10248 25872 10260
rect 25280 10220 25872 10248
rect 25280 10208 25286 10220
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 24075 10152 24348 10180
rect 24412 10152 25084 10180
rect 24075 10149 24087 10152
rect 24029 10143 24087 10149
rect 8110 10112 8116 10124
rect 7024 10084 8116 10112
rect 8110 10072 8116 10084
rect 8168 10112 8174 10124
rect 9306 10112 9312 10124
rect 8168 10084 9312 10112
rect 8168 10072 8174 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10778 10112 10784 10124
rect 10739 10084 10784 10112
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 16850 10112 16856 10124
rect 16811 10084 16856 10112
rect 16850 10072 16856 10084
rect 16908 10072 16914 10124
rect 19426 10072 19432 10124
rect 19484 10112 19490 10124
rect 19610 10112 19616 10124
rect 19484 10084 19616 10112
rect 19484 10072 19490 10084
rect 19610 10072 19616 10084
rect 19668 10072 19674 10124
rect 20806 10072 20812 10124
rect 20864 10112 20870 10124
rect 21266 10112 21272 10124
rect 20864 10084 21272 10112
rect 20864 10072 20870 10084
rect 21266 10072 21272 10084
rect 21324 10072 21330 10124
rect 21634 10072 21640 10124
rect 21692 10112 21698 10124
rect 24412 10112 24440 10152
rect 21692 10084 24440 10112
rect 24949 10115 25007 10121
rect 21692 10072 21698 10084
rect 24949 10081 24961 10115
rect 24995 10112 25007 10115
rect 26513 10115 26571 10121
rect 24995 10084 25084 10112
rect 24995 10081 25007 10084
rect 24949 10075 25007 10081
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2958 10044 2964 10056
rect 2639 10016 2964 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 1949 9979 2007 9985
rect 1949 9945 1961 9979
rect 1995 9976 2007 9979
rect 2608 9976 2636 10007
rect 2958 10004 2964 10016
rect 3016 10004 3022 10056
rect 3970 10004 3976 10056
rect 4028 10044 4034 10056
rect 4065 10047 4123 10053
rect 4065 10044 4077 10047
rect 4028 10016 4077 10044
rect 4028 10004 4034 10016
rect 4065 10013 4077 10016
rect 4111 10013 4123 10047
rect 4065 10007 4123 10013
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 1995 9948 2636 9976
rect 1995 9945 2007 9948
rect 1949 9939 2007 9945
rect 5810 9936 5816 9988
rect 5868 9976 5874 9988
rect 6089 9979 6147 9985
rect 6089 9976 6101 9979
rect 5868 9948 6101 9976
rect 5868 9936 5874 9948
rect 6089 9945 6101 9948
rect 6135 9976 6147 9979
rect 6457 9979 6515 9985
rect 6457 9976 6469 9979
rect 6135 9948 6469 9976
rect 6135 9945 6147 9948
rect 6089 9939 6147 9945
rect 6457 9945 6469 9948
rect 6503 9976 6515 9979
rect 7116 9976 7144 10007
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 8665 10047 8723 10053
rect 8665 10044 8677 10047
rect 7800 10016 8677 10044
rect 7800 10004 7806 10016
rect 8665 10013 8677 10016
rect 8711 10013 8723 10047
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 8665 10007 8723 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17126 10044 17132 10056
rect 17087 10016 17132 10044
rect 17126 10004 17132 10016
rect 17184 10004 17190 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 19153 10047 19211 10053
rect 19153 10044 19165 10047
rect 18380 10016 19165 10044
rect 18380 10004 18386 10016
rect 19153 10013 19165 10016
rect 19199 10044 19211 10047
rect 19889 10047 19947 10053
rect 19889 10044 19901 10047
rect 19199 10016 19901 10044
rect 19199 10013 19211 10016
rect 19153 10007 19211 10013
rect 19889 10013 19901 10016
rect 19935 10044 19947 10047
rect 20162 10044 20168 10056
rect 19935 10016 20168 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20162 10004 20168 10016
rect 20220 10044 20226 10056
rect 21545 10047 21603 10053
rect 21545 10044 21557 10047
rect 20220 10016 21557 10044
rect 20220 10004 20226 10016
rect 21545 10013 21557 10016
rect 21591 10044 21603 10047
rect 21726 10044 21732 10056
rect 21591 10016 21732 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21726 10004 21732 10016
rect 21784 10004 21790 10056
rect 6503 9948 7144 9976
rect 6503 9945 6515 9948
rect 6457 9939 6515 9945
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2222 9908 2228 9920
rect 2087 9880 2228 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 3697 9911 3755 9917
rect 3697 9877 3709 9911
rect 3743 9908 3755 9911
rect 4062 9908 4068 9920
rect 3743 9880 4068 9908
rect 3743 9877 3755 9880
rect 3697 9871 3755 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 5718 9868 5724 9920
rect 5776 9908 5782 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 5776 9880 6561 9908
rect 5776 9868 5782 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 6549 9871 6607 9877
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7432 9880 7573 9908
rect 7432 9868 7438 9880
rect 7561 9877 7573 9880
rect 7607 9877 7619 9911
rect 7561 9871 7619 9877
rect 8297 9911 8355 9917
rect 8297 9877 8309 9911
rect 8343 9908 8355 9911
rect 8386 9908 8392 9920
rect 8343 9880 8392 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 16482 9908 16488 9920
rect 16443 9880 16488 9908
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 20714 9868 20720 9920
rect 20772 9908 20778 9920
rect 21913 9911 21971 9917
rect 21913 9908 21925 9911
rect 20772 9880 21925 9908
rect 20772 9868 20778 9880
rect 21913 9877 21925 9880
rect 21959 9908 21971 9911
rect 22370 9908 22376 9920
rect 21959 9880 22376 9908
rect 21959 9877 21971 9880
rect 21913 9871 21971 9877
rect 22370 9868 22376 9880
rect 22428 9868 22434 9920
rect 24946 9868 24952 9920
rect 25004 9908 25010 9920
rect 25056 9908 25084 10084
rect 26513 10081 26525 10115
rect 26559 10112 26571 10115
rect 26602 10112 26608 10124
rect 26559 10084 26608 10112
rect 26559 10081 26571 10084
rect 26513 10075 26571 10081
rect 26602 10072 26608 10084
rect 26660 10072 26666 10124
rect 25225 10047 25283 10053
rect 25225 10013 25237 10047
rect 25271 10044 25283 10047
rect 25590 10044 25596 10056
rect 25271 10016 25596 10044
rect 25271 10013 25283 10016
rect 25225 10007 25283 10013
rect 25590 10004 25596 10016
rect 25648 10044 25654 10056
rect 26694 10044 26700 10056
rect 25648 10016 26700 10044
rect 25648 10004 25654 10016
rect 26694 10004 26700 10016
rect 26752 10044 26758 10056
rect 27065 10047 27123 10053
rect 27065 10044 27077 10047
rect 26752 10016 27077 10044
rect 26752 10004 26758 10016
rect 27065 10013 27077 10016
rect 27111 10013 27123 10047
rect 27065 10007 27123 10013
rect 26237 9979 26295 9985
rect 26237 9945 26249 9979
rect 26283 9976 26295 9979
rect 26510 9976 26516 9988
rect 26283 9948 26516 9976
rect 26283 9945 26295 9948
rect 26237 9939 26295 9945
rect 26510 9936 26516 9948
rect 26568 9936 26574 9988
rect 25004 9880 25084 9908
rect 26697 9911 26755 9917
rect 25004 9868 25010 9880
rect 26697 9877 26709 9911
rect 26743 9908 26755 9911
rect 26970 9908 26976 9920
rect 26743 9880 26976 9908
rect 26743 9877 26755 9880
rect 26697 9871 26755 9877
rect 26970 9868 26976 9880
rect 27028 9868 27034 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 2924 9676 3372 9704
rect 2924 9664 2930 9676
rect 2133 9639 2191 9645
rect 2133 9605 2145 9639
rect 2179 9636 2191 9639
rect 2498 9636 2504 9648
rect 2179 9608 2504 9636
rect 2179 9605 2191 9608
rect 2133 9599 2191 9605
rect 2498 9596 2504 9608
rect 2556 9596 2562 9648
rect 2958 9636 2964 9648
rect 2884 9608 2964 9636
rect 2884 9580 2912 9608
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 3344 9636 3372 9676
rect 3878 9664 3884 9716
rect 3936 9704 3942 9716
rect 6641 9707 6699 9713
rect 3936 9676 4108 9704
rect 3936 9664 3942 9676
rect 3602 9636 3608 9648
rect 3344 9608 3608 9636
rect 3602 9596 3608 9608
rect 3660 9596 3666 9648
rect 4080 9636 4108 9676
rect 6641 9673 6653 9707
rect 6687 9704 6699 9707
rect 7006 9704 7012 9716
rect 6687 9676 7012 9704
rect 6687 9673 6699 9676
rect 6641 9667 6699 9673
rect 7006 9664 7012 9676
rect 7064 9664 7070 9716
rect 8110 9704 8116 9716
rect 8071 9676 8116 9704
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 16942 9704 16948 9716
rect 16500 9676 16948 9704
rect 4157 9639 4215 9645
rect 4157 9636 4169 9639
rect 4080 9608 4169 9636
rect 4157 9605 4169 9608
rect 4203 9605 4215 9639
rect 4157 9599 4215 9605
rect 5629 9639 5687 9645
rect 5629 9605 5641 9639
rect 5675 9636 5687 9639
rect 6825 9639 6883 9645
rect 6825 9636 6837 9639
rect 5675 9608 6837 9636
rect 5675 9605 5687 9608
rect 5629 9599 5687 9605
rect 6825 9605 6837 9608
rect 6871 9605 6883 9639
rect 6825 9599 6883 9605
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 1394 9500 1400 9512
rect 1355 9472 1400 9500
rect 1394 9460 1400 9472
rect 1452 9460 1458 9512
rect 3050 9432 3056 9444
rect 3011 9404 3056 9432
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3160 9432 3188 9531
rect 3234 9528 3240 9580
rect 3292 9568 3298 9580
rect 3697 9571 3755 9577
rect 3292 9540 3464 9568
rect 3292 9528 3298 9540
rect 3436 9512 3464 9540
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 4706 9568 4712 9580
rect 3743 9540 4712 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 3418 9460 3424 9512
rect 3476 9460 3482 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5644 9500 5672 9599
rect 8938 9596 8944 9648
rect 8996 9636 9002 9648
rect 9122 9636 9128 9648
rect 8996 9608 9128 9636
rect 8996 9596 9002 9608
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 15654 9596 15660 9648
rect 15712 9636 15718 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15712 9608 15945 9636
rect 15712 9596 15718 9608
rect 15933 9605 15945 9608
rect 15979 9636 15991 9639
rect 16500 9636 16528 9676
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 19426 9704 19432 9716
rect 19076 9676 19432 9704
rect 15979 9608 16528 9636
rect 18601 9639 18659 9645
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 18601 9605 18613 9639
rect 18647 9636 18659 9639
rect 19076 9636 19104 9676
rect 19426 9664 19432 9676
rect 19484 9664 19490 9716
rect 21085 9707 21143 9713
rect 21085 9673 21097 9707
rect 21131 9704 21143 9707
rect 21358 9704 21364 9716
rect 21131 9676 21364 9704
rect 21131 9673 21143 9676
rect 21085 9667 21143 9673
rect 21358 9664 21364 9676
rect 21416 9664 21422 9716
rect 21726 9704 21732 9716
rect 21687 9676 21732 9704
rect 21726 9664 21732 9676
rect 21784 9664 21790 9716
rect 25222 9704 25228 9716
rect 25183 9676 25228 9704
rect 25222 9664 25228 9676
rect 25280 9664 25286 9716
rect 26602 9664 26608 9716
rect 26660 9704 26666 9716
rect 26973 9707 27031 9713
rect 26973 9704 26985 9707
rect 26660 9676 26985 9704
rect 26660 9664 26666 9676
rect 26973 9673 26985 9676
rect 27019 9673 27031 9707
rect 26973 9667 27031 9673
rect 18647 9608 19104 9636
rect 24397 9639 24455 9645
rect 18647 9605 18659 9608
rect 18601 9599 18659 9605
rect 24397 9605 24409 9639
rect 24443 9636 24455 9639
rect 24762 9636 24768 9648
rect 24443 9608 24768 9636
rect 24443 9605 24455 9608
rect 24397 9599 24455 9605
rect 24762 9596 24768 9608
rect 24820 9596 24826 9648
rect 25498 9636 25504 9648
rect 25459 9608 25504 9636
rect 25498 9596 25504 9608
rect 25556 9596 25562 9648
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6181 9571 6239 9577
rect 6181 9568 6193 9571
rect 5868 9540 6193 9568
rect 5868 9528 5874 9540
rect 6181 9537 6193 9540
rect 6227 9537 6239 9571
rect 7374 9568 7380 9580
rect 7335 9540 7380 9568
rect 6181 9531 6239 9537
rect 4571 9472 5672 9500
rect 6196 9500 6224 9531
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 15562 9568 15568 9580
rect 15475 9540 15568 9568
rect 15562 9528 15568 9540
rect 15620 9568 15626 9580
rect 16758 9568 16764 9580
rect 15620 9540 16764 9568
rect 15620 9528 15626 9540
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 17037 9571 17095 9577
rect 17037 9537 17049 9571
rect 17083 9568 17095 9571
rect 17126 9568 17132 9580
rect 17083 9540 17132 9568
rect 17083 9537 17095 9540
rect 17037 9531 17095 9537
rect 17126 9528 17132 9540
rect 17184 9568 17190 9580
rect 17184 9540 17908 9568
rect 17184 9528 17190 9540
rect 6822 9500 6828 9512
rect 6196 9472 6828 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 6822 9460 6828 9472
rect 6880 9460 6886 9512
rect 16298 9500 16304 9512
rect 16259 9472 16304 9500
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 3234 9432 3240 9444
rect 3160 9404 3240 9432
rect 3234 9392 3240 9404
rect 3292 9432 3298 9444
rect 3694 9432 3700 9444
rect 3292 9404 3700 9432
rect 3292 9392 3298 9404
rect 3694 9392 3700 9404
rect 3752 9392 3758 9444
rect 3970 9392 3976 9444
rect 4028 9432 4034 9444
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 4028 9404 4077 9432
rect 4028 9392 4034 9404
rect 4065 9401 4077 9404
rect 4111 9432 4123 9435
rect 4890 9432 4896 9444
rect 4111 9404 4896 9432
rect 4111 9401 4123 9404
rect 4065 9395 4123 9401
rect 4890 9392 4896 9404
rect 4948 9392 4954 9444
rect 5721 9435 5779 9441
rect 5721 9401 5733 9435
rect 5767 9432 5779 9435
rect 7190 9432 7196 9444
rect 5767 9404 7196 9432
rect 5767 9401 5779 9404
rect 5721 9395 5779 9401
rect 7190 9392 7196 9404
rect 7248 9392 7254 9444
rect 15286 9392 15292 9444
rect 15344 9432 15350 9444
rect 17880 9441 17908 9540
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21361 9571 21419 9577
rect 21361 9568 21373 9571
rect 21324 9540 21373 9568
rect 21324 9528 21330 9540
rect 21361 9537 21373 9540
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 19061 9503 19119 9509
rect 19061 9469 19073 9503
rect 19107 9500 19119 9503
rect 19150 9500 19156 9512
rect 19107 9472 19156 9500
rect 19107 9469 19119 9472
rect 19061 9463 19119 9469
rect 19150 9460 19156 9472
rect 19208 9460 19214 9512
rect 23934 9460 23940 9512
rect 23992 9500 23998 9512
rect 24029 9503 24087 9509
rect 24029 9500 24041 9503
rect 23992 9472 24041 9500
rect 23992 9460 23998 9472
rect 24029 9469 24041 9472
rect 24075 9500 24087 9503
rect 24213 9503 24271 9509
rect 24213 9500 24225 9503
rect 24075 9472 24225 9500
rect 24075 9469 24087 9472
rect 24029 9463 24087 9469
rect 24213 9469 24225 9472
rect 24259 9469 24271 9503
rect 25314 9500 25320 9512
rect 25275 9472 25320 9500
rect 24213 9463 24271 9469
rect 25314 9460 25320 9472
rect 25372 9500 25378 9512
rect 25869 9503 25927 9509
rect 25869 9500 25881 9503
rect 25372 9472 25881 9500
rect 25372 9460 25378 9472
rect 25869 9469 25881 9472
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 26329 9503 26387 9509
rect 26329 9469 26341 9503
rect 26375 9500 26387 9503
rect 26418 9500 26424 9512
rect 26375 9472 26424 9500
rect 26375 9469 26387 9472
rect 26329 9463 26387 9469
rect 26418 9460 26424 9472
rect 26476 9460 26482 9512
rect 27522 9500 27528 9512
rect 27483 9472 27528 9500
rect 27522 9460 27528 9472
rect 27580 9500 27586 9512
rect 28077 9503 28135 9509
rect 28077 9500 28089 9503
rect 27580 9472 28089 9500
rect 27580 9460 27586 9472
rect 28077 9469 28089 9472
rect 28123 9469 28135 9503
rect 28077 9463 28135 9469
rect 16761 9435 16819 9441
rect 16761 9432 16773 9435
rect 15344 9404 16773 9432
rect 15344 9392 15350 9404
rect 16761 9401 16773 9404
rect 16807 9432 16819 9435
rect 17405 9435 17463 9441
rect 17405 9432 17417 9435
rect 16807 9404 17417 9432
rect 16807 9401 16819 9404
rect 16761 9395 16819 9401
rect 17405 9401 17417 9404
rect 17451 9401 17463 9435
rect 17405 9395 17463 9401
rect 17865 9435 17923 9441
rect 17865 9401 17877 9435
rect 17911 9432 17923 9435
rect 19328 9435 19386 9441
rect 17911 9404 19012 9432
rect 17911 9401 17923 9404
rect 17865 9395 17923 9401
rect 1581 9367 1639 9373
rect 1581 9333 1593 9367
rect 1627 9364 1639 9367
rect 1670 9364 1676 9376
rect 1627 9336 1676 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2593 9367 2651 9373
rect 2593 9364 2605 9367
rect 1912 9336 2605 9364
rect 1912 9324 1918 9336
rect 2593 9333 2605 9336
rect 2639 9333 2651 9367
rect 2593 9327 2651 9333
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 2958 9364 2964 9376
rect 2832 9336 2964 9364
rect 2832 9324 2838 9336
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3068 9364 3096 9392
rect 3602 9364 3608 9376
rect 3068 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 4614 9364 4620 9376
rect 4527 9336 4620 9364
rect 4614 9324 4620 9336
rect 4672 9364 4678 9376
rect 5169 9367 5227 9373
rect 5169 9364 5181 9367
rect 4672 9336 5181 9364
rect 4672 9324 4678 9336
rect 5169 9333 5181 9336
rect 5215 9333 5227 9367
rect 5169 9327 5227 9333
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7285 9367 7343 9373
rect 7285 9364 7297 9367
rect 7064 9336 7297 9364
rect 7064 9324 7070 9336
rect 7285 9333 7297 9336
rect 7331 9333 7343 9367
rect 16390 9364 16396 9376
rect 16351 9336 16396 9364
rect 7285 9327 7343 9333
rect 16390 9324 16396 9336
rect 16448 9324 16454 9376
rect 16850 9364 16856 9376
rect 16811 9336 16856 9364
rect 16850 9324 16856 9336
rect 16908 9324 16914 9376
rect 18874 9364 18880 9376
rect 18835 9336 18880 9364
rect 18874 9324 18880 9336
rect 18932 9324 18938 9376
rect 18984 9364 19012 9404
rect 19328 9401 19340 9435
rect 19374 9432 19386 9435
rect 20622 9432 20628 9444
rect 19374 9404 20628 9432
rect 19374 9401 19386 9404
rect 19328 9395 19386 9401
rect 20622 9392 20628 9404
rect 20680 9392 20686 9444
rect 20438 9364 20444 9376
rect 18984 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 24854 9364 24860 9376
rect 24815 9336 24860 9364
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 26605 9367 26663 9373
rect 26605 9333 26617 9367
rect 26651 9364 26663 9367
rect 26694 9364 26700 9376
rect 26651 9336 26700 9364
rect 26651 9333 26663 9336
rect 26605 9327 26663 9333
rect 26694 9324 26700 9336
rect 26752 9324 26758 9376
rect 27709 9367 27767 9373
rect 27709 9333 27721 9367
rect 27755 9364 27767 9367
rect 27798 9364 27804 9376
rect 27755 9336 27804 9364
rect 27755 9333 27767 9336
rect 27709 9327 27767 9333
rect 27798 9324 27804 9336
rect 27856 9324 27862 9376
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1581 9163 1639 9169
rect 1581 9160 1593 9163
rect 1452 9132 1593 9160
rect 1452 9120 1458 9132
rect 1581 9129 1593 9132
rect 1627 9129 1639 9163
rect 1581 9123 1639 9129
rect 2038 9120 2044 9172
rect 2096 9160 2102 9172
rect 2317 9163 2375 9169
rect 2317 9160 2329 9163
rect 2096 9132 2329 9160
rect 2096 9120 2102 9132
rect 2317 9129 2329 9132
rect 2363 9129 2375 9163
rect 2866 9160 2872 9172
rect 2827 9132 2872 9160
rect 2317 9123 2375 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3602 9160 3608 9172
rect 3563 9132 3608 9160
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 7190 9160 7196 9172
rect 7151 9132 7196 9160
rect 7190 9120 7196 9132
rect 7248 9120 7254 9172
rect 15286 9160 15292 9172
rect 15247 9132 15292 9160
rect 15286 9120 15292 9132
rect 15344 9120 15350 9172
rect 19150 9160 19156 9172
rect 19111 9132 19156 9160
rect 19150 9120 19156 9132
rect 19208 9120 19214 9172
rect 19702 9160 19708 9172
rect 19663 9132 19708 9160
rect 19702 9120 19708 9132
rect 19760 9120 19766 9172
rect 24670 9160 24676 9172
rect 24631 9132 24676 9160
rect 24670 9120 24676 9132
rect 24728 9120 24734 9172
rect 2222 9092 2228 9104
rect 2183 9064 2228 9092
rect 2222 9052 2228 9064
rect 2280 9092 2286 9104
rect 2682 9092 2688 9104
rect 2280 9064 2688 9092
rect 2280 9052 2286 9064
rect 2682 9052 2688 9064
rect 2740 9052 2746 9104
rect 5160 9095 5218 9101
rect 5160 9061 5172 9095
rect 5206 9092 5218 9095
rect 5350 9092 5356 9104
rect 5206 9064 5356 9092
rect 5206 9061 5218 9064
rect 5160 9055 5218 9061
rect 5350 9052 5356 9064
rect 5408 9092 5414 9104
rect 7374 9092 7380 9104
rect 5408 9064 7380 9092
rect 5408 9052 5414 9064
rect 7374 9052 7380 9064
rect 7432 9092 7438 9104
rect 16574 9101 16580 9104
rect 16209 9095 16267 9101
rect 7432 9064 7880 9092
rect 7432 9052 7438 9064
rect 1854 8984 1860 9036
rect 1912 9024 1918 9036
rect 2866 9024 2872 9036
rect 1912 8996 2872 9024
rect 1912 8984 1918 8996
rect 2866 8984 2872 8996
rect 2924 8984 2930 9036
rect 7558 8984 7564 9036
rect 7616 9024 7622 9036
rect 7745 9027 7803 9033
rect 7745 9024 7757 9027
rect 7616 8996 7757 9024
rect 7616 8984 7622 8996
rect 7745 8993 7757 8996
rect 7791 8993 7803 9027
rect 7852 9024 7880 9064
rect 16209 9061 16221 9095
rect 16255 9092 16267 9095
rect 16568 9092 16580 9101
rect 16255 9064 16580 9092
rect 16255 9061 16267 9064
rect 16209 9055 16267 9061
rect 16568 9055 16580 9064
rect 16632 9092 16638 9104
rect 17126 9092 17132 9104
rect 16632 9064 17132 9092
rect 16574 9052 16580 9055
rect 16632 9052 16638 9064
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 19613 9095 19671 9101
rect 19613 9061 19625 9095
rect 19659 9092 19671 9095
rect 20530 9092 20536 9104
rect 19659 9064 20536 9092
rect 19659 9061 19671 9064
rect 19613 9055 19671 9061
rect 20530 9052 20536 9064
rect 20588 9052 20594 9104
rect 16298 9024 16304 9036
rect 7852 8996 7972 9024
rect 16259 8996 16304 9024
rect 7745 8987 7803 8993
rect 2501 8959 2559 8965
rect 2501 8956 2513 8959
rect 2424 8928 2513 8956
rect 2424 8900 2452 8928
rect 2501 8925 2513 8928
rect 2547 8956 2559 8959
rect 3234 8956 3240 8968
rect 2547 8928 3240 8956
rect 2547 8925 2559 8928
rect 2501 8919 2559 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4890 8956 4896 8968
rect 4851 8928 4896 8956
rect 4890 8916 4896 8928
rect 4948 8916 4954 8968
rect 6914 8916 6920 8968
rect 6972 8956 6978 8968
rect 7834 8956 7840 8968
rect 6972 8928 7840 8956
rect 6972 8916 6978 8928
rect 7834 8916 7840 8928
rect 7892 8916 7898 8968
rect 7944 8965 7972 8996
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 25314 9024 25320 9036
rect 25275 8996 25320 9024
rect 25314 8984 25320 8996
rect 25372 8984 25378 9036
rect 26510 9024 26516 9036
rect 26471 8996 26516 9024
rect 26510 8984 26516 8996
rect 26568 8984 26574 9036
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8202 8956 8208 8968
rect 7975 8928 8208 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8202 8916 8208 8928
rect 8260 8916 8266 8968
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8956 19947 8959
rect 20162 8956 20168 8968
rect 19935 8928 20168 8956
rect 19935 8925 19947 8928
rect 19889 8919 19947 8925
rect 2406 8848 2412 8900
rect 2464 8848 2470 8900
rect 4341 8891 4399 8897
rect 4341 8857 4353 8891
rect 4387 8888 4399 8891
rect 4706 8888 4712 8900
rect 4387 8860 4712 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 4706 8848 4712 8860
rect 4764 8888 4770 8900
rect 4764 8860 4936 8888
rect 4764 8848 4770 8860
rect 1854 8820 1860 8832
rect 1815 8792 1860 8820
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 4798 8820 4804 8832
rect 4759 8792 4804 8820
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4908 8820 4936 8860
rect 18598 8848 18604 8900
rect 18656 8888 18662 8900
rect 18785 8891 18843 8897
rect 18785 8888 18797 8891
rect 18656 8860 18797 8888
rect 18656 8848 18662 8860
rect 18785 8857 18797 8860
rect 18831 8888 18843 8891
rect 19904 8888 19932 8919
rect 20162 8916 20168 8928
rect 20220 8956 20226 8968
rect 20622 8956 20628 8968
rect 20220 8928 20628 8956
rect 20220 8916 20226 8928
rect 20622 8916 20628 8928
rect 20680 8916 20686 8968
rect 18831 8860 19932 8888
rect 18831 8857 18843 8860
rect 18785 8851 18843 8857
rect 5626 8820 5632 8832
rect 4908 8792 5632 8820
rect 5626 8780 5632 8792
rect 5684 8820 5690 8832
rect 6273 8823 6331 8829
rect 6273 8820 6285 8823
rect 5684 8792 6285 8820
rect 5684 8780 5690 8792
rect 6273 8789 6285 8792
rect 6319 8789 6331 8823
rect 6914 8820 6920 8832
rect 6875 8792 6920 8820
rect 6273 8783 6331 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7374 8820 7380 8832
rect 7335 8792 7380 8820
rect 7374 8780 7380 8792
rect 7432 8780 7438 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17000 8792 17693 8820
rect 17000 8780 17006 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 19150 8780 19156 8832
rect 19208 8820 19214 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 19208 8792 19257 8820
rect 19208 8780 19214 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 25498 8820 25504 8832
rect 25459 8792 25504 8820
rect 19245 8783 19303 8789
rect 25498 8780 25504 8792
rect 25556 8780 25562 8832
rect 25866 8780 25872 8832
rect 25924 8820 25930 8832
rect 26697 8823 26755 8829
rect 26697 8820 26709 8823
rect 25924 8792 26709 8820
rect 25924 8780 25930 8792
rect 26697 8789 26709 8792
rect 26743 8789 26755 8823
rect 26697 8783 26755 8789
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 1946 8616 1952 8628
rect 1907 8588 1952 8616
rect 1946 8576 1952 8588
rect 2004 8576 2010 8628
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3329 8619 3387 8625
rect 3329 8616 3341 8619
rect 3016 8588 3341 8616
rect 3016 8576 3022 8588
rect 3329 8585 3341 8588
rect 3375 8585 3387 8619
rect 3694 8616 3700 8628
rect 3655 8588 3700 8616
rect 3329 8579 3387 8585
rect 3694 8576 3700 8588
rect 3752 8576 3758 8628
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4212 8588 4813 8616
rect 4212 8576 4218 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 9125 8619 9183 8625
rect 9125 8616 9137 8619
rect 7892 8588 9137 8616
rect 7892 8576 7898 8588
rect 9125 8585 9137 8588
rect 9171 8585 9183 8619
rect 9125 8579 9183 8585
rect 16209 8619 16267 8625
rect 16209 8585 16221 8619
rect 16255 8616 16267 8619
rect 16298 8616 16304 8628
rect 16255 8588 16304 8616
rect 16255 8585 16267 8588
rect 16209 8579 16267 8585
rect 16298 8576 16304 8588
rect 16356 8616 16362 8628
rect 16666 8616 16672 8628
rect 16356 8588 16672 8616
rect 16356 8576 16362 8588
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 18598 8616 18604 8628
rect 18559 8588 18604 8616
rect 18598 8576 18604 8588
rect 18656 8576 18662 8628
rect 19702 8616 19708 8628
rect 19663 8588 19708 8616
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20530 8616 20536 8628
rect 20211 8588 20536 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 25130 8616 25136 8628
rect 25091 8588 25136 8616
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25314 8576 25320 8628
rect 25372 8616 25378 8628
rect 25869 8619 25927 8625
rect 25869 8616 25881 8619
rect 25372 8588 25881 8616
rect 25372 8576 25378 8588
rect 25869 8585 25881 8588
rect 25915 8585 25927 8619
rect 25869 8579 25927 8585
rect 26510 8576 26516 8628
rect 26568 8616 26574 8628
rect 27341 8619 27399 8625
rect 27341 8616 27353 8619
rect 26568 8588 27353 8616
rect 26568 8576 26574 8588
rect 27341 8585 27353 8588
rect 27387 8585 27399 8619
rect 27706 8616 27712 8628
rect 27667 8588 27712 8616
rect 27341 8579 27399 8585
rect 27706 8576 27712 8588
rect 27764 8576 27770 8628
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28077 8619 28135 8625
rect 28077 8616 28089 8619
rect 28040 8588 28089 8616
rect 28040 8576 28046 8588
rect 28077 8585 28089 8588
rect 28123 8585 28135 8619
rect 28077 8579 28135 8585
rect 1780 8480 1808 8576
rect 8202 8548 8208 8560
rect 8163 8520 8208 8548
rect 8202 8508 8208 8520
rect 8260 8548 8266 8560
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8260 8520 8769 8548
rect 8260 8508 8266 8520
rect 8757 8517 8769 8520
rect 8803 8517 8815 8551
rect 8757 8511 8815 8517
rect 15841 8551 15899 8557
rect 15841 8517 15853 8551
rect 15887 8548 15899 8551
rect 19720 8548 19748 8576
rect 25501 8551 25559 8557
rect 15887 8520 16896 8548
rect 19720 8520 20668 8548
rect 15887 8517 15899 8520
rect 15841 8511 15899 8517
rect 16868 8492 16896 8520
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 1780 8452 2513 8480
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3326 8480 3332 8492
rect 3099 8452 3332 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4430 8480 4436 8492
rect 4203 8452 4436 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2314 8412 2320 8424
rect 1912 8384 2320 8412
rect 1912 8372 1918 8384
rect 2314 8372 2320 8384
rect 2372 8372 2378 8424
rect 3513 8415 3571 8421
rect 3513 8381 3525 8415
rect 3559 8412 3571 8415
rect 4172 8412 4200 8443
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 5166 8480 5172 8492
rect 4856 8452 5172 8480
rect 4856 8440 4862 8452
rect 5166 8440 5172 8452
rect 5224 8480 5230 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 5224 8452 5273 8480
rect 5224 8440 5230 8452
rect 5261 8449 5273 8452
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5626 8480 5632 8492
rect 5491 8452 5632 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5626 8440 5632 8452
rect 5684 8440 5690 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 16482 8480 16488 8492
rect 15519 8452 16488 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 16482 8440 16488 8452
rect 16540 8480 16546 8492
rect 16761 8483 16819 8489
rect 16761 8480 16773 8483
rect 16540 8452 16773 8480
rect 16540 8440 16546 8452
rect 16761 8449 16773 8452
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 16850 8440 16856 8492
rect 16908 8480 16914 8492
rect 17865 8483 17923 8489
rect 16908 8452 17001 8480
rect 16908 8440 16914 8452
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 19150 8480 19156 8492
rect 17911 8452 19156 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 19702 8480 19708 8492
rect 19383 8452 19708 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 19702 8440 19708 8452
rect 19760 8480 19766 8492
rect 20438 8480 20444 8492
rect 19760 8452 20444 8480
rect 19760 8440 19766 8452
rect 20438 8440 20444 8452
rect 20496 8440 20502 8492
rect 20640 8480 20668 8520
rect 25501 8517 25513 8551
rect 25547 8548 25559 8551
rect 25590 8548 25596 8560
rect 25547 8520 25596 8548
rect 25547 8517 25559 8520
rect 25501 8511 25559 8517
rect 25590 8508 25596 8520
rect 25648 8508 25654 8560
rect 26602 8548 26608 8560
rect 26563 8520 26608 8548
rect 26602 8508 26608 8520
rect 26660 8508 26666 8560
rect 20640 8452 21956 8480
rect 3559 8384 4200 8412
rect 4709 8415 4767 8421
rect 3559 8381 3571 8384
rect 3513 8375 3571 8381
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4890 8412 4896 8424
rect 4755 8384 4896 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 4890 8372 4896 8384
rect 4948 8412 4954 8424
rect 6362 8412 6368 8424
rect 4948 8384 6368 8412
rect 4948 8372 4954 8384
rect 6362 8372 6368 8384
rect 6420 8412 6426 8424
rect 6546 8412 6552 8424
rect 6420 8384 6552 8412
rect 6420 8372 6426 8384
rect 6546 8372 6552 8384
rect 6604 8412 6610 8424
rect 6825 8415 6883 8421
rect 6825 8412 6837 8415
rect 6604 8384 6837 8412
rect 6604 8372 6610 8384
rect 6825 8381 6837 8384
rect 6871 8381 6883 8415
rect 6825 8375 6883 8381
rect 16390 8372 16396 8424
rect 16448 8412 16454 8424
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 16448 8384 16681 8412
rect 16448 8372 16454 8384
rect 16669 8381 16681 8384
rect 16715 8412 16727 8415
rect 17313 8415 17371 8421
rect 17313 8412 17325 8415
rect 16715 8384 17325 8412
rect 16715 8381 16727 8384
rect 16669 8375 16727 8381
rect 17313 8381 17325 8384
rect 17359 8381 17371 8415
rect 17313 8375 17371 8381
rect 5169 8347 5227 8353
rect 5169 8313 5181 8347
rect 5215 8344 5227 8347
rect 5258 8344 5264 8356
rect 5215 8316 5264 8344
rect 5215 8313 5227 8316
rect 5169 8307 5227 8313
rect 5258 8304 5264 8316
rect 5316 8304 5322 8356
rect 6273 8347 6331 8353
rect 6273 8313 6285 8347
rect 6319 8344 6331 8347
rect 7092 8347 7150 8353
rect 7092 8344 7104 8347
rect 6319 8316 7104 8344
rect 6319 8313 6331 8316
rect 6273 8307 6331 8313
rect 7092 8313 7104 8316
rect 7138 8344 7150 8347
rect 7282 8344 7288 8356
rect 7138 8316 7288 8344
rect 7138 8313 7150 8316
rect 7092 8307 7150 8313
rect 7282 8304 7288 8316
rect 7340 8304 7346 8356
rect 19061 8347 19119 8353
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 20441 8347 20499 8353
rect 20441 8344 20453 8347
rect 19107 8316 20453 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 20441 8313 20453 8316
rect 20487 8344 20499 8347
rect 20714 8344 20720 8356
rect 20487 8316 20720 8344
rect 20487 8313 20499 8316
rect 20441 8307 20499 8313
rect 20714 8304 20720 8316
rect 20772 8304 20778 8356
rect 2409 8279 2467 8285
rect 2409 8245 2421 8279
rect 2455 8276 2467 8279
rect 2866 8276 2872 8288
rect 2455 8248 2872 8276
rect 2455 8245 2467 8248
rect 2409 8239 2467 8245
rect 2866 8236 2872 8248
rect 2924 8236 2930 8288
rect 5350 8236 5356 8288
rect 5408 8276 5414 8288
rect 5813 8279 5871 8285
rect 5813 8276 5825 8279
rect 5408 8248 5825 8276
rect 5408 8236 5414 8248
rect 5813 8245 5825 8248
rect 5859 8245 5871 8279
rect 16298 8276 16304 8288
rect 16259 8248 16304 8276
rect 5813 8239 5871 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 18690 8276 18696 8288
rect 18651 8248 18696 8276
rect 18690 8236 18696 8248
rect 18748 8236 18754 8288
rect 21928 8276 21956 8452
rect 25130 8372 25136 8424
rect 25188 8412 25194 8424
rect 25317 8415 25375 8421
rect 25317 8412 25329 8415
rect 25188 8384 25329 8412
rect 25188 8372 25194 8384
rect 25317 8381 25329 8384
rect 25363 8381 25375 8415
rect 26418 8412 26424 8424
rect 26379 8384 26424 8412
rect 25317 8375 25375 8381
rect 26418 8372 26424 8384
rect 26476 8412 26482 8424
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26476 8384 26985 8412
rect 26476 8372 26482 8384
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 26973 8375 27031 8381
rect 27525 8415 27583 8421
rect 27525 8381 27537 8415
rect 27571 8412 27583 8415
rect 27982 8412 27988 8424
rect 27571 8384 27988 8412
rect 27571 8381 27583 8384
rect 27525 8375 27583 8381
rect 27982 8372 27988 8384
rect 28040 8372 28046 8424
rect 27062 8276 27068 8288
rect 21928 8248 27068 8276
rect 27062 8236 27068 8248
rect 27120 8236 27126 8288
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 2038 8032 2044 8084
rect 2096 8072 2102 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 2096 8044 2329 8072
rect 2096 8032 2102 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2317 8035 2375 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2924 8044 3433 8072
rect 2924 8032 2930 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 4614 8072 4620 8084
rect 4575 8044 4620 8072
rect 3421 8035 3479 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 4982 8072 4988 8084
rect 4943 8044 4988 8072
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5626 8072 5632 8084
rect 5587 8044 5632 8072
rect 5626 8032 5632 8044
rect 5684 8032 5690 8084
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6641 8075 6699 8081
rect 6641 8072 6653 8075
rect 6512 8044 6653 8072
rect 6512 8032 6518 8044
rect 6641 8041 6653 8044
rect 6687 8041 6699 8075
rect 6641 8035 6699 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7834 8072 7840 8084
rect 7524 8044 7840 8072
rect 7524 8032 7530 8044
rect 7834 8032 7840 8044
rect 7892 8072 7898 8084
rect 8205 8075 8263 8081
rect 8205 8072 8217 8075
rect 7892 8044 8217 8072
rect 7892 8032 7898 8044
rect 8205 8041 8217 8044
rect 8251 8041 8263 8075
rect 8205 8035 8263 8041
rect 16393 8075 16451 8081
rect 16393 8041 16405 8075
rect 16439 8072 16451 8075
rect 16482 8072 16488 8084
rect 16439 8044 16488 8072
rect 16439 8041 16451 8044
rect 16393 8035 16451 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 20162 8072 20168 8084
rect 20123 8044 20168 8072
rect 20162 8032 20168 8044
rect 20220 8032 20226 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 20901 8075 20959 8081
rect 20901 8072 20913 8075
rect 20772 8044 20913 8072
rect 20772 8032 20778 8044
rect 20901 8041 20913 8044
rect 20947 8041 20959 8075
rect 21266 8072 21272 8084
rect 21179 8044 21272 8072
rect 20901 8035 20959 8041
rect 21266 8032 21272 8044
rect 21324 8072 21330 8084
rect 21634 8072 21640 8084
rect 21324 8044 21640 8072
rect 21324 8032 21330 8044
rect 21634 8032 21640 8044
rect 21692 8032 21698 8084
rect 25498 8072 25504 8084
rect 25459 8044 25504 8072
rect 25498 8032 25504 8044
rect 25556 8032 25562 8084
rect 2222 7964 2228 8016
rect 2280 8004 2286 8016
rect 2280 7976 2544 8004
rect 2280 7964 2286 7976
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2041 7939 2099 7945
rect 2041 7905 2053 7939
rect 2087 7936 2099 7939
rect 2406 7936 2412 7948
rect 2087 7908 2412 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 2406 7896 2412 7908
rect 2464 7896 2470 7948
rect 2516 7945 2544 7976
rect 2774 7964 2780 8016
rect 2832 8004 2838 8016
rect 3053 8007 3111 8013
rect 3053 8004 3065 8007
rect 2832 7976 3065 8004
rect 2832 7964 2838 7976
rect 3053 7973 3065 7976
rect 3099 7973 3111 8007
rect 3053 7967 3111 7973
rect 4525 8007 4583 8013
rect 4525 7973 4537 8007
rect 4571 8004 4583 8007
rect 5258 8004 5264 8016
rect 4571 7976 5264 8004
rect 4571 7973 4583 7976
rect 4525 7967 4583 7973
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 8110 8004 8116 8016
rect 5368 7976 8116 8004
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7936 2559 7939
rect 2590 7936 2596 7948
rect 2547 7908 2596 7936
rect 2547 7905 2559 7908
rect 2501 7899 2559 7905
rect 2590 7896 2596 7908
rect 2648 7896 2654 7948
rect 5368 7936 5396 7976
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 16850 7964 16856 8016
rect 16908 8013 16914 8016
rect 16908 8007 16972 8013
rect 16908 7973 16926 8007
rect 16960 7973 16972 8007
rect 16908 7967 16972 7973
rect 16908 7964 16914 7967
rect 4172 7908 5396 7936
rect 1302 7828 1308 7880
rect 1360 7868 1366 7880
rect 4172 7868 4200 7908
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6328 7908 6561 7936
rect 6328 7896 6334 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 16666 7936 16672 7948
rect 16627 7908 16672 7936
rect 6549 7899 6607 7905
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 19058 7896 19064 7948
rect 19116 7936 19122 7948
rect 19521 7939 19579 7945
rect 19521 7936 19533 7939
rect 19116 7908 19533 7936
rect 19116 7896 19122 7908
rect 19521 7905 19533 7908
rect 19567 7905 19579 7939
rect 25314 7936 25320 7948
rect 25275 7908 25320 7936
rect 19521 7899 19579 7905
rect 25314 7896 25320 7908
rect 25372 7896 25378 7948
rect 26513 7939 26571 7945
rect 26513 7905 26525 7939
rect 26559 7936 26571 7939
rect 26786 7936 26792 7948
rect 26559 7908 26792 7936
rect 26559 7905 26571 7908
rect 26513 7899 26571 7905
rect 26786 7896 26792 7908
rect 26844 7896 26850 7948
rect 1360 7840 4200 7868
rect 5077 7871 5135 7877
rect 1360 7828 1366 7840
rect 5077 7837 5089 7871
rect 5123 7837 5135 7871
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 5077 7831 5135 7837
rect 5092 7744 5120 7831
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 6089 7871 6147 7877
rect 6089 7837 6101 7871
rect 6135 7868 6147 7871
rect 6825 7871 6883 7877
rect 6825 7868 6837 7871
rect 6135 7840 6837 7868
rect 6135 7837 6147 7840
rect 6089 7831 6147 7837
rect 6825 7837 6837 7840
rect 6871 7868 6883 7871
rect 7282 7868 7288 7880
rect 6871 7840 7288 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7282 7828 7288 7840
rect 7340 7828 7346 7880
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7558 7868 7564 7880
rect 7515 7840 7564 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 8294 7868 8300 7880
rect 8255 7840 8300 7868
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 19610 7868 19616 7880
rect 19571 7840 19616 7868
rect 19610 7828 19616 7840
rect 19668 7828 19674 7880
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 21358 7868 21364 7880
rect 19760 7840 19805 7868
rect 21319 7840 21364 7868
rect 19760 7828 19766 7840
rect 21358 7828 21364 7840
rect 21416 7828 21422 7880
rect 21453 7871 21511 7877
rect 21453 7837 21465 7871
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 5810 7760 5816 7812
rect 5868 7800 5874 7812
rect 6181 7803 6239 7809
rect 6181 7800 6193 7803
rect 5868 7772 6193 7800
rect 5868 7760 5874 7772
rect 6181 7769 6193 7772
rect 6227 7769 6239 7803
rect 9122 7800 9128 7812
rect 6181 7763 6239 7769
rect 6288 7772 9128 7800
rect 1394 7692 1400 7744
rect 1452 7732 1458 7744
rect 1581 7735 1639 7741
rect 1581 7732 1593 7735
rect 1452 7704 1593 7732
rect 1452 7692 1458 7704
rect 1581 7701 1593 7704
rect 1627 7701 1639 7735
rect 5074 7732 5080 7744
rect 4987 7704 5080 7732
rect 1581 7695 1639 7701
rect 5074 7692 5080 7704
rect 5132 7732 5138 7744
rect 6288 7732 6316 7772
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 18785 7803 18843 7809
rect 18785 7769 18797 7803
rect 18831 7800 18843 7803
rect 19242 7800 19248 7812
rect 18831 7772 19248 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 19242 7760 19248 7772
rect 19300 7800 19306 7812
rect 19720 7800 19748 7828
rect 19300 7772 19748 7800
rect 19300 7760 19306 7772
rect 20162 7760 20168 7812
rect 20220 7800 20226 7812
rect 21468 7800 21496 7831
rect 21634 7800 21640 7812
rect 20220 7772 21640 7800
rect 20220 7760 20226 7772
rect 21634 7760 21640 7772
rect 21692 7760 21698 7812
rect 7742 7732 7748 7744
rect 5132 7704 6316 7732
rect 7703 7704 7748 7732
rect 5132 7692 5138 7704
rect 7742 7692 7748 7704
rect 7800 7692 7806 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 17092 7704 18061 7732
rect 17092 7692 17098 7704
rect 18049 7701 18061 7704
rect 18095 7732 18107 7735
rect 18598 7732 18604 7744
rect 18095 7704 18604 7732
rect 18095 7701 18107 7704
rect 18049 7695 18107 7701
rect 18598 7692 18604 7704
rect 18656 7692 18662 7744
rect 19150 7732 19156 7744
rect 19111 7704 19156 7732
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 26697 7735 26755 7741
rect 26697 7701 26709 7735
rect 26743 7732 26755 7735
rect 26786 7732 26792 7744
rect 26743 7704 26792 7732
rect 26743 7701 26755 7704
rect 26697 7695 26755 7701
rect 26786 7692 26792 7704
rect 26844 7692 26850 7744
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 1578 7488 1584 7540
rect 1636 7528 1642 7540
rect 1949 7531 2007 7537
rect 1949 7528 1961 7531
rect 1636 7500 1961 7528
rect 1636 7488 1642 7500
rect 1949 7497 1961 7500
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 2409 7531 2467 7537
rect 2409 7497 2421 7531
rect 2455 7528 2467 7531
rect 2590 7528 2596 7540
rect 2455 7500 2596 7528
rect 2455 7497 2467 7500
rect 2409 7491 2467 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 4246 7528 4252 7540
rect 4207 7500 4252 7528
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4709 7531 4767 7537
rect 4709 7497 4721 7531
rect 4755 7528 4767 7531
rect 4982 7528 4988 7540
rect 4755 7500 4988 7528
rect 4755 7497 4767 7500
rect 4709 7491 4767 7497
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5166 7528 5172 7540
rect 5127 7500 5172 7528
rect 5166 7488 5172 7500
rect 5224 7488 5230 7540
rect 6273 7531 6331 7537
rect 6273 7497 6285 7531
rect 6319 7528 6331 7531
rect 6454 7528 6460 7540
rect 6319 7500 6460 7528
rect 6319 7497 6331 7500
rect 6273 7491 6331 7497
rect 6454 7488 6460 7500
rect 6512 7488 6518 7540
rect 6822 7528 6828 7540
rect 6783 7500 6828 7528
rect 6822 7488 6828 7500
rect 6880 7488 6886 7540
rect 7834 7528 7840 7540
rect 7795 7500 7840 7528
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 8168 7500 8217 7528
rect 8168 7488 8174 7500
rect 8205 7497 8217 7500
rect 8251 7497 8263 7531
rect 8205 7491 8263 7497
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 17034 7528 17040 7540
rect 16347 7500 17040 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 17034 7488 17040 7500
rect 17092 7488 17098 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 19153 7531 19211 7537
rect 19153 7528 19165 7531
rect 19116 7500 19165 7528
rect 19116 7488 19122 7500
rect 19153 7497 19165 7500
rect 19199 7497 19211 7531
rect 19153 7491 19211 7497
rect 20993 7531 21051 7537
rect 20993 7497 21005 7531
rect 21039 7528 21051 7531
rect 21358 7528 21364 7540
rect 21039 7500 21364 7528
rect 21039 7497 21051 7500
rect 20993 7491 21051 7497
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 21634 7528 21640 7540
rect 21595 7500 21640 7528
rect 21634 7488 21640 7500
rect 21692 7488 21698 7540
rect 25314 7528 25320 7540
rect 25275 7500 25320 7528
rect 25314 7488 25320 7500
rect 25372 7488 25378 7540
rect 27062 7528 27068 7540
rect 27023 7500 27068 7528
rect 27062 7488 27068 7500
rect 27120 7488 27126 7540
rect 2682 7460 2688 7472
rect 2643 7432 2688 7460
rect 2682 7420 2688 7432
rect 2740 7420 2746 7472
rect 5074 7460 5080 7472
rect 5035 7432 5080 7460
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 18049 7463 18107 7469
rect 18049 7460 18061 7463
rect 16868 7432 18061 7460
rect 3142 7392 3148 7404
rect 2516 7364 3148 7392
rect 1397 7327 1455 7333
rect 1397 7293 1409 7327
rect 1443 7324 1455 7327
rect 1578 7324 1584 7336
rect 1443 7296 1584 7324
rect 1443 7293 1455 7296
rect 1397 7287 1455 7293
rect 1578 7284 1584 7296
rect 1636 7284 1642 7336
rect 2516 7333 2544 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 5258 7352 5264 7404
rect 5316 7392 5322 7404
rect 5721 7395 5779 7401
rect 5721 7392 5733 7395
rect 5316 7364 5733 7392
rect 5316 7352 5322 7364
rect 5721 7361 5733 7364
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 7282 7352 7288 7404
rect 7340 7392 7346 7404
rect 7469 7395 7527 7401
rect 7469 7392 7481 7395
rect 7340 7364 7481 7392
rect 7340 7352 7346 7364
rect 7469 7361 7481 7364
rect 7515 7392 7527 7395
rect 8294 7392 8300 7404
rect 7515 7364 8300 7392
rect 7515 7361 7527 7364
rect 7469 7355 7527 7361
rect 8294 7352 8300 7364
rect 8352 7352 8358 7404
rect 16868 7401 16896 7432
rect 18049 7429 18061 7432
rect 18095 7429 18107 7463
rect 21266 7460 21272 7472
rect 21227 7432 21272 7460
rect 18049 7423 18107 7429
rect 21266 7420 21272 7432
rect 21324 7420 21330 7472
rect 26878 7420 26884 7472
rect 26936 7460 26942 7472
rect 27341 7463 27399 7469
rect 27341 7460 27353 7463
rect 26936 7432 27353 7460
rect 26936 7420 26942 7432
rect 27341 7429 27353 7432
rect 27387 7429 27399 7463
rect 27341 7423 27399 7429
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16853 7395 16911 7401
rect 16853 7392 16865 7395
rect 15979 7364 16865 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16853 7361 16865 7364
rect 16899 7361 16911 7395
rect 17034 7392 17040 7404
rect 16995 7364 17040 7392
rect 16853 7355 16911 7361
rect 17034 7352 17040 7364
rect 17092 7352 17098 7404
rect 18601 7395 18659 7401
rect 18601 7392 18613 7395
rect 17788 7364 18613 7392
rect 2507 7327 2565 7333
rect 2507 7293 2519 7327
rect 2553 7293 2565 7327
rect 2507 7287 2565 7293
rect 3605 7327 3663 7333
rect 3605 7293 3617 7327
rect 3651 7324 3663 7327
rect 4246 7324 4252 7336
rect 3651 7296 4252 7324
rect 3651 7293 3663 7296
rect 3605 7287 3663 7293
rect 4246 7284 4252 7296
rect 4304 7284 4310 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7324 5687 7327
rect 5810 7324 5816 7336
rect 5675 7296 5816 7324
rect 5675 7293 5687 7296
rect 5629 7287 5687 7293
rect 5810 7284 5816 7296
rect 5868 7284 5874 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7324 6699 7327
rect 6730 7324 6736 7336
rect 6687 7296 6736 7324
rect 6687 7293 6699 7296
rect 6641 7287 6699 7293
rect 6730 7284 6736 7296
rect 6788 7324 6794 7336
rect 7374 7324 7380 7336
rect 6788 7296 7380 7324
rect 6788 7284 6794 7296
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7324 15623 7327
rect 16298 7324 16304 7336
rect 15611 7296 16304 7324
rect 15611 7293 15623 7296
rect 15565 7287 15623 7293
rect 16298 7284 16304 7296
rect 16356 7324 16362 7336
rect 16761 7327 16819 7333
rect 16761 7324 16773 7327
rect 16356 7296 16773 7324
rect 16356 7284 16362 7296
rect 16761 7293 16773 7296
rect 16807 7293 16819 7327
rect 16761 7287 16819 7293
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 5537 7259 5595 7265
rect 5537 7256 5549 7259
rect 5500 7228 5549 7256
rect 5500 7216 5506 7228
rect 5537 7225 5549 7228
rect 5583 7256 5595 7259
rect 7742 7256 7748 7268
rect 5583 7228 7748 7256
rect 5583 7225 5595 7228
rect 5537 7219 5595 7225
rect 7742 7216 7748 7228
rect 7800 7216 7806 7268
rect 16850 7216 16856 7268
rect 16908 7256 16914 7268
rect 17788 7265 17816 7364
rect 18601 7361 18613 7364
rect 18647 7361 18659 7395
rect 20162 7392 20168 7404
rect 20123 7364 20168 7392
rect 18601 7355 18659 7361
rect 20162 7352 20168 7364
rect 20220 7352 20226 7404
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7324 18475 7327
rect 18506 7324 18512 7336
rect 18463 7296 18512 7324
rect 18463 7293 18475 7296
rect 18417 7287 18475 7293
rect 18506 7284 18512 7296
rect 18564 7324 18570 7336
rect 19150 7324 19156 7336
rect 18564 7296 19156 7324
rect 18564 7284 18570 7296
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 19978 7324 19984 7336
rect 19939 7296 19984 7324
rect 19978 7284 19984 7296
rect 20036 7284 20042 7336
rect 26421 7327 26479 7333
rect 26421 7293 26433 7327
rect 26467 7324 26479 7327
rect 27062 7324 27068 7336
rect 26467 7296 27068 7324
rect 26467 7293 26479 7296
rect 26421 7287 26479 7293
rect 27062 7284 27068 7296
rect 27120 7284 27126 7336
rect 27154 7284 27160 7336
rect 27212 7324 27218 7336
rect 27525 7327 27583 7333
rect 27525 7324 27537 7327
rect 27212 7296 27537 7324
rect 27212 7284 27218 7296
rect 27525 7293 27537 7296
rect 27571 7324 27583 7327
rect 28077 7327 28135 7333
rect 28077 7324 28089 7327
rect 27571 7296 28089 7324
rect 27571 7293 27583 7296
rect 27525 7287 27583 7293
rect 28077 7293 28089 7296
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 17773 7259 17831 7265
rect 17773 7256 17785 7259
rect 16908 7228 17785 7256
rect 16908 7216 16914 7228
rect 17773 7225 17785 7228
rect 17819 7225 17831 7259
rect 17773 7219 17831 7225
rect 19702 7216 19708 7268
rect 19760 7256 19766 7268
rect 20073 7259 20131 7265
rect 20073 7256 20085 7259
rect 19760 7228 20085 7256
rect 19760 7216 19766 7228
rect 20073 7225 20085 7228
rect 20119 7225 20131 7259
rect 20073 7219 20131 7225
rect 1578 7188 1584 7200
rect 1539 7160 1584 7188
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3786 7188 3792 7200
rect 3747 7160 3792 7188
rect 3786 7148 3792 7160
rect 3844 7148 3850 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 7064 7160 7205 7188
rect 7064 7148 7070 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7374 7188 7380 7200
rect 7331 7160 7380 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8573 7191 8631 7197
rect 8573 7188 8585 7191
rect 8352 7160 8585 7188
rect 8352 7148 8358 7160
rect 8573 7157 8585 7160
rect 8619 7157 8631 7191
rect 16390 7188 16396 7200
rect 16351 7160 16396 7188
rect 8573 7151 8631 7157
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 17405 7191 17463 7197
rect 17405 7188 17417 7191
rect 16724 7160 17417 7188
rect 16724 7148 16730 7160
rect 17405 7157 17417 7160
rect 17451 7157 17463 7191
rect 17405 7151 17463 7157
rect 18509 7191 18567 7197
rect 18509 7157 18521 7191
rect 18555 7188 18567 7191
rect 18690 7188 18696 7200
rect 18555 7160 18696 7188
rect 18555 7157 18567 7160
rect 18509 7151 18567 7157
rect 18690 7148 18696 7160
rect 18748 7148 18754 7200
rect 19610 7188 19616 7200
rect 19571 7160 19616 7188
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 26605 7191 26663 7197
rect 26605 7157 26617 7191
rect 26651 7188 26663 7191
rect 26878 7188 26884 7200
rect 26651 7160 26884 7188
rect 26651 7157 26663 7160
rect 26605 7151 26663 7157
rect 26878 7148 26884 7160
rect 26936 7148 26942 7200
rect 27706 7188 27712 7200
rect 27667 7160 27712 7188
rect 27706 7148 27712 7160
rect 27764 7148 27770 7200
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 2038 6984 2044 6996
rect 1999 6956 2044 6984
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 4709 6987 4767 6993
rect 4709 6953 4721 6987
rect 4755 6984 4767 6987
rect 5169 6987 5227 6993
rect 5169 6984 5181 6987
rect 4755 6956 5181 6984
rect 4755 6953 4767 6956
rect 4709 6947 4767 6953
rect 5169 6953 5181 6956
rect 5215 6984 5227 6987
rect 5258 6984 5264 6996
rect 5215 6956 5264 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 5629 6987 5687 6993
rect 5629 6953 5641 6987
rect 5675 6984 5687 6987
rect 5810 6984 5816 6996
rect 5675 6956 5816 6984
rect 5675 6953 5687 6956
rect 5629 6947 5687 6953
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 6270 6984 6276 6996
rect 6231 6956 6276 6984
rect 6270 6944 6276 6956
rect 6328 6944 6334 6996
rect 7282 6984 7288 6996
rect 7243 6956 7288 6984
rect 7282 6944 7288 6956
rect 7340 6944 7346 6996
rect 16761 6987 16819 6993
rect 16761 6953 16773 6987
rect 16807 6984 16819 6987
rect 16850 6984 16856 6996
rect 16807 6956 16856 6984
rect 16807 6953 16819 6956
rect 16761 6947 16819 6953
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 18506 6984 18512 6996
rect 18467 6956 18512 6984
rect 18506 6944 18512 6956
rect 18564 6944 18570 6996
rect 19242 6984 19248 6996
rect 19203 6956 19248 6984
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 19702 6984 19708 6996
rect 19663 6956 19708 6984
rect 19702 6944 19708 6956
rect 19760 6944 19766 6996
rect 19978 6984 19984 6996
rect 19939 6956 19984 6984
rect 19978 6944 19984 6956
rect 20036 6944 20042 6996
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6916 18199 6919
rect 18690 6916 18696 6928
rect 18187 6888 18696 6916
rect 18187 6885 18199 6888
rect 18141 6879 18199 6885
rect 18690 6876 18696 6888
rect 18748 6876 18754 6928
rect 19610 6916 19616 6928
rect 19260 6888 19616 6916
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2038 6848 2044 6860
rect 1443 6820 2044 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2498 6848 2504 6860
rect 2459 6820 2504 6848
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 15289 6851 15347 6857
rect 15289 6817 15301 6851
rect 15335 6848 15347 6851
rect 15378 6848 15384 6860
rect 15335 6820 15384 6848
rect 15335 6817 15347 6820
rect 15289 6811 15347 6817
rect 15378 6808 15384 6820
rect 15436 6848 15442 6860
rect 16390 6848 16396 6860
rect 15436 6820 16396 6848
rect 15436 6808 15442 6820
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 18877 6851 18935 6857
rect 18877 6817 18889 6851
rect 18923 6848 18935 6851
rect 19260 6848 19288 6888
rect 19610 6876 19616 6888
rect 19668 6876 19674 6928
rect 26510 6848 26516 6860
rect 18923 6820 19288 6848
rect 26471 6820 26516 6848
rect 18923 6817 18935 6820
rect 18877 6811 18935 6817
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 2130 6672 2136 6724
rect 2188 6712 2194 6724
rect 2685 6715 2743 6721
rect 2685 6712 2697 6715
rect 2188 6684 2697 6712
rect 2188 6672 2194 6684
rect 2685 6681 2697 6684
rect 2731 6681 2743 6715
rect 2685 6675 2743 6681
rect 1578 6644 1584 6656
rect 1539 6616 1584 6644
rect 1578 6604 1584 6616
rect 1636 6604 1642 6656
rect 6914 6644 6920 6656
rect 6875 6616 6920 6644
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 26694 6644 26700 6656
rect 26655 6616 26700 6644
rect 26694 6604 26700 6616
rect 26752 6604 26758 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 1544 6412 1593 6440
rect 1544 6400 1550 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 2406 6440 2412 6452
rect 2367 6412 2412 6440
rect 1581 6403 1639 6409
rect 2406 6400 2412 6412
rect 2464 6400 2470 6452
rect 3142 6440 3148 6452
rect 3103 6412 3148 6440
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 5261 6443 5319 6449
rect 5261 6409 5273 6443
rect 5307 6440 5319 6443
rect 5442 6440 5448 6452
rect 5307 6412 5448 6440
rect 5307 6409 5319 6412
rect 5261 6403 5319 6409
rect 5442 6400 5448 6412
rect 5500 6400 5506 6452
rect 15378 6440 15384 6452
rect 15339 6412 15384 6440
rect 15378 6400 15384 6412
rect 15436 6400 15442 6452
rect 26510 6440 26516 6452
rect 26471 6412 26516 6440
rect 26510 6400 26516 6412
rect 26568 6400 26574 6452
rect 2038 6372 2044 6384
rect 1951 6344 2044 6372
rect 2038 6332 2044 6344
rect 2096 6372 2102 6384
rect 5074 6372 5080 6384
rect 2096 6344 5080 6372
rect 2096 6332 2102 6344
rect 5074 6332 5080 6344
rect 5132 6332 5138 6384
rect 1397 6239 1455 6245
rect 1397 6205 1409 6239
rect 1443 6236 1455 6239
rect 2406 6236 2412 6248
rect 1443 6208 2412 6236
rect 1443 6205 1455 6208
rect 1397 6199 1455 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2501 6239 2559 6245
rect 2501 6205 2513 6239
rect 2547 6236 2559 6239
rect 3142 6236 3148 6248
rect 2547 6208 3148 6236
rect 2547 6205 2559 6208
rect 2501 6199 2559 6205
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 2498 5896 2504 5908
rect 2459 5868 2504 5896
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 1360 5732 1409 5760
rect 1360 5720 1366 5732
rect 1397 5729 1409 5732
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 1394 5516 1400 5568
rect 1452 5556 1458 5568
rect 1581 5559 1639 5565
rect 1581 5556 1593 5559
rect 1452 5528 1593 5556
rect 1452 5516 1458 5528
rect 1581 5525 1593 5528
rect 1627 5525 1639 5559
rect 1581 5519 1639 5525
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1360 5324 1593 5352
rect 1360 5312 1366 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 26418 5148 26424 5160
rect 26379 5120 26424 5148
rect 26418 5108 26424 5120
rect 26476 5148 26482 5160
rect 26973 5151 27031 5157
rect 26973 5148 26985 5151
rect 26476 5120 26985 5148
rect 26476 5108 26482 5120
rect 26973 5117 26985 5120
rect 27019 5117 27031 5151
rect 26973 5111 27031 5117
rect 26602 5012 26608 5024
rect 26563 4984 26608 5012
rect 26602 4972 26608 4984
rect 26660 4972 26666 5024
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 1397 2975 1455 2981
rect 1397 2941 1409 2975
rect 1443 2972 1455 2975
rect 2038 2972 2044 2984
rect 1443 2944 2044 2972
rect 1443 2941 1455 2944
rect 1397 2935 1455 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 26418 2972 26424 2984
rect 26379 2944 26424 2972
rect 26418 2932 26424 2944
rect 26476 2972 26482 2984
rect 26973 2975 27031 2981
rect 26973 2972 26985 2975
rect 26476 2944 26985 2972
rect 26476 2932 26482 2944
rect 26973 2941 26985 2944
rect 27019 2941 27031 2975
rect 26973 2935 27031 2941
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 26602 2836 26608 2848
rect 26563 2808 26608 2836
rect 26602 2796 26608 2808
rect 26660 2796 26666 2848
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 6365 2635 6423 2641
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6546 2632 6552 2644
rect 6411 2604 6552 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 8294 2632 8300 2644
rect 8255 2604 8300 2632
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 7190 2505 7196 2508
rect 6733 2499 6791 2505
rect 6733 2465 6745 2499
rect 6779 2496 6791 2499
rect 7184 2496 7196 2505
rect 6779 2468 7196 2496
rect 6779 2465 6791 2468
rect 6733 2459 6791 2465
rect 7184 2459 7196 2468
rect 7190 2456 7196 2459
rect 7248 2456 7254 2508
rect 6546 2388 6552 2440
rect 6604 2428 6610 2440
rect 6917 2431 6975 2437
rect 6917 2428 6929 2431
rect 6604 2400 6929 2428
rect 6604 2388 6610 2400
rect 6917 2397 6929 2400
rect 6963 2397 6975 2431
rect 6917 2391 6975 2397
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 3332 22788 3384 22840
rect 10600 22788 10652 22840
rect 3516 22516 3568 22568
rect 7380 22516 7432 22568
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 14004 21088 14056 21140
rect 19616 21088 19668 21140
rect 17960 21020 18012 21072
rect 12164 20995 12216 21004
rect 12164 20961 12173 20995
rect 12173 20961 12207 20995
rect 12207 20961 12216 20995
rect 12164 20952 12216 20961
rect 16580 20952 16632 21004
rect 18972 20952 19024 21004
rect 18512 20884 18564 20936
rect 4068 20816 4120 20868
rect 5632 20816 5684 20868
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 19248 20816 19300 20868
rect 21732 20816 21784 20868
rect 25044 20816 25096 20868
rect 4988 20791 5040 20800
rect 4988 20757 4997 20791
rect 4997 20757 5031 20791
rect 5031 20757 5040 20791
rect 4988 20748 5040 20757
rect 12716 20791 12768 20800
rect 12716 20757 12725 20791
rect 12725 20757 12759 20791
rect 12759 20757 12768 20791
rect 12716 20748 12768 20757
rect 18328 20791 18380 20800
rect 18328 20757 18337 20791
rect 18337 20757 18371 20791
rect 18371 20757 18380 20791
rect 18328 20748 18380 20757
rect 20168 20791 20220 20800
rect 20168 20757 20177 20791
rect 20177 20757 20211 20791
rect 20211 20757 20220 20791
rect 20168 20748 20220 20757
rect 22192 20748 22244 20800
rect 24860 20748 24912 20800
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 940 20544 992 20596
rect 2688 20544 2740 20596
rect 8208 20544 8260 20596
rect 10232 20544 10284 20596
rect 15844 20544 15896 20596
rect 17776 20544 17828 20596
rect 20168 20544 20220 20596
rect 12164 20476 12216 20528
rect 17960 20476 18012 20528
rect 19340 20476 19392 20528
rect 4988 20408 5040 20460
rect 2136 20340 2188 20392
rect 4712 20340 4764 20392
rect 12716 20408 12768 20460
rect 1952 20247 2004 20256
rect 1952 20213 1961 20247
rect 1961 20213 1995 20247
rect 1995 20213 2004 20247
rect 1952 20204 2004 20213
rect 4160 20204 4212 20256
rect 17592 20408 17644 20460
rect 25228 20544 25280 20596
rect 26608 20587 26660 20596
rect 26608 20553 26617 20587
rect 26617 20553 26651 20587
rect 26651 20553 26660 20587
rect 26608 20544 26660 20553
rect 25412 20519 25464 20528
rect 25412 20485 25421 20519
rect 25421 20485 25455 20519
rect 25455 20485 25464 20519
rect 25412 20476 25464 20485
rect 13636 20340 13688 20392
rect 13820 20340 13872 20392
rect 16764 20383 16816 20392
rect 16764 20349 16773 20383
rect 16773 20349 16807 20383
rect 16807 20349 16816 20383
rect 16764 20340 16816 20349
rect 20168 20340 20220 20392
rect 12808 20315 12860 20324
rect 12808 20281 12817 20315
rect 12817 20281 12851 20315
rect 12851 20281 12860 20315
rect 12808 20272 12860 20281
rect 19984 20315 20036 20324
rect 19984 20281 19993 20315
rect 19993 20281 20027 20315
rect 20027 20281 20036 20315
rect 19984 20272 20036 20281
rect 4896 20247 4948 20256
rect 4896 20213 4905 20247
rect 4905 20213 4939 20247
rect 4939 20213 4948 20247
rect 4896 20204 4948 20213
rect 7472 20204 7524 20256
rect 9772 20247 9824 20256
rect 9772 20213 9781 20247
rect 9781 20213 9815 20247
rect 9815 20213 9824 20247
rect 9772 20204 9824 20213
rect 12256 20204 12308 20256
rect 16580 20247 16632 20256
rect 16580 20213 16589 20247
rect 16589 20213 16623 20247
rect 16623 20213 16632 20247
rect 16580 20204 16632 20213
rect 18604 20204 18656 20256
rect 18696 20204 18748 20256
rect 19340 20204 19392 20256
rect 24768 20204 24820 20256
rect 26608 20340 26660 20392
rect 25872 20204 25924 20256
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 4436 20043 4488 20052
rect 4436 20009 4445 20043
rect 4445 20009 4479 20043
rect 4479 20009 4488 20043
rect 4436 20000 4488 20009
rect 4988 20000 5040 20052
rect 5632 20043 5684 20052
rect 5632 20009 5641 20043
rect 5641 20009 5675 20043
rect 5675 20009 5684 20043
rect 5632 20000 5684 20009
rect 12716 20000 12768 20052
rect 16764 20043 16816 20052
rect 16764 20009 16773 20043
rect 16773 20009 16807 20043
rect 16807 20009 16816 20043
rect 16764 20000 16816 20009
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 21548 20000 21600 20052
rect 23388 20000 23440 20052
rect 12256 19932 12308 19984
rect 4068 19864 4120 19916
rect 12348 19864 12400 19916
rect 15200 19864 15252 19916
rect 15752 19907 15804 19916
rect 15752 19873 15761 19907
rect 15761 19873 15795 19907
rect 15795 19873 15804 19907
rect 17776 19907 17828 19916
rect 15752 19864 15804 19873
rect 17776 19873 17785 19907
rect 17785 19873 17819 19907
rect 17819 19873 17828 19907
rect 17776 19864 17828 19873
rect 19616 19864 19668 19916
rect 20904 19907 20956 19916
rect 20904 19873 20913 19907
rect 20913 19873 20947 19907
rect 20947 19873 20956 19907
rect 20904 19864 20956 19873
rect 21916 19907 21968 19916
rect 21916 19873 21925 19907
rect 21925 19873 21959 19907
rect 21959 19873 21968 19907
rect 21916 19864 21968 19873
rect 5724 19839 5776 19848
rect 5724 19805 5733 19839
rect 5733 19805 5767 19839
rect 5767 19805 5776 19839
rect 5724 19796 5776 19805
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 19156 19796 19208 19848
rect 18788 19728 18840 19780
rect 20720 19796 20772 19848
rect 27436 19796 27488 19848
rect 3884 19660 3936 19712
rect 5264 19660 5316 19712
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 14924 19703 14976 19712
rect 14924 19669 14933 19703
rect 14933 19669 14967 19703
rect 14967 19669 14976 19703
rect 14924 19660 14976 19669
rect 15292 19703 15344 19712
rect 15292 19669 15301 19703
rect 15301 19669 15335 19703
rect 15335 19669 15344 19703
rect 15292 19660 15344 19669
rect 18236 19660 18288 19712
rect 18696 19660 18748 19712
rect 20168 19703 20220 19712
rect 20168 19669 20177 19703
rect 20177 19669 20211 19703
rect 20211 19669 20220 19703
rect 20168 19660 20220 19669
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 5632 19456 5684 19508
rect 6368 19456 6420 19508
rect 13636 19456 13688 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 17684 19456 17736 19508
rect 14556 19388 14608 19440
rect 14924 19388 14976 19440
rect 3700 19320 3752 19372
rect 4896 19320 4948 19372
rect 5264 19320 5316 19372
rect 5724 19252 5776 19304
rect 12164 19320 12216 19372
rect 10876 19252 10928 19304
rect 1676 19159 1728 19168
rect 1676 19125 1685 19159
rect 1685 19125 1719 19159
rect 1719 19125 1728 19159
rect 1676 19116 1728 19125
rect 1952 19159 2004 19168
rect 1952 19125 1961 19159
rect 1961 19125 1995 19159
rect 1995 19125 2004 19159
rect 1952 19116 2004 19125
rect 4068 19184 4120 19236
rect 4896 19227 4948 19236
rect 4896 19193 4905 19227
rect 4905 19193 4939 19227
rect 4939 19193 4948 19227
rect 4896 19184 4948 19193
rect 11336 19184 11388 19236
rect 3884 19159 3936 19168
rect 3884 19125 3893 19159
rect 3893 19125 3927 19159
rect 3927 19125 3936 19159
rect 3884 19116 3936 19125
rect 4988 19159 5040 19168
rect 4988 19125 4997 19159
rect 4997 19125 5031 19159
rect 5031 19125 5040 19159
rect 4988 19116 5040 19125
rect 5448 19159 5500 19168
rect 5448 19125 5457 19159
rect 5457 19125 5491 19159
rect 5491 19125 5500 19159
rect 5448 19116 5500 19125
rect 6828 19159 6880 19168
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 10784 19159 10836 19168
rect 10784 19125 10793 19159
rect 10793 19125 10827 19159
rect 10827 19125 10836 19159
rect 10784 19116 10836 19125
rect 11888 19116 11940 19168
rect 12532 19252 12584 19304
rect 15200 19320 15252 19372
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 17776 19252 17828 19304
rect 18880 19295 18932 19304
rect 18880 19261 18889 19295
rect 18889 19261 18923 19295
rect 18923 19261 18932 19295
rect 18880 19252 18932 19261
rect 26516 19320 26568 19372
rect 17868 19184 17920 19236
rect 14924 19159 14976 19168
rect 14924 19125 14933 19159
rect 14933 19125 14967 19159
rect 14967 19125 14976 19159
rect 14924 19116 14976 19125
rect 15016 19116 15068 19168
rect 15752 19116 15804 19168
rect 18420 19184 18472 19236
rect 19248 19184 19300 19236
rect 20168 19252 20220 19304
rect 22284 19252 22336 19304
rect 20352 19184 20404 19236
rect 20904 19184 20956 19236
rect 18696 19116 18748 19168
rect 19340 19116 19392 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 22100 19116 22152 19168
rect 22560 19116 22612 19168
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 24676 19184 24728 19236
rect 25964 19159 26016 19168
rect 25964 19125 25973 19159
rect 25973 19125 26007 19159
rect 26007 19125 26016 19159
rect 25964 19116 26016 19125
rect 26516 19159 26568 19168
rect 26516 19125 26525 19159
rect 26525 19125 26559 19159
rect 26559 19125 26568 19159
rect 26516 19116 26568 19125
rect 26884 19159 26936 19168
rect 26884 19125 26893 19159
rect 26893 19125 26927 19159
rect 26927 19125 26936 19159
rect 26884 19116 26936 19125
rect 27068 19159 27120 19168
rect 27068 19125 27077 19159
rect 27077 19125 27111 19159
rect 27111 19125 27120 19159
rect 27068 19116 27120 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 2688 18955 2740 18964
rect 2688 18921 2697 18955
rect 2697 18921 2731 18955
rect 2731 18921 2740 18955
rect 2688 18912 2740 18921
rect 4068 18912 4120 18964
rect 4712 18955 4764 18964
rect 4712 18921 4721 18955
rect 4721 18921 4755 18955
rect 4755 18921 4764 18955
rect 4712 18912 4764 18921
rect 6184 18955 6236 18964
rect 6184 18921 6193 18955
rect 6193 18921 6227 18955
rect 6227 18921 6236 18955
rect 6184 18912 6236 18921
rect 7288 18955 7340 18964
rect 7288 18921 7297 18955
rect 7297 18921 7331 18955
rect 7331 18921 7340 18955
rect 7288 18912 7340 18921
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 9864 18955 9916 18964
rect 9864 18921 9873 18955
rect 9873 18921 9907 18955
rect 9907 18921 9916 18955
rect 9864 18912 9916 18921
rect 11336 18912 11388 18964
rect 13820 18912 13872 18964
rect 14280 18912 14332 18964
rect 15292 18912 15344 18964
rect 15844 18912 15896 18964
rect 18880 18955 18932 18964
rect 18880 18921 18889 18955
rect 18889 18921 18923 18955
rect 18923 18921 18932 18955
rect 18880 18912 18932 18921
rect 19156 18912 19208 18964
rect 24768 18955 24820 18964
rect 24768 18921 24777 18955
rect 24777 18921 24811 18955
rect 24811 18921 24820 18955
rect 24768 18912 24820 18921
rect 2872 18844 2924 18896
rect 2044 18819 2096 18828
rect 2044 18785 2053 18819
rect 2053 18785 2087 18819
rect 2087 18785 2096 18819
rect 2044 18776 2096 18785
rect 2504 18819 2556 18828
rect 2504 18785 2513 18819
rect 2513 18785 2547 18819
rect 2547 18785 2556 18819
rect 2504 18776 2556 18785
rect 5540 18844 5592 18896
rect 18788 18844 18840 18896
rect 6460 18776 6512 18828
rect 7656 18819 7708 18828
rect 7656 18785 7665 18819
rect 7665 18785 7699 18819
rect 7699 18785 7708 18819
rect 7656 18776 7708 18785
rect 9680 18819 9732 18828
rect 9680 18785 9689 18819
rect 9689 18785 9723 18819
rect 9723 18785 9732 18819
rect 9680 18776 9732 18785
rect 11428 18819 11480 18828
rect 11428 18785 11462 18819
rect 11462 18785 11480 18819
rect 11428 18776 11480 18785
rect 13912 18776 13964 18828
rect 16764 18819 16816 18828
rect 16764 18785 16798 18819
rect 16798 18785 16816 18819
rect 16764 18776 16816 18785
rect 19064 18776 19116 18828
rect 19432 18819 19484 18828
rect 19432 18785 19441 18819
rect 19441 18785 19475 18819
rect 19475 18785 19484 18819
rect 19432 18776 19484 18785
rect 23112 18776 23164 18828
rect 4804 18751 4856 18760
rect 4804 18717 4813 18751
rect 4813 18717 4847 18751
rect 4847 18717 4856 18751
rect 4804 18708 4856 18717
rect 7840 18751 7892 18760
rect 7840 18717 7849 18751
rect 7849 18717 7883 18751
rect 7883 18717 7892 18751
rect 7840 18708 7892 18717
rect 3240 18640 3292 18692
rect 9036 18640 9088 18692
rect 2228 18572 2280 18624
rect 3884 18572 3936 18624
rect 5448 18572 5500 18624
rect 7012 18572 7064 18624
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 10784 18615 10836 18624
rect 10784 18581 10793 18615
rect 10793 18581 10827 18615
rect 10827 18581 10836 18615
rect 10784 18572 10836 18581
rect 13636 18708 13688 18760
rect 14096 18751 14148 18760
rect 14096 18717 14105 18751
rect 14105 18717 14139 18751
rect 14139 18717 14148 18751
rect 14096 18708 14148 18717
rect 16488 18751 16540 18760
rect 12532 18683 12584 18692
rect 12532 18649 12541 18683
rect 12541 18649 12575 18683
rect 12575 18649 12584 18683
rect 12532 18640 12584 18649
rect 13084 18640 13136 18692
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 18880 18708 18932 18760
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 25228 18751 25280 18760
rect 25228 18717 25237 18751
rect 25237 18717 25271 18751
rect 25271 18717 25280 18751
rect 25228 18708 25280 18717
rect 25412 18751 25464 18760
rect 25412 18717 25421 18751
rect 25421 18717 25455 18751
rect 25455 18717 25464 18751
rect 25412 18708 25464 18717
rect 25964 18708 26016 18760
rect 19984 18683 20036 18692
rect 19984 18649 19993 18683
rect 19993 18649 20027 18683
rect 20027 18649 20036 18683
rect 19984 18640 20036 18649
rect 24584 18640 24636 18692
rect 26332 18776 26384 18828
rect 27068 18844 27120 18896
rect 26976 18819 27028 18828
rect 26976 18785 26985 18819
rect 26985 18785 27019 18819
rect 27019 18785 27028 18819
rect 26976 18776 27028 18785
rect 27068 18751 27120 18760
rect 27068 18717 27077 18751
rect 27077 18717 27111 18751
rect 27111 18717 27120 18751
rect 27068 18708 27120 18717
rect 11888 18572 11940 18624
rect 17868 18615 17920 18624
rect 17868 18581 17877 18615
rect 17877 18581 17911 18615
rect 17911 18581 17920 18615
rect 17868 18572 17920 18581
rect 23388 18572 23440 18624
rect 24676 18615 24728 18624
rect 24676 18581 24685 18615
rect 24685 18581 24719 18615
rect 24719 18581 24728 18615
rect 24676 18572 24728 18581
rect 25780 18615 25832 18624
rect 25780 18581 25789 18615
rect 25789 18581 25823 18615
rect 25823 18581 25832 18615
rect 25780 18572 25832 18581
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 3976 18368 4028 18420
rect 5448 18368 5500 18420
rect 10600 18411 10652 18420
rect 10600 18377 10609 18411
rect 10609 18377 10643 18411
rect 10643 18377 10652 18411
rect 10600 18368 10652 18377
rect 10876 18368 10928 18420
rect 12256 18368 12308 18420
rect 17776 18368 17828 18420
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 19616 18411 19668 18420
rect 19616 18377 19625 18411
rect 19625 18377 19659 18411
rect 19659 18377 19668 18411
rect 19616 18368 19668 18377
rect 23112 18411 23164 18420
rect 23112 18377 23121 18411
rect 23121 18377 23155 18411
rect 23155 18377 23164 18411
rect 23112 18368 23164 18377
rect 25412 18368 25464 18420
rect 27068 18411 27120 18420
rect 7656 18300 7708 18352
rect 8116 18300 8168 18352
rect 16764 18300 16816 18352
rect 1676 18232 1728 18284
rect 2228 18275 2280 18284
rect 1952 18207 2004 18216
rect 1952 18173 1961 18207
rect 1961 18173 1995 18207
rect 1995 18173 2004 18207
rect 1952 18164 2004 18173
rect 2228 18241 2237 18275
rect 2237 18241 2271 18275
rect 2271 18241 2280 18275
rect 2228 18232 2280 18241
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 4160 18232 4212 18284
rect 4344 18232 4396 18284
rect 7288 18232 7340 18284
rect 8668 18232 8720 18284
rect 10876 18232 10928 18284
rect 11428 18275 11480 18284
rect 11428 18241 11437 18275
rect 11437 18241 11471 18275
rect 11471 18241 11480 18275
rect 13084 18275 13136 18284
rect 11428 18232 11480 18241
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 18328 18232 18380 18284
rect 18880 18300 18932 18352
rect 19248 18300 19300 18352
rect 21272 18300 21324 18352
rect 21640 18300 21692 18352
rect 22560 18300 22612 18352
rect 25228 18300 25280 18352
rect 18788 18232 18840 18284
rect 20168 18275 20220 18284
rect 20168 18241 20177 18275
rect 20177 18241 20211 18275
rect 20211 18241 20220 18275
rect 20168 18232 20220 18241
rect 22192 18275 22244 18284
rect 2412 18164 2464 18216
rect 3700 18207 3752 18216
rect 3700 18173 3709 18207
rect 3709 18173 3743 18207
rect 3743 18173 3752 18207
rect 3700 18164 3752 18173
rect 4896 18164 4948 18216
rect 2136 18096 2188 18148
rect 2688 18071 2740 18080
rect 2688 18037 2697 18071
rect 2697 18037 2731 18071
rect 2731 18037 2740 18071
rect 2688 18028 2740 18037
rect 3976 18028 4028 18080
rect 4896 18028 4948 18080
rect 5080 18028 5132 18080
rect 5724 18028 5776 18080
rect 6920 18096 6972 18148
rect 7840 18139 7892 18148
rect 7840 18105 7849 18139
rect 7849 18105 7883 18139
rect 7883 18105 7892 18139
rect 7840 18096 7892 18105
rect 7012 18028 7064 18080
rect 9312 18164 9364 18216
rect 9680 18207 9732 18216
rect 9680 18173 9689 18207
rect 9689 18173 9723 18207
rect 9723 18173 9732 18207
rect 9680 18164 9732 18173
rect 10600 18164 10652 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 14280 18207 14332 18216
rect 14280 18173 14314 18207
rect 14314 18173 14332 18207
rect 8300 18096 8352 18148
rect 8944 18139 8996 18148
rect 8944 18105 8953 18139
rect 8953 18105 8987 18139
rect 8987 18105 8996 18139
rect 8944 18096 8996 18105
rect 11888 18139 11940 18148
rect 11888 18105 11897 18139
rect 11897 18105 11931 18139
rect 11931 18105 11940 18139
rect 11888 18096 11940 18105
rect 12532 18096 12584 18148
rect 14280 18164 14332 18173
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 18696 18164 18748 18216
rect 14648 18096 14700 18148
rect 16488 18139 16540 18148
rect 16488 18105 16497 18139
rect 16497 18105 16531 18139
rect 16531 18105 16540 18139
rect 16488 18096 16540 18105
rect 19064 18139 19116 18148
rect 19064 18105 19073 18139
rect 19073 18105 19107 18139
rect 19107 18105 19116 18139
rect 19064 18096 19116 18105
rect 19616 18096 19668 18148
rect 22192 18241 22201 18275
rect 22201 18241 22235 18275
rect 22235 18241 22244 18275
rect 22192 18232 22244 18241
rect 22376 18275 22428 18284
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 24676 18232 24728 18284
rect 27068 18377 27077 18411
rect 27077 18377 27111 18411
rect 27111 18377 27120 18411
rect 27068 18368 27120 18377
rect 22284 18164 22336 18216
rect 21640 18139 21692 18148
rect 21640 18105 21649 18139
rect 21649 18105 21683 18139
rect 21683 18105 21692 18139
rect 21640 18096 21692 18105
rect 25780 18164 25832 18216
rect 26516 18164 26568 18216
rect 27160 18164 27212 18216
rect 26976 18096 27028 18148
rect 8668 18028 8720 18080
rect 9036 18071 9088 18080
rect 9036 18037 9045 18071
rect 9045 18037 9079 18071
rect 9079 18037 9088 18071
rect 9036 18028 9088 18037
rect 9588 18028 9640 18080
rect 10048 18028 10100 18080
rect 10784 18028 10836 18080
rect 11336 18028 11388 18080
rect 12992 18028 13044 18080
rect 13636 18071 13688 18080
rect 13636 18037 13645 18071
rect 13645 18037 13679 18071
rect 13679 18037 13688 18071
rect 13636 18028 13688 18037
rect 15476 18028 15528 18080
rect 19984 18028 20036 18080
rect 21548 18028 21600 18080
rect 24492 18071 24544 18080
rect 24492 18037 24501 18071
rect 24501 18037 24535 18071
rect 24535 18037 24544 18071
rect 24492 18028 24544 18037
rect 24584 18071 24636 18080
rect 24584 18037 24593 18071
rect 24593 18037 24627 18071
rect 24627 18037 24636 18071
rect 25504 18071 25556 18080
rect 24584 18028 24636 18037
rect 25504 18037 25513 18071
rect 25513 18037 25547 18071
rect 25547 18037 25556 18071
rect 25504 18028 25556 18037
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 2504 17824 2556 17876
rect 2688 17867 2740 17876
rect 2688 17833 2697 17867
rect 2697 17833 2731 17867
rect 2731 17833 2740 17867
rect 2688 17824 2740 17833
rect 3700 17824 3752 17876
rect 4344 17867 4396 17876
rect 4344 17833 4353 17867
rect 4353 17833 4387 17867
rect 4387 17833 4396 17867
rect 4344 17824 4396 17833
rect 4804 17867 4856 17876
rect 4804 17833 4813 17867
rect 4813 17833 4847 17867
rect 4847 17833 4856 17867
rect 4804 17824 4856 17833
rect 5540 17824 5592 17876
rect 6828 17824 6880 17876
rect 7656 17867 7708 17876
rect 7656 17833 7665 17867
rect 7665 17833 7699 17867
rect 7699 17833 7708 17867
rect 7656 17824 7708 17833
rect 10876 17867 10928 17876
rect 10876 17833 10885 17867
rect 10885 17833 10919 17867
rect 10919 17833 10928 17867
rect 10876 17824 10928 17833
rect 13084 17824 13136 17876
rect 13728 17824 13780 17876
rect 14280 17824 14332 17876
rect 14924 17824 14976 17876
rect 15200 17824 15252 17876
rect 17592 17824 17644 17876
rect 18972 17824 19024 17876
rect 20168 17867 20220 17876
rect 20168 17833 20177 17867
rect 20177 17833 20211 17867
rect 20211 17833 20220 17867
rect 20168 17824 20220 17833
rect 21916 17824 21968 17876
rect 22376 17867 22428 17876
rect 22376 17833 22385 17867
rect 22385 17833 22419 17867
rect 22419 17833 22428 17867
rect 22376 17824 22428 17833
rect 25228 17867 25280 17876
rect 25228 17833 25237 17867
rect 25237 17833 25271 17867
rect 25271 17833 25280 17867
rect 25228 17824 25280 17833
rect 25412 17824 25464 17876
rect 26332 17867 26384 17876
rect 26332 17833 26341 17867
rect 26341 17833 26375 17867
rect 26375 17833 26384 17867
rect 26332 17824 26384 17833
rect 26976 17824 27028 17876
rect 4160 17756 4212 17808
rect 5264 17799 5316 17808
rect 5264 17765 5276 17799
rect 5276 17765 5316 17799
rect 5264 17756 5316 17765
rect 7288 17756 7340 17808
rect 7748 17756 7800 17808
rect 13912 17756 13964 17808
rect 14648 17799 14700 17808
rect 14648 17765 14657 17799
rect 14657 17765 14691 17799
rect 14691 17765 14700 17799
rect 14648 17756 14700 17765
rect 21456 17799 21508 17808
rect 21456 17765 21465 17799
rect 21465 17765 21499 17799
rect 21499 17765 21508 17799
rect 21456 17756 21508 17765
rect 2136 17663 2188 17672
rect 2136 17629 2145 17663
rect 2145 17629 2179 17663
rect 2179 17629 2188 17663
rect 2136 17620 2188 17629
rect 2320 17663 2372 17672
rect 2320 17629 2329 17663
rect 2329 17629 2363 17663
rect 2363 17629 2372 17663
rect 2320 17620 2372 17629
rect 2688 17620 2740 17672
rect 4804 17688 4856 17740
rect 8300 17688 8352 17740
rect 12072 17688 12124 17740
rect 13820 17688 13872 17740
rect 16488 17688 16540 17740
rect 16948 17731 17000 17740
rect 16948 17697 16982 17731
rect 16982 17697 17000 17731
rect 16948 17688 17000 17697
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 21364 17731 21416 17740
rect 21364 17697 21373 17731
rect 21373 17697 21407 17731
rect 21407 17697 21416 17731
rect 21364 17688 21416 17697
rect 8484 17663 8536 17672
rect 8484 17629 8493 17663
rect 8493 17629 8527 17663
rect 8527 17629 8536 17663
rect 8484 17620 8536 17629
rect 8668 17663 8720 17672
rect 8668 17629 8677 17663
rect 8677 17629 8711 17663
rect 8711 17629 8720 17663
rect 8668 17620 8720 17629
rect 11612 17620 11664 17672
rect 10600 17552 10652 17604
rect 12164 17620 12216 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 18604 17620 18656 17672
rect 19064 17552 19116 17604
rect 21088 17620 21140 17672
rect 22560 17731 22612 17740
rect 22560 17697 22569 17731
rect 22569 17697 22603 17731
rect 22603 17697 22612 17731
rect 22560 17688 22612 17697
rect 23388 17688 23440 17740
rect 26884 17731 26936 17740
rect 26884 17697 26893 17731
rect 26893 17697 26927 17731
rect 26927 17697 26936 17731
rect 26884 17688 26936 17697
rect 26792 17620 26844 17672
rect 27160 17663 27212 17672
rect 27160 17629 27169 17663
rect 27169 17629 27203 17663
rect 27203 17629 27212 17663
rect 27160 17620 27212 17629
rect 24768 17552 24820 17604
rect 4068 17484 4120 17536
rect 7840 17484 7892 17536
rect 9956 17527 10008 17536
rect 9956 17493 9965 17527
rect 9965 17493 9999 17527
rect 9999 17493 10008 17527
rect 9956 17484 10008 17493
rect 11428 17527 11480 17536
rect 11428 17493 11437 17527
rect 11437 17493 11471 17527
rect 11471 17493 11480 17527
rect 11428 17484 11480 17493
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 18788 17527 18840 17536
rect 18788 17493 18797 17527
rect 18797 17493 18831 17527
rect 18831 17493 18840 17527
rect 18788 17484 18840 17493
rect 22284 17484 22336 17536
rect 23848 17484 23900 17536
rect 24860 17527 24912 17536
rect 24860 17493 24869 17527
rect 24869 17493 24903 17527
rect 24903 17493 24912 17527
rect 24860 17484 24912 17493
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2136 17280 2188 17332
rect 5264 17280 5316 17332
rect 7932 17280 7984 17332
rect 10600 17323 10652 17332
rect 8116 17212 8168 17264
rect 2320 17076 2372 17128
rect 4344 17076 4396 17128
rect 7840 17076 7892 17128
rect 10600 17289 10609 17323
rect 10609 17289 10643 17323
rect 10643 17289 10652 17323
rect 10600 17280 10652 17289
rect 11980 17280 12032 17332
rect 12440 17323 12492 17332
rect 12440 17289 12449 17323
rect 12449 17289 12483 17323
rect 12483 17289 12492 17323
rect 12440 17280 12492 17289
rect 13084 17280 13136 17332
rect 14188 17280 14240 17332
rect 16948 17280 17000 17332
rect 17592 17280 17644 17332
rect 20168 17323 20220 17332
rect 9128 17144 9180 17196
rect 4804 17008 4856 17060
rect 8484 17008 8536 17060
rect 11428 17144 11480 17196
rect 14648 17212 14700 17264
rect 11980 17008 12032 17060
rect 15108 17187 15160 17196
rect 15108 17153 15117 17187
rect 15117 17153 15151 17187
rect 15151 17153 15160 17187
rect 15108 17144 15160 17153
rect 16488 17144 16540 17196
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 21088 17323 21140 17332
rect 21088 17289 21097 17323
rect 21097 17289 21131 17323
rect 21131 17289 21140 17323
rect 21088 17280 21140 17289
rect 22560 17280 22612 17332
rect 23204 17280 23256 17332
rect 23388 17323 23440 17332
rect 23388 17289 23397 17323
rect 23397 17289 23431 17323
rect 23431 17289 23440 17323
rect 23388 17280 23440 17289
rect 23940 17323 23992 17332
rect 23940 17289 23949 17323
rect 23949 17289 23983 17323
rect 23983 17289 23992 17323
rect 23940 17280 23992 17289
rect 24492 17280 24544 17332
rect 24860 17280 24912 17332
rect 26792 17280 26844 17332
rect 25504 17255 25556 17264
rect 25504 17221 25513 17255
rect 25513 17221 25547 17255
rect 25547 17221 25556 17255
rect 25504 17212 25556 17221
rect 26884 17212 26936 17264
rect 18788 17119 18840 17128
rect 18788 17085 18797 17119
rect 18797 17085 18831 17119
rect 18831 17085 18840 17119
rect 18788 17076 18840 17085
rect 23020 17144 23072 17196
rect 24768 17187 24820 17196
rect 24768 17153 24777 17187
rect 24777 17153 24811 17187
rect 24811 17153 24820 17187
rect 24768 17144 24820 17153
rect 25688 17187 25740 17196
rect 25688 17153 25697 17187
rect 25697 17153 25731 17187
rect 25731 17153 25740 17187
rect 25688 17144 25740 17153
rect 27988 17144 28040 17196
rect 19064 17119 19116 17128
rect 19064 17085 19087 17119
rect 19087 17085 19116 17119
rect 19064 17076 19116 17085
rect 23940 17076 23992 17128
rect 16672 17008 16724 17060
rect 22468 17051 22520 17060
rect 1676 16983 1728 16992
rect 1676 16949 1685 16983
rect 1685 16949 1719 16983
rect 1719 16949 1728 16983
rect 1676 16940 1728 16949
rect 7932 16940 7984 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 11612 16940 11664 16992
rect 12072 16940 12124 16992
rect 12716 16940 12768 16992
rect 14556 16983 14608 16992
rect 14556 16949 14565 16983
rect 14565 16949 14599 16983
rect 14599 16949 14608 16983
rect 14556 16940 14608 16949
rect 18604 16983 18656 16992
rect 18604 16949 18613 16983
rect 18613 16949 18647 16983
rect 18647 16949 18656 16983
rect 18604 16940 18656 16949
rect 20812 16940 20864 16992
rect 22468 17017 22477 17051
rect 22477 17017 22511 17051
rect 22511 17017 22520 17051
rect 22468 17008 22520 17017
rect 25412 17008 25464 17060
rect 22008 16983 22060 16992
rect 22008 16949 22017 16983
rect 22017 16949 22051 16983
rect 22051 16949 22060 16983
rect 22008 16940 22060 16949
rect 22284 16940 22336 16992
rect 24584 16983 24636 16992
rect 24584 16949 24593 16983
rect 24593 16949 24627 16983
rect 24627 16949 24636 16983
rect 24584 16940 24636 16949
rect 26424 16940 26476 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16736 1728 16788
rect 2320 16736 2372 16788
rect 4804 16736 4856 16788
rect 7932 16779 7984 16788
rect 2228 16668 2280 16720
rect 3056 16668 3108 16720
rect 7932 16745 7941 16779
rect 7941 16745 7975 16779
rect 7975 16745 7984 16779
rect 7932 16736 7984 16745
rect 8484 16736 8536 16788
rect 9128 16736 9180 16788
rect 9680 16779 9732 16788
rect 5356 16668 5408 16720
rect 8116 16668 8168 16720
rect 8300 16668 8352 16720
rect 9680 16745 9689 16779
rect 9689 16745 9723 16779
rect 9723 16745 9732 16779
rect 9680 16736 9732 16745
rect 9956 16736 10008 16788
rect 13084 16736 13136 16788
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 13912 16736 13964 16788
rect 14280 16779 14332 16788
rect 14280 16745 14289 16779
rect 14289 16745 14323 16779
rect 14323 16745 14332 16779
rect 14280 16736 14332 16745
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 18512 16779 18564 16788
rect 18512 16745 18521 16779
rect 18521 16745 18555 16779
rect 18555 16745 18564 16779
rect 18512 16736 18564 16745
rect 21456 16736 21508 16788
rect 22560 16779 22612 16788
rect 22560 16745 22569 16779
rect 22569 16745 22603 16779
rect 22603 16745 22612 16779
rect 22560 16736 22612 16745
rect 23112 16736 23164 16788
rect 24768 16736 24820 16788
rect 25872 16779 25924 16788
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 9588 16668 9640 16720
rect 10324 16668 10376 16720
rect 10784 16643 10836 16652
rect 3516 16532 3568 16584
rect 8116 16532 8168 16584
rect 8852 16532 8904 16584
rect 10784 16609 10793 16643
rect 10793 16609 10827 16643
rect 10827 16609 10836 16643
rect 10784 16600 10836 16609
rect 11888 16668 11940 16720
rect 15844 16668 15896 16720
rect 18972 16711 19024 16720
rect 12164 16600 12216 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 18972 16677 18981 16711
rect 18981 16677 19015 16711
rect 19015 16677 19024 16711
rect 18972 16668 19024 16677
rect 25872 16745 25881 16779
rect 25881 16745 25915 16779
rect 25915 16745 25924 16779
rect 25872 16736 25924 16745
rect 18880 16643 18932 16652
rect 9864 16532 9916 16584
rect 3608 16396 3660 16448
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 6276 16396 6328 16448
rect 15108 16532 15160 16584
rect 17776 16532 17828 16584
rect 18880 16609 18889 16643
rect 18889 16609 18923 16643
rect 18923 16609 18932 16643
rect 18880 16600 18932 16609
rect 19524 16643 19576 16652
rect 19524 16609 19533 16643
rect 19533 16609 19567 16643
rect 19567 16609 19576 16643
rect 19524 16600 19576 16609
rect 21180 16643 21232 16652
rect 21180 16609 21189 16643
rect 21189 16609 21223 16643
rect 21223 16609 21232 16643
rect 21180 16600 21232 16609
rect 21272 16600 21324 16652
rect 22376 16600 22428 16652
rect 23112 16600 23164 16652
rect 23848 16600 23900 16652
rect 19064 16575 19116 16584
rect 19064 16541 19073 16575
rect 19073 16541 19107 16575
rect 19107 16541 19116 16575
rect 19064 16532 19116 16541
rect 23204 16532 23256 16584
rect 23756 16532 23808 16584
rect 25412 16532 25464 16584
rect 11428 16396 11480 16448
rect 18144 16439 18196 16448
rect 18144 16405 18153 16439
rect 18153 16405 18187 16439
rect 18187 16405 18196 16439
rect 18144 16396 18196 16405
rect 26516 16600 26568 16652
rect 26884 16643 26936 16652
rect 26884 16609 26893 16643
rect 26893 16609 26927 16643
rect 26927 16609 26936 16643
rect 26884 16600 26936 16609
rect 27160 16575 27212 16584
rect 27160 16541 27169 16575
rect 27169 16541 27203 16575
rect 27203 16541 27212 16575
rect 27160 16532 27212 16541
rect 27160 16396 27212 16448
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 3056 16235 3108 16244
rect 3056 16201 3065 16235
rect 3065 16201 3099 16235
rect 3099 16201 3108 16235
rect 3056 16192 3108 16201
rect 4160 16235 4212 16244
rect 3608 16167 3660 16176
rect 3608 16133 3617 16167
rect 3617 16133 3651 16167
rect 3651 16133 3660 16167
rect 3608 16124 3660 16133
rect 4160 16201 4169 16235
rect 4169 16201 4203 16235
rect 4203 16201 4212 16235
rect 4160 16192 4212 16201
rect 5172 16235 5224 16244
rect 5172 16201 5181 16235
rect 5181 16201 5215 16235
rect 5215 16201 5224 16235
rect 5172 16192 5224 16201
rect 5540 16235 5592 16244
rect 5540 16201 5549 16235
rect 5549 16201 5583 16235
rect 5583 16201 5592 16235
rect 5540 16192 5592 16201
rect 7380 16192 7432 16244
rect 8116 16235 8168 16244
rect 8116 16201 8125 16235
rect 8125 16201 8159 16235
rect 8159 16201 8168 16235
rect 8116 16192 8168 16201
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 9864 16192 9916 16244
rect 12164 16235 12216 16244
rect 12164 16201 12173 16235
rect 12173 16201 12207 16235
rect 12207 16201 12216 16235
rect 12164 16192 12216 16201
rect 15016 16235 15068 16244
rect 15016 16201 15025 16235
rect 15025 16201 15059 16235
rect 15059 16201 15068 16235
rect 15016 16192 15068 16201
rect 17592 16192 17644 16244
rect 19984 16235 20036 16244
rect 19984 16201 19993 16235
rect 19993 16201 20027 16235
rect 20027 16201 20036 16235
rect 19984 16192 20036 16201
rect 21180 16235 21232 16244
rect 21180 16201 21189 16235
rect 21189 16201 21223 16235
rect 21223 16201 21232 16235
rect 21180 16192 21232 16201
rect 21364 16192 21416 16244
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 23204 16192 23256 16244
rect 24400 16235 24452 16244
rect 24400 16201 24409 16235
rect 24409 16201 24443 16235
rect 24443 16201 24452 16235
rect 24400 16192 24452 16201
rect 24584 16235 24636 16244
rect 24584 16201 24593 16235
rect 24593 16201 24627 16235
rect 24627 16201 24636 16235
rect 24584 16192 24636 16201
rect 25688 16192 25740 16244
rect 13912 16124 13964 16176
rect 15108 16124 15160 16176
rect 21272 16124 21324 16176
rect 7288 16099 7340 16108
rect 7288 16065 7297 16099
rect 7297 16065 7331 16099
rect 7331 16065 7340 16099
rect 7288 16056 7340 16065
rect 11428 16099 11480 16108
rect 11428 16065 11437 16099
rect 11437 16065 11471 16099
rect 11471 16065 11480 16099
rect 11428 16056 11480 16065
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 8300 16031 8352 16040
rect 8300 15997 8309 16031
rect 8309 15997 8343 16031
rect 8343 15997 8352 16031
rect 8300 15988 8352 15997
rect 11152 16031 11204 16040
rect 11152 15997 11161 16031
rect 11161 15997 11195 16031
rect 11195 15997 11204 16031
rect 11152 15988 11204 15997
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 14740 16056 14792 16108
rect 15844 16056 15896 16108
rect 18052 16099 18104 16108
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22560 16099 22612 16108
rect 22008 16056 22060 16065
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 25412 16056 25464 16108
rect 27160 16192 27212 16244
rect 15476 15988 15528 16040
rect 18144 15988 18196 16040
rect 21548 15988 21600 16040
rect 23572 15988 23624 16040
rect 24952 16031 25004 16040
rect 24952 15997 24961 16031
rect 24961 15997 24995 16031
rect 24995 15997 25004 16031
rect 24952 15988 25004 15997
rect 2688 15920 2740 15972
rect 4528 15963 4580 15972
rect 4528 15929 4537 15963
rect 4537 15929 4571 15963
rect 4571 15929 4580 15963
rect 4528 15920 4580 15929
rect 8668 15920 8720 15972
rect 9496 15920 9548 15972
rect 26424 15963 26476 15972
rect 26424 15929 26458 15963
rect 26458 15929 26476 15963
rect 26424 15920 26476 15929
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 8852 15852 8904 15904
rect 10324 15895 10376 15904
rect 10324 15861 10333 15895
rect 10333 15861 10367 15895
rect 10367 15861 10376 15895
rect 10324 15852 10376 15861
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 11520 15852 11572 15904
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 11888 15852 11940 15861
rect 13360 15895 13412 15904
rect 13360 15861 13369 15895
rect 13369 15861 13403 15895
rect 13403 15861 13412 15895
rect 13360 15852 13412 15861
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 15568 15852 15620 15904
rect 17776 15895 17828 15904
rect 17776 15861 17785 15895
rect 17785 15861 17819 15895
rect 17819 15861 17828 15895
rect 17776 15852 17828 15861
rect 18604 15852 18656 15904
rect 22192 15852 22244 15904
rect 25412 15852 25464 15904
rect 27252 15852 27304 15904
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 2044 15691 2096 15700
rect 2044 15657 2053 15691
rect 2053 15657 2087 15691
rect 2087 15657 2096 15691
rect 2044 15648 2096 15657
rect 3516 15691 3568 15700
rect 3516 15657 3525 15691
rect 3525 15657 3559 15691
rect 3559 15657 3568 15691
rect 3516 15648 3568 15657
rect 3608 15648 3660 15700
rect 5816 15648 5868 15700
rect 8208 15648 8260 15700
rect 8392 15691 8444 15700
rect 8392 15657 8401 15691
rect 8401 15657 8435 15691
rect 8435 15657 8444 15691
rect 8392 15648 8444 15657
rect 9956 15648 10008 15700
rect 10876 15648 10928 15700
rect 11428 15648 11480 15700
rect 14740 15691 14792 15700
rect 14740 15657 14749 15691
rect 14749 15657 14783 15691
rect 14783 15657 14792 15691
rect 14740 15648 14792 15657
rect 15844 15648 15896 15700
rect 18052 15691 18104 15700
rect 18052 15657 18061 15691
rect 18061 15657 18095 15691
rect 18095 15657 18104 15691
rect 18052 15648 18104 15657
rect 21456 15648 21508 15700
rect 22192 15691 22244 15700
rect 22192 15657 22201 15691
rect 22201 15657 22235 15691
rect 22235 15657 22244 15691
rect 22192 15648 22244 15657
rect 23204 15691 23256 15700
rect 23204 15657 23213 15691
rect 23213 15657 23247 15691
rect 23247 15657 23256 15691
rect 23204 15648 23256 15657
rect 23480 15648 23532 15700
rect 23756 15648 23808 15700
rect 26884 15648 26936 15700
rect 5264 15580 5316 15632
rect 4712 15512 4764 15564
rect 5172 15512 5224 15564
rect 5448 15512 5500 15564
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 2688 15487 2740 15496
rect 2688 15453 2697 15487
rect 2697 15453 2731 15487
rect 2731 15453 2740 15487
rect 2688 15444 2740 15453
rect 1676 15351 1728 15360
rect 1676 15317 1685 15351
rect 1685 15317 1719 15351
rect 1719 15317 1728 15351
rect 1676 15308 1728 15317
rect 3056 15308 3108 15360
rect 8576 15444 8628 15496
rect 15476 15580 15528 15632
rect 8392 15376 8444 15428
rect 10416 15444 10468 15496
rect 12532 15512 12584 15564
rect 15108 15512 15160 15564
rect 20720 15623 20772 15632
rect 20720 15589 20729 15623
rect 20729 15589 20763 15623
rect 20763 15589 20772 15623
rect 20720 15580 20772 15589
rect 24768 15623 24820 15632
rect 24768 15589 24777 15623
rect 24777 15589 24811 15623
rect 24811 15589 24820 15623
rect 24768 15580 24820 15589
rect 25872 15580 25924 15632
rect 18420 15512 18472 15564
rect 18604 15555 18656 15564
rect 18604 15521 18638 15555
rect 18638 15521 18656 15555
rect 18604 15512 18656 15521
rect 21548 15555 21600 15564
rect 21548 15521 21557 15555
rect 21557 15521 21591 15555
rect 21591 15521 21600 15555
rect 21548 15512 21600 15521
rect 23112 15555 23164 15564
rect 23112 15521 23121 15555
rect 23121 15521 23155 15555
rect 23155 15521 23164 15555
rect 23112 15512 23164 15521
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 21732 15487 21784 15496
rect 21732 15453 21741 15487
rect 21741 15453 21775 15487
rect 21775 15453 21784 15487
rect 21732 15444 21784 15453
rect 22008 15444 22060 15496
rect 22376 15376 22428 15428
rect 24584 15444 24636 15496
rect 26608 15512 26660 15564
rect 26884 15555 26936 15564
rect 26884 15521 26893 15555
rect 26893 15521 26927 15555
rect 26927 15521 26936 15555
rect 26884 15512 26936 15521
rect 25412 15487 25464 15496
rect 25412 15453 25421 15487
rect 25421 15453 25455 15487
rect 25455 15453 25464 15487
rect 26976 15487 27028 15496
rect 25412 15444 25464 15453
rect 26976 15453 26985 15487
rect 26985 15453 27019 15487
rect 27019 15453 27028 15487
rect 26976 15444 27028 15453
rect 24492 15376 24544 15428
rect 26424 15376 26476 15428
rect 27528 15444 27580 15496
rect 4344 15308 4396 15360
rect 4620 15351 4672 15360
rect 4620 15317 4629 15351
rect 4629 15317 4663 15351
rect 4663 15317 4672 15351
rect 4620 15308 4672 15317
rect 5264 15351 5316 15360
rect 5264 15317 5273 15351
rect 5273 15317 5307 15351
rect 5307 15317 5316 15351
rect 5264 15308 5316 15317
rect 8300 15308 8352 15360
rect 9036 15351 9088 15360
rect 9036 15317 9045 15351
rect 9045 15317 9079 15351
rect 9079 15317 9088 15351
rect 9036 15308 9088 15317
rect 11428 15351 11480 15360
rect 11428 15317 11437 15351
rect 11437 15317 11471 15351
rect 11471 15317 11480 15351
rect 11428 15308 11480 15317
rect 12256 15308 12308 15360
rect 13820 15351 13872 15360
rect 13820 15317 13829 15351
rect 13829 15317 13863 15351
rect 13863 15317 13872 15351
rect 13820 15308 13872 15317
rect 14372 15308 14424 15360
rect 15568 15308 15620 15360
rect 19708 15351 19760 15360
rect 19708 15317 19717 15351
rect 19717 15317 19751 15351
rect 19751 15317 19760 15351
rect 19708 15308 19760 15317
rect 27160 15308 27212 15360
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 2044 15147 2096 15156
rect 2044 15113 2053 15147
rect 2053 15113 2087 15147
rect 2087 15113 2096 15147
rect 2044 15104 2096 15113
rect 2412 15104 2464 15156
rect 7932 15147 7984 15156
rect 7932 15113 7941 15147
rect 7941 15113 7975 15147
rect 7975 15113 7984 15147
rect 7932 15104 7984 15113
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 12532 15104 12584 15156
rect 13728 15104 13780 15156
rect 18420 15147 18472 15156
rect 18420 15113 18429 15147
rect 18429 15113 18463 15147
rect 18463 15113 18472 15147
rect 18420 15104 18472 15113
rect 20628 15104 20680 15156
rect 13820 15036 13872 15088
rect 14740 15036 14792 15088
rect 16028 15079 16080 15088
rect 16028 15045 16037 15079
rect 16037 15045 16071 15079
rect 16071 15045 16080 15079
rect 16028 15036 16080 15045
rect 21272 15104 21324 15156
rect 22376 15104 22428 15156
rect 23480 15147 23532 15156
rect 23480 15113 23489 15147
rect 23489 15113 23523 15147
rect 23523 15113 23532 15147
rect 23480 15104 23532 15113
rect 24584 15104 24636 15156
rect 27620 15104 27672 15156
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 3608 14968 3660 15020
rect 5264 14968 5316 15020
rect 6276 14968 6328 15020
rect 10416 15011 10468 15020
rect 10416 14977 10425 15011
rect 10425 14977 10459 15011
rect 10459 14977 10468 15011
rect 10416 14968 10468 14977
rect 11336 15011 11388 15020
rect 11336 14977 11345 15011
rect 11345 14977 11379 15011
rect 11379 14977 11388 15011
rect 11336 14968 11388 14977
rect 13728 15011 13780 15020
rect 13728 14977 13737 15011
rect 13737 14977 13771 15011
rect 13771 14977 13780 15011
rect 13728 14968 13780 14977
rect 13912 14968 13964 15020
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 15476 14968 15528 15020
rect 20628 14968 20680 15020
rect 26884 15036 26936 15088
rect 27712 15079 27764 15088
rect 27712 15045 27721 15079
rect 27721 15045 27755 15079
rect 27755 15045 27764 15079
rect 27712 15036 27764 15045
rect 23756 14968 23808 15020
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 2504 14900 2556 14952
rect 4620 14900 4672 14952
rect 5632 14943 5684 14952
rect 3516 14875 3568 14884
rect 3516 14841 3525 14875
rect 3525 14841 3559 14875
rect 3559 14841 3568 14875
rect 3516 14832 3568 14841
rect 5632 14909 5641 14943
rect 5641 14909 5675 14943
rect 5675 14909 5684 14943
rect 5632 14900 5684 14909
rect 8208 14900 8260 14952
rect 8392 14943 8444 14952
rect 8392 14909 8426 14943
rect 8426 14909 8444 14943
rect 8392 14900 8444 14909
rect 12256 14900 12308 14952
rect 13820 14900 13872 14952
rect 16028 14900 16080 14952
rect 16948 14900 17000 14952
rect 26792 14900 26844 14952
rect 27160 14943 27212 14952
rect 27160 14909 27169 14943
rect 27169 14909 27203 14943
rect 27203 14909 27212 14943
rect 27160 14900 27212 14909
rect 5264 14832 5316 14884
rect 8484 14832 8536 14884
rect 11520 14832 11572 14884
rect 11888 14875 11940 14884
rect 11888 14841 11897 14875
rect 11897 14841 11931 14875
rect 11931 14841 11940 14875
rect 11888 14832 11940 14841
rect 13728 14832 13780 14884
rect 14556 14832 14608 14884
rect 16580 14875 16632 14884
rect 16580 14841 16589 14875
rect 16589 14841 16623 14875
rect 16623 14841 16632 14875
rect 16580 14832 16632 14841
rect 18144 14832 18196 14884
rect 18604 14832 18656 14884
rect 2412 14807 2464 14816
rect 2412 14773 2421 14807
rect 2421 14773 2455 14807
rect 2455 14773 2464 14807
rect 2412 14764 2464 14773
rect 2964 14764 3016 14816
rect 4712 14807 4764 14816
rect 4712 14773 4721 14807
rect 4721 14773 4755 14807
rect 4755 14773 4764 14807
rect 4712 14764 4764 14773
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 5632 14764 5684 14816
rect 6736 14764 6788 14816
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 11428 14764 11480 14816
rect 11796 14764 11848 14816
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 13544 14764 13596 14773
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 15016 14807 15068 14816
rect 14464 14764 14516 14773
rect 15016 14773 15025 14807
rect 15025 14773 15059 14807
rect 15059 14773 15068 14807
rect 15016 14764 15068 14773
rect 15660 14807 15712 14816
rect 15660 14773 15669 14807
rect 15669 14773 15703 14807
rect 15703 14773 15712 14807
rect 15660 14764 15712 14773
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 19892 14807 19944 14816
rect 19892 14773 19901 14807
rect 19901 14773 19935 14807
rect 19935 14773 19944 14807
rect 19892 14764 19944 14773
rect 20076 14764 20128 14816
rect 20444 14764 20496 14816
rect 24492 14875 24544 14884
rect 24492 14841 24526 14875
rect 24526 14841 24544 14875
rect 24492 14832 24544 14841
rect 26976 14832 27028 14884
rect 23112 14807 23164 14816
rect 23112 14773 23121 14807
rect 23121 14773 23155 14807
rect 23155 14773 23164 14807
rect 23112 14764 23164 14773
rect 25596 14807 25648 14816
rect 25596 14773 25605 14807
rect 25605 14773 25639 14807
rect 25639 14773 25648 14807
rect 25596 14764 25648 14773
rect 26700 14807 26752 14816
rect 26700 14773 26709 14807
rect 26709 14773 26743 14807
rect 26743 14773 26752 14807
rect 26700 14764 26752 14773
rect 26792 14764 26844 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 1860 14603 1912 14612
rect 1860 14569 1869 14603
rect 1869 14569 1903 14603
rect 1903 14569 1912 14603
rect 1860 14560 1912 14569
rect 3056 14560 3108 14612
rect 3608 14603 3660 14612
rect 3608 14569 3617 14603
rect 3617 14569 3651 14603
rect 3651 14569 3660 14603
rect 3608 14560 3660 14569
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 8392 14560 8444 14612
rect 8944 14560 8996 14612
rect 10784 14560 10836 14612
rect 12532 14560 12584 14612
rect 13544 14560 13596 14612
rect 16212 14560 16264 14612
rect 21548 14560 21600 14612
rect 26332 14560 26384 14612
rect 11152 14492 11204 14544
rect 13912 14492 13964 14544
rect 14464 14492 14516 14544
rect 15476 14492 15528 14544
rect 15844 14492 15896 14544
rect 17408 14535 17460 14544
rect 17408 14501 17442 14535
rect 17442 14501 17460 14535
rect 17408 14492 17460 14501
rect 21732 14492 21784 14544
rect 24584 14492 24636 14544
rect 25596 14492 25648 14544
rect 756 14424 808 14476
rect 2044 14424 2096 14476
rect 4068 14467 4120 14476
rect 4068 14433 4077 14467
rect 4077 14433 4111 14467
rect 4111 14433 4120 14467
rect 4068 14424 4120 14433
rect 5448 14424 5500 14476
rect 5632 14424 5684 14476
rect 5816 14467 5868 14476
rect 5816 14433 5850 14467
rect 5850 14433 5868 14467
rect 5816 14424 5868 14433
rect 8300 14424 8352 14476
rect 10876 14467 10928 14476
rect 10876 14433 10885 14467
rect 10885 14433 10919 14467
rect 10919 14433 10928 14467
rect 10876 14424 10928 14433
rect 11428 14424 11480 14476
rect 15108 14467 15160 14476
rect 15108 14433 15117 14467
rect 15117 14433 15151 14467
rect 15151 14433 15160 14467
rect 15108 14424 15160 14433
rect 20904 14424 20956 14476
rect 23756 14424 23808 14476
rect 26884 14467 26936 14476
rect 26884 14433 26893 14467
rect 26893 14433 26927 14467
rect 26927 14433 26936 14467
rect 26884 14424 26936 14433
rect 1492 14220 1544 14272
rect 2688 14356 2740 14408
rect 2964 14399 3016 14408
rect 2964 14365 2973 14399
rect 2973 14365 3007 14399
rect 3007 14365 3016 14399
rect 2964 14356 3016 14365
rect 4712 14356 4764 14408
rect 8668 14399 8720 14408
rect 8668 14365 8677 14399
rect 8677 14365 8711 14399
rect 8711 14365 8720 14399
rect 8668 14356 8720 14365
rect 9680 14356 9732 14408
rect 10232 14399 10284 14408
rect 5264 14288 5316 14340
rect 9772 14331 9824 14340
rect 9772 14297 9781 14331
rect 9781 14297 9815 14331
rect 9815 14297 9824 14331
rect 9772 14288 9824 14297
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 13728 14356 13780 14408
rect 15200 14356 15252 14408
rect 15752 14356 15804 14408
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 21732 14399 21784 14408
rect 21732 14365 21741 14399
rect 21741 14365 21775 14399
rect 21775 14365 21784 14399
rect 21732 14356 21784 14365
rect 11152 14288 11204 14340
rect 19340 14288 19392 14340
rect 19892 14331 19944 14340
rect 19892 14297 19901 14331
rect 19901 14297 19935 14331
rect 19935 14297 19944 14331
rect 19892 14288 19944 14297
rect 20628 14288 20680 14340
rect 22376 14356 22428 14408
rect 22928 14399 22980 14408
rect 22928 14365 22937 14399
rect 22937 14365 22971 14399
rect 22971 14365 22980 14399
rect 22928 14356 22980 14365
rect 26700 14356 26752 14408
rect 2320 14220 2372 14272
rect 3056 14220 3108 14272
rect 4160 14220 4212 14272
rect 4804 14263 4856 14272
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 6920 14263 6972 14272
rect 6920 14229 6929 14263
rect 6929 14229 6963 14263
rect 6963 14229 6972 14263
rect 6920 14220 6972 14229
rect 8024 14263 8076 14272
rect 8024 14229 8033 14263
rect 8033 14229 8067 14263
rect 8067 14229 8076 14263
rect 8024 14220 8076 14229
rect 9956 14220 10008 14272
rect 11336 14220 11388 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 18052 14220 18104 14272
rect 19156 14263 19208 14272
rect 19156 14229 19165 14263
rect 19165 14229 19199 14263
rect 19199 14229 19208 14263
rect 19156 14220 19208 14229
rect 20076 14220 20128 14272
rect 20536 14220 20588 14272
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 23480 14263 23532 14272
rect 23480 14229 23489 14263
rect 23489 14229 23523 14263
rect 23523 14229 23532 14263
rect 23480 14220 23532 14229
rect 23848 14263 23900 14272
rect 23848 14229 23857 14263
rect 23857 14229 23891 14263
rect 23891 14229 23900 14263
rect 23848 14220 23900 14229
rect 25688 14220 25740 14272
rect 27160 14220 27212 14272
rect 27252 14220 27304 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 4068 14016 4120 14068
rect 4620 14016 4672 14068
rect 5632 14016 5684 14068
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 8300 14016 8352 14068
rect 8944 14059 8996 14068
rect 8944 14025 8953 14059
rect 8953 14025 8987 14059
rect 8987 14025 8996 14059
rect 8944 14016 8996 14025
rect 11152 14016 11204 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 14740 14059 14792 14068
rect 14740 14025 14749 14059
rect 14749 14025 14783 14059
rect 14783 14025 14792 14059
rect 14740 14016 14792 14025
rect 15752 14016 15804 14068
rect 16304 14059 16356 14068
rect 16304 14025 16313 14059
rect 16313 14025 16347 14059
rect 16347 14025 16356 14059
rect 16304 14016 16356 14025
rect 16580 14016 16632 14068
rect 17408 14016 17460 14068
rect 4804 13880 4856 13932
rect 6276 13880 6328 13932
rect 11336 13880 11388 13932
rect 15844 13948 15896 14000
rect 19524 13991 19576 14000
rect 19524 13957 19533 13991
rect 19533 13957 19567 13991
rect 19567 13957 19576 13991
rect 19524 13948 19576 13957
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15384 13880 15436 13889
rect 15476 13923 15528 13932
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 20628 13991 20680 14000
rect 20628 13957 20637 13991
rect 20637 13957 20671 13991
rect 20671 13957 20680 13991
rect 20628 13948 20680 13957
rect 20904 13991 20956 14000
rect 20904 13957 20913 13991
rect 20913 13957 20947 13991
rect 20947 13957 20956 13991
rect 20904 13948 20956 13957
rect 22100 13948 22152 14000
rect 23756 14016 23808 14068
rect 24032 14059 24084 14068
rect 24032 14025 24041 14059
rect 24041 14025 24075 14059
rect 24075 14025 24084 14059
rect 24032 14016 24084 14025
rect 25412 14016 25464 14068
rect 27160 14016 27212 14068
rect 26884 13948 26936 14000
rect 2320 13812 2372 13864
rect 4620 13855 4672 13864
rect 4620 13821 4629 13855
rect 4629 13821 4663 13855
rect 4663 13821 4672 13855
rect 4620 13812 4672 13821
rect 2504 13787 2556 13796
rect 2504 13753 2538 13787
rect 2538 13753 2556 13787
rect 2504 13744 2556 13753
rect 5632 13744 5684 13796
rect 6552 13812 6604 13864
rect 6828 13812 6880 13864
rect 8668 13812 8720 13864
rect 5908 13744 5960 13796
rect 9036 13744 9088 13796
rect 9956 13812 10008 13864
rect 10600 13812 10652 13864
rect 19984 13855 20036 13864
rect 11428 13744 11480 13796
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 20076 13812 20128 13864
rect 23848 13880 23900 13932
rect 13268 13744 13320 13796
rect 2044 13676 2096 13728
rect 6184 13719 6236 13728
rect 6184 13685 6193 13719
rect 6193 13685 6227 13719
rect 6227 13685 6236 13719
rect 6184 13676 6236 13685
rect 7012 13676 7064 13728
rect 7104 13676 7156 13728
rect 8392 13719 8444 13728
rect 8392 13685 8401 13719
rect 8401 13685 8435 13719
rect 8435 13685 8444 13719
rect 8392 13676 8444 13685
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 15108 13676 15160 13728
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 18236 13719 18288 13728
rect 18236 13685 18245 13719
rect 18245 13685 18279 13719
rect 18279 13685 18288 13719
rect 18236 13676 18288 13685
rect 19156 13676 19208 13728
rect 19892 13719 19944 13728
rect 19892 13685 19901 13719
rect 19901 13685 19935 13719
rect 19935 13685 19944 13719
rect 19892 13676 19944 13685
rect 21180 13812 21232 13864
rect 23480 13812 23532 13864
rect 24400 13855 24452 13864
rect 24400 13821 24409 13855
rect 24409 13821 24443 13855
rect 24443 13821 24452 13855
rect 24400 13812 24452 13821
rect 24584 13923 24636 13932
rect 24584 13889 24593 13923
rect 24593 13889 24627 13923
rect 24627 13889 24636 13923
rect 25596 13923 25648 13932
rect 24584 13880 24636 13889
rect 24768 13812 24820 13864
rect 23756 13744 23808 13796
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 26700 13880 26752 13932
rect 25688 13812 25740 13864
rect 21272 13676 21324 13728
rect 27068 13676 27120 13728
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 4988 13472 5040 13524
rect 5632 13515 5684 13524
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 5908 13472 5960 13524
rect 6644 13472 6696 13524
rect 10232 13472 10284 13524
rect 11336 13515 11388 13524
rect 11336 13481 11345 13515
rect 11345 13481 11379 13515
rect 11379 13481 11388 13515
rect 11336 13472 11388 13481
rect 11796 13515 11848 13524
rect 11796 13481 11805 13515
rect 11805 13481 11839 13515
rect 11839 13481 11848 13515
rect 11796 13472 11848 13481
rect 12256 13515 12308 13524
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 12808 13472 12860 13524
rect 13728 13472 13780 13524
rect 15844 13515 15896 13524
rect 15844 13481 15853 13515
rect 15853 13481 15887 13515
rect 15887 13481 15896 13515
rect 15844 13472 15896 13481
rect 19248 13515 19300 13524
rect 19248 13481 19257 13515
rect 19257 13481 19291 13515
rect 19291 13481 19300 13515
rect 19248 13472 19300 13481
rect 21732 13472 21784 13524
rect 24216 13515 24268 13524
rect 24216 13481 24225 13515
rect 24225 13481 24259 13515
rect 24259 13481 24268 13515
rect 24216 13472 24268 13481
rect 25688 13472 25740 13524
rect 3608 13404 3660 13456
rect 5816 13404 5868 13456
rect 6920 13404 6972 13456
rect 7196 13404 7248 13456
rect 9588 13404 9640 13456
rect 13268 13447 13320 13456
rect 13268 13413 13277 13447
rect 13277 13413 13311 13447
rect 13311 13413 13320 13447
rect 13268 13404 13320 13413
rect 13544 13404 13596 13456
rect 1584 13336 1636 13388
rect 1768 13379 1820 13388
rect 1768 13345 1802 13379
rect 1802 13345 1820 13379
rect 1768 13336 1820 13345
rect 3056 13336 3108 13388
rect 4252 13336 4304 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 7656 13336 7708 13388
rect 11060 13336 11112 13388
rect 12164 13379 12216 13388
rect 12164 13345 12173 13379
rect 12173 13345 12207 13379
rect 12207 13345 12216 13379
rect 12164 13336 12216 13345
rect 14096 13379 14148 13388
rect 14096 13345 14105 13379
rect 14105 13345 14139 13379
rect 14139 13345 14148 13379
rect 14096 13336 14148 13345
rect 17132 13404 17184 13456
rect 16856 13379 16908 13388
rect 16856 13345 16890 13379
rect 16890 13345 16908 13379
rect 16856 13336 16908 13345
rect 17868 13336 17920 13388
rect 18972 13336 19024 13388
rect 20444 13336 20496 13388
rect 2504 13268 2556 13320
rect 4804 13268 4856 13320
rect 5448 13268 5500 13320
rect 6184 13268 6236 13320
rect 6736 13268 6788 13320
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 10600 13311 10652 13320
rect 10600 13277 10609 13311
rect 10609 13277 10643 13311
rect 10643 13277 10652 13311
rect 10600 13268 10652 13277
rect 11888 13200 11940 13252
rect 14464 13268 14516 13320
rect 19708 13311 19760 13320
rect 19708 13277 19717 13311
rect 19717 13277 19751 13311
rect 19751 13277 19760 13311
rect 19708 13268 19760 13277
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 20628 13268 20680 13320
rect 13268 13200 13320 13252
rect 15292 13200 15344 13252
rect 20996 13268 21048 13320
rect 21824 13379 21876 13388
rect 21824 13345 21833 13379
rect 21833 13345 21867 13379
rect 21867 13345 21876 13379
rect 21824 13336 21876 13345
rect 23020 13336 23072 13388
rect 24124 13379 24176 13388
rect 24124 13345 24133 13379
rect 24133 13345 24167 13379
rect 24167 13345 24176 13379
rect 24124 13336 24176 13345
rect 25320 13379 25372 13388
rect 25320 13345 25329 13379
rect 25329 13345 25363 13379
rect 25363 13345 25372 13379
rect 25320 13336 25372 13345
rect 25504 13336 25556 13388
rect 28172 13336 28224 13388
rect 22100 13268 22152 13320
rect 26424 13268 26476 13320
rect 27068 13311 27120 13320
rect 27068 13277 27077 13311
rect 27077 13277 27111 13311
rect 27111 13277 27120 13311
rect 27068 13268 27120 13277
rect 4160 13132 4212 13184
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 5264 13132 5316 13141
rect 7104 13132 7156 13184
rect 8484 13175 8536 13184
rect 8484 13141 8493 13175
rect 8493 13141 8527 13175
rect 8527 13141 8536 13175
rect 8484 13132 8536 13141
rect 15108 13132 15160 13184
rect 16488 13175 16540 13184
rect 16488 13141 16497 13175
rect 16497 13141 16531 13175
rect 16531 13141 16540 13175
rect 16488 13132 16540 13141
rect 17960 13175 18012 13184
rect 17960 13141 17969 13175
rect 17969 13141 18003 13175
rect 18003 13141 18012 13175
rect 17960 13132 18012 13141
rect 21088 13175 21140 13184
rect 21088 13141 21097 13175
rect 21097 13141 21131 13175
rect 21131 13141 21140 13175
rect 21088 13132 21140 13141
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 23480 13132 23532 13184
rect 23756 13175 23808 13184
rect 23756 13141 23765 13175
rect 23765 13141 23799 13175
rect 23799 13141 23808 13175
rect 23756 13132 23808 13141
rect 25044 13132 25096 13184
rect 25136 13175 25188 13184
rect 25136 13141 25145 13175
rect 25145 13141 25179 13175
rect 25179 13141 25188 13175
rect 25136 13132 25188 13141
rect 25412 13132 25464 13184
rect 26332 13175 26384 13184
rect 26332 13141 26341 13175
rect 26341 13141 26375 13175
rect 26375 13141 26384 13175
rect 26332 13132 26384 13141
rect 26516 13175 26568 13184
rect 26516 13141 26525 13175
rect 26525 13141 26559 13175
rect 26559 13141 26568 13175
rect 26516 13132 26568 13141
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 3056 12971 3108 12980
rect 3056 12937 3065 12971
rect 3065 12937 3099 12971
rect 3099 12937 3108 12971
rect 3056 12928 3108 12937
rect 4252 12928 4304 12980
rect 4988 12971 5040 12980
rect 4988 12937 4997 12971
rect 4997 12937 5031 12971
rect 5031 12937 5040 12971
rect 4988 12928 5040 12937
rect 6460 12928 6512 12980
rect 6644 12928 6696 12980
rect 6736 12928 6788 12980
rect 6552 12903 6604 12912
rect 6552 12869 6561 12903
rect 6561 12869 6595 12903
rect 6595 12869 6604 12903
rect 6552 12860 6604 12869
rect 5264 12792 5316 12844
rect 6368 12792 6420 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 5172 12724 5224 12776
rect 7012 12792 7064 12844
rect 7656 12792 7708 12844
rect 10416 12928 10468 12980
rect 11336 12928 11388 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12256 12928 12308 12980
rect 12440 12971 12492 12980
rect 12440 12937 12449 12971
rect 12449 12937 12483 12971
rect 12483 12937 12492 12971
rect 12440 12928 12492 12937
rect 13544 12928 13596 12980
rect 13820 12928 13872 12980
rect 14096 12971 14148 12980
rect 14096 12937 14105 12971
rect 14105 12937 14139 12971
rect 14139 12937 14148 12971
rect 14096 12928 14148 12937
rect 16396 12971 16448 12980
rect 16396 12937 16405 12971
rect 16405 12937 16439 12971
rect 16439 12937 16448 12971
rect 16396 12928 16448 12937
rect 19800 12928 19852 12980
rect 20076 12928 20128 12980
rect 23020 12971 23072 12980
rect 23020 12937 23029 12971
rect 23029 12937 23063 12971
rect 23063 12937 23072 12971
rect 23020 12928 23072 12937
rect 23940 12971 23992 12980
rect 23940 12937 23949 12971
rect 23949 12937 23983 12971
rect 23983 12937 23992 12971
rect 23940 12928 23992 12937
rect 24124 12928 24176 12980
rect 25320 12971 25372 12980
rect 25320 12937 25329 12971
rect 25329 12937 25363 12971
rect 25363 12937 25372 12971
rect 25320 12928 25372 12937
rect 25780 12928 25832 12980
rect 26424 12928 26476 12980
rect 11060 12903 11112 12912
rect 11060 12869 11069 12903
rect 11069 12869 11103 12903
rect 11103 12869 11112 12903
rect 11060 12860 11112 12869
rect 11980 12860 12032 12912
rect 12164 12860 12216 12912
rect 10600 12792 10652 12844
rect 13268 12792 13320 12844
rect 15292 12835 15344 12844
rect 15292 12801 15301 12835
rect 15301 12801 15335 12835
rect 15335 12801 15344 12835
rect 15292 12792 15344 12801
rect 16764 12860 16816 12912
rect 20352 12860 20404 12912
rect 20628 12860 20680 12912
rect 20996 12860 21048 12912
rect 24216 12860 24268 12912
rect 16488 12792 16540 12844
rect 7380 12724 7432 12776
rect 8484 12724 8536 12776
rect 12808 12767 12860 12776
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 17408 12792 17460 12844
rect 17960 12792 18012 12844
rect 19984 12835 20036 12844
rect 19984 12801 19993 12835
rect 19993 12801 20027 12835
rect 20027 12801 20036 12835
rect 19984 12792 20036 12801
rect 23296 12792 23348 12844
rect 24860 12860 24912 12912
rect 28172 12903 28224 12912
rect 28172 12869 28181 12903
rect 28181 12869 28215 12903
rect 28215 12869 28224 12903
rect 28172 12860 28224 12869
rect 25044 12792 25096 12844
rect 25596 12792 25648 12844
rect 26148 12835 26200 12844
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 2872 12656 2924 12708
rect 3332 12656 3384 12708
rect 8300 12656 8352 12708
rect 12164 12699 12216 12708
rect 12164 12665 12173 12699
rect 12173 12665 12207 12699
rect 12207 12665 12216 12699
rect 12164 12656 12216 12665
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 5356 12588 5408 12640
rect 6736 12588 6788 12640
rect 10232 12588 10284 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 20628 12656 20680 12708
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 15844 12631 15896 12640
rect 15844 12597 15853 12631
rect 15853 12597 15887 12631
rect 15887 12597 15896 12631
rect 15844 12588 15896 12597
rect 17132 12588 17184 12640
rect 18972 12631 19024 12640
rect 18972 12597 18981 12631
rect 18981 12597 19015 12631
rect 19015 12597 19024 12631
rect 18972 12588 19024 12597
rect 19708 12588 19760 12640
rect 20260 12588 20312 12640
rect 20352 12588 20404 12640
rect 21088 12724 21140 12776
rect 23664 12724 23716 12776
rect 25136 12724 25188 12776
rect 21272 12699 21324 12708
rect 21272 12665 21306 12699
rect 21306 12665 21324 12699
rect 21272 12656 21324 12665
rect 26240 12656 26292 12708
rect 27528 12631 27580 12640
rect 27528 12597 27537 12631
rect 27537 12597 27571 12631
rect 27571 12597 27580 12631
rect 27528 12588 27580 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 1676 12427 1728 12436
rect 1676 12393 1685 12427
rect 1685 12393 1719 12427
rect 1719 12393 1728 12427
rect 1676 12384 1728 12393
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 5264 12384 5316 12436
rect 5448 12384 5500 12436
rect 3516 12359 3568 12368
rect 3516 12325 3525 12359
rect 3525 12325 3559 12359
rect 3559 12325 3568 12359
rect 8392 12384 8444 12436
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 16488 12384 16540 12436
rect 3516 12316 3568 12325
rect 5816 12316 5868 12368
rect 10232 12316 10284 12368
rect 4068 12248 4120 12300
rect 12716 12248 12768 12300
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 15384 12248 15436 12300
rect 4804 12112 4856 12164
rect 2596 12044 2648 12096
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 4068 12087 4120 12096
rect 4068 12053 4077 12087
rect 4077 12053 4111 12087
rect 4111 12053 4120 12087
rect 4068 12044 4120 12053
rect 7196 12180 7248 12232
rect 7656 12155 7708 12164
rect 7656 12121 7665 12155
rect 7665 12121 7699 12155
rect 7699 12121 7708 12155
rect 7656 12112 7708 12121
rect 8668 12112 8720 12164
rect 9772 12180 9824 12232
rect 12164 12180 12216 12232
rect 14832 12180 14884 12232
rect 15844 12180 15896 12232
rect 16764 12384 16816 12436
rect 19984 12384 20036 12436
rect 26148 12427 26200 12436
rect 26148 12393 26157 12427
rect 26157 12393 26191 12427
rect 26191 12393 26200 12427
rect 26148 12384 26200 12393
rect 26516 12384 26568 12436
rect 17408 12291 17460 12300
rect 17408 12257 17442 12291
rect 17442 12257 17460 12291
rect 17408 12248 17460 12257
rect 20168 12248 20220 12300
rect 23480 12248 23532 12300
rect 24492 12248 24544 12300
rect 26148 12248 26200 12300
rect 26608 12248 26660 12300
rect 17132 12223 17184 12232
rect 14464 12112 14516 12164
rect 15660 12112 15712 12164
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 20628 12180 20680 12232
rect 20904 12223 20956 12232
rect 20904 12189 20913 12223
rect 20913 12189 20947 12223
rect 20947 12189 20956 12223
rect 20904 12180 20956 12189
rect 23296 12112 23348 12164
rect 27528 12180 27580 12232
rect 6368 12044 6420 12096
rect 6552 12044 6604 12096
rect 8300 12044 8352 12096
rect 8760 12087 8812 12096
rect 8760 12053 8769 12087
rect 8769 12053 8803 12087
rect 8803 12053 8812 12087
rect 8760 12044 8812 12053
rect 11428 12087 11480 12096
rect 11428 12053 11437 12087
rect 11437 12053 11471 12087
rect 11471 12053 11480 12087
rect 11428 12044 11480 12053
rect 11888 12044 11940 12096
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 14556 12087 14608 12096
rect 14556 12053 14565 12087
rect 14565 12053 14599 12087
rect 14599 12053 14608 12087
rect 14556 12044 14608 12053
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 18420 12044 18472 12096
rect 20260 12087 20312 12096
rect 20260 12053 20269 12087
rect 20269 12053 20303 12087
rect 20303 12053 20312 12087
rect 20260 12044 20312 12053
rect 20444 12044 20496 12096
rect 21272 12044 21324 12096
rect 24308 12044 24360 12096
rect 25780 12044 25832 12096
rect 25872 12044 25924 12096
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 1676 11840 1728 11892
rect 1768 11704 1820 11756
rect 4528 11772 4580 11824
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 7196 11840 7248 11892
rect 2412 11636 2464 11688
rect 3516 11568 3568 11620
rect 5816 11568 5868 11620
rect 7564 11840 7616 11892
rect 9772 11883 9824 11892
rect 9772 11849 9781 11883
rect 9781 11849 9815 11883
rect 9815 11849 9824 11883
rect 9772 11840 9824 11849
rect 10876 11840 10928 11892
rect 14832 11883 14884 11892
rect 14832 11849 14841 11883
rect 14841 11849 14875 11883
rect 14875 11849 14884 11883
rect 14832 11840 14884 11849
rect 20536 11840 20588 11892
rect 22836 11840 22888 11892
rect 11704 11772 11756 11824
rect 12164 11772 12216 11824
rect 12716 11815 12768 11824
rect 12716 11781 12725 11815
rect 12725 11781 12759 11815
rect 12759 11781 12768 11815
rect 12716 11772 12768 11781
rect 20352 11772 20404 11824
rect 20904 11772 20956 11824
rect 23296 11772 23348 11824
rect 23480 11815 23532 11824
rect 23480 11781 23489 11815
rect 23489 11781 23523 11815
rect 23523 11781 23532 11815
rect 23480 11772 23532 11781
rect 8668 11704 8720 11756
rect 11428 11704 11480 11756
rect 12900 11704 12952 11756
rect 12992 11704 13044 11756
rect 14464 11704 14516 11756
rect 14924 11704 14976 11756
rect 15752 11704 15804 11756
rect 16488 11704 16540 11756
rect 17040 11747 17092 11756
rect 17040 11713 17049 11747
rect 17049 11713 17083 11747
rect 17083 11713 17092 11747
rect 17040 11704 17092 11713
rect 17132 11704 17184 11756
rect 8392 11636 8444 11688
rect 10508 11636 10560 11688
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 15292 11636 15344 11688
rect 15844 11679 15896 11688
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 16948 11636 17000 11688
rect 17776 11636 17828 11688
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 18420 11679 18472 11688
rect 18420 11645 18454 11679
rect 18454 11645 18472 11679
rect 18420 11636 18472 11645
rect 19984 11636 20036 11688
rect 20536 11636 20588 11688
rect 21824 11679 21876 11688
rect 21824 11645 21833 11679
rect 21833 11645 21867 11679
rect 21867 11645 21876 11679
rect 21824 11636 21876 11645
rect 24860 11840 24912 11892
rect 26792 11883 26844 11892
rect 26792 11849 26801 11883
rect 26801 11849 26835 11883
rect 26835 11849 26844 11883
rect 26792 11840 26844 11849
rect 27160 11840 27212 11892
rect 25780 11772 25832 11824
rect 24492 11747 24544 11756
rect 24492 11713 24501 11747
rect 24501 11713 24535 11747
rect 24535 11713 24544 11747
rect 24492 11704 24544 11713
rect 25872 11747 25924 11756
rect 25320 11636 25372 11688
rect 25872 11713 25881 11747
rect 25881 11713 25915 11747
rect 25915 11713 25924 11747
rect 25872 11704 25924 11713
rect 26608 11747 26660 11756
rect 26608 11713 26617 11747
rect 26617 11713 26651 11747
rect 26651 11713 26660 11747
rect 26608 11704 26660 11713
rect 27436 11747 27488 11756
rect 27436 11713 27445 11747
rect 27445 11713 27479 11747
rect 27479 11713 27488 11747
rect 27436 11704 27488 11713
rect 27528 11747 27580 11756
rect 27528 11713 27537 11747
rect 27537 11713 27571 11747
rect 27571 11713 27580 11747
rect 27528 11704 27580 11713
rect 20352 11568 20404 11620
rect 20812 11568 20864 11620
rect 21640 11568 21692 11620
rect 24952 11568 25004 11620
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4804 11500 4856 11552
rect 5172 11543 5224 11552
rect 5172 11509 5181 11543
rect 5181 11509 5215 11543
rect 5215 11509 5224 11543
rect 5172 11500 5224 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 6368 11500 6420 11552
rect 7104 11500 7156 11552
rect 8208 11500 8260 11552
rect 8392 11543 8444 11552
rect 8392 11509 8401 11543
rect 8401 11509 8435 11543
rect 8435 11509 8444 11543
rect 8392 11500 8444 11509
rect 10324 11500 10376 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 15292 11543 15344 11552
rect 15292 11509 15301 11543
rect 15301 11509 15335 11543
rect 15335 11509 15344 11543
rect 15292 11500 15344 11509
rect 16212 11543 16264 11552
rect 16212 11509 16221 11543
rect 16221 11509 16255 11543
rect 16255 11509 16264 11543
rect 16212 11500 16264 11509
rect 16396 11543 16448 11552
rect 16396 11509 16405 11543
rect 16405 11509 16439 11543
rect 16439 11509 16448 11543
rect 16396 11500 16448 11509
rect 20168 11543 20220 11552
rect 20168 11509 20177 11543
rect 20177 11509 20211 11543
rect 20211 11509 20220 11543
rect 20168 11500 20220 11509
rect 21272 11543 21324 11552
rect 21272 11509 21281 11543
rect 21281 11509 21315 11543
rect 21315 11509 21324 11543
rect 21272 11500 21324 11509
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 26424 11543 26476 11552
rect 26424 11509 26433 11543
rect 26433 11509 26467 11543
rect 26467 11509 26476 11543
rect 27160 11568 27212 11620
rect 26424 11500 26476 11509
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 2136 11339 2188 11348
rect 2136 11305 2145 11339
rect 2145 11305 2179 11339
rect 2179 11305 2188 11339
rect 2136 11296 2188 11305
rect 3148 11296 3200 11348
rect 3516 11339 3568 11348
rect 3516 11305 3525 11339
rect 3525 11305 3559 11339
rect 3559 11305 3568 11339
rect 3516 11296 3568 11305
rect 4068 11296 4120 11348
rect 5816 11296 5868 11348
rect 6920 11339 6972 11348
rect 6920 11305 6929 11339
rect 6929 11305 6963 11339
rect 6963 11305 6972 11339
rect 6920 11296 6972 11305
rect 7012 11296 7064 11348
rect 8024 11296 8076 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 11336 11296 11388 11348
rect 12532 11296 12584 11348
rect 12992 11296 13044 11348
rect 14556 11296 14608 11348
rect 15200 11296 15252 11348
rect 16488 11296 16540 11348
rect 17408 11296 17460 11348
rect 18144 11339 18196 11348
rect 18144 11305 18153 11339
rect 18153 11305 18187 11339
rect 18187 11305 18196 11339
rect 18144 11296 18196 11305
rect 18420 11296 18472 11348
rect 20260 11296 20312 11348
rect 20720 11296 20772 11348
rect 23664 11339 23716 11348
rect 23664 11305 23673 11339
rect 23673 11305 23707 11339
rect 23707 11305 23716 11339
rect 23664 11296 23716 11305
rect 24952 11296 25004 11348
rect 25872 11296 25924 11348
rect 26516 11339 26568 11348
rect 26516 11305 26525 11339
rect 26525 11305 26559 11339
rect 26559 11305 26568 11339
rect 26516 11296 26568 11305
rect 26884 11339 26936 11348
rect 26884 11305 26893 11339
rect 26893 11305 26927 11339
rect 26927 11305 26936 11339
rect 26884 11296 26936 11305
rect 27344 11296 27396 11348
rect 27528 11339 27580 11348
rect 27528 11305 27537 11339
rect 27537 11305 27571 11339
rect 27571 11305 27580 11339
rect 27528 11296 27580 11305
rect 10232 11228 10284 11280
rect 14924 11271 14976 11280
rect 3056 11160 3108 11212
rect 4068 11160 4120 11212
rect 5264 11203 5316 11212
rect 5264 11169 5298 11203
rect 5298 11169 5316 11203
rect 5264 11160 5316 11169
rect 8208 11160 8260 11212
rect 10600 11203 10652 11212
rect 10600 11169 10609 11203
rect 10609 11169 10643 11203
rect 10643 11169 10652 11203
rect 10600 11160 10652 11169
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 2320 11092 2372 11144
rect 2964 11135 3016 11144
rect 2688 11024 2740 11076
rect 2964 11101 2973 11135
rect 2973 11101 3007 11135
rect 3007 11101 3016 11135
rect 2964 11092 3016 11101
rect 3516 11092 3568 11144
rect 8300 11092 8352 11144
rect 8760 11092 8812 11144
rect 10140 11092 10192 11144
rect 10692 11135 10744 11144
rect 10692 11101 10701 11135
rect 10701 11101 10735 11135
rect 10735 11101 10744 11135
rect 10692 11092 10744 11101
rect 14924 11237 14933 11271
rect 14933 11237 14967 11271
rect 14967 11237 14976 11271
rect 14924 11228 14976 11237
rect 15660 11271 15712 11280
rect 15660 11237 15669 11271
rect 15669 11237 15703 11271
rect 15703 11237 15712 11271
rect 15660 11228 15712 11237
rect 17776 11228 17828 11280
rect 18512 11228 18564 11280
rect 19892 11228 19944 11280
rect 22100 11228 22152 11280
rect 23480 11228 23532 11280
rect 23756 11228 23808 11280
rect 27620 11228 27672 11280
rect 11888 11160 11940 11212
rect 11704 11092 11756 11144
rect 15568 11160 15620 11212
rect 16304 11160 16356 11212
rect 19248 11160 19300 11212
rect 20812 11160 20864 11212
rect 21916 11160 21968 11212
rect 22560 11203 22612 11212
rect 22560 11169 22569 11203
rect 22569 11169 22603 11203
rect 22603 11169 22612 11203
rect 22560 11160 22612 11169
rect 25596 11160 25648 11212
rect 3884 10999 3936 11008
rect 3884 10965 3893 10999
rect 3893 10965 3927 10999
rect 3927 10965 3936 10999
rect 3884 10956 3936 10965
rect 3976 10956 4028 11008
rect 12164 11024 12216 11076
rect 16672 11135 16724 11144
rect 16672 11101 16681 11135
rect 16681 11101 16715 11135
rect 16715 11101 16724 11135
rect 18328 11135 18380 11144
rect 16672 11092 16724 11101
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 16488 11024 16540 11076
rect 4988 10956 5040 11008
rect 7012 10956 7064 11008
rect 7656 10956 7708 11008
rect 18972 10956 19024 11008
rect 20444 11092 20496 11144
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 23480 11092 23532 11144
rect 23848 11092 23900 11144
rect 24308 11135 24360 11144
rect 24308 11101 24317 11135
rect 24317 11101 24351 11135
rect 24351 11101 24360 11135
rect 24308 11092 24360 11101
rect 22744 11067 22796 11076
rect 22744 11033 22753 11067
rect 22753 11033 22787 11067
rect 22787 11033 22796 11067
rect 22744 11024 22796 11033
rect 25688 11024 25740 11076
rect 27252 11092 27304 11144
rect 21732 10956 21784 11008
rect 23296 10956 23348 11008
rect 23664 10956 23716 11008
rect 26700 10956 26752 11008
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 3148 10795 3200 10804
rect 3148 10761 3157 10795
rect 3157 10761 3191 10795
rect 3191 10761 3200 10795
rect 3148 10752 3200 10761
rect 3608 10795 3660 10804
rect 3608 10761 3617 10795
rect 3617 10761 3651 10795
rect 3651 10761 3660 10795
rect 3608 10752 3660 10761
rect 4160 10752 4212 10804
rect 7472 10752 7524 10804
rect 8208 10752 8260 10804
rect 10140 10795 10192 10804
rect 10140 10761 10149 10795
rect 10149 10761 10183 10795
rect 10183 10761 10192 10795
rect 10140 10752 10192 10761
rect 10324 10795 10376 10804
rect 10324 10761 10333 10795
rect 10333 10761 10367 10795
rect 10367 10761 10376 10795
rect 10324 10752 10376 10761
rect 3792 10684 3844 10736
rect 8300 10727 8352 10736
rect 8300 10693 8309 10727
rect 8309 10693 8343 10727
rect 8343 10693 8352 10727
rect 8300 10684 8352 10693
rect 1584 10616 1636 10668
rect 2136 10616 2188 10668
rect 2964 10616 3016 10668
rect 5264 10616 5316 10668
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 8116 10616 8168 10668
rect 11336 10616 11388 10668
rect 11704 10752 11756 10804
rect 11888 10795 11940 10804
rect 11888 10761 11897 10795
rect 11897 10761 11931 10795
rect 11931 10761 11940 10795
rect 11888 10752 11940 10761
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 12532 10752 12584 10804
rect 15292 10752 15344 10804
rect 17776 10795 17828 10804
rect 17776 10761 17785 10795
rect 17785 10761 17819 10795
rect 17819 10761 17828 10795
rect 17776 10752 17828 10761
rect 18972 10795 19024 10804
rect 18972 10761 18981 10795
rect 18981 10761 19015 10795
rect 19015 10761 19024 10795
rect 18972 10752 19024 10761
rect 15384 10684 15436 10736
rect 15568 10727 15620 10736
rect 15568 10693 15577 10727
rect 15577 10693 15611 10727
rect 15611 10693 15620 10727
rect 15568 10684 15620 10693
rect 16580 10616 16632 10668
rect 17868 10616 17920 10668
rect 19340 10616 19392 10668
rect 20352 10752 20404 10804
rect 21456 10795 21508 10804
rect 21456 10761 21465 10795
rect 21465 10761 21499 10795
rect 21499 10761 21508 10795
rect 21456 10752 21508 10761
rect 22560 10752 22612 10804
rect 24768 10752 24820 10804
rect 27344 10752 27396 10804
rect 27620 10795 27672 10804
rect 27620 10761 27629 10795
rect 27629 10761 27663 10795
rect 27663 10761 27672 10795
rect 27620 10752 27672 10761
rect 21732 10616 21784 10668
rect 24952 10684 25004 10736
rect 25228 10684 25280 10736
rect 26700 10659 26752 10668
rect 2780 10548 2832 10600
rect 3884 10548 3936 10600
rect 7748 10591 7800 10600
rect 7748 10557 7757 10591
rect 7757 10557 7791 10591
rect 7791 10557 7800 10591
rect 7748 10548 7800 10557
rect 4252 10480 4304 10532
rect 6920 10480 6972 10532
rect 10600 10548 10652 10600
rect 10784 10548 10836 10600
rect 16856 10591 16908 10600
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 21824 10591 21876 10600
rect 21824 10557 21833 10591
rect 21833 10557 21867 10591
rect 21867 10557 21876 10591
rect 21824 10548 21876 10557
rect 22376 10591 22428 10600
rect 22376 10557 22385 10591
rect 22385 10557 22419 10591
rect 22419 10557 22428 10591
rect 22376 10548 22428 10557
rect 23572 10548 23624 10600
rect 23664 10591 23716 10600
rect 23664 10557 23673 10591
rect 23673 10557 23707 10591
rect 23707 10557 23716 10591
rect 23664 10548 23716 10557
rect 24308 10548 24360 10600
rect 25596 10591 25648 10600
rect 25596 10557 25605 10591
rect 25605 10557 25639 10591
rect 25639 10557 25648 10591
rect 25596 10548 25648 10557
rect 26700 10625 26709 10659
rect 26709 10625 26743 10659
rect 26743 10625 26752 10659
rect 26700 10616 26752 10625
rect 16764 10523 16816 10532
rect 16764 10489 16773 10523
rect 16773 10489 16807 10523
rect 16807 10489 16816 10523
rect 16764 10480 16816 10489
rect 20352 10480 20404 10532
rect 25780 10480 25832 10532
rect 2044 10455 2096 10464
rect 2044 10421 2053 10455
rect 2053 10421 2087 10455
rect 2087 10421 2096 10455
rect 2044 10412 2096 10421
rect 4068 10455 4120 10464
rect 4068 10421 4077 10455
rect 4077 10421 4111 10455
rect 4111 10421 4120 10455
rect 4068 10412 4120 10421
rect 5540 10455 5592 10464
rect 5540 10421 5549 10455
rect 5549 10421 5583 10455
rect 5583 10421 5592 10455
rect 5540 10412 5592 10421
rect 6368 10412 6420 10464
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 7656 10455 7708 10464
rect 7656 10421 7665 10455
rect 7665 10421 7699 10455
rect 7699 10421 7708 10455
rect 7656 10412 7708 10421
rect 9036 10455 9088 10464
rect 9036 10421 9045 10455
rect 9045 10421 9079 10455
rect 9079 10421 9088 10455
rect 9036 10412 9088 10421
rect 10324 10412 10376 10464
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 20628 10412 20680 10464
rect 21916 10455 21968 10464
rect 21916 10421 21925 10455
rect 21925 10421 21959 10455
rect 21959 10421 21968 10455
rect 21916 10412 21968 10421
rect 26516 10412 26568 10464
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 1400 10208 1452 10260
rect 2412 10251 2464 10260
rect 2412 10217 2421 10251
rect 2421 10217 2455 10251
rect 2455 10217 2464 10251
rect 2412 10208 2464 10217
rect 2504 10251 2556 10260
rect 2504 10217 2513 10251
rect 2513 10217 2547 10251
rect 2547 10217 2556 10251
rect 2504 10208 2556 10217
rect 2964 10208 3016 10260
rect 5264 10208 5316 10260
rect 6552 10208 6604 10260
rect 7012 10251 7064 10260
rect 7012 10217 7021 10251
rect 7021 10217 7055 10251
rect 7055 10217 7064 10251
rect 7012 10208 7064 10217
rect 8024 10251 8076 10260
rect 8024 10217 8033 10251
rect 8033 10217 8067 10251
rect 8067 10217 8076 10251
rect 8024 10208 8076 10217
rect 10324 10251 10376 10260
rect 10324 10217 10333 10251
rect 10333 10217 10367 10251
rect 10367 10217 10376 10251
rect 10324 10208 10376 10217
rect 11336 10208 11388 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 16396 10208 16448 10260
rect 17684 10251 17736 10260
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 19248 10251 19300 10260
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 19524 10208 19576 10260
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 20812 10208 20864 10260
rect 21364 10251 21416 10260
rect 21364 10217 21373 10251
rect 21373 10217 21407 10251
rect 21407 10217 21416 10251
rect 21364 10208 21416 10217
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 24124 10208 24176 10260
rect 24308 10208 24360 10260
rect 24584 10251 24636 10260
rect 24584 10217 24593 10251
rect 24593 10217 24627 10251
rect 24627 10217 24636 10251
rect 24584 10208 24636 10217
rect 4804 10140 4856 10192
rect 4712 10072 4764 10124
rect 6920 10115 6972 10124
rect 6920 10081 6929 10115
rect 6929 10081 6963 10115
rect 6963 10081 6972 10115
rect 6920 10072 6972 10081
rect 7656 10140 7708 10192
rect 21916 10140 21968 10192
rect 23388 10140 23440 10192
rect 25228 10208 25280 10260
rect 25872 10208 25924 10260
rect 8116 10115 8168 10124
rect 8116 10081 8125 10115
rect 8125 10081 8159 10115
rect 8159 10081 8168 10115
rect 8116 10072 8168 10081
rect 9312 10072 9364 10124
rect 10784 10115 10836 10124
rect 10784 10081 10793 10115
rect 10793 10081 10827 10115
rect 10827 10081 10836 10115
rect 10784 10072 10836 10081
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 19432 10072 19484 10124
rect 19616 10115 19668 10124
rect 19616 10081 19625 10115
rect 19625 10081 19659 10115
rect 19659 10081 19668 10115
rect 19616 10072 19668 10081
rect 20812 10072 20864 10124
rect 21272 10115 21324 10124
rect 21272 10081 21281 10115
rect 21281 10081 21315 10115
rect 21315 10081 21324 10115
rect 21272 10072 21324 10081
rect 21640 10072 21692 10124
rect 2964 10004 3016 10056
rect 3976 10004 4028 10056
rect 5816 9936 5868 9988
rect 7748 10004 7800 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 17132 10047 17184 10056
rect 17132 10013 17141 10047
rect 17141 10013 17175 10047
rect 17175 10013 17184 10047
rect 17132 10004 17184 10013
rect 18328 10004 18380 10056
rect 20168 10004 20220 10056
rect 21732 10004 21784 10056
rect 2228 9868 2280 9920
rect 4068 9868 4120 9920
rect 5724 9868 5776 9920
rect 7380 9868 7432 9920
rect 8392 9868 8444 9920
rect 16488 9911 16540 9920
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 20720 9868 20772 9920
rect 22376 9868 22428 9920
rect 24952 9868 25004 9920
rect 26608 10072 26660 10124
rect 25596 10004 25648 10056
rect 26700 10004 26752 10056
rect 26516 9936 26568 9988
rect 26976 9868 27028 9920
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 2872 9664 2924 9716
rect 2504 9596 2556 9648
rect 2964 9596 3016 9648
rect 3884 9664 3936 9716
rect 3608 9596 3660 9648
rect 7012 9664 7064 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 2872 9528 2924 9580
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 3240 9528 3292 9580
rect 4712 9571 4764 9580
rect 4712 9537 4721 9571
rect 4721 9537 4755 9571
rect 4755 9537 4764 9571
rect 4712 9528 4764 9537
rect 3424 9460 3476 9512
rect 8944 9596 8996 9648
rect 9128 9596 9180 9648
rect 15660 9596 15712 9648
rect 16948 9664 17000 9716
rect 19432 9664 19484 9716
rect 21364 9664 21416 9716
rect 21732 9707 21784 9716
rect 21732 9673 21741 9707
rect 21741 9673 21775 9707
rect 21775 9673 21784 9707
rect 21732 9664 21784 9673
rect 25228 9707 25280 9716
rect 25228 9673 25237 9707
rect 25237 9673 25271 9707
rect 25271 9673 25280 9707
rect 25228 9664 25280 9673
rect 26608 9664 26660 9716
rect 24768 9596 24820 9648
rect 25504 9639 25556 9648
rect 25504 9605 25513 9639
rect 25513 9605 25547 9639
rect 25547 9605 25556 9639
rect 25504 9596 25556 9605
rect 5816 9528 5868 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 16764 9528 16816 9580
rect 17132 9528 17184 9580
rect 6828 9460 6880 9512
rect 16304 9503 16356 9512
rect 16304 9469 16313 9503
rect 16313 9469 16347 9503
rect 16347 9469 16356 9503
rect 16304 9460 16356 9469
rect 3240 9392 3292 9444
rect 3700 9392 3752 9444
rect 3976 9392 4028 9444
rect 4896 9392 4948 9444
rect 7196 9435 7248 9444
rect 7196 9401 7205 9435
rect 7205 9401 7239 9435
rect 7239 9401 7248 9435
rect 7196 9392 7248 9401
rect 15292 9392 15344 9444
rect 21272 9528 21324 9580
rect 19156 9460 19208 9512
rect 23940 9460 23992 9512
rect 25320 9503 25372 9512
rect 25320 9469 25329 9503
rect 25329 9469 25363 9503
rect 25363 9469 25372 9503
rect 25320 9460 25372 9469
rect 26424 9503 26476 9512
rect 26424 9469 26433 9503
rect 26433 9469 26467 9503
rect 26467 9469 26476 9503
rect 26424 9460 26476 9469
rect 27528 9503 27580 9512
rect 27528 9469 27537 9503
rect 27537 9469 27571 9503
rect 27571 9469 27580 9503
rect 27528 9460 27580 9469
rect 1676 9324 1728 9376
rect 1860 9324 1912 9376
rect 2780 9324 2832 9376
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3608 9324 3660 9376
rect 4620 9367 4672 9376
rect 4620 9333 4629 9367
rect 4629 9333 4663 9367
rect 4663 9333 4672 9367
rect 4620 9324 4672 9333
rect 7012 9324 7064 9376
rect 16396 9367 16448 9376
rect 16396 9333 16405 9367
rect 16405 9333 16439 9367
rect 16439 9333 16448 9367
rect 16396 9324 16448 9333
rect 16856 9367 16908 9376
rect 16856 9333 16865 9367
rect 16865 9333 16899 9367
rect 16899 9333 16908 9367
rect 16856 9324 16908 9333
rect 18880 9367 18932 9376
rect 18880 9333 18889 9367
rect 18889 9333 18923 9367
rect 18923 9333 18932 9367
rect 18880 9324 18932 9333
rect 20628 9392 20680 9444
rect 20444 9367 20496 9376
rect 20444 9333 20453 9367
rect 20453 9333 20487 9367
rect 20487 9333 20496 9367
rect 20444 9324 20496 9333
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 26700 9324 26752 9376
rect 27804 9324 27856 9376
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 1400 9120 1452 9172
rect 2044 9120 2096 9172
rect 2872 9163 2924 9172
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3608 9163 3660 9172
rect 3608 9129 3617 9163
rect 3617 9129 3651 9163
rect 3651 9129 3660 9163
rect 3608 9120 3660 9129
rect 7196 9163 7248 9172
rect 7196 9129 7205 9163
rect 7205 9129 7239 9163
rect 7239 9129 7248 9163
rect 7196 9120 7248 9129
rect 15292 9163 15344 9172
rect 15292 9129 15301 9163
rect 15301 9129 15335 9163
rect 15335 9129 15344 9163
rect 15292 9120 15344 9129
rect 19156 9163 19208 9172
rect 19156 9129 19165 9163
rect 19165 9129 19199 9163
rect 19199 9129 19208 9163
rect 19156 9120 19208 9129
rect 19708 9163 19760 9172
rect 19708 9129 19717 9163
rect 19717 9129 19751 9163
rect 19751 9129 19760 9163
rect 19708 9120 19760 9129
rect 24676 9163 24728 9172
rect 24676 9129 24685 9163
rect 24685 9129 24719 9163
rect 24719 9129 24728 9163
rect 24676 9120 24728 9129
rect 2228 9095 2280 9104
rect 2228 9061 2237 9095
rect 2237 9061 2271 9095
rect 2271 9061 2280 9095
rect 2228 9052 2280 9061
rect 2688 9052 2740 9104
rect 5356 9052 5408 9104
rect 7380 9052 7432 9104
rect 1860 8984 1912 9036
rect 2872 8984 2924 9036
rect 7564 8984 7616 9036
rect 16580 9095 16632 9104
rect 16580 9061 16614 9095
rect 16614 9061 16632 9095
rect 16580 9052 16632 9061
rect 17132 9052 17184 9104
rect 20536 9052 20588 9104
rect 16304 9027 16356 9036
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 6920 8916 6972 8968
rect 7840 8959 7892 8968
rect 7840 8925 7849 8959
rect 7849 8925 7883 8959
rect 7883 8925 7892 8959
rect 7840 8916 7892 8925
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 26516 9027 26568 9036
rect 26516 8993 26525 9027
rect 26525 8993 26559 9027
rect 26559 8993 26568 9027
rect 26516 8984 26568 8993
rect 8208 8916 8260 8968
rect 2412 8848 2464 8900
rect 4712 8848 4764 8900
rect 1860 8823 1912 8832
rect 1860 8789 1869 8823
rect 1869 8789 1903 8823
rect 1903 8789 1912 8823
rect 1860 8780 1912 8789
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 18604 8848 18656 8900
rect 20168 8916 20220 8968
rect 20628 8916 20680 8968
rect 5632 8780 5684 8832
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 6920 8780 6972 8789
rect 7380 8823 7432 8832
rect 7380 8789 7389 8823
rect 7389 8789 7423 8823
rect 7423 8789 7432 8823
rect 7380 8780 7432 8789
rect 16948 8780 17000 8832
rect 19156 8780 19208 8832
rect 25504 8823 25556 8832
rect 25504 8789 25513 8823
rect 25513 8789 25547 8823
rect 25547 8789 25556 8823
rect 25504 8780 25556 8789
rect 25872 8780 25924 8832
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 1952 8619 2004 8628
rect 1952 8585 1961 8619
rect 1961 8585 1995 8619
rect 1995 8585 2004 8619
rect 1952 8576 2004 8585
rect 2964 8576 3016 8628
rect 3700 8619 3752 8628
rect 3700 8585 3709 8619
rect 3709 8585 3743 8619
rect 3743 8585 3752 8619
rect 3700 8576 3752 8585
rect 4160 8576 4212 8628
rect 7840 8576 7892 8628
rect 16304 8576 16356 8628
rect 16672 8576 16724 8628
rect 18604 8619 18656 8628
rect 18604 8585 18613 8619
rect 18613 8585 18647 8619
rect 18647 8585 18656 8619
rect 18604 8576 18656 8585
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20536 8576 20588 8628
rect 25136 8619 25188 8628
rect 25136 8585 25145 8619
rect 25145 8585 25179 8619
rect 25179 8585 25188 8619
rect 25136 8576 25188 8585
rect 25320 8576 25372 8628
rect 26516 8576 26568 8628
rect 27712 8619 27764 8628
rect 27712 8585 27721 8619
rect 27721 8585 27755 8619
rect 27755 8585 27764 8619
rect 27712 8576 27764 8585
rect 27988 8576 28040 8628
rect 8208 8551 8260 8560
rect 8208 8517 8217 8551
rect 8217 8517 8251 8551
rect 8251 8517 8260 8551
rect 8208 8508 8260 8517
rect 3332 8440 3384 8492
rect 1860 8372 1912 8424
rect 2320 8415 2372 8424
rect 2320 8381 2329 8415
rect 2329 8381 2363 8415
rect 2363 8381 2372 8415
rect 2320 8372 2372 8381
rect 4436 8440 4488 8492
rect 4804 8440 4856 8492
rect 5172 8440 5224 8492
rect 5632 8440 5684 8492
rect 16488 8440 16540 8492
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 19156 8483 19208 8492
rect 19156 8449 19165 8483
rect 19165 8449 19199 8483
rect 19199 8449 19208 8483
rect 19156 8440 19208 8449
rect 19708 8440 19760 8492
rect 20444 8440 20496 8492
rect 25596 8508 25648 8560
rect 26608 8551 26660 8560
rect 26608 8517 26617 8551
rect 26617 8517 26651 8551
rect 26651 8517 26660 8551
rect 26608 8508 26660 8517
rect 4896 8372 4948 8424
rect 6368 8372 6420 8424
rect 6552 8415 6604 8424
rect 6552 8381 6561 8415
rect 6561 8381 6595 8415
rect 6595 8381 6604 8415
rect 6552 8372 6604 8381
rect 16396 8372 16448 8424
rect 5264 8304 5316 8356
rect 7288 8304 7340 8356
rect 20720 8304 20772 8356
rect 2872 8236 2924 8288
rect 5356 8236 5408 8288
rect 16304 8279 16356 8288
rect 16304 8245 16313 8279
rect 16313 8245 16347 8279
rect 16347 8245 16356 8279
rect 16304 8236 16356 8245
rect 18696 8279 18748 8288
rect 18696 8245 18705 8279
rect 18705 8245 18739 8279
rect 18739 8245 18748 8279
rect 18696 8236 18748 8245
rect 25136 8372 25188 8424
rect 26424 8415 26476 8424
rect 26424 8381 26433 8415
rect 26433 8381 26467 8415
rect 26467 8381 26476 8415
rect 26424 8372 26476 8381
rect 27988 8372 28040 8424
rect 27068 8236 27120 8288
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 2044 8032 2096 8084
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 2872 8032 2924 8084
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 5632 8075 5684 8084
rect 5632 8041 5641 8075
rect 5641 8041 5675 8075
rect 5675 8041 5684 8075
rect 5632 8032 5684 8041
rect 6460 8032 6512 8084
rect 7472 8032 7524 8084
rect 7840 8032 7892 8084
rect 16488 8032 16540 8084
rect 20168 8075 20220 8084
rect 20168 8041 20177 8075
rect 20177 8041 20211 8075
rect 20211 8041 20220 8075
rect 20168 8032 20220 8041
rect 20720 8032 20772 8084
rect 21272 8075 21324 8084
rect 21272 8041 21281 8075
rect 21281 8041 21315 8075
rect 21315 8041 21324 8075
rect 21272 8032 21324 8041
rect 21640 8032 21692 8084
rect 25504 8075 25556 8084
rect 25504 8041 25513 8075
rect 25513 8041 25547 8075
rect 25547 8041 25556 8075
rect 25504 8032 25556 8041
rect 2228 7964 2280 8016
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2412 7896 2464 7948
rect 2780 7964 2832 8016
rect 5264 7964 5316 8016
rect 8116 8007 8168 8016
rect 2596 7896 2648 7948
rect 8116 7973 8125 8007
rect 8125 7973 8159 8007
rect 8159 7973 8168 8007
rect 8116 7964 8168 7973
rect 16856 7964 16908 8016
rect 1308 7828 1360 7880
rect 6276 7896 6328 7948
rect 16672 7939 16724 7948
rect 16672 7905 16681 7939
rect 16681 7905 16715 7939
rect 16715 7905 16724 7939
rect 16672 7896 16724 7905
rect 19064 7896 19116 7948
rect 25320 7939 25372 7948
rect 25320 7905 25329 7939
rect 25329 7905 25363 7939
rect 25363 7905 25372 7939
rect 25320 7896 25372 7905
rect 26792 7896 26844 7948
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 7288 7828 7340 7880
rect 7564 7828 7616 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 21364 7871 21416 7880
rect 19708 7828 19760 7837
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 5816 7760 5868 7812
rect 1400 7692 1452 7744
rect 5080 7692 5132 7744
rect 9128 7760 9180 7812
rect 19248 7760 19300 7812
rect 20168 7760 20220 7812
rect 21640 7760 21692 7812
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 17040 7692 17092 7744
rect 18604 7692 18656 7744
rect 19156 7735 19208 7744
rect 19156 7701 19165 7735
rect 19165 7701 19199 7735
rect 19199 7701 19208 7735
rect 19156 7692 19208 7701
rect 26792 7692 26844 7744
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 1584 7488 1636 7540
rect 2596 7488 2648 7540
rect 4252 7531 4304 7540
rect 4252 7497 4261 7531
rect 4261 7497 4295 7531
rect 4295 7497 4304 7531
rect 4252 7488 4304 7497
rect 4988 7488 5040 7540
rect 5172 7531 5224 7540
rect 5172 7497 5181 7531
rect 5181 7497 5215 7531
rect 5215 7497 5224 7531
rect 5172 7488 5224 7497
rect 6460 7488 6512 7540
rect 6828 7531 6880 7540
rect 6828 7497 6837 7531
rect 6837 7497 6871 7531
rect 6871 7497 6880 7531
rect 6828 7488 6880 7497
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 7840 7488 7892 7497
rect 8116 7488 8168 7540
rect 17040 7488 17092 7540
rect 19064 7488 19116 7540
rect 21364 7488 21416 7540
rect 21640 7531 21692 7540
rect 21640 7497 21649 7531
rect 21649 7497 21683 7531
rect 21683 7497 21692 7531
rect 21640 7488 21692 7497
rect 25320 7531 25372 7540
rect 25320 7497 25329 7531
rect 25329 7497 25363 7531
rect 25363 7497 25372 7531
rect 25320 7488 25372 7497
rect 27068 7531 27120 7540
rect 27068 7497 27077 7531
rect 27077 7497 27111 7531
rect 27111 7497 27120 7531
rect 27068 7488 27120 7497
rect 2688 7463 2740 7472
rect 2688 7429 2697 7463
rect 2697 7429 2731 7463
rect 2731 7429 2740 7463
rect 2688 7420 2740 7429
rect 5080 7463 5132 7472
rect 5080 7429 5089 7463
rect 5089 7429 5123 7463
rect 5123 7429 5132 7463
rect 5080 7420 5132 7429
rect 3148 7395 3200 7404
rect 1584 7284 1636 7336
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 5264 7352 5316 7404
rect 7288 7352 7340 7404
rect 8300 7352 8352 7404
rect 21272 7463 21324 7472
rect 21272 7429 21281 7463
rect 21281 7429 21315 7463
rect 21315 7429 21324 7463
rect 21272 7420 21324 7429
rect 26884 7420 26936 7472
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 4252 7284 4304 7336
rect 5816 7284 5868 7336
rect 6736 7284 6788 7336
rect 7380 7284 7432 7336
rect 16304 7284 16356 7336
rect 5448 7216 5500 7268
rect 7748 7216 7800 7268
rect 16856 7216 16908 7268
rect 20168 7395 20220 7404
rect 20168 7361 20177 7395
rect 20177 7361 20211 7395
rect 20211 7361 20220 7395
rect 20168 7352 20220 7361
rect 18512 7284 18564 7336
rect 19156 7284 19208 7336
rect 19984 7327 20036 7336
rect 19984 7293 19993 7327
rect 19993 7293 20027 7327
rect 20027 7293 20036 7327
rect 19984 7284 20036 7293
rect 27068 7284 27120 7336
rect 27160 7284 27212 7336
rect 19708 7216 19760 7268
rect 1584 7191 1636 7200
rect 1584 7157 1593 7191
rect 1593 7157 1627 7191
rect 1627 7157 1636 7191
rect 1584 7148 1636 7157
rect 3792 7191 3844 7200
rect 3792 7157 3801 7191
rect 3801 7157 3835 7191
rect 3835 7157 3844 7191
rect 3792 7148 3844 7157
rect 7012 7148 7064 7200
rect 7380 7148 7432 7200
rect 8300 7148 8352 7200
rect 16396 7191 16448 7200
rect 16396 7157 16405 7191
rect 16405 7157 16439 7191
rect 16439 7157 16448 7191
rect 16396 7148 16448 7157
rect 16672 7148 16724 7200
rect 18696 7148 18748 7200
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 26884 7148 26936 7200
rect 27712 7191 27764 7200
rect 27712 7157 27721 7191
rect 27721 7157 27755 7191
rect 27755 7157 27764 7191
rect 27712 7148 27764 7157
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 2044 6987 2096 6996
rect 2044 6953 2053 6987
rect 2053 6953 2087 6987
rect 2087 6953 2096 6987
rect 2044 6944 2096 6953
rect 5264 6944 5316 6996
rect 5816 6944 5868 6996
rect 6276 6987 6328 6996
rect 6276 6953 6285 6987
rect 6285 6953 6319 6987
rect 6319 6953 6328 6987
rect 6276 6944 6328 6953
rect 7288 6987 7340 6996
rect 7288 6953 7297 6987
rect 7297 6953 7331 6987
rect 7331 6953 7340 6987
rect 7288 6944 7340 6953
rect 16856 6944 16908 6996
rect 18512 6987 18564 6996
rect 18512 6953 18521 6987
rect 18521 6953 18555 6987
rect 18555 6953 18564 6987
rect 18512 6944 18564 6953
rect 19248 6987 19300 6996
rect 19248 6953 19257 6987
rect 19257 6953 19291 6987
rect 19291 6953 19300 6987
rect 19248 6944 19300 6953
rect 19708 6987 19760 6996
rect 19708 6953 19717 6987
rect 19717 6953 19751 6987
rect 19751 6953 19760 6987
rect 19708 6944 19760 6953
rect 19984 6987 20036 6996
rect 19984 6953 19993 6987
rect 19993 6953 20027 6987
rect 20027 6953 20036 6987
rect 19984 6944 20036 6953
rect 18696 6876 18748 6928
rect 2044 6808 2096 6860
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 2504 6851 2556 6860
rect 2504 6817 2513 6851
rect 2513 6817 2547 6851
rect 2547 6817 2556 6851
rect 2504 6808 2556 6817
rect 15384 6808 15436 6860
rect 16396 6808 16448 6860
rect 19616 6876 19668 6928
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 2136 6672 2188 6724
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 26700 6647 26752 6656
rect 26700 6613 26709 6647
rect 26709 6613 26743 6647
rect 26743 6613 26752 6647
rect 26700 6604 26752 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 1492 6400 1544 6452
rect 2412 6443 2464 6452
rect 2412 6409 2421 6443
rect 2421 6409 2455 6443
rect 2455 6409 2464 6443
rect 2412 6400 2464 6409
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 5448 6400 5500 6452
rect 15384 6443 15436 6452
rect 15384 6409 15393 6443
rect 15393 6409 15427 6443
rect 15427 6409 15436 6443
rect 15384 6400 15436 6409
rect 26516 6443 26568 6452
rect 26516 6409 26525 6443
rect 26525 6409 26559 6443
rect 26559 6409 26568 6443
rect 26516 6400 26568 6409
rect 2044 6375 2096 6384
rect 2044 6341 2053 6375
rect 2053 6341 2087 6375
rect 2087 6341 2096 6375
rect 2044 6332 2096 6341
rect 5080 6332 5132 6384
rect 2412 6196 2464 6248
rect 3148 6196 3200 6248
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 1308 5720 1360 5772
rect 1400 5516 1452 5568
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 1308 5312 1360 5364
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 26608 5015 26660 5024
rect 26608 4981 26617 5015
rect 26617 4981 26651 5015
rect 26651 4981 26660 5015
rect 26608 4972 26660 4981
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2044 2932 2096 2984
rect 26424 2975 26476 2984
rect 26424 2941 26433 2975
rect 26433 2941 26467 2975
rect 26467 2941 26476 2975
rect 26424 2932 26476 2941
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 26608 2839 26660 2848
rect 26608 2805 26617 2839
rect 26617 2805 26651 2839
rect 26651 2805 26660 2839
rect 26608 2796 26660 2805
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 6552 2592 6604 2644
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 7196 2499 7248 2508
rect 7196 2465 7230 2499
rect 7230 2465 7248 2499
rect 7196 2456 7248 2465
rect 6552 2388 6604 2440
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 938 23520 994 24000
rect 2778 23520 2834 24000
rect 3330 23624 3386 23633
rect 3330 23559 3386 23568
rect 952 20602 980 23520
rect 2792 20618 2820 23520
rect 3344 22846 3372 23559
rect 4618 23520 4674 24000
rect 6550 23520 6606 24000
rect 8390 23520 8446 24000
rect 10230 23520 10286 24000
rect 12162 23520 12218 24000
rect 14002 23520 14058 24000
rect 15934 23520 15990 24000
rect 17774 23520 17830 24000
rect 19614 23520 19670 24000
rect 21546 23520 21602 24000
rect 23386 23520 23442 24000
rect 25042 23624 25098 23633
rect 25042 23559 25098 23568
rect 3514 23080 3570 23089
rect 3514 23015 3570 23024
rect 3332 22840 3384 22846
rect 3332 22782 3384 22788
rect 3528 22574 3556 23015
rect 3516 22568 3568 22574
rect 3516 22510 3568 22516
rect 2870 22400 2926 22409
rect 2870 22335 2926 22344
rect 2700 20602 2820 20618
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 2688 20596 2820 20602
rect 2740 20590 2820 20596
rect 2688 20538 2740 20544
rect 2136 20392 2188 20398
rect 2136 20334 2188 20340
rect 1952 20256 2004 20262
rect 1950 20224 1952 20233
rect 2004 20224 2006 20233
rect 1950 20159 2006 20168
rect 1676 19168 1728 19174
rect 1676 19110 1728 19116
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1688 18290 1716 19110
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1964 18222 1992 19110
rect 2042 18864 2098 18873
rect 2042 18799 2044 18808
rect 2096 18799 2098 18808
rect 2044 18770 2096 18776
rect 2148 18578 2176 20334
rect 2686 19408 2742 19417
rect 2686 19343 2742 19352
rect 2700 18970 2728 19343
rect 2688 18964 2740 18970
rect 2688 18906 2740 18912
rect 2884 18902 2912 22335
rect 3330 21856 3386 21865
rect 3330 21791 3386 21800
rect 2962 20632 3018 20641
rect 2962 20567 3018 20576
rect 2872 18896 2924 18902
rect 2792 18856 2872 18884
rect 2504 18828 2556 18834
rect 2504 18770 2556 18776
rect 2056 18550 2176 18578
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 1952 18216 2004 18222
rect 1952 18158 2004 18164
rect 1964 17898 1992 18158
rect 1872 17870 1992 17898
rect 1676 16992 1728 16998
rect 1676 16934 1728 16940
rect 1688 16794 1716 16934
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1688 16046 1716 16730
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 754 15872 810 15881
rect 754 15807 810 15816
rect 768 14482 796 15807
rect 1688 15366 1716 15982
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1872 14618 1900 17870
rect 2056 17762 2084 18550
rect 2240 18290 2268 18566
rect 2228 18284 2280 18290
rect 2228 18226 2280 18232
rect 2136 18148 2188 18154
rect 2136 18090 2188 18096
rect 1964 17734 2084 17762
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 756 14476 808 14482
rect 756 14418 808 14424
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10266 1440 11086
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1504 10010 1532 14214
rect 1584 13388 1636 13394
rect 1768 13388 1820 13394
rect 1636 13348 1716 13376
rect 1584 13330 1636 13336
rect 1688 12782 1716 13348
rect 1768 13330 1820 13336
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 1688 11898 1716 12378
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1780 11762 1808 13330
rect 1768 11756 1820 11762
rect 1768 11698 1820 11704
rect 1584 10668 1636 10674
rect 1584 10610 1636 10616
rect 1412 9982 1532 10010
rect 1412 9738 1440 9982
rect 1490 9888 1546 9897
rect 1490 9823 1546 9832
rect 1320 9710 1440 9738
rect 1320 7886 1348 9710
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1412 9518 1440 9551
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 1412 9178 1440 9454
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1398 7984 1454 7993
rect 1398 7919 1400 7928
rect 1452 7919 1454 7928
rect 1400 7890 1452 7896
rect 1308 7880 1360 7886
rect 1308 7822 1360 7828
rect 1320 5778 1348 7822
rect 1400 7744 1452 7750
rect 1400 7686 1452 7692
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1320 5370 1348 5714
rect 1412 5681 1440 7686
rect 1504 6458 1532 9823
rect 1596 7546 1624 10610
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1596 7342 1624 7482
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 1596 6361 1624 6598
rect 1582 6352 1638 6361
rect 1582 6287 1638 6296
rect 1398 5672 1454 5681
rect 1398 5607 1454 5616
rect 1400 5568 1452 5574
rect 1400 5510 1452 5516
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1412 1465 1440 5510
rect 1688 4457 1716 9318
rect 1780 8634 1808 11698
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1872 9042 1900 9318
rect 1860 9036 1912 9042
rect 1860 8978 1912 8984
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1872 8430 1900 8774
rect 1964 8634 1992 17734
rect 2148 17678 2176 18090
rect 2136 17672 2188 17678
rect 2136 17614 2188 17620
rect 2148 17338 2176 17614
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2240 16726 2268 18226
rect 2412 18216 2464 18222
rect 2412 18158 2464 18164
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2332 17134 2360 17614
rect 2320 17128 2372 17134
rect 2320 17070 2372 17076
rect 2332 16794 2360 17070
rect 2320 16788 2372 16794
rect 2320 16730 2372 16736
rect 2228 16720 2280 16726
rect 2228 16662 2280 16668
rect 2042 15872 2098 15881
rect 2042 15807 2098 15816
rect 2056 15706 2084 15807
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2042 15600 2098 15609
rect 2042 15535 2098 15544
rect 2056 15162 2084 15535
rect 2424 15162 2452 18158
rect 2516 17882 2544 18770
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2700 17882 2728 18022
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2700 17678 2728 17818
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2688 15972 2740 15978
rect 2688 15914 2740 15920
rect 2700 15502 2728 15914
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2412 15156 2464 15162
rect 2412 15098 2464 15104
rect 2516 14958 2544 15438
rect 2700 15026 2728 15438
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2504 14952 2556 14958
rect 2504 14894 2556 14900
rect 2412 14816 2464 14822
rect 2410 14784 2412 14793
rect 2464 14784 2466 14793
rect 2410 14719 2466 14728
rect 2516 14634 2544 14894
rect 2424 14606 2544 14634
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2056 13734 2084 14418
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2332 13870 2360 14214
rect 2320 13864 2372 13870
rect 2320 13806 2372 13812
rect 2044 13728 2096 13734
rect 2044 13670 2096 13676
rect 2056 13297 2084 13670
rect 2042 13288 2098 13297
rect 2042 13223 2098 13232
rect 2134 11792 2190 11801
rect 2134 11727 2190 11736
rect 2320 11756 2372 11762
rect 2148 11354 2176 11727
rect 2320 11698 2372 11704
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 2148 10674 2176 11290
rect 2332 11150 2360 11698
rect 2424 11694 2452 14606
rect 2700 14414 2728 14962
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2504 13796 2556 13802
rect 2504 13738 2556 13744
rect 2516 13326 2544 13738
rect 2504 13320 2556 13326
rect 2504 13262 2556 13268
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 11144 2372 11150
rect 2320 11086 2372 11092
rect 2424 10996 2452 11630
rect 2332 10968 2452 10996
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2134 10432 2190 10441
rect 2056 9178 2084 10406
rect 2134 10367 2190 10376
rect 2044 9172 2096 9178
rect 2044 9114 2096 9120
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2056 8090 2084 9114
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2042 7984 2098 7993
rect 2042 7919 2098 7928
rect 2056 7002 2084 7919
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2056 6390 2084 6802
rect 2148 6730 2176 10367
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2240 9110 2268 9862
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2332 8956 2360 10968
rect 2502 10568 2558 10577
rect 2502 10503 2558 10512
rect 2516 10266 2544 10503
rect 2412 10260 2464 10266
rect 2412 10202 2464 10208
rect 2504 10260 2556 10266
rect 2504 10202 2556 10208
rect 2424 9722 2452 10202
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2516 9654 2544 10202
rect 2504 9648 2556 9654
rect 2504 9590 2556 9596
rect 2240 8928 2360 8956
rect 2240 8022 2268 8928
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 2320 8424 2372 8430
rect 2320 8366 2372 8372
rect 2228 8016 2280 8022
rect 2228 7958 2280 7964
rect 2332 6866 2360 8366
rect 2424 7954 2452 8842
rect 2412 7948 2464 7954
rect 2412 7890 2464 7896
rect 2410 6896 2466 6905
rect 2320 6860 2372 6866
rect 2516 6866 2544 9590
rect 2608 9489 2636 12038
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 2700 9568 2728 11018
rect 2792 10606 2820 18856
rect 2872 18838 2924 18844
rect 2976 18680 3004 20567
rect 2884 18652 3004 18680
rect 3240 18692 3292 18698
rect 2884 14793 2912 18652
rect 3240 18634 3292 18640
rect 2962 18592 3018 18601
rect 2962 18527 3018 18536
rect 2976 15586 3004 18527
rect 3146 18320 3202 18329
rect 3146 18255 3202 18264
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 3068 16250 3096 16662
rect 3056 16244 3108 16250
rect 3056 16186 3108 16192
rect 3160 15745 3188 18255
rect 3146 15736 3202 15745
rect 3146 15671 3202 15680
rect 2976 15558 3188 15586
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2964 14816 3016 14822
rect 2870 14784 2926 14793
rect 2964 14758 3016 14764
rect 2870 14719 2926 14728
rect 2976 14414 3004 14758
rect 3068 14618 3096 15302
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 3068 14278 3096 14554
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3068 12986 3096 13330
rect 3056 12980 3108 12986
rect 3056 12922 3108 12928
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2884 9722 2912 12650
rect 3160 11354 3188 15558
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10674 3004 11086
rect 3068 10690 3096 11154
rect 3160 10810 3188 11290
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2964 10668 3016 10674
rect 3068 10662 3188 10690
rect 2964 10610 3016 10616
rect 2976 10266 3004 10610
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2976 10062 3004 10202
rect 2964 10056 3016 10062
rect 2964 9998 3016 10004
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2976 9654 3004 9998
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2872 9580 2924 9586
rect 2700 9540 2820 9568
rect 2594 9480 2650 9489
rect 2594 9415 2650 9424
rect 2792 9382 2820 9540
rect 2872 9522 2924 9528
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2884 9178 2912 9522
rect 3160 9489 3188 10662
rect 3252 9586 3280 18634
rect 3344 12714 3372 21791
rect 4066 21312 4122 21321
rect 4066 21247 4122 21256
rect 4080 20874 4108 21247
rect 4068 20868 4120 20874
rect 4068 20810 4120 20816
rect 4160 20256 4212 20262
rect 3422 20224 3478 20233
rect 3422 20159 3478 20168
rect 3988 20204 4160 20210
rect 3988 20198 4212 20204
rect 3988 20182 4200 20198
rect 3436 13274 3464 20159
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3712 19281 3740 19314
rect 3698 19272 3754 19281
rect 3698 19207 3754 19216
rect 3896 19174 3924 19654
rect 3884 19168 3936 19174
rect 3882 19136 3884 19145
rect 3936 19136 3938 19145
rect 3882 19071 3938 19080
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3698 18320 3754 18329
rect 3896 18290 3924 18566
rect 3988 18426 4016 20182
rect 4434 20088 4490 20097
rect 4434 20023 4436 20032
rect 4488 20023 4490 20032
rect 4436 19994 4488 20000
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4080 19242 4108 19858
rect 4632 19417 4660 23520
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 5632 20868 5684 20874
rect 5632 20810 5684 20816
rect 4988 20800 5040 20806
rect 4988 20742 5040 20748
rect 5000 20466 5028 20742
rect 4988 20460 5040 20466
rect 4988 20402 5040 20408
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4618 19408 4674 19417
rect 4618 19343 4674 19352
rect 4068 19236 4120 19242
rect 4068 19178 4120 19184
rect 4080 18970 4108 19178
rect 4724 18970 4752 20334
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4908 19378 4936 20198
rect 5000 20058 5028 20402
rect 5644 20058 5672 20810
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 6564 20097 6592 23520
rect 8404 23474 8432 23520
rect 8312 23446 8432 23474
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 6550 20088 6606 20097
rect 4988 20052 5040 20058
rect 4988 19994 5040 20000
rect 5632 20052 5684 20058
rect 6550 20023 6606 20032
rect 5632 19994 5684 20000
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 5276 19378 5304 19654
rect 5644 19514 5672 19994
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 4908 18816 4936 19178
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 5000 19009 5028 19110
rect 4986 19000 5042 19009
rect 4986 18935 5042 18944
rect 4908 18788 5028 18816
rect 4804 18760 4856 18766
rect 4804 18702 4856 18708
rect 3976 18420 4028 18426
rect 3976 18362 4028 18368
rect 3698 18255 3754 18264
rect 3884 18284 3936 18290
rect 3712 18222 3740 18255
rect 3884 18226 3936 18232
rect 4160 18284 4212 18290
rect 4160 18226 4212 18232
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 3700 18216 3752 18222
rect 3700 18158 3752 18164
rect 3712 17882 3740 18158
rect 3976 18080 4028 18086
rect 3976 18022 4028 18028
rect 3700 17876 3752 17882
rect 3700 17818 3752 17824
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3528 15706 3556 16526
rect 3608 16448 3660 16454
rect 3608 16390 3660 16396
rect 3620 16182 3648 16390
rect 3608 16176 3660 16182
rect 3608 16118 3660 16124
rect 3620 15706 3648 16118
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3620 15026 3648 15642
rect 3790 15328 3846 15337
rect 3790 15263 3846 15272
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3516 14884 3568 14890
rect 3516 14826 3568 14832
rect 3528 13433 3556 14826
rect 3620 14618 3648 14962
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3620 14074 3648 14554
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3620 13462 3648 14010
rect 3608 13456 3660 13462
rect 3514 13424 3570 13433
rect 3608 13398 3660 13404
rect 3514 13359 3570 13368
rect 3436 13246 3648 13274
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3528 11626 3556 12310
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3422 11384 3478 11393
rect 3528 11354 3556 11562
rect 3422 11319 3478 11328
rect 3516 11348 3568 11354
rect 3436 9636 3464 11319
rect 3516 11290 3568 11296
rect 3528 11150 3556 11290
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3620 10810 3648 13246
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 11558 3740 12582
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3608 9648 3660 9654
rect 3436 9608 3556 9636
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3424 9512 3476 9518
rect 2962 9480 3018 9489
rect 3146 9480 3202 9489
rect 3018 9450 3096 9466
rect 3018 9444 3108 9450
rect 3018 9438 3056 9444
rect 2962 9415 3018 9424
rect 3330 9480 3386 9489
rect 3146 9415 3202 9424
rect 3240 9444 3292 9450
rect 3056 9386 3108 9392
rect 3424 9454 3476 9460
rect 3330 9415 3386 9424
rect 3240 9386 3292 9392
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2688 9104 2740 9110
rect 2688 9046 2740 9052
rect 2700 8956 2728 9046
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2700 8928 2820 8956
rect 2686 8664 2742 8673
rect 2686 8599 2742 8608
rect 2700 8090 2728 8599
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 8022 2820 8928
rect 2884 8294 2912 8978
rect 2976 8634 3004 9318
rect 3252 8974 3280 9386
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3344 8498 3372 9415
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 8090 2912 8230
rect 3436 8129 3464 9454
rect 3422 8120 3478 8129
rect 2872 8084 2924 8090
rect 3422 8055 3478 8064
rect 2872 8026 2924 8032
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 2608 7546 2636 7890
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2688 7472 2740 7478
rect 2686 7440 2688 7449
rect 2740 7440 2742 7449
rect 2686 7375 2742 7384
rect 3146 7440 3202 7449
rect 3146 7375 3148 7384
rect 3200 7375 3202 7384
rect 3148 7346 3200 7352
rect 2410 6831 2466 6840
rect 2504 6860 2556 6866
rect 2320 6802 2372 6808
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2424 6458 2452 6831
rect 2504 6802 2556 6808
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2044 6384 2096 6390
rect 2044 6326 2096 6332
rect 2424 6254 2452 6394
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2516 5914 2544 6802
rect 3146 6760 3202 6769
rect 3146 6695 3202 6704
rect 3160 6458 3188 6695
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3160 6254 3188 6394
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 1674 4448 1730 4457
rect 1674 4383 1730 4392
rect 2042 4040 2098 4049
rect 2042 3975 2098 3984
rect 2056 3194 2084 3975
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 2056 2990 2084 3130
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 2689 1624 2790
rect 1582 2680 1638 2689
rect 1582 2615 1638 2624
rect 1398 1456 1454 1465
rect 1398 1391 1454 1400
rect 2700 377 2728 6054
rect 3528 5137 3556 9608
rect 3608 9590 3660 9596
rect 3620 9489 3648 9590
rect 3606 9480 3662 9489
rect 3712 9450 3740 11494
rect 3804 10742 3832 15263
rect 3988 13569 4016 18022
rect 4172 17814 4200 18226
rect 4356 17882 4384 18226
rect 4816 17882 4844 18702
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 18086 4936 18158
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4344 17876 4396 17882
rect 4344 17818 4396 17824
rect 4804 17876 4856 17882
rect 4804 17818 4856 17824
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4068 17536 4120 17542
rect 4120 17496 4200 17524
rect 4068 17478 4120 17484
rect 4172 16250 4200 17496
rect 4356 17134 4384 17818
rect 4816 17746 4844 17818
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4816 17066 4844 17682
rect 4804 17060 4856 17066
rect 4804 17002 4856 17008
rect 4816 16794 4844 17002
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4528 15972 4580 15978
rect 4528 15914 4580 15920
rect 4540 15881 4568 15914
rect 4632 15910 4660 16390
rect 4620 15904 4672 15910
rect 4526 15872 4582 15881
rect 4620 15846 4672 15852
rect 4526 15807 4582 15816
rect 4632 15609 4660 15846
rect 4618 15600 4674 15609
rect 4618 15535 4674 15544
rect 4712 15564 4764 15570
rect 4712 15506 4764 15512
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4620 15360 4672 15366
rect 4620 15302 4672 15308
rect 4066 15056 4122 15065
rect 4066 14991 4122 15000
rect 4080 14482 4108 14991
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4080 14074 4108 14418
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3974 13560 4030 13569
rect 3974 13495 4030 13504
rect 4172 13410 4200 14214
rect 4250 13696 4306 13705
rect 4250 13631 4306 13640
rect 3988 13382 4200 13410
rect 4264 13394 4292 13631
rect 4252 13388 4304 13394
rect 3884 12096 3936 12102
rect 3882 12064 3884 12073
rect 3936 12064 3938 12073
rect 3882 11999 3938 12008
rect 3988 11665 4016 13382
rect 4252 13330 4304 13336
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4080 12102 4108 12242
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 4080 11354 4108 12038
rect 4172 11393 4200 13126
rect 4264 12986 4292 13330
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4158 11384 4214 11393
rect 4068 11348 4120 11354
rect 4158 11319 4214 11328
rect 4068 11290 4120 11296
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3976 11008 4028 11014
rect 3976 10950 4028 10956
rect 3792 10736 3844 10742
rect 3792 10678 3844 10684
rect 3896 10606 3924 10950
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3896 9722 3924 10542
rect 3988 10062 4016 10950
rect 4080 10792 4108 11154
rect 4160 10804 4212 10810
rect 4080 10764 4160 10792
rect 4160 10746 4212 10752
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4068 10464 4120 10470
rect 4068 10406 4120 10412
rect 3976 10056 4028 10062
rect 3976 9998 4028 10004
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3988 9450 4016 9998
rect 4080 9926 4108 10406
rect 4068 9920 4120 9926
rect 4120 9868 4200 9874
rect 4068 9862 4200 9868
rect 4080 9846 4200 9862
rect 3606 9415 3662 9424
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3698 9344 3754 9353
rect 3620 9178 3648 9318
rect 3698 9279 3754 9288
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3712 8634 3740 9279
rect 4172 8634 4200 9846
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4264 7546 4292 10474
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 4264 7342 4292 7482
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 3792 7200 3844 7206
rect 3792 7142 3844 7148
rect 3514 5128 3570 5137
rect 3514 5063 3570 5072
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 3712 480 3740 3431
rect 3804 3369 3832 7142
rect 4356 3913 4384 15302
rect 4632 14958 4660 15302
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4632 14074 4660 14894
rect 4724 14822 4752 15506
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 14414 4752 14758
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4620 14068 4672 14074
rect 4620 14010 4672 14016
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4434 13560 4490 13569
rect 4434 13495 4490 13504
rect 4448 12617 4476 13495
rect 4434 12608 4490 12617
rect 4434 12543 4490 12552
rect 4448 8498 4476 12543
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4540 11830 4568 12378
rect 4632 12345 4660 13806
rect 4724 13433 4752 14350
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4816 13938 4844 14214
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4710 13424 4766 13433
rect 4710 13359 4766 13368
rect 4816 13326 4844 13874
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4908 12730 4936 18022
rect 5000 17785 5028 18788
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4986 17776 5042 17785
rect 4986 17711 5042 17720
rect 5000 14113 5028 17711
rect 4986 14104 5042 14113
rect 4986 14039 5042 14048
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 5000 12986 5028 13466
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4986 12744 5042 12753
rect 4908 12702 4986 12730
rect 4986 12679 5042 12688
rect 4618 12336 4674 12345
rect 4618 12271 4674 12280
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4816 11558 4844 12106
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 10198 4844 11494
rect 5000 11014 5028 12679
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4712 10124 4764 10130
rect 4712 10066 4764 10072
rect 4724 9586 4752 10066
rect 5092 9761 5120 18022
rect 5276 17814 5304 19314
rect 5736 19310 5764 19790
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 5724 19304 5776 19310
rect 5354 19272 5410 19281
rect 5724 19246 5776 19252
rect 6182 19272 6238 19281
rect 5354 19207 5410 19216
rect 5264 17808 5316 17814
rect 5264 17750 5316 17756
rect 5276 17338 5304 17750
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5368 16726 5396 19207
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5460 18630 5488 19110
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 18426 5488 18566
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5552 17882 5580 18838
rect 5736 18193 5764 19246
rect 6182 19207 6238 19216
rect 6196 18970 6224 19207
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5722 18184 5778 18193
rect 5722 18119 5778 18128
rect 5724 18080 5776 18086
rect 5724 18022 5776 18028
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5356 16720 5408 16726
rect 5408 16668 5580 16674
rect 5356 16662 5580 16668
rect 5172 16652 5224 16658
rect 5368 16646 5580 16662
rect 5172 16594 5224 16600
rect 5184 16250 5212 16594
rect 5552 16250 5580 16646
rect 5736 16425 5764 18022
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 6276 16448 6328 16454
rect 5722 16416 5778 16425
rect 6276 16390 6328 16396
rect 5722 16351 5778 16360
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5184 15570 5212 16186
rect 5816 15700 5868 15706
rect 5816 15642 5868 15648
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5276 15366 5304 15574
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5264 15360 5316 15366
rect 5264 15302 5316 15308
rect 5276 15026 5304 15302
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 12782 5212 14758
rect 5276 14618 5304 14826
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5276 14346 5304 14554
rect 5460 14482 5488 15506
rect 5632 14952 5684 14958
rect 5630 14920 5632 14929
rect 5684 14920 5686 14929
rect 5630 14855 5686 14864
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14482 5672 14758
rect 5828 14482 5856 15642
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 6288 15026 6316 16390
rect 6276 15020 6328 15026
rect 6276 14962 6328 14968
rect 5448 14476 5500 14482
rect 5448 14418 5500 14424
rect 5632 14476 5684 14482
rect 5632 14418 5684 14424
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5264 14340 5316 14346
rect 5264 14282 5316 14288
rect 5354 14104 5410 14113
rect 5644 14074 5672 14418
rect 5354 14039 5410 14048
rect 5632 14068 5684 14074
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5276 12850 5304 13126
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5172 12776 5224 12782
rect 5170 12744 5172 12753
rect 5224 12744 5226 12753
rect 5368 12730 5396 14039
rect 5632 14010 5684 14016
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5644 13569 5672 13738
rect 5630 13560 5686 13569
rect 5630 13495 5632 13504
rect 5684 13495 5686 13504
rect 5632 13466 5684 13472
rect 5828 13462 5856 14418
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 6288 13938 6316 14962
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 5920 13530 5948 13738
rect 6184 13728 6236 13734
rect 6288 13716 6316 13874
rect 6236 13688 6316 13716
rect 6184 13670 6236 13676
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 6196 13326 6224 13670
rect 6274 13560 6330 13569
rect 6380 13546 6408 19450
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 7286 19136 7342 19145
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6472 17513 6500 18770
rect 6840 18329 6868 19110
rect 7286 19071 7342 19080
rect 7300 18970 7328 19071
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6826 18320 6882 18329
rect 6826 18255 6882 18264
rect 6920 18148 6972 18154
rect 6840 18108 6920 18136
rect 6840 17882 6868 18108
rect 6920 18090 6972 18096
rect 7024 18086 7052 18566
rect 7288 18284 7340 18290
rect 7288 18226 7340 18232
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 7300 17814 7328 18226
rect 7288 17808 7340 17814
rect 7288 17750 7340 17756
rect 6458 17504 6514 17513
rect 6458 17439 6514 17448
rect 6458 17096 6514 17105
rect 6458 17031 6514 17040
rect 6472 13682 6500 17031
rect 7286 16416 7342 16425
rect 7286 16351 7342 16360
rect 7300 16114 7328 16351
rect 7392 16250 7420 22510
rect 8208 20596 8260 20602
rect 8312 20584 8340 23446
rect 10244 20602 10272 23520
rect 12176 23474 12204 23520
rect 12084 23446 12204 23474
rect 10600 22840 10652 22846
rect 10600 22782 10652 22788
rect 8260 20556 8340 20584
rect 10232 20596 10284 20602
rect 8208 20538 8260 20544
rect 10232 20538 10284 20544
rect 7472 20256 7524 20262
rect 7472 20198 7524 20204
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 6642 15056 6698 15065
rect 6642 14991 6698 15000
rect 6550 14648 6606 14657
rect 6550 14583 6606 14592
rect 6564 14074 6592 14583
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6564 13870 6592 14010
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6472 13654 6592 13682
rect 6380 13518 6500 13546
rect 6274 13495 6330 13504
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 6184 13320 6236 13326
rect 6184 13262 6236 13268
rect 5170 12679 5226 12688
rect 5276 12702 5396 12730
rect 5276 12442 5304 12702
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5368 11642 5396 12582
rect 5460 12442 5488 13262
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 5448 12436 5500 12442
rect 5448 12378 5500 12384
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5722 12064 5778 12073
rect 5722 11999 5778 12008
rect 5368 11614 5672 11642
rect 5644 11558 5672 11614
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5540 11552 5592 11558
rect 5632 11552 5684 11558
rect 5540 11494 5592 11500
rect 5630 11520 5632 11529
rect 5684 11520 5686 11529
rect 5184 10713 5212 11494
rect 5552 11393 5580 11494
rect 5630 11455 5686 11464
rect 5538 11384 5594 11393
rect 5538 11319 5594 11328
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5170 10704 5226 10713
rect 5276 10674 5304 11154
rect 5170 10639 5226 10648
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5276 10266 5304 10610
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5552 10169 5580 10406
rect 5644 10305 5672 10610
rect 5630 10296 5686 10305
rect 5630 10231 5686 10240
rect 5538 10160 5594 10169
rect 5538 10095 5594 10104
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5078 9752 5134 9761
rect 5078 9687 5134 9696
rect 5644 9625 5672 9959
rect 5736 9926 5764 11999
rect 5828 11626 5856 12310
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5828 11354 5856 11562
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5828 10674 5856 11290
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5828 9994 5856 10610
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5724 9920 5776 9926
rect 5724 9862 5776 9868
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5814 9752 5870 9761
rect 5956 9744 6252 9764
rect 5814 9687 5870 9696
rect 5630 9616 5686 9625
rect 4712 9580 4764 9586
rect 5828 9586 5856 9687
rect 5630 9551 5686 9560
rect 5816 9580 5868 9586
rect 4712 9522 4764 9528
rect 5816 9522 5868 9528
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4632 8090 4660 9318
rect 4724 8906 4752 9522
rect 4986 9480 5042 9489
rect 4896 9444 4948 9450
rect 4986 9415 5042 9424
rect 4896 9386 4948 9392
rect 4908 8974 4936 9386
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 4816 8498 4844 8774
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4908 8430 4936 8910
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 5000 8090 5028 9415
rect 5356 9104 5408 9110
rect 5356 9046 5408 9052
rect 5172 8492 5224 8498
rect 5172 8434 5224 8440
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5000 7546 5028 8026
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5092 7478 5120 7686
rect 5184 7546 5212 8434
rect 5262 8392 5318 8401
rect 5262 8327 5264 8336
rect 5316 8327 5318 8336
rect 5264 8298 5316 8304
rect 5276 8022 5304 8298
rect 5368 8294 5396 9046
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 5644 8498 5672 8774
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5356 8288 5408 8294
rect 5356 8230 5408 8236
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5264 7880 5316 7886
rect 5368 7834 5396 8230
rect 5644 8090 5672 8434
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 6288 7954 6316 13495
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6380 12850 6408 13330
rect 6472 13161 6500 13518
rect 6458 13152 6514 13161
rect 6458 13087 6514 13096
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6380 11558 6408 12038
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 10470 6408 11494
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 8430 6408 10406
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6472 8090 6500 12922
rect 6564 12918 6592 13654
rect 6656 13530 6684 14991
rect 7286 14920 7342 14929
rect 7286 14855 7342 14864
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6656 12986 6684 13466
rect 6748 13326 6776 14758
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12986 6776 13262
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 6748 12730 6776 12922
rect 6564 12702 6776 12730
rect 6564 12102 6592 12702
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6748 11393 6776 12582
rect 6734 11384 6790 11393
rect 6734 11319 6790 11328
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10266 6592 10406
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6840 10146 6868 13806
rect 6932 13462 6960 14214
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 7024 12850 7052 13670
rect 7116 13190 7144 13670
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6918 12744 6974 12753
rect 6918 12679 6974 12688
rect 6932 11354 6960 12679
rect 7024 11354 7052 12786
rect 7116 11642 7144 13126
rect 7208 12238 7236 13398
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 11898 7236 12174
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7116 11614 7236 11642
rect 7104 11552 7156 11558
rect 7104 11494 7156 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 7116 11121 7144 11494
rect 7102 11112 7158 11121
rect 7102 11047 7158 11056
rect 7012 11008 7064 11014
rect 7208 10962 7236 11614
rect 7012 10950 7064 10956
rect 7024 10849 7052 10950
rect 7116 10934 7236 10962
rect 7010 10840 7066 10849
rect 7010 10775 7066 10784
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6748 10118 6868 10146
rect 6932 10130 6960 10474
rect 7024 10266 7052 10775
rect 7012 10260 7064 10266
rect 7012 10202 7064 10208
rect 6920 10124 6972 10130
rect 6552 8424 6604 8430
rect 6552 8366 6604 8372
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 5316 7828 5396 7834
rect 5264 7822 5396 7828
rect 5276 7806 5396 7822
rect 5816 7812 5868 7818
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5092 6390 5120 7414
rect 5276 7410 5304 7806
rect 5816 7754 5868 7760
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 7002 5304 7346
rect 5828 7342 5856 7754
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 5816 7336 5868 7342
rect 5816 7278 5868 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5460 6458 5488 7210
rect 5828 7002 5856 7278
rect 6288 7002 6316 7890
rect 6472 7546 6500 8026
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6288 6769 6316 6938
rect 6274 6760 6330 6769
rect 6274 6695 6330 6704
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5080 6384 5132 6390
rect 5080 6326 5132 6332
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 3790 3360 3846 3369
rect 3790 3295 3846 3304
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 6564 2650 6592 8366
rect 6748 7342 6776 10118
rect 6920 10066 6972 10072
rect 6932 10010 6960 10066
rect 6840 9982 6960 10010
rect 6840 9518 6868 9982
rect 7024 9722 7052 10202
rect 7012 9716 7064 9722
rect 7012 9658 7064 9664
rect 7010 9616 7066 9625
rect 7010 9551 7066 9560
rect 6828 9512 6880 9518
rect 6828 9454 6880 9460
rect 7024 9382 7052 9551
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 8968 6972 8974
rect 6840 8928 6920 8956
rect 6840 7546 6868 8928
rect 6920 8910 6972 8916
rect 6920 8832 6972 8838
rect 7024 8786 7052 9318
rect 6972 8780 7052 8786
rect 6920 8774 7052 8780
rect 6932 8758 7052 8774
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 6932 6905 6960 8758
rect 7116 7528 7144 10934
rect 7196 9444 7248 9450
rect 7196 9386 7248 9392
rect 7208 9178 7236 9386
rect 7196 9172 7248 9178
rect 7196 9114 7248 9120
rect 7300 8922 7328 14855
rect 7378 13016 7434 13025
rect 7378 12951 7434 12960
rect 7392 12782 7420 12951
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7484 10810 7512 20198
rect 7746 19000 7802 19009
rect 7746 18935 7748 18944
rect 7800 18935 7802 18944
rect 7748 18906 7800 18912
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7668 18358 7696 18770
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7668 17882 7696 18294
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7760 17814 7788 18906
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 7852 18154 7880 18702
rect 9036 18692 9088 18698
rect 9036 18634 9088 18640
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 7930 18184 7986 18193
rect 7840 18148 7892 18154
rect 7930 18119 7986 18128
rect 7840 18090 7892 18096
rect 7748 17808 7800 17814
rect 7748 17750 7800 17756
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 17134 7880 17478
rect 7944 17338 7972 18119
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 8128 17270 8156 18294
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8300 18148 8352 18154
rect 8220 18108 8300 18136
rect 8116 17264 8168 17270
rect 8116 17206 8168 17212
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7944 16794 7972 16934
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 8128 16726 8156 17206
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8116 16584 8168 16590
rect 8116 16526 8168 16532
rect 8128 16250 8156 16526
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 7562 15872 7618 15881
rect 7562 15807 7618 15816
rect 7576 11898 7604 15807
rect 7930 15736 7986 15745
rect 7930 15671 7986 15680
rect 7944 15162 7972 15671
rect 8128 15609 8156 16186
rect 8220 15706 8248 18108
rect 8300 18090 8352 18096
rect 8680 18086 8708 18226
rect 8956 18154 8984 18566
rect 8944 18148 8996 18154
rect 8944 18090 8996 18096
rect 9048 18086 9076 18634
rect 9692 18222 9720 18770
rect 9312 18216 9364 18222
rect 9680 18216 9732 18222
rect 9312 18158 9364 18164
rect 9678 18184 9680 18193
rect 9732 18184 9734 18193
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 8300 17740 8352 17746
rect 8300 17682 8352 17688
rect 8312 16726 8340 17682
rect 8680 17678 8708 18022
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8668 17672 8720 17678
rect 8668 17614 8720 17620
rect 8496 17066 8524 17614
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8496 16794 8524 17002
rect 8680 16998 8708 17614
rect 8942 17232 8998 17241
rect 8942 17167 8998 17176
rect 9128 17196 9180 17202
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8300 16040 8352 16046
rect 8300 15982 8352 15988
rect 8208 15700 8260 15706
rect 8208 15642 8260 15648
rect 8114 15600 8170 15609
rect 8114 15535 8170 15544
rect 8312 15366 8340 15982
rect 8680 15978 8708 16934
rect 8852 16584 8904 16590
rect 8852 16526 8904 16532
rect 8668 15972 8720 15978
rect 8668 15914 8720 15920
rect 8864 15910 8892 16526
rect 8852 15904 8904 15910
rect 8852 15846 8904 15852
rect 8390 15736 8446 15745
rect 8390 15671 8392 15680
rect 8444 15671 8446 15680
rect 8392 15642 8444 15648
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8392 15428 8444 15434
rect 8392 15370 8444 15376
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 7932 15156 7984 15162
rect 7760 15116 7932 15144
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 12850 7696 13330
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7668 12170 7696 12786
rect 7656 12164 7708 12170
rect 7656 12106 7708 12112
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7760 11098 7788 15116
rect 7932 15098 7984 15104
rect 8312 15042 8340 15302
rect 8220 15014 8340 15042
rect 8220 14958 8248 15014
rect 8404 14958 8432 15370
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 8392 14952 8444 14958
rect 8588 14906 8616 15438
rect 8392 14894 8444 14900
rect 8298 14784 8354 14793
rect 8298 14719 8354 14728
rect 8312 14482 8340 14719
rect 8404 14618 8432 14894
rect 8496 14890 8616 14906
rect 8484 14884 8616 14890
rect 8536 14878 8616 14884
rect 8484 14826 8536 14832
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 11354 8064 14214
rect 8312 14074 8340 14418
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8312 13841 8340 14010
rect 8298 13832 8354 13841
rect 8298 13767 8354 13776
rect 8392 13728 8444 13734
rect 8392 13670 8444 13676
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8312 12102 8340 12650
rect 8404 12442 8432 13670
rect 8484 13184 8536 13190
rect 8484 13126 8536 13132
rect 8496 12782 8524 13126
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8300 12096 8352 12102
rect 8128 12044 8300 12050
rect 8128 12038 8352 12044
rect 8128 12022 8340 12038
rect 8024 11348 8076 11354
rect 8024 11290 8076 11296
rect 7576 11070 7788 11098
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 7392 9586 7420 9862
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 9110 7420 9522
rect 7380 9104 7432 9110
rect 7380 9046 7432 9052
rect 7576 9042 7604 11070
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10470 7696 10950
rect 7746 10704 7802 10713
rect 7746 10639 7802 10648
rect 7760 10606 7788 10639
rect 7748 10600 7800 10606
rect 7748 10542 7800 10548
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10198 7696 10406
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7760 10062 7788 10542
rect 8036 10266 8064 11290
rect 8128 10674 8156 12022
rect 8404 11694 8432 12378
rect 8588 12209 8616 14878
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13870 8708 14350
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8574 12200 8630 12209
rect 8680 12170 8708 13806
rect 8864 13546 8892 15846
rect 8956 14618 8984 17167
rect 9128 17138 9180 17144
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9048 15366 9076 16934
rect 9140 16794 9168 17138
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 9324 16289 9352 18158
rect 9678 18119 9734 18128
rect 9588 18080 9640 18086
rect 9640 18040 9720 18068
rect 9588 18022 9640 18028
rect 9692 16794 9720 18040
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9588 16720 9640 16726
rect 9640 16668 9720 16674
rect 9588 16662 9720 16668
rect 9600 16646 9720 16662
rect 9310 16280 9366 16289
rect 9692 16250 9720 16646
rect 9310 16215 9366 16224
rect 9680 16244 9732 16250
rect 9036 15360 9088 15366
rect 9036 15302 9088 15308
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 8956 14074 8984 14554
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 8956 13705 8984 14010
rect 9048 13802 9076 15302
rect 9036 13796 9088 13802
rect 9036 13738 9088 13744
rect 8942 13696 8998 13705
rect 8942 13631 8998 13640
rect 8864 13518 8984 13546
rect 8574 12135 8630 12144
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8680 11762 8708 12106
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8482 11520 8538 11529
rect 8220 11218 8248 11494
rect 8404 11257 8432 11494
rect 8482 11455 8538 11464
rect 8496 11354 8524 11455
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8390 11248 8446 11257
rect 8208 11212 8260 11218
rect 8390 11183 8446 11192
rect 8208 11154 8260 11160
rect 8220 10810 8248 11154
rect 8772 11150 8800 12038
rect 8850 11384 8906 11393
rect 8850 11319 8852 11328
rect 8904 11319 8906 11328
rect 8852 11290 8904 11296
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8312 10742 8340 11086
rect 8300 10736 8352 10742
rect 8300 10678 8352 10684
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8128 9722 8156 10066
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7300 8894 7512 8922
rect 7380 8832 7432 8838
rect 7380 8774 7432 8780
rect 7392 8401 7420 8774
rect 7378 8392 7434 8401
rect 7288 8356 7340 8362
rect 7378 8327 7434 8336
rect 7288 8298 7340 8304
rect 7300 7886 7328 8298
rect 7484 8090 7512 8894
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7576 7886 7604 8978
rect 7840 8968 7892 8974
rect 7840 8910 7892 8916
rect 8208 8968 8260 8974
rect 8208 8910 8260 8916
rect 7852 8634 7880 8910
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8220 8566 8248 8910
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7288 7880 7340 7886
rect 7564 7880 7616 7886
rect 7288 7822 7340 7828
rect 7562 7848 7564 7857
rect 7616 7848 7618 7857
rect 7024 7500 7144 7528
rect 7024 7449 7052 7500
rect 7010 7440 7066 7449
rect 7300 7410 7328 7822
rect 7562 7783 7618 7792
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7010 7375 7066 7384
rect 7288 7404 7340 7410
rect 7024 7206 7052 7375
rect 7288 7346 7340 7352
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 6918 6896 6974 6905
rect 6918 6831 6974 6840
rect 7024 6746 7052 7142
rect 7300 7002 7328 7346
rect 7392 7342 7420 7373
rect 7380 7336 7432 7342
rect 7378 7304 7380 7313
rect 7432 7304 7434 7313
rect 7760 7274 7788 7686
rect 7852 7546 7880 8026
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 8128 7546 8156 7958
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8312 7410 8340 7822
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 7378 7239 7434 7248
rect 7748 7268 7800 7274
rect 7392 7206 7420 7239
rect 7748 7210 7800 7216
rect 8312 7206 8340 7346
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 6932 6718 7052 6746
rect 6932 6662 6960 6718
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 4049 6960 6598
rect 6918 4040 6974 4049
rect 6918 3975 6974 3984
rect 8312 2650 8340 7142
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 6564 2446 6592 2586
rect 8404 2553 8432 9862
rect 8956 9654 8984 13518
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8390 2544 8446 2553
rect 7196 2508 7248 2514
rect 8390 2479 8446 2488
rect 7196 2450 7248 2456
rect 6552 2440 6604 2446
rect 7208 2417 7236 2450
rect 6552 2382 6604 2388
rect 7194 2408 7250 2417
rect 7194 2343 7250 2352
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 9048 921 9076 10406
rect 9324 10130 9352 16215
rect 9680 16186 9732 16192
rect 9496 15972 9548 15978
rect 9496 15914 9548 15920
rect 9508 15162 9536 15914
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9680 14408 9732 14414
rect 9600 14368 9680 14396
rect 9600 13462 9628 14368
rect 9680 14350 9732 14356
rect 9784 14346 9812 20198
rect 9862 19408 9918 19417
rect 9862 19343 9918 19352
rect 9876 18970 9904 19343
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 10612 18426 10640 22782
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 10782 19952 10838 19961
rect 10782 19887 10838 19896
rect 10796 19174 10824 19887
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19310 10916 19654
rect 12084 19417 12112 23446
rect 14016 21146 14044 23520
rect 15948 23474 15976 23520
rect 15856 23446 15976 23474
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 12164 21004 12216 21010
rect 12164 20946 12216 20952
rect 12176 20534 12204 20946
rect 12716 20800 12768 20806
rect 12716 20742 12768 20748
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12728 20466 12756 20742
rect 15856 20602 15884 23446
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 16580 21004 16632 21010
rect 16580 20946 16632 20952
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19990 12296 20198
rect 12728 20058 12756 20402
rect 13636 20392 13688 20398
rect 13820 20392 13872 20398
rect 13636 20334 13688 20340
rect 13740 20340 13820 20346
rect 13740 20334 13872 20340
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12256 19984 12308 19990
rect 12820 19961 12848 20266
rect 12256 19926 12308 19932
rect 12806 19952 12862 19961
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12070 19408 12126 19417
rect 12176 19378 12204 19790
rect 12070 19343 12126 19352
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 10876 19304 10928 19310
rect 10876 19246 10928 19252
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 10784 18624 10836 18630
rect 10784 18566 10836 18572
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10612 18222 10640 18362
rect 10796 18329 10824 18566
rect 10888 18426 10916 19246
rect 11336 19236 11388 19242
rect 11336 19178 11388 19184
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 11348 18970 11376 19178
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11334 18728 11390 18737
rect 11334 18663 11390 18672
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10782 18320 10838 18329
rect 10782 18255 10838 18264
rect 10876 18284 10928 18290
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10796 18086 10824 18255
rect 10876 18226 10928 18232
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 9862 17640 9918 17649
rect 9862 17575 9918 17584
rect 9876 16697 9904 17575
rect 9956 17536 10008 17542
rect 9956 17478 10008 17484
rect 9968 16794 9996 17478
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9862 16688 9918 16697
rect 9862 16623 9918 16632
rect 9864 16584 9916 16590
rect 9864 16526 9916 16532
rect 9876 16250 9904 16526
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9968 15706 9996 16730
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 9956 14272 10008 14278
rect 9956 14214 10008 14220
rect 9968 13870 9996 14214
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9692 12220 9720 13670
rect 9772 12232 9824 12238
rect 9692 12192 9772 12220
rect 9772 12174 9824 12180
rect 9784 11898 9812 12174
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 10060 11801 10088 18022
rect 10888 17882 10916 18226
rect 11152 18216 11204 18222
rect 11150 18184 11152 18193
rect 11204 18184 11206 18193
rect 11150 18119 11206 18128
rect 11348 18086 11376 18663
rect 11440 18290 11468 18770
rect 11900 18630 11928 19110
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11428 18284 11480 18290
rect 11428 18226 11480 18232
rect 11900 18154 11928 18566
rect 12268 18426 12296 19926
rect 12348 19916 12400 19922
rect 12806 19887 12862 19896
rect 12348 19858 12400 19864
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12360 18306 12388 19858
rect 13648 19514 13676 20334
rect 13740 20318 13860 20334
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18698 12572 19246
rect 13636 18760 13688 18766
rect 13636 18702 13688 18708
rect 12532 18692 12584 18698
rect 12532 18634 12584 18640
rect 13084 18692 13136 18698
rect 13084 18634 13136 18640
rect 12360 18278 12480 18306
rect 13096 18290 13124 18634
rect 11888 18148 11940 18154
rect 11888 18090 11940 18096
rect 11336 18080 11388 18086
rect 11336 18022 11388 18028
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 11612 17672 11664 17678
rect 11612 17614 11664 17620
rect 10600 17604 10652 17610
rect 10600 17546 10652 17552
rect 10612 17338 10640 17546
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 11440 17202 11468 17478
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 11624 16998 11652 17614
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10324 16720 10376 16726
rect 10324 16662 10376 16668
rect 10506 16688 10562 16697
rect 10336 15910 10364 16662
rect 10506 16623 10562 16632
rect 10784 16652 10836 16658
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 14929 10364 15846
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15065 10456 15438
rect 10414 15056 10470 15065
rect 10414 14991 10416 15000
rect 10468 14991 10470 15000
rect 10416 14962 10468 14968
rect 10322 14920 10378 14929
rect 10322 14855 10378 14864
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10244 13530 10272 14350
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 10244 12374 10272 12582
rect 10232 12368 10284 12374
rect 10232 12310 10284 12316
rect 10046 11792 10102 11801
rect 10046 11727 10102 11736
rect 10244 11286 10272 12310
rect 10520 11694 10548 16623
rect 10784 16594 10836 16600
rect 10796 16425 10824 16594
rect 11428 16448 11480 16454
rect 10782 16416 10838 16425
rect 10782 16351 10838 16360
rect 11150 16416 11206 16425
rect 11428 16390 11480 16396
rect 11150 16351 11206 16360
rect 11164 16046 11192 16351
rect 11440 16114 11468 16390
rect 11518 16144 11574 16153
rect 11428 16108 11480 16114
rect 11518 16079 11574 16088
rect 11428 16050 11480 16056
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 10600 15904 10652 15910
rect 10598 15872 10600 15881
rect 10652 15872 10654 15881
rect 10598 15807 10654 15816
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 11440 15706 11468 16050
rect 11532 15910 11560 16079
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14618 10824 14758
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10888 14521 10916 15642
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 11152 14544 11204 14550
rect 10874 14512 10930 14521
rect 11152 14486 11204 14492
rect 10874 14447 10876 14456
rect 10928 14447 10930 14456
rect 10876 14418 10928 14424
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10612 13326 10640 13806
rect 10782 13560 10838 13569
rect 10888 13546 10916 14418
rect 11164 14346 11192 14486
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11164 14074 11192 14282
rect 11348 14278 11376 14962
rect 11440 14822 11468 15302
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11428 14476 11480 14482
rect 11532 14464 11560 14826
rect 11480 14436 11560 14464
rect 11428 14418 11480 14424
rect 11336 14272 11388 14278
rect 11334 14240 11336 14249
rect 11388 14240 11390 14249
rect 11334 14175 11390 14184
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11164 13716 11192 14010
rect 11348 13938 11376 14175
rect 11336 13932 11388 13938
rect 11336 13874 11388 13880
rect 11440 13802 11468 14418
rect 11428 13796 11480 13802
rect 11428 13738 11480 13744
rect 11164 13688 11376 13716
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 10838 13518 10916 13546
rect 11348 13530 11376 13688
rect 11336 13524 11388 13530
rect 10782 13495 10838 13504
rect 11336 13466 11388 13472
rect 11060 13388 11112 13394
rect 11060 13330 11112 13336
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10612 12850 10640 13262
rect 11072 12918 11100 13330
rect 11336 12980 11388 12986
rect 11336 12922 11388 12928
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11060 12912 11112 12918
rect 10888 12860 11060 12866
rect 10888 12854 11112 12860
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10888 12838 11100 12854
rect 10888 11898 10916 12838
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10232 11280 10284 11286
rect 10232 11222 10284 11228
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 10152 10849 10180 11086
rect 10138 10840 10194 10849
rect 10336 10810 10364 11494
rect 10612 11218 10640 11591
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 11348 11354 11376 12922
rect 11428 12096 11480 12102
rect 11428 12038 11480 12044
rect 11440 11762 11468 12038
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10690 11248 10746 11257
rect 10600 11212 10652 11218
rect 10690 11183 10746 11192
rect 10600 11154 10652 11160
rect 10138 10775 10140 10784
rect 10192 10775 10194 10784
rect 10324 10804 10376 10810
rect 10140 10746 10192 10752
rect 10324 10746 10376 10752
rect 10612 10606 10640 11154
rect 10704 11150 10732 11183
rect 10692 11144 10744 11150
rect 10692 11086 10744 11092
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 10600 10600 10652 10606
rect 10322 10568 10378 10577
rect 10600 10542 10652 10548
rect 10784 10600 10836 10606
rect 10784 10542 10836 10548
rect 10322 10503 10378 10512
rect 10336 10470 10364 10503
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 10305 10364 10406
rect 10322 10296 10378 10305
rect 10322 10231 10324 10240
rect 10376 10231 10378 10240
rect 10324 10202 10376 10208
rect 10796 10169 10824 10542
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 11348 10266 11376 10610
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10782 10160 10838 10169
rect 9312 10124 9364 10130
rect 10782 10095 10784 10104
rect 9312 10066 9364 10072
rect 10836 10095 10838 10104
rect 10784 10066 10836 10072
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9140 8809 9168 9590
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 9126 8800 9182 8809
rect 9126 8735 9182 8744
rect 9140 7818 9168 8735
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 11532 7993 11560 12922
rect 11624 11257 11652 16934
rect 11900 16726 11928 18090
rect 11978 17776 12034 17785
rect 11978 17711 12034 17720
rect 12072 17740 12124 17746
rect 11992 17338 12020 17711
rect 12072 17682 12124 17688
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11992 17066 12020 17274
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 12084 16998 12112 17682
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11900 15910 11928 16662
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15502 11928 15846
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 14890 11928 15438
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 13530 11836 14758
rect 11796 13524 11848 13530
rect 11796 13466 11848 13472
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11900 12102 11928 13194
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11704 11824 11756 11830
rect 11704 11766 11756 11772
rect 11610 11248 11666 11257
rect 11610 11183 11666 11192
rect 11716 11150 11744 11766
rect 11900 11218 11928 12038
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11716 10810 11744 11086
rect 11900 10810 11928 11154
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11992 10713 12020 12854
rect 12084 11665 12112 16934
rect 12176 16658 12204 17614
rect 12452 17338 12480 18278
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12544 17542 12572 18090
rect 12992 18080 13044 18086
rect 12990 18048 12992 18057
rect 13044 18048 13046 18057
rect 12990 17983 13046 17992
rect 13096 17882 13124 18226
rect 13648 18086 13676 18702
rect 13636 18080 13688 18086
rect 13636 18022 13688 18028
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12176 16250 12204 16594
rect 12346 16280 12402 16289
rect 12164 16244 12216 16250
rect 12544 16266 12572 17478
rect 13096 17338 13124 17818
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12402 16238 12572 16266
rect 12346 16215 12402 16224
rect 12164 16186 12216 16192
rect 12544 15881 12572 16238
rect 12530 15872 12586 15881
rect 12530 15807 12586 15816
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15178 12296 15302
rect 12268 15150 12480 15178
rect 12544 15162 12572 15506
rect 12268 14958 12296 15150
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12254 13560 12310 13569
rect 12254 13495 12256 13504
rect 12308 13495 12310 13504
rect 12256 13466 12308 13472
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 12176 13161 12204 13330
rect 12162 13152 12218 13161
rect 12162 13087 12218 13096
rect 12176 12918 12204 13087
rect 12268 12986 12296 13466
rect 12452 12986 12480 15150
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12544 14618 12572 15098
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12162 12744 12218 12753
rect 12162 12679 12164 12688
rect 12216 12679 12218 12688
rect 12164 12650 12216 12656
rect 12728 12306 12756 16934
rect 13096 16794 13124 17274
rect 13542 17232 13598 17241
rect 13542 17167 13598 17176
rect 13556 16794 13584 17167
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13360 15904 13412 15910
rect 12898 15872 12954 15881
rect 13360 15846 13412 15852
rect 12898 15807 12954 15816
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 12782 12848 13466
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12912 12442 12940 15807
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13280 13802 13308 14214
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13280 13462 13308 13738
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13280 13258 13308 13398
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13280 12850 13308 13194
rect 13372 13161 13400 15846
rect 13648 15201 13676 18022
rect 13740 17882 13768 20318
rect 16592 20262 16620 20946
rect 17788 20602 17816 23520
rect 19628 21146 19656 23520
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 17960 21072 18012 21078
rect 17960 21014 18012 21020
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17972 20534 18000 21014
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18512 20936 18564 20942
rect 18512 20878 18564 20884
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 16764 20392 16816 20398
rect 16764 20334 16816 20340
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 15752 19916 15804 19922
rect 16592 19904 16620 20198
rect 16776 20058 16804 20334
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 15752 19858 15804 19864
rect 16408 19876 16620 19904
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13832 18970 13860 19450
rect 14936 19446 14964 19654
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14924 19440 14976 19446
rect 14924 19382 14976 19388
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14280 18964 14332 18970
rect 14280 18906 14332 18912
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13924 17814 13952 18770
rect 14096 18760 14148 18766
rect 14094 18728 14096 18737
rect 14148 18728 14150 18737
rect 14094 18663 14150 18672
rect 14292 18222 14320 18906
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 13820 17740 13872 17746
rect 13820 17682 13872 17688
rect 13832 16658 13860 17682
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 17338 14228 17614
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14292 16794 14320 17818
rect 14568 16998 14596 19382
rect 15212 19378 15240 19858
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14924 19168 14976 19174
rect 14924 19110 14976 19116
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14648 18148 14700 18154
rect 14648 18090 14700 18096
rect 14660 17814 14688 18090
rect 14936 17882 14964 19110
rect 14924 17876 14976 17882
rect 14924 17818 14976 17824
rect 14648 17808 14700 17814
rect 14648 17750 14700 17756
rect 14660 17270 14688 17750
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14556 16992 14608 16998
rect 14556 16934 14608 16940
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 13820 16652 13872 16658
rect 13740 16612 13820 16640
rect 13634 15192 13690 15201
rect 13740 15162 13768 16612
rect 13820 16594 13872 16600
rect 13924 16538 13952 16730
rect 13832 16510 13952 16538
rect 13832 16046 13860 16510
rect 13912 16176 13964 16182
rect 13912 16118 13964 16124
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13634 15127 13690 15136
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13832 15094 13860 15302
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13740 14890 13768 14962
rect 13832 14958 13860 15030
rect 13924 15026 13952 16118
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13728 14884 13780 14890
rect 13728 14826 13780 14832
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14618 13584 14758
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13924 14550 13952 14962
rect 13912 14544 13964 14550
rect 13912 14486 13964 14492
rect 13728 14408 13780 14414
rect 13728 14350 13780 14356
rect 13542 13832 13598 13841
rect 13542 13767 13598 13776
rect 13556 13462 13584 13767
rect 13740 13530 13768 14350
rect 13818 14240 13874 14249
rect 13818 14175 13874 14184
rect 13832 14074 13860 14175
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13544 13456 13596 13462
rect 13544 13398 13596 13404
rect 14094 13424 14150 13433
rect 13358 13152 13414 13161
rect 13358 13087 13414 13096
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12716 12300 12768 12306
rect 12716 12242 12768 12248
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12176 11830 12204 12174
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 12544 11354 12572 12038
rect 12728 11830 12756 12242
rect 12716 11824 12768 11830
rect 12716 11766 12768 11772
rect 12912 11762 12940 12378
rect 12990 12336 13046 12345
rect 12990 12271 12992 12280
rect 13044 12271 13046 12280
rect 12992 12242 13044 12248
rect 12990 12200 13046 12209
rect 12990 12135 13046 12144
rect 13004 11762 13032 12135
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13004 11354 13032 11698
rect 13268 11552 13320 11558
rect 13266 11520 13268 11529
rect 13320 11520 13322 11529
rect 13266 11455 13322 11464
rect 12532 11348 12584 11354
rect 12532 11290 12584 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12164 11076 12216 11082
rect 12164 11018 12216 11024
rect 12176 10810 12204 11018
rect 12544 10810 12572 11290
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 11978 10704 12034 10713
rect 11978 10639 12034 10648
rect 11518 7984 11574 7993
rect 11518 7919 11574 7928
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 13372 5137 13400 13087
rect 13556 12986 13584 13398
rect 14094 13359 14096 13368
rect 14148 13359 14150 13368
rect 14096 13330 14148 13336
rect 14108 12986 14136 13330
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 13634 12880 13690 12889
rect 13634 12815 13690 12824
rect 13648 11694 13676 12815
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13832 9081 13860 12922
rect 13818 9072 13874 9081
rect 13818 9007 13874 9016
rect 14384 7585 14412 15302
rect 14568 14890 14596 16934
rect 15028 16250 15056 19110
rect 15212 17882 15240 19314
rect 15304 19310 15332 19654
rect 15292 19304 15344 19310
rect 15764 19281 15792 19858
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15292 19246 15344 19252
rect 15750 19272 15806 19281
rect 15304 18970 15332 19246
rect 15750 19207 15806 19216
rect 15764 19174 15792 19207
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15476 18080 15528 18086
rect 15476 18022 15528 18028
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 15120 16590 15148 17138
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15120 16182 15148 16526
rect 15108 16176 15160 16182
rect 15108 16118 15160 16124
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14752 15706 14780 16050
rect 14740 15700 14792 15706
rect 14740 15642 14792 15648
rect 14752 15094 14780 15642
rect 15120 15570 15148 16118
rect 15488 16046 15516 18022
rect 15764 16153 15792 19110
rect 15856 18970 15884 19790
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 15844 18964 15896 18970
rect 15844 18906 15896 18912
rect 15856 16726 15884 18906
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15750 16144 15806 16153
rect 15856 16114 15884 16662
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15750 16079 15806 16088
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15566 16008 15622 16017
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15609 15424 15846
rect 15488 15638 15516 15982
rect 15566 15943 15622 15952
rect 15580 15910 15608 15943
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15476 15632 15528 15638
rect 15382 15600 15438 15609
rect 15108 15564 15160 15570
rect 15476 15574 15528 15580
rect 15382 15535 15438 15544
rect 15108 15506 15160 15512
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14738 14920 14794 14929
rect 14556 14884 14608 14890
rect 14738 14855 14794 14864
rect 14556 14826 14608 14832
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14657 14504 14758
rect 14462 14648 14518 14657
rect 14462 14583 14518 14592
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 14476 14074 14504 14486
rect 14752 14074 14780 14855
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 14385 15056 14758
rect 15120 14482 15148 15506
rect 15488 15026 15516 15574
rect 15580 15366 15608 15846
rect 15856 15706 15884 16050
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16028 15088 16080 15094
rect 16026 15056 16028 15065
rect 16080 15056 16082 15065
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15476 15020 15528 15026
rect 16026 14991 16082 15000
rect 15476 14962 15528 14968
rect 15108 14476 15160 14482
rect 15108 14418 15160 14424
rect 15212 14414 15240 14962
rect 15488 14550 15516 14962
rect 16040 14958 16068 14991
rect 16028 14952 16080 14958
rect 16028 14894 16080 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 15476 14544 15528 14550
rect 15672 14521 15700 14758
rect 16224 14618 16252 14758
rect 16212 14612 16264 14618
rect 16264 14572 16344 14600
rect 16212 14554 16264 14560
rect 15844 14544 15896 14550
rect 15476 14486 15528 14492
rect 15658 14512 15714 14521
rect 15200 14408 15252 14414
rect 15014 14376 15070 14385
rect 15200 14350 15252 14356
rect 15014 14311 15070 14320
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 15488 13938 15516 14486
rect 15844 14486 15896 14492
rect 15658 14447 15714 14456
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15764 14074 15792 14350
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15856 14006 15884 14486
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 16316 14074 16344 14572
rect 16304 14068 16356 14074
rect 16304 14010 16356 14016
rect 15844 14000 15896 14006
rect 15844 13942 15896 13948
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15108 13728 15160 13734
rect 15108 13670 15160 13676
rect 14464 13320 14516 13326
rect 14464 13262 14516 13268
rect 14476 12646 14504 13262
rect 15120 13190 15148 13670
rect 15292 13252 15344 13258
rect 15292 13194 15344 13200
rect 15108 13184 15160 13190
rect 15108 13126 15160 13132
rect 14464 12640 14516 12646
rect 15120 12617 15148 13126
rect 15304 12850 15332 13194
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15200 12640 15252 12646
rect 14464 12582 14516 12588
rect 14922 12608 14978 12617
rect 14476 12170 14504 12582
rect 14922 12543 14978 12552
rect 15106 12608 15162 12617
rect 15200 12582 15252 12588
rect 15106 12543 15162 12552
rect 14832 12232 14884 12238
rect 14936 12209 14964 12543
rect 14832 12174 14884 12180
rect 14922 12200 14978 12209
rect 14464 12164 14516 12170
rect 14464 12106 14516 12112
rect 14476 11762 14504 12106
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14568 11354 14596 12038
rect 14844 11898 14872 12174
rect 14922 12135 14978 12144
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14936 11286 14964 11698
rect 15212 11354 15240 12582
rect 15396 12424 15424 13874
rect 15856 13530 15884 13942
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 16302 13288 16358 13297
rect 16302 13223 16358 13232
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15844 12640 15896 12646
rect 15844 12582 15896 12588
rect 15304 12396 15424 12424
rect 15304 12209 15332 12396
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15290 12200 15346 12209
rect 15290 12135 15346 12144
rect 15304 11694 15332 12135
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15292 11552 15344 11558
rect 15396 11529 15424 12242
rect 15856 12238 15884 12582
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15292 11494 15344 11500
rect 15382 11520 15438 11529
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 15304 10810 15332 11494
rect 15382 11455 15438 11464
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15396 10742 15424 11455
rect 15672 11286 15700 12106
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15660 11280 15712 11286
rect 15660 11222 15712 11228
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15580 10742 15608 11154
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15764 10266 15792 11698
rect 15844 11688 15896 11694
rect 15842 11656 15844 11665
rect 15896 11656 15898 11665
rect 15842 11591 15898 11600
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11257 16252 11494
rect 16210 11248 16266 11257
rect 16316 11218 16344 13223
rect 16408 12986 16436 19876
rect 16764 18828 16816 18834
rect 16764 18770 16816 18776
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 16500 18154 16528 18702
rect 16776 18358 16804 18770
rect 16764 18352 16816 18358
rect 16764 18294 16816 18300
rect 16488 18148 16540 18154
rect 16488 18090 16540 18096
rect 16500 17746 16528 18090
rect 17604 17882 17632 20402
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17696 19514 17724 19994
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17684 19508 17736 19514
rect 17684 19450 17736 19456
rect 17788 19310 17816 19858
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17788 18426 17816 19246
rect 17880 19242 17908 19790
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 17868 19236 17920 19242
rect 17868 19178 17920 19184
rect 17880 18630 17908 19178
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17880 17898 17908 18566
rect 18248 18170 18276 19654
rect 18340 18290 18368 20742
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18432 18222 18460 19178
rect 18420 18216 18472 18222
rect 18248 18142 18368 18170
rect 18420 18158 18472 18164
rect 17592 17876 17644 17882
rect 17880 17870 18184 17898
rect 17592 17818 17644 17824
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16500 17202 16528 17682
rect 16960 17338 16988 17682
rect 17604 17338 17632 17818
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 16684 16794 16712 17002
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 17038 16552 17094 16561
rect 17038 16487 17094 16496
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16592 14226 16620 14826
rect 16592 14198 16712 14226
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16488 13184 16540 13190
rect 16488 13126 16540 13132
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16500 12850 16528 13126
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16500 12442 16528 12786
rect 16488 12436 16540 12442
rect 16488 12378 16540 12384
rect 16592 11778 16620 14010
rect 16500 11762 16620 11778
rect 16488 11756 16620 11762
rect 16540 11750 16620 11756
rect 16488 11698 16540 11704
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16592 11506 16620 11750
rect 16684 11642 16712 14198
rect 16856 13388 16908 13394
rect 16776 13348 16856 13376
rect 16776 12918 16804 13348
rect 16856 13330 16908 13336
rect 16960 13002 16988 14894
rect 16868 12974 16988 13002
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16776 12442 16804 12854
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16684 11614 16804 11642
rect 16408 11393 16436 11494
rect 16592 11478 16712 11506
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 16500 11257 16528 11290
rect 16486 11248 16542 11257
rect 16210 11183 16266 11192
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16408 11206 16486 11234
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16408 10266 16436 11206
rect 16486 11183 16542 11192
rect 16684 11150 16712 11478
rect 16672 11144 16724 11150
rect 16776 11121 16804 11614
rect 16672 11086 16724 11092
rect 16762 11112 16818 11121
rect 16488 11076 16540 11082
rect 16540 11036 16620 11064
rect 16762 11047 16818 11056
rect 16488 11018 16540 11024
rect 16592 10674 16620 11036
rect 16580 10668 16632 10674
rect 16580 10610 16632 10616
rect 16776 10538 16804 11047
rect 16868 10606 16896 12974
rect 17052 12186 17080 16487
rect 17604 16250 17632 17274
rect 17776 16584 17828 16590
rect 17776 16526 17828 16532
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17788 15910 17816 16526
rect 18156 16454 18184 17870
rect 18340 17649 18368 18142
rect 18326 17640 18382 17649
rect 18326 17575 18382 17584
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17406 14648 17462 14657
rect 17406 14583 17462 14592
rect 17420 14550 17448 14583
rect 17408 14544 17460 14550
rect 17408 14486 17460 14492
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17144 13734 17172 14350
rect 17420 14074 17448 14486
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13462 17172 13670
rect 17132 13456 17184 13462
rect 17132 13398 17184 13404
rect 17144 12646 17172 13398
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 17132 12640 17184 12646
rect 17132 12582 17184 12588
rect 17144 12238 17172 12582
rect 17420 12306 17448 12786
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 16960 12158 17080 12186
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 16960 11694 16988 12158
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 11762 17080 12038
rect 17144 11762 17172 12174
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 17420 11354 17448 12242
rect 17788 11694 17816 15846
rect 18064 15706 18092 16050
rect 18156 16046 18184 16390
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 17868 13388 17920 13394
rect 18064 13376 18092 14214
rect 17920 13348 18092 13376
rect 17868 13330 17920 13336
rect 17960 13184 18012 13190
rect 17960 13126 18012 13132
rect 17972 12850 18000 13126
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 18156 11506 18184 14826
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18248 13297 18276 13670
rect 18340 13569 18368 17575
rect 18524 16794 18552 20878
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18696 20256 18748 20262
rect 18696 20198 18748 20204
rect 18616 18034 18644 20198
rect 18708 19718 18736 20198
rect 18788 19780 18840 19786
rect 18788 19722 18840 19728
rect 18696 19712 18748 19718
rect 18696 19654 18748 19660
rect 18696 19168 18748 19174
rect 18696 19110 18748 19116
rect 18708 18222 18736 19110
rect 18800 18902 18828 19722
rect 18892 19310 18920 20878
rect 18880 19304 18932 19310
rect 18880 19246 18932 19252
rect 18892 18970 18920 19246
rect 18880 18964 18932 18970
rect 18880 18906 18932 18912
rect 18788 18896 18840 18902
rect 18788 18838 18840 18844
rect 18800 18290 18828 18838
rect 18892 18766 18920 18906
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18880 18352 18932 18358
rect 18880 18294 18932 18300
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18696 18216 18748 18222
rect 18696 18158 18748 18164
rect 18616 18006 18736 18034
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18616 16998 18644 17614
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18512 16788 18564 16794
rect 18512 16730 18564 16736
rect 18616 15994 18644 16934
rect 18708 16697 18736 18006
rect 18788 17536 18840 17542
rect 18892 17524 18920 18294
rect 18984 17882 19012 20946
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19260 20516 19288 20810
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 20180 20602 20208 20742
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 19340 20528 19392 20534
rect 19260 20488 19340 20516
rect 19340 20470 19392 20476
rect 20168 20392 20220 20398
rect 19982 20360 20038 20369
rect 20168 20334 20220 20340
rect 19982 20295 19984 20304
rect 20036 20295 20038 20304
rect 19984 20266 20036 20272
rect 19340 20256 19392 20262
rect 19340 20198 19392 20204
rect 19156 19848 19208 19854
rect 19156 19790 19208 19796
rect 19168 18970 19196 19790
rect 19352 19258 19380 20198
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19260 19242 19380 19258
rect 19248 19236 19380 19242
rect 19300 19230 19380 19236
rect 19248 19178 19300 19184
rect 19340 19168 19392 19174
rect 19260 19116 19340 19122
rect 19260 19110 19392 19116
rect 19260 19094 19380 19110
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19064 18828 19116 18834
rect 19064 18770 19116 18776
rect 19076 18193 19104 18770
rect 19260 18358 19288 19094
rect 19430 18864 19486 18873
rect 19430 18799 19432 18808
rect 19484 18799 19486 18808
rect 19432 18770 19484 18776
rect 19444 18426 19472 18770
rect 19628 18426 19656 19858
rect 20180 19718 20208 20334
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 21560 20058 21588 23520
rect 21732 20868 21784 20874
rect 21732 20810 21784 20816
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 20904 19916 20956 19922
rect 20904 19858 20956 19864
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20168 19712 20220 19718
rect 20168 19654 20220 19660
rect 20180 19310 20208 19654
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 19982 18728 20038 18737
rect 19982 18663 19984 18672
rect 20036 18663 20038 18672
rect 19984 18634 20036 18640
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19248 18352 19300 18358
rect 19248 18294 19300 18300
rect 19996 18193 20024 18634
rect 20180 18290 20208 19246
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20168 18284 20220 18290
rect 20168 18226 20220 18232
rect 19062 18184 19118 18193
rect 19982 18184 20038 18193
rect 19062 18119 19064 18128
rect 19116 18119 19118 18128
rect 19616 18148 19668 18154
rect 19064 18090 19116 18096
rect 19982 18119 20038 18128
rect 19616 18090 19668 18096
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19064 17604 19116 17610
rect 19064 17546 19116 17552
rect 18840 17496 18920 17524
rect 18788 17478 18840 17484
rect 18800 17134 18828 17478
rect 19076 17134 19104 17546
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18970 16960 19026 16969
rect 18970 16895 19026 16904
rect 18984 16726 19012 16895
rect 18972 16720 19024 16726
rect 18694 16688 18750 16697
rect 18972 16662 19024 16668
rect 18694 16623 18750 16632
rect 18880 16652 18932 16658
rect 18524 15966 18644 15994
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 15162 18460 15506
rect 18524 15337 18552 15966
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15570 18644 15846
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18510 15328 18566 15337
rect 18510 15263 18566 15272
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18326 13560 18382 13569
rect 18326 13495 18382 13504
rect 18234 13288 18290 13297
rect 18234 13223 18290 13232
rect 18524 12345 18552 15263
rect 18616 14890 18644 15506
rect 18604 14884 18656 14890
rect 18604 14826 18656 14832
rect 18602 13016 18658 13025
rect 18602 12951 18658 12960
rect 18616 12753 18644 12951
rect 18602 12744 18658 12753
rect 18602 12679 18658 12688
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18432 11694 18460 12038
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 17880 11478 18184 11506
rect 17682 11384 17738 11393
rect 17408 11348 17460 11354
rect 17682 11319 17738 11328
rect 17408 11290 17460 11296
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16764 10532 16816 10538
rect 16764 10474 16816 10480
rect 16868 10305 16896 10542
rect 16854 10296 16910 10305
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 16396 10260 16448 10266
rect 17696 10266 17724 11319
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17788 10810 17816 11222
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17880 10674 17908 11478
rect 18142 11384 18198 11393
rect 18432 11354 18460 11630
rect 18142 11319 18144 11328
rect 18196 11319 18198 11328
rect 18420 11348 18472 11354
rect 18144 11290 18196 11296
rect 18420 11290 18472 11296
rect 18524 11286 18552 12271
rect 18512 11280 18564 11286
rect 18512 11222 18564 11228
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 18340 10470 18368 11086
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 16854 10231 16910 10240
rect 17684 10260 17736 10266
rect 16396 10202 16448 10208
rect 17684 10202 17736 10208
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 15660 9648 15712 9654
rect 15566 9616 15622 9625
rect 15660 9590 15712 9596
rect 15566 9551 15568 9560
rect 15620 9551 15622 9560
rect 15568 9522 15620 9528
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15304 9178 15332 9386
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15672 8809 15700 9590
rect 16304 9512 16356 9518
rect 16302 9480 16304 9489
rect 16356 9480 16358 9489
rect 16302 9415 16358 9424
rect 16396 9376 16448 9382
rect 16396 9318 16448 9324
rect 16302 9208 16358 9217
rect 16302 9143 16358 9152
rect 16316 9042 16344 9143
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 15658 8800 15714 8809
rect 15658 8735 15714 8744
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16316 8634 16344 8978
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16408 8430 16436 9318
rect 16500 8498 16528 9862
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16776 9330 16804 9522
rect 16868 9489 16896 10066
rect 18340 10062 18368 10406
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17132 10056 17184 10062
rect 17132 9998 17184 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 16960 9897 16988 9998
rect 16946 9888 17002 9897
rect 16946 9823 17002 9832
rect 16960 9722 16988 9823
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 17144 9586 17172 9998
rect 18708 9625 18736 16623
rect 18880 16594 18932 16600
rect 18892 16561 18920 16594
rect 19076 16590 19104 17070
rect 19536 16658 19564 17682
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19064 16584 19116 16590
rect 18878 16552 18934 16561
rect 19064 16526 19116 16532
rect 18878 16487 18934 16496
rect 19430 16416 19486 16425
rect 19430 16351 19486 16360
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19156 14272 19208 14278
rect 19352 14226 19380 14282
rect 19156 14214 19208 14220
rect 19168 13734 19196 14214
rect 19260 14198 19380 14226
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19260 13530 19288 14198
rect 19338 14104 19394 14113
rect 19338 14039 19394 14048
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18984 12646 19012 13330
rect 18972 12640 19024 12646
rect 18970 12608 18972 12617
rect 19024 12608 19026 12617
rect 18970 12543 19026 12552
rect 19352 12481 19380 14039
rect 19338 12472 19394 12481
rect 19338 12407 19394 12416
rect 19248 11212 19300 11218
rect 19248 11154 19300 11160
rect 18972 11008 19024 11014
rect 18972 10950 19024 10956
rect 18984 10810 19012 10950
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19260 10266 19288 11154
rect 19340 10668 19392 10674
rect 19340 10610 19392 10616
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19352 9738 19380 10610
rect 19444 10130 19472 16351
rect 19536 15881 19564 16594
rect 19522 15872 19578 15881
rect 19522 15807 19578 15816
rect 19536 15473 19564 15807
rect 19522 15464 19578 15473
rect 19522 15399 19578 15408
rect 19536 14113 19564 15399
rect 19522 14104 19578 14113
rect 19522 14039 19578 14048
rect 19524 14000 19576 14006
rect 19522 13968 19524 13977
rect 19576 13968 19578 13977
rect 19522 13903 19578 13912
rect 19628 13546 19656 18090
rect 19996 18086 20024 18119
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 20180 17882 20208 18226
rect 20168 17876 20220 17882
rect 20168 17818 20220 17824
rect 20180 17338 20208 17818
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 19982 16552 20038 16561
rect 19982 16487 20038 16496
rect 19996 16250 20024 16487
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19996 16153 20024 16186
rect 19982 16144 20038 16153
rect 19982 16079 20038 16088
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19720 14657 19748 15302
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19706 14648 19762 14657
rect 19706 14583 19762 14592
rect 19904 14346 19932 14758
rect 19982 14512 20038 14521
rect 19982 14447 20038 14456
rect 19892 14340 19944 14346
rect 19892 14282 19944 14288
rect 19996 13870 20024 14447
rect 20088 14278 20116 14758
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19892 13728 19944 13734
rect 19892 13670 19944 13676
rect 19536 13518 19656 13546
rect 19536 12594 19564 13518
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 19720 12646 19748 13262
rect 19812 12986 19840 13262
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 19904 12753 19932 13670
rect 20088 12986 20116 13806
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19984 12844 20036 12850
rect 20088 12832 20116 12922
rect 20364 12918 20392 19178
rect 20732 19174 20760 19790
rect 20916 19242 20944 19858
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21652 18358 21680 18702
rect 21272 18352 21324 18358
rect 21272 18294 21324 18300
rect 21640 18352 21692 18358
rect 21640 18294 21692 18300
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21100 17338 21128 17614
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20812 16992 20864 16998
rect 20810 16960 20812 16969
rect 20864 16960 20866 16969
rect 20810 16895 20866 16904
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 21284 16776 21312 18294
rect 21640 18148 21692 18154
rect 21744 18136 21772 20810
rect 22192 20800 22244 20806
rect 22192 20742 22244 20748
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21928 19156 21956 19858
rect 22100 19168 22152 19174
rect 21928 19128 22100 19156
rect 21744 18108 21864 18136
rect 21640 18090 21692 18096
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21456 17808 21508 17814
rect 21456 17750 21508 17756
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 21192 16748 21312 16776
rect 21192 16658 21220 16748
rect 21180 16652 21232 16658
rect 21180 16594 21232 16600
rect 21272 16652 21324 16658
rect 21272 16594 21324 16600
rect 21192 16250 21220 16594
rect 21180 16244 21232 16250
rect 21180 16186 21232 16192
rect 21284 16182 21312 16594
rect 21376 16250 21404 17682
rect 21468 16794 21496 17750
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21364 16244 21416 16250
rect 21364 16186 21416 16192
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 21468 15706 21496 16730
rect 21560 16046 21588 18022
rect 21652 17864 21680 18090
rect 21652 17836 21772 17864
rect 21744 17660 21772 17836
rect 21652 17632 21772 17660
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20628 15156 20680 15162
rect 20732 15144 20760 15574
rect 21548 15564 21600 15570
rect 21548 15506 21600 15512
rect 20680 15116 20760 15144
rect 21272 15156 21324 15162
rect 20628 15098 20680 15104
rect 21272 15098 21324 15104
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 13394 20484 14758
rect 20640 14346 20668 14962
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20904 14476 20956 14482
rect 20904 14418 20956 14424
rect 20916 14385 20944 14418
rect 20902 14376 20958 14385
rect 20628 14340 20680 14346
rect 20902 14311 20958 14320
rect 20628 14282 20680 14288
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20444 13388 20496 13394
rect 20444 13330 20496 13336
rect 20352 12912 20404 12918
rect 20352 12854 20404 12860
rect 20036 12804 20116 12832
rect 19984 12786 20036 12792
rect 19890 12744 19946 12753
rect 19890 12679 19946 12688
rect 19708 12640 19760 12646
rect 19536 12566 19656 12594
rect 19708 12582 19760 12588
rect 19522 12472 19578 12481
rect 19522 12407 19578 12416
rect 19536 10266 19564 12407
rect 19628 11937 19656 12566
rect 19720 12209 19748 12582
rect 19996 12442 20024 12786
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20352 12640 20404 12646
rect 20352 12582 20404 12588
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20168 12300 20220 12306
rect 20168 12242 20220 12248
rect 19706 12200 19762 12209
rect 19706 12135 19762 12144
rect 19890 12200 19946 12209
rect 19890 12135 19946 12144
rect 19614 11928 19670 11937
rect 19614 11863 19670 11872
rect 19904 11286 19932 12135
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 19996 11121 20024 11630
rect 20180 11558 20208 12242
rect 20272 12102 20300 12582
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 19982 11112 20038 11121
rect 19982 11047 20038 11056
rect 19706 10976 19762 10985
rect 19706 10911 19762 10920
rect 19720 10305 19748 10911
rect 19706 10296 19762 10305
rect 19524 10260 19576 10266
rect 19706 10231 19762 10240
rect 19524 10202 19576 10208
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19536 9738 19564 10202
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19168 9710 19380 9738
rect 19444 9722 19564 9738
rect 19432 9716 19564 9722
rect 18694 9616 18750 9625
rect 17132 9580 17184 9586
rect 18694 9551 18750 9560
rect 17132 9522 17184 9528
rect 16854 9480 16910 9489
rect 16854 9415 16910 9424
rect 16856 9376 16908 9382
rect 16776 9324 16856 9330
rect 16776 9318 16908 9324
rect 16776 9302 16896 9318
rect 16580 9104 16632 9110
rect 16580 9046 16632 9052
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16396 8424 16448 8430
rect 16592 8378 16620 9046
rect 16868 8945 16896 9302
rect 17144 9110 17172 9522
rect 19168 9518 19196 9710
rect 19484 9710 19564 9716
rect 19432 9658 19484 9664
rect 19156 9512 19208 9518
rect 19156 9454 19208 9460
rect 18880 9376 18932 9382
rect 18880 9318 18932 9324
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 16948 8832 17000 8838
rect 16868 8780 16948 8786
rect 16868 8774 17000 8780
rect 16868 8758 16988 8774
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16396 8366 16448 8372
rect 16500 8350 16620 8378
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 14370 7576 14426 7585
rect 15956 7568 16252 7588
rect 14370 7511 14426 7520
rect 16316 7342 16344 8230
rect 16500 8090 16528 8350
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16684 7954 16712 8570
rect 16868 8498 16896 8758
rect 18616 8634 18644 8842
rect 18604 8628 18656 8634
rect 18604 8570 18656 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 8022 16896 8434
rect 18892 8401 18920 9318
rect 19168 9217 19196 9454
rect 19154 9208 19210 9217
rect 19154 9143 19156 9152
rect 19208 9143 19210 9152
rect 19156 9114 19208 9120
rect 19168 9083 19196 9114
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8498 19196 8774
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19628 8401 19656 10066
rect 19720 9178 19748 10231
rect 20180 10062 20208 11494
rect 20272 11354 20300 12038
rect 20364 11830 20392 12582
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20364 11626 20392 11766
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20260 11348 20312 11354
rect 20260 11290 20312 11296
rect 20364 10810 20392 11562
rect 20456 11150 20484 12038
rect 20548 11898 20576 14214
rect 20640 14006 20668 14282
rect 20916 14006 20944 14311
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20904 14000 20956 14006
rect 20904 13942 20956 13948
rect 21192 13870 21220 14214
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21284 13734 21312 15098
rect 21560 14618 21588 15506
rect 21548 14612 21600 14618
rect 21548 14554 21600 14560
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21362 13696 21418 13705
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 20628 13320 20680 13326
rect 20996 13320 21048 13326
rect 20680 13280 20760 13308
rect 20628 13262 20680 13268
rect 20628 12912 20680 12918
rect 20626 12880 20628 12889
rect 20680 12880 20682 12889
rect 20626 12815 20682 12824
rect 20628 12708 20680 12714
rect 20732 12696 20760 13280
rect 20996 13262 21048 13268
rect 21008 12918 21036 13262
rect 21088 13184 21140 13190
rect 21284 13172 21312 13670
rect 21362 13631 21418 13640
rect 21140 13144 21312 13172
rect 21088 13126 21140 13132
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 21100 12782 21128 13126
rect 21376 13025 21404 13631
rect 21362 13016 21418 13025
rect 21362 12951 21418 12960
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 20680 12668 20760 12696
rect 20628 12650 20680 12656
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 20444 11144 20496 11150
rect 20444 11086 20496 11092
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20350 10704 20406 10713
rect 20350 10639 20406 10648
rect 20364 10538 20392 10639
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 20364 10266 20392 10474
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 19708 9172 19760 9178
rect 19708 9114 19760 9120
rect 19720 8634 19748 9114
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19708 8492 19760 8498
rect 19708 8434 19760 8440
rect 18878 8392 18934 8401
rect 18878 8327 18934 8336
rect 19614 8392 19670 8401
rect 19614 8327 19670 8336
rect 18696 8288 18748 8294
rect 18696 8230 18748 8236
rect 16856 8016 16908 8022
rect 16856 7958 16908 7964
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 16684 7206 16712 7890
rect 16868 7274 16896 7958
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 17052 7546 17080 7686
rect 17040 7540 17092 7546
rect 17040 7482 17092 7488
rect 17052 7410 17080 7482
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 16856 7268 16908 7274
rect 16856 7210 16908 7216
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16408 6866 16436 7142
rect 16868 7002 16896 7210
rect 18524 7002 18552 7278
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15396 6458 15424 6802
rect 18616 6746 18644 7686
rect 18708 7206 18736 8230
rect 19064 7948 19116 7954
rect 19064 7890 19116 7896
rect 19076 7857 19104 7890
rect 19720 7886 19748 8434
rect 20180 8090 20208 8910
rect 20456 8498 20484 9318
rect 20548 9110 20576 11630
rect 20640 11064 20668 12174
rect 20732 11354 20760 12668
rect 21272 12708 21324 12714
rect 21272 12650 21324 12656
rect 20810 12608 20866 12617
rect 20810 12543 20866 12552
rect 20824 11626 20852 12543
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20904 12232 20956 12238
rect 20904 12174 20956 12180
rect 20916 11830 20944 12174
rect 21284 12102 21312 12650
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 20904 11824 20956 11830
rect 20904 11766 20956 11772
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 20720 11348 20772 11354
rect 20720 11290 20772 11296
rect 20812 11212 20864 11218
rect 20812 11154 20864 11160
rect 20640 11036 20760 11064
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 9450 20668 10406
rect 20732 10146 20760 11036
rect 20824 10266 20852 11154
rect 21284 10985 21312 11494
rect 21270 10976 21326 10985
rect 21270 10911 21326 10920
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 21376 10266 21404 12951
rect 21652 11778 21680 17632
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21744 14550 21772 15438
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21732 14408 21784 14414
rect 21732 14350 21784 14356
rect 21744 13530 21772 14350
rect 21836 13705 21864 18108
rect 21928 17882 21956 19128
rect 22100 19110 22152 19116
rect 22204 18290 22232 20742
rect 23400 20058 23428 23520
rect 24858 21584 24914 21593
rect 24858 21519 24914 21528
rect 24872 20806 24900 21519
rect 25056 21434 25084 23559
rect 25226 23520 25282 24000
rect 27158 23520 27214 24000
rect 28998 23520 29054 24000
rect 24964 21406 25084 21434
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 23938 20360 23994 20369
rect 23938 20295 23994 20304
rect 23388 20052 23440 20058
rect 23388 19994 23440 20000
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22192 18284 22244 18290
rect 22192 18226 22244 18232
rect 22296 18222 22324 19246
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22572 18358 22600 19110
rect 23112 18828 23164 18834
rect 23112 18770 23164 18776
rect 23124 18426 23152 18770
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 22560 18352 22612 18358
rect 22560 18294 22612 18300
rect 22834 18320 22890 18329
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22284 18216 22336 18222
rect 22284 18158 22336 18164
rect 22388 17882 22416 18226
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22296 16998 22324 17478
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22020 16833 22048 16934
rect 22006 16824 22062 16833
rect 22006 16759 22062 16768
rect 22296 16153 22324 16934
rect 22388 16658 22416 17818
rect 22572 17746 22600 18294
rect 22834 18255 22890 18264
rect 22560 17740 22612 17746
rect 22560 17682 22612 17688
rect 22572 17338 22600 17682
rect 22560 17332 22612 17338
rect 22560 17274 22612 17280
rect 22468 17060 22520 17066
rect 22468 17002 22520 17008
rect 22480 16697 22508 17002
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22466 16688 22522 16697
rect 22376 16652 22428 16658
rect 22466 16623 22522 16632
rect 22376 16594 22428 16600
rect 22282 16144 22338 16153
rect 22008 16108 22060 16114
rect 22282 16079 22338 16088
rect 22008 16050 22060 16056
rect 22020 15502 22048 16050
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22204 15706 22232 15846
rect 22192 15700 22244 15706
rect 22192 15642 22244 15648
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22388 15434 22416 16594
rect 22572 16114 22600 16730
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22558 15600 22614 15609
rect 22558 15535 22614 15544
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22388 15162 22416 15370
rect 22376 15156 22428 15162
rect 22376 15098 22428 15104
rect 22388 14414 22416 15098
rect 22376 14408 22428 14414
rect 22006 14376 22062 14385
rect 22376 14350 22428 14356
rect 22006 14311 22062 14320
rect 21822 13696 21878 13705
rect 21822 13631 21878 13640
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21822 13424 21878 13433
rect 21822 13359 21824 13368
rect 21876 13359 21878 13368
rect 21824 13330 21876 13336
rect 21822 12336 21878 12345
rect 21822 12271 21878 12280
rect 21560 11750 21680 11778
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21468 10810 21496 11086
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 20732 10130 20852 10146
rect 20732 10124 20864 10130
rect 20732 10118 20812 10124
rect 20812 10066 20864 10072
rect 21272 10124 21324 10130
rect 21272 10066 21324 10072
rect 20718 10024 20774 10033
rect 20718 9959 20774 9968
rect 20732 9926 20760 9959
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 21284 9586 21312 10066
rect 21376 9722 21404 10202
rect 21364 9716 21416 9722
rect 21364 9658 21416 9664
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 20628 9444 20680 9450
rect 20628 9386 20680 9392
rect 20536 9104 20588 9110
rect 20536 9046 20588 9052
rect 20548 8634 20576 9046
rect 20640 8974 20668 9386
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20628 8968 20680 8974
rect 21560 8945 21588 11750
rect 21836 11694 21864 12271
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21652 10130 21680 11562
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 21744 10674 21772 10950
rect 21822 10840 21878 10849
rect 21822 10775 21878 10784
rect 21732 10668 21784 10674
rect 21732 10610 21784 10616
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 20628 8910 20680 8916
rect 21546 8936 21602 8945
rect 21546 8871 21602 8880
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20444 8492 20496 8498
rect 20444 8434 20496 8440
rect 20720 8356 20772 8362
rect 20720 8298 20772 8304
rect 20732 8090 20760 8298
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 21652 8090 21680 10066
rect 21744 10062 21772 10610
rect 21836 10606 21864 10775
rect 21824 10600 21876 10606
rect 21824 10542 21876 10548
rect 21928 10470 21956 11154
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 10198 21956 10406
rect 21916 10192 21968 10198
rect 21916 10134 21968 10140
rect 21732 10056 21784 10062
rect 21732 9998 21784 10004
rect 21744 9722 21772 9998
rect 21732 9716 21784 9722
rect 21732 9658 21784 9664
rect 22020 9217 22048 14311
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22112 13326 22140 13942
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22112 11762 22140 13262
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 22006 9208 22062 9217
rect 22006 9143 22062 9152
rect 20168 8084 20220 8090
rect 20168 8026 20220 8032
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 21272 8084 21324 8090
rect 21272 8026 21324 8032
rect 21640 8084 21692 8090
rect 21640 8026 21692 8032
rect 19616 7880 19668 7886
rect 19062 7848 19118 7857
rect 19616 7822 19668 7828
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19062 7783 19118 7792
rect 19248 7812 19300 7818
rect 19076 7546 19104 7783
rect 19248 7754 19300 7760
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19168 7342 19196 7686
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 18696 7200 18748 7206
rect 18696 7142 18748 7148
rect 18708 6934 18736 7142
rect 19260 7002 19288 7754
rect 19628 7206 19656 7822
rect 20180 7818 20208 8026
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 19982 7440 20038 7449
rect 20180 7410 20208 7754
rect 21284 7478 21312 8026
rect 21364 7880 21416 7886
rect 21362 7848 21364 7857
rect 22112 7857 22140 11222
rect 22572 11218 22600 15535
rect 22848 11898 22876 18255
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23032 16674 23060 17138
rect 23124 16794 23152 18362
rect 23400 17746 23428 18566
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23400 17338 23428 17682
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23112 16788 23164 16794
rect 23112 16730 23164 16736
rect 23032 16658 23152 16674
rect 23032 16652 23164 16658
rect 23032 16646 23112 16652
rect 23112 16594 23164 16600
rect 23124 16250 23152 16594
rect 23216 16590 23244 17274
rect 23860 16658 23888 17478
rect 23952 17338 23980 20295
rect 24768 20256 24820 20262
rect 24768 20198 24820 20204
rect 24676 19236 24728 19242
rect 24676 19178 24728 19184
rect 24584 18692 24636 18698
rect 24584 18634 24636 18640
rect 24214 18184 24270 18193
rect 24214 18119 24270 18128
rect 23940 17332 23992 17338
rect 23940 17274 23992 17280
rect 23952 17134 23980 17274
rect 23940 17128 23992 17134
rect 23940 17070 23992 17076
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23204 16584 23256 16590
rect 23204 16526 23256 16532
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 23216 16250 23244 16526
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23204 16244 23256 16250
rect 23204 16186 23256 16192
rect 23572 16040 23624 16046
rect 23202 16008 23258 16017
rect 23572 15982 23624 15988
rect 23202 15943 23258 15952
rect 23216 15706 23244 15943
rect 23204 15700 23256 15706
rect 23204 15642 23256 15648
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 23124 14822 23152 15506
rect 23492 15162 23520 15642
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 22928 14408 22980 14414
rect 22928 14350 22980 14356
rect 22836 11892 22888 11898
rect 22836 11834 22888 11840
rect 22940 11529 22968 14350
rect 23020 13388 23072 13394
rect 23020 13330 23072 13336
rect 23032 13161 23060 13330
rect 23018 13152 23074 13161
rect 23018 13087 23074 13096
rect 23032 12986 23060 13087
rect 23020 12980 23072 12986
rect 23020 12922 23072 12928
rect 22926 11520 22982 11529
rect 22926 11455 22982 11464
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22572 10810 22600 11154
rect 22742 11112 22798 11121
rect 22742 11047 22744 11056
rect 22796 11047 22798 11056
rect 22744 11018 22796 11024
rect 22560 10804 22612 10810
rect 22560 10746 22612 10752
rect 22376 10600 22428 10606
rect 22376 10542 22428 10548
rect 22388 9926 22416 10542
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 23124 9489 23152 14758
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23492 13870 23520 14214
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23308 12850 23336 13126
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23492 12306 23520 13126
rect 23480 12300 23532 12306
rect 23480 12242 23532 12248
rect 23296 12164 23348 12170
rect 23296 12106 23348 12112
rect 23308 11830 23336 12106
rect 23478 11928 23534 11937
rect 23478 11863 23534 11872
rect 23492 11830 23520 11863
rect 23296 11824 23348 11830
rect 23296 11766 23348 11772
rect 23480 11824 23532 11830
rect 23480 11766 23532 11772
rect 23308 11014 23336 11766
rect 23480 11280 23532 11286
rect 23400 11228 23480 11234
rect 23400 11222 23532 11228
rect 23400 11206 23520 11222
rect 23296 11008 23348 11014
rect 23296 10950 23348 10956
rect 23400 10198 23428 11206
rect 23480 11144 23532 11150
rect 23480 11086 23532 11092
rect 23492 10266 23520 11086
rect 23584 10606 23612 15982
rect 23768 15706 23796 16526
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23768 15026 23796 15642
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14482 23796 14962
rect 23756 14476 23808 14482
rect 23756 14418 23808 14424
rect 23768 14074 23796 14418
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23768 13802 23796 14010
rect 23860 13938 23888 14214
rect 23952 13954 23980 17070
rect 24030 14376 24086 14385
rect 24030 14311 24086 14320
rect 24044 14074 24072 14311
rect 24032 14068 24084 14074
rect 24032 14010 24084 14016
rect 23848 13932 23900 13938
rect 23952 13926 24072 13954
rect 23848 13874 23900 13880
rect 23756 13796 23808 13802
rect 23756 13738 23808 13744
rect 23938 13696 23994 13705
rect 23938 13631 23994 13640
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23664 12776 23716 12782
rect 23664 12718 23716 12724
rect 23676 11354 23704 12718
rect 23664 11348 23716 11354
rect 23664 11290 23716 11296
rect 23768 11286 23796 13126
rect 23952 12986 23980 13631
rect 23940 12980 23992 12986
rect 23940 12922 23992 12928
rect 23848 11552 23900 11558
rect 23848 11494 23900 11500
rect 23756 11280 23808 11286
rect 23756 11222 23808 11228
rect 23860 11150 23888 11494
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23676 10606 23704 10950
rect 23572 10600 23624 10606
rect 23572 10542 23624 10548
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23388 10192 23440 10198
rect 23388 10134 23440 10140
rect 23940 9512 23992 9518
rect 23110 9480 23166 9489
rect 23110 9415 23166 9424
rect 23938 9480 23940 9489
rect 23992 9480 23994 9489
rect 23938 9415 23994 9424
rect 24044 7993 24072 13926
rect 24228 13530 24256 18119
rect 24596 18086 24624 18634
rect 24688 18630 24716 19178
rect 24780 18970 24808 20198
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24676 18624 24728 18630
rect 24676 18566 24728 18572
rect 24688 18290 24716 18566
rect 24676 18284 24728 18290
rect 24676 18226 24728 18232
rect 24964 18193 24992 21406
rect 25042 21312 25098 21321
rect 25042 21247 25098 21256
rect 25056 20874 25084 21247
rect 25044 20868 25096 20874
rect 25044 20810 25096 20816
rect 25240 20602 25268 23520
rect 25778 23080 25834 23089
rect 25778 23015 25834 23024
rect 25228 20596 25280 20602
rect 25228 20538 25280 20544
rect 25412 20528 25464 20534
rect 25410 20496 25412 20505
rect 25464 20496 25466 20505
rect 25792 20482 25820 23015
rect 25870 22400 25926 22409
rect 25870 22335 25926 22344
rect 25410 20431 25466 20440
rect 25700 20454 25820 20482
rect 25042 19408 25098 19417
rect 25042 19343 25098 19352
rect 24950 18184 25006 18193
rect 24950 18119 25006 18128
rect 24492 18080 24544 18086
rect 24584 18080 24636 18086
rect 24492 18022 24544 18028
rect 24582 18048 24584 18057
rect 24636 18048 24638 18057
rect 24504 17338 24532 18022
rect 24582 17983 24638 17992
rect 24768 17604 24820 17610
rect 24768 17546 24820 17552
rect 24492 17332 24544 17338
rect 24492 17274 24544 17280
rect 24780 17202 24808 17546
rect 24860 17536 24912 17542
rect 24860 17478 24912 17484
rect 24872 17338 24900 17478
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24768 17196 24820 17202
rect 24768 17138 24820 17144
rect 24584 16992 24636 16998
rect 24584 16934 24636 16940
rect 24398 16416 24454 16425
rect 24398 16351 24454 16360
rect 24412 16250 24440 16351
rect 24596 16250 24624 16934
rect 24780 16794 24808 17138
rect 24768 16788 24820 16794
rect 24768 16730 24820 16736
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24950 16144 25006 16153
rect 24950 16079 25006 16088
rect 24964 16046 24992 16079
rect 24952 16040 25004 16046
rect 25056 16017 25084 19343
rect 25700 19281 25728 20454
rect 25884 20346 25912 22335
rect 25956 21788 26252 21808
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 26606 20632 26662 20641
rect 26606 20567 26608 20576
rect 26660 20567 26662 20576
rect 26608 20538 26660 20544
rect 27172 20505 27200 23520
rect 29012 20641 29040 23520
rect 28998 20632 29054 20641
rect 28998 20567 29054 20576
rect 27158 20496 27214 20505
rect 27158 20431 27214 20440
rect 25792 20318 25912 20346
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 25686 19272 25742 19281
rect 25686 19207 25742 19216
rect 25792 19145 25820 20318
rect 25872 20256 25924 20262
rect 25872 20198 25924 20204
rect 25778 19136 25834 19145
rect 25778 19071 25834 19080
rect 25228 18760 25280 18766
rect 25228 18702 25280 18708
rect 25412 18760 25464 18766
rect 25412 18702 25464 18708
rect 25240 18358 25268 18702
rect 25424 18426 25452 18702
rect 25780 18624 25832 18630
rect 25780 18566 25832 18572
rect 25412 18420 25464 18426
rect 25412 18362 25464 18368
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 25240 17882 25268 18294
rect 25424 17882 25452 18362
rect 25792 18222 25820 18566
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25228 17876 25280 17882
rect 25228 17818 25280 17824
rect 25412 17876 25464 17882
rect 25412 17818 25464 17824
rect 25424 17066 25452 17818
rect 25516 17270 25544 18022
rect 25504 17264 25556 17270
rect 25504 17206 25556 17212
rect 25884 17218 25912 20198
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 26516 19372 26568 19378
rect 26516 19314 26568 19320
rect 26528 19174 26556 19314
rect 25964 19168 26016 19174
rect 25964 19110 26016 19116
rect 26516 19168 26568 19174
rect 26516 19110 26568 19116
rect 25976 18766 26004 19110
rect 26332 18828 26384 18834
rect 26332 18770 26384 18776
rect 25964 18760 26016 18766
rect 25964 18702 26016 18708
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 26344 17882 26372 18770
rect 26528 18222 26556 19110
rect 26516 18216 26568 18222
rect 26516 18158 26568 18164
rect 26514 18048 26570 18057
rect 26514 17983 26570 17992
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25688 17196 25740 17202
rect 25884 17190 26004 17218
rect 25688 17138 25740 17144
rect 25412 17060 25464 17066
rect 25412 17002 25464 17008
rect 25412 16584 25464 16590
rect 25412 16526 25464 16532
rect 25424 16114 25452 16526
rect 25502 16280 25558 16289
rect 25700 16250 25728 17138
rect 25870 16824 25926 16833
rect 25870 16759 25872 16768
rect 25924 16759 25926 16768
rect 25872 16730 25924 16736
rect 25778 16688 25834 16697
rect 25778 16623 25834 16632
rect 25502 16215 25558 16224
rect 25688 16244 25740 16250
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 24952 15982 25004 15988
rect 25042 16008 25098 16017
rect 25042 15943 25098 15952
rect 25424 15910 25452 16050
rect 25412 15904 25464 15910
rect 24858 15872 24914 15881
rect 25412 15846 25464 15852
rect 24858 15807 24914 15816
rect 24768 15632 24820 15638
rect 24768 15574 24820 15580
rect 24584 15496 24636 15502
rect 24780 15473 24808 15574
rect 24584 15438 24636 15444
rect 24766 15464 24822 15473
rect 24492 15428 24544 15434
rect 24492 15370 24544 15376
rect 24504 14929 24532 15370
rect 24596 15337 24624 15438
rect 24766 15399 24822 15408
rect 24582 15328 24638 15337
rect 24582 15263 24638 15272
rect 24596 15162 24624 15263
rect 24584 15156 24636 15162
rect 24584 15098 24636 15104
rect 24490 14920 24546 14929
rect 24490 14855 24492 14864
rect 24544 14855 24546 14864
rect 24492 14826 24544 14832
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24596 13938 24624 14486
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24400 13864 24452 13870
rect 24400 13806 24452 13812
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24136 12986 24164 13330
rect 24124 12980 24176 12986
rect 24124 12922 24176 12928
rect 24136 10266 24164 12922
rect 24228 12918 24256 13466
rect 24216 12912 24268 12918
rect 24216 12854 24268 12860
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24320 11150 24348 12038
rect 24412 11393 24440 13806
rect 24582 12744 24638 12753
rect 24582 12679 24638 12688
rect 24492 12300 24544 12306
rect 24492 12242 24544 12248
rect 24504 11762 24532 12242
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24398 11384 24454 11393
rect 24398 11319 24454 11328
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24320 10606 24348 11086
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24320 10266 24348 10542
rect 24596 10266 24624 12679
rect 24780 10810 24808 13806
rect 24872 13161 24900 15807
rect 25424 15502 25452 15846
rect 25412 15496 25464 15502
rect 24950 15464 25006 15473
rect 25412 15438 25464 15444
rect 24950 15399 25006 15408
rect 24858 13152 24914 13161
rect 24858 13087 24914 13096
rect 24860 12912 24912 12918
rect 24860 12854 24912 12860
rect 24872 11898 24900 12854
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24858 11792 24914 11801
rect 24964 11778 24992 15399
rect 25226 14648 25282 14657
rect 25226 14583 25282 14592
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25136 13184 25188 13190
rect 25136 13126 25188 13132
rect 25056 12850 25084 13126
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25056 11914 25084 12786
rect 25148 12782 25176 13126
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25240 12050 25268 14583
rect 25424 14074 25452 15438
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25516 13394 25544 16215
rect 25688 16186 25740 16192
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25608 14550 25636 14758
rect 25596 14544 25648 14550
rect 25596 14486 25648 14492
rect 25688 14272 25740 14278
rect 25688 14214 25740 14220
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25320 13388 25372 13394
rect 25320 13330 25372 13336
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25332 12986 25360 13330
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25424 12186 25452 13126
rect 25608 12850 25636 13874
rect 25700 13870 25728 14214
rect 25688 13864 25740 13870
rect 25688 13806 25740 13812
rect 25700 13530 25728 13806
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 25686 13424 25742 13433
rect 25686 13359 25742 13368
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25424 12158 25544 12186
rect 25240 12022 25452 12050
rect 25056 11886 25268 11914
rect 24964 11750 25084 11778
rect 24858 11727 24914 11736
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 24308 10260 24360 10266
rect 24308 10202 24360 10208
rect 24584 10260 24636 10266
rect 24584 10202 24636 10208
rect 24872 10044 24900 11727
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24964 11354 24992 11562
rect 24952 11348 25004 11354
rect 24952 11290 25004 11296
rect 24952 10736 25004 10742
rect 24950 10704 24952 10713
rect 25004 10704 25006 10713
rect 24950 10639 25006 10648
rect 25056 10169 25084 11750
rect 25134 10840 25190 10849
rect 25134 10775 25190 10784
rect 25042 10160 25098 10169
rect 25042 10095 25098 10104
rect 24872 10016 25084 10044
rect 24952 9920 25004 9926
rect 24858 9888 24914 9897
rect 24952 9862 25004 9868
rect 24858 9823 24914 9832
rect 24674 9752 24730 9761
rect 24674 9687 24730 9696
rect 24688 9178 24716 9687
rect 24768 9648 24820 9654
rect 24872 9602 24900 9823
rect 24820 9596 24900 9602
rect 24768 9590 24900 9596
rect 24780 9574 24900 9590
rect 24964 9466 24992 9862
rect 24872 9438 24992 9466
rect 24872 9382 24900 9438
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24030 7984 24086 7993
rect 24030 7919 24086 7928
rect 21416 7848 21418 7857
rect 22098 7848 22154 7857
rect 21362 7783 21418 7792
rect 21640 7812 21692 7818
rect 21376 7546 21404 7783
rect 22098 7783 22154 7792
rect 21640 7754 21692 7760
rect 21652 7546 21680 7754
rect 24872 7721 24900 9318
rect 24858 7712 24914 7721
rect 24858 7647 24914 7656
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21640 7540 21692 7546
rect 21640 7482 21692 7488
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 19982 7375 20038 7384
rect 20168 7404 20220 7410
rect 19996 7342 20024 7375
rect 20168 7346 20220 7352
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19616 7200 19668 7206
rect 19720 7177 19748 7210
rect 19616 7142 19668 7148
rect 19706 7168 19762 7177
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19628 6934 19656 7142
rect 19706 7103 19762 7112
rect 19720 7002 19748 7103
rect 19996 7002 20024 7278
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 24872 7041 24900 7647
rect 24858 7032 24914 7041
rect 19708 6996 19760 7002
rect 19708 6938 19760 6944
rect 19984 6996 20036 7002
rect 24858 6967 24914 6976
rect 19984 6938 20036 6944
rect 18696 6928 18748 6934
rect 18696 6870 18748 6876
rect 19616 6928 19668 6934
rect 19616 6870 19668 6876
rect 18616 6718 18736 6746
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15384 6452 15436 6458
rect 15384 6394 15436 6400
rect 13358 5128 13414 5137
rect 13358 5063 13414 5072
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 15488 3505 15516 6598
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 15474 3496 15530 3505
rect 15474 3431 15530 3440
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 11150 2408 11206 2417
rect 11150 2343 11206 2352
rect 9034 912 9090 921
rect 9034 847 9090 856
rect 11164 480 11192 2343
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 18708 480 18736 6718
rect 19720 4049 19748 6938
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 19706 4040 19762 4049
rect 19706 3975 19762 3984
rect 25056 3913 25084 10016
rect 25148 8634 25176 10775
rect 25240 10742 25268 11886
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25228 10736 25280 10742
rect 25228 10678 25280 10684
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25240 9722 25268 10202
rect 25228 9716 25280 9722
rect 25228 9658 25280 9664
rect 25332 9518 25360 11630
rect 25320 9512 25372 9518
rect 25320 9454 25372 9460
rect 25318 9072 25374 9081
rect 25318 9007 25320 9016
rect 25372 9007 25374 9016
rect 25320 8978 25372 8984
rect 25332 8634 25360 8978
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25148 8430 25176 8570
rect 25136 8424 25188 8430
rect 25136 8366 25188 8372
rect 25318 7984 25374 7993
rect 25318 7919 25320 7928
rect 25372 7919 25374 7928
rect 25320 7890 25372 7896
rect 25332 7546 25360 7890
rect 25320 7540 25372 7546
rect 25320 7482 25372 7488
rect 25424 7449 25452 12022
rect 25516 11801 25544 12158
rect 25502 11792 25558 11801
rect 25502 11727 25558 11736
rect 25502 11656 25558 11665
rect 25502 11591 25558 11600
rect 25516 9654 25544 11591
rect 25596 11212 25648 11218
rect 25700 11200 25728 13359
rect 25792 12986 25820 16623
rect 25976 16538 26004 17190
rect 26424 16992 26476 16998
rect 26424 16934 26476 16940
rect 25976 16510 26372 16538
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25872 15632 25924 15638
rect 25872 15574 25924 15580
rect 25884 13841 25912 15574
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 26344 14618 26372 16510
rect 26436 15978 26464 16934
rect 26528 16658 26556 17983
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26620 16538 26648 20334
rect 26790 20088 26846 20097
rect 26790 20023 26846 20032
rect 26804 18873 26832 20023
rect 27436 19848 27488 19854
rect 27436 19790 27488 19796
rect 27448 19310 27476 19790
rect 27436 19304 27488 19310
rect 27342 19272 27398 19281
rect 27436 19246 27488 19252
rect 27342 19207 27398 19216
rect 26884 19168 26936 19174
rect 26882 19136 26884 19145
rect 27068 19168 27120 19174
rect 26936 19136 26938 19145
rect 27068 19110 27120 19116
rect 26882 19071 26938 19080
rect 27080 18902 27108 19110
rect 27068 18896 27120 18902
rect 26790 18864 26846 18873
rect 27068 18838 27120 18844
rect 26790 18799 26846 18808
rect 26976 18828 27028 18834
rect 26804 17678 26832 18799
rect 26976 18770 27028 18776
rect 26988 18154 27016 18770
rect 27068 18760 27120 18766
rect 27068 18702 27120 18708
rect 27080 18426 27108 18702
rect 27068 18420 27120 18426
rect 27068 18362 27120 18368
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 26976 18148 27028 18154
rect 26976 18090 27028 18096
rect 26988 17882 27016 18090
rect 26976 17876 27028 17882
rect 26976 17818 27028 17824
rect 26882 17776 26938 17785
rect 26882 17711 26884 17720
rect 26936 17711 26938 17720
rect 26884 17682 26936 17688
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26804 17338 26832 17614
rect 26792 17332 26844 17338
rect 26792 17274 26844 17280
rect 26896 17270 26924 17682
rect 27172 17678 27200 18158
rect 27160 17672 27212 17678
rect 27160 17614 27212 17620
rect 26884 17264 26936 17270
rect 26884 17206 26936 17212
rect 26884 16652 26936 16658
rect 26884 16594 26936 16600
rect 26528 16510 26648 16538
rect 26424 15972 26476 15978
rect 26424 15914 26476 15920
rect 26436 15434 26464 15914
rect 26424 15428 26476 15434
rect 26424 15370 26476 15376
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 25870 13832 25926 13841
rect 25870 13767 25926 13776
rect 25780 12980 25832 12986
rect 25780 12922 25832 12928
rect 25884 12209 25912 13767
rect 26528 13705 26556 16510
rect 26896 15706 26924 16594
rect 27172 16590 27200 17614
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27172 16454 27200 16526
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27172 16250 27200 16390
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27252 15904 27304 15910
rect 27252 15846 27304 15852
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26884 15564 26936 15570
rect 26884 15506 26936 15512
rect 26514 13696 26570 13705
rect 26514 13631 26570 13640
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26332 13184 26384 13190
rect 26332 13126 26384 13132
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 26344 12866 26372 13126
rect 26436 12986 26464 13262
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26424 12980 26476 12986
rect 26424 12922 26476 12928
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26252 12838 26372 12866
rect 26160 12442 26188 12786
rect 26252 12714 26280 12838
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26148 12436 26200 12442
rect 26148 12378 26200 12384
rect 26252 12322 26280 12650
rect 26160 12306 26280 12322
rect 26148 12300 26280 12306
rect 26200 12294 26280 12300
rect 26148 12242 26200 12248
rect 25870 12200 25926 12209
rect 25870 12135 25926 12144
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 25792 11830 25820 12038
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 25884 11762 25912 12038
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26436 11778 26464 12922
rect 26528 12442 26556 13126
rect 26516 12436 26568 12442
rect 26516 12378 26568 12384
rect 26620 12306 26648 15506
rect 26896 15094 26924 15506
rect 26976 15496 27028 15502
rect 26976 15438 27028 15444
rect 26884 15088 26936 15094
rect 26884 15030 26936 15036
rect 26792 14952 26844 14958
rect 26792 14894 26844 14900
rect 26804 14822 26832 14894
rect 26988 14890 27016 15438
rect 27160 15360 27212 15366
rect 27160 15302 27212 15308
rect 27172 14958 27200 15302
rect 27264 15026 27292 15846
rect 27252 15020 27304 15026
rect 27252 14962 27304 14968
rect 27160 14952 27212 14958
rect 27264 14929 27292 14962
rect 27160 14894 27212 14900
rect 27250 14920 27306 14929
rect 26976 14884 27028 14890
rect 27250 14855 27306 14864
rect 26976 14826 27028 14832
rect 26700 14816 26752 14822
rect 26700 14758 26752 14764
rect 26792 14816 26844 14822
rect 26792 14758 26844 14764
rect 26712 14521 26740 14758
rect 26698 14512 26754 14521
rect 26698 14447 26754 14456
rect 26700 14408 26752 14414
rect 26700 14350 26752 14356
rect 26712 13977 26740 14350
rect 26698 13968 26754 13977
rect 26698 13903 26700 13912
rect 26752 13903 26754 13912
rect 26700 13874 26752 13880
rect 26712 13843 26740 13874
rect 26804 13784 26832 14758
rect 26884 14476 26936 14482
rect 26884 14418 26936 14424
rect 26896 14385 26924 14418
rect 26882 14376 26938 14385
rect 26882 14311 26938 14320
rect 26896 14006 26924 14311
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26804 13756 26924 13784
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 25872 11756 25924 11762
rect 26436 11750 26556 11778
rect 26620 11762 26648 12242
rect 26790 11928 26846 11937
rect 26790 11863 26792 11872
rect 26844 11863 26846 11872
rect 26792 11834 26844 11840
rect 26896 11778 26924 13756
rect 25872 11698 25924 11704
rect 25884 11354 25912 11698
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26528 11506 26556 11750
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26804 11750 26924 11778
rect 25872 11348 25924 11354
rect 25872 11290 25924 11296
rect 25700 11172 25912 11200
rect 25596 11154 25648 11160
rect 25608 10606 25636 11154
rect 25688 11076 25740 11082
rect 25688 11018 25740 11024
rect 25596 10600 25648 10606
rect 25594 10568 25596 10577
rect 25648 10568 25650 10577
rect 25594 10503 25650 10512
rect 25596 10056 25648 10062
rect 25596 9998 25648 10004
rect 25608 9761 25636 9998
rect 25594 9752 25650 9761
rect 25594 9687 25650 9696
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25594 9344 25650 9353
rect 25594 9279 25650 9288
rect 25504 8832 25556 8838
rect 25504 8774 25556 8780
rect 25516 8537 25544 8774
rect 25608 8566 25636 9279
rect 25596 8560 25648 8566
rect 25502 8528 25558 8537
rect 25596 8502 25648 8508
rect 25502 8463 25558 8472
rect 25502 8120 25558 8129
rect 25502 8055 25504 8064
rect 25556 8055 25558 8064
rect 25504 8026 25556 8032
rect 25410 7440 25466 7449
rect 25410 7375 25466 7384
rect 25042 3904 25098 3913
rect 20956 3836 21252 3856
rect 25042 3839 25098 3848
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 25700 3505 25728 11018
rect 25780 10532 25832 10538
rect 25780 10474 25832 10480
rect 25686 3496 25742 3505
rect 25686 3431 25742 3440
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 25792 1306 25820 10474
rect 25884 10266 25912 11172
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 26436 9518 26464 11494
rect 26528 11478 26648 11506
rect 26514 11384 26570 11393
rect 26514 11319 26516 11328
rect 26568 11319 26570 11328
rect 26516 11290 26568 11296
rect 26514 10704 26570 10713
rect 26514 10639 26570 10648
rect 26528 10470 26556 10639
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26528 10033 26556 10406
rect 26620 10130 26648 11478
rect 26700 11008 26752 11014
rect 26700 10950 26752 10956
rect 26712 10674 26740 10950
rect 26700 10668 26752 10674
rect 26700 10610 26752 10616
rect 26608 10124 26660 10130
rect 26608 10066 26660 10072
rect 26514 10024 26570 10033
rect 26514 9959 26516 9968
rect 26568 9959 26570 9968
rect 26516 9930 26568 9936
rect 26620 9722 26648 10066
rect 26712 10062 26740 10610
rect 26700 10056 26752 10062
rect 26700 9998 26752 10004
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 26424 9512 26476 9518
rect 26424 9454 26476 9460
rect 26700 9376 26752 9382
rect 26700 9318 26752 9324
rect 26422 9208 26478 9217
rect 26422 9143 26478 9152
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 25884 4593 25912 8774
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 26436 8430 26464 9143
rect 26516 9036 26568 9042
rect 26516 8978 26568 8984
rect 26528 8634 26556 8978
rect 26516 8628 26568 8634
rect 26516 8570 26568 8576
rect 26424 8424 26476 8430
rect 26528 8401 26556 8570
rect 26608 8560 26660 8566
rect 26608 8502 26660 8508
rect 26424 8366 26476 8372
rect 26514 8392 26570 8401
rect 26514 8327 26570 8336
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 26620 7449 26648 8502
rect 26606 7440 26662 7449
rect 26606 7375 26662 7384
rect 26514 7032 26570 7041
rect 26514 6967 26570 6976
rect 26528 6866 26556 6967
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 26528 6458 26556 6802
rect 26712 6746 26740 9318
rect 26804 7954 26832 11750
rect 26882 11520 26938 11529
rect 26882 11455 26938 11464
rect 26896 11354 26924 11455
rect 26884 11348 26936 11354
rect 26884 11290 26936 11296
rect 26988 10010 27016 14826
rect 27264 14278 27292 14855
rect 27160 14272 27212 14278
rect 27160 14214 27212 14220
rect 27252 14272 27304 14278
rect 27252 14214 27304 14220
rect 27172 14074 27200 14214
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27068 13728 27120 13734
rect 27068 13670 27120 13676
rect 27080 13326 27108 13670
rect 27068 13320 27120 13326
rect 27068 13262 27120 13268
rect 27160 11892 27212 11898
rect 27160 11834 27212 11840
rect 27172 11626 27200 11834
rect 27160 11620 27212 11626
rect 27160 11562 27212 11568
rect 26988 9982 27108 10010
rect 26976 9920 27028 9926
rect 26976 9862 27028 9868
rect 26792 7948 26844 7954
rect 26792 7890 26844 7896
rect 26804 7857 26832 7890
rect 26790 7848 26846 7857
rect 26846 7806 26924 7834
rect 26790 7783 26846 7792
rect 26792 7744 26844 7750
rect 26792 7686 26844 7692
rect 26620 6718 26740 6746
rect 26516 6452 26568 6458
rect 26516 6394 26568 6400
rect 26620 5545 26648 6718
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26712 6361 26740 6598
rect 26698 6352 26754 6361
rect 26698 6287 26754 6296
rect 26606 5536 26662 5545
rect 25956 5468 26252 5488
rect 26606 5471 26662 5480
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 26424 5160 26476 5166
rect 26422 5128 26424 5137
rect 26476 5128 26478 5137
rect 26422 5063 26478 5072
rect 26606 5128 26662 5137
rect 26606 5063 26662 5072
rect 26620 5030 26648 5063
rect 26608 5024 26660 5030
rect 26608 4966 26660 4972
rect 25870 4584 25926 4593
rect 25870 4519 25926 4528
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 26422 4040 26478 4049
rect 26422 3975 26478 3984
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 26436 2990 26464 3975
rect 26424 2984 26476 2990
rect 26424 2926 26476 2932
rect 26608 2848 26660 2854
rect 26606 2816 26608 2825
rect 26660 2816 26662 2825
rect 26606 2751 26662 2760
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 26804 1465 26832 7686
rect 26896 7478 26924 7806
rect 26884 7472 26936 7478
rect 26884 7414 26936 7420
rect 26884 7200 26936 7206
rect 26884 7142 26936 7148
rect 26790 1456 26846 1465
rect 26790 1391 26846 1400
rect 25792 1278 26188 1306
rect 26160 480 26188 1278
rect 2686 368 2742 377
rect 2686 303 2742 312
rect 3698 0 3754 480
rect 11150 0 11206 480
rect 18694 0 18750 480
rect 26146 0 26202 480
rect 26896 377 26924 7142
rect 26988 6338 27016 9862
rect 27080 8294 27108 9982
rect 27068 8288 27120 8294
rect 27068 8230 27120 8236
rect 27080 7546 27108 8230
rect 27068 7540 27120 7546
rect 27068 7482 27120 7488
rect 27080 7342 27108 7482
rect 27172 7342 27200 11562
rect 27264 11150 27292 14214
rect 27356 11354 27384 19207
rect 29366 17232 29422 17241
rect 27988 17196 28040 17202
rect 29366 17167 29422 17176
rect 27988 17138 28040 17144
rect 27528 15496 27580 15502
rect 27580 15456 27660 15484
rect 27528 15438 27580 15444
rect 27632 15162 27660 15456
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27712 15088 27764 15094
rect 27712 15030 27764 15036
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 27540 12238 27568 12582
rect 27724 12345 27752 15030
rect 27710 12336 27766 12345
rect 27710 12271 27766 12280
rect 27528 12232 27580 12238
rect 27434 12200 27490 12209
rect 27528 12174 27580 12180
rect 27434 12135 27490 12144
rect 27448 11762 27476 12135
rect 27540 11762 27568 12174
rect 27436 11756 27488 11762
rect 27436 11698 27488 11704
rect 27528 11756 27580 11762
rect 27528 11698 27580 11704
rect 27540 11354 27568 11698
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27528 11348 27580 11354
rect 27528 11290 27580 11296
rect 27252 11144 27304 11150
rect 27252 11086 27304 11092
rect 27356 10810 27384 11290
rect 27620 11280 27672 11286
rect 27620 11222 27672 11228
rect 27632 10810 27660 11222
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27710 10432 27766 10441
rect 27710 10367 27766 10376
rect 27526 9616 27582 9625
rect 27526 9551 27582 9560
rect 27540 9518 27568 9551
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27724 8634 27752 10367
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27712 7200 27764 7206
rect 27712 7142 27764 7148
rect 27724 7041 27752 7142
rect 27710 7032 27766 7041
rect 27710 6967 27766 6976
rect 26988 6310 27108 6338
rect 26974 5536 27030 5545
rect 26974 5471 27030 5480
rect 26988 2145 27016 5471
rect 26974 2136 27030 2145
rect 26974 2071 27030 2080
rect 27080 921 27108 6310
rect 27816 5681 27844 9318
rect 28000 8634 28028 17138
rect 29380 17105 29408 17167
rect 29366 17096 29422 17105
rect 29366 17031 29422 17040
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 28184 12918 28212 13330
rect 28172 12912 28224 12918
rect 28170 12880 28172 12889
rect 28224 12880 28226 12889
rect 28170 12815 28226 12824
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 28000 8430 28028 8570
rect 27988 8424 28040 8430
rect 27988 8366 28040 8372
rect 27802 5672 27858 5681
rect 27802 5607 27858 5616
rect 27066 912 27122 921
rect 27066 847 27122 856
rect 26882 368 26938 377
rect 26882 303 26938 312
<< via2 >>
rect 3330 23568 3386 23624
rect 25042 23568 25098 23624
rect 3514 23024 3570 23080
rect 2870 22344 2926 22400
rect 1950 20204 1952 20224
rect 1952 20204 2004 20224
rect 2004 20204 2006 20224
rect 1950 20168 2006 20204
rect 2042 18828 2098 18864
rect 2042 18808 2044 18828
rect 2044 18808 2096 18828
rect 2096 18808 2098 18828
rect 2686 19352 2742 19408
rect 3330 21800 3386 21856
rect 2962 20576 3018 20632
rect 754 15816 810 15872
rect 1490 9832 1546 9888
rect 1398 9560 1454 9616
rect 1398 7948 1454 7984
rect 1398 7928 1400 7948
rect 1400 7928 1452 7948
rect 1452 7928 1454 7948
rect 1582 6840 1638 6896
rect 1582 6296 1638 6352
rect 1398 5616 1454 5672
rect 2042 15816 2098 15872
rect 2042 15544 2098 15600
rect 2410 14764 2412 14784
rect 2412 14764 2464 14784
rect 2464 14764 2466 14784
rect 2410 14728 2466 14764
rect 2042 13232 2098 13288
rect 2134 11736 2190 11792
rect 2134 10376 2190 10432
rect 2042 7928 2098 7984
rect 2502 10512 2558 10568
rect 2410 6840 2466 6896
rect 2962 18536 3018 18592
rect 3146 18264 3202 18320
rect 3146 15680 3202 15736
rect 2870 14728 2926 14784
rect 2594 9424 2650 9480
rect 4066 21256 4122 21312
rect 3422 20168 3478 20224
rect 3698 19216 3754 19272
rect 3882 19116 3884 19136
rect 3884 19116 3936 19136
rect 3936 19116 3938 19136
rect 3882 19080 3938 19116
rect 3698 18264 3754 18320
rect 4434 20052 4490 20088
rect 4434 20032 4436 20052
rect 4436 20032 4488 20052
rect 4488 20032 4490 20052
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 4618 19352 4674 19408
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 6550 20032 6606 20088
rect 4986 18944 5042 19000
rect 3790 15272 3846 15328
rect 3514 13368 3570 13424
rect 3422 11328 3478 11384
rect 2962 9424 3018 9480
rect 3146 9424 3202 9480
rect 3330 9424 3386 9480
rect 2686 8608 2742 8664
rect 3422 8064 3478 8120
rect 2686 7420 2688 7440
rect 2688 7420 2740 7440
rect 2740 7420 2742 7440
rect 2686 7384 2742 7420
rect 3146 7404 3202 7440
rect 3146 7384 3148 7404
rect 3148 7384 3200 7404
rect 3200 7384 3202 7404
rect 3146 6704 3202 6760
rect 1674 4392 1730 4448
rect 2042 3984 2098 4040
rect 1582 2624 1638 2680
rect 1398 1400 1454 1456
rect 3606 9424 3662 9480
rect 4526 15816 4582 15872
rect 4618 15544 4674 15600
rect 4066 15000 4122 15056
rect 3974 13504 4030 13560
rect 4250 13640 4306 13696
rect 3882 12044 3884 12064
rect 3884 12044 3936 12064
rect 3936 12044 3938 12064
rect 3882 12008 3938 12044
rect 3974 11600 4030 11656
rect 4158 11328 4214 11384
rect 3698 9288 3754 9344
rect 3514 5072 3570 5128
rect 3698 3440 3754 3496
rect 4434 13504 4490 13560
rect 4434 12552 4490 12608
rect 4710 13368 4766 13424
rect 4986 17720 5042 17776
rect 4986 14048 5042 14104
rect 4986 12688 5042 12744
rect 4618 12280 4674 12336
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 5354 19216 5410 19272
rect 6182 19216 6238 19272
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5722 18128 5778 18184
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 5722 16360 5778 16416
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 5630 14900 5632 14920
rect 5632 14900 5684 14920
rect 5684 14900 5686 14920
rect 5630 14864 5686 14900
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5354 14048 5410 14104
rect 5170 12724 5172 12744
rect 5172 12724 5224 12744
rect 5224 12724 5226 12744
rect 5630 13524 5686 13560
rect 5630 13504 5632 13524
rect 5632 13504 5684 13524
rect 5684 13504 5686 13524
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 6274 13504 6330 13560
rect 7286 19080 7342 19136
rect 6826 18264 6882 18320
rect 6458 17448 6514 17504
rect 6458 17040 6514 17096
rect 7286 16360 7342 16416
rect 6642 15000 6698 15056
rect 6550 14592 6606 14648
rect 5170 12688 5226 12724
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5722 12008 5778 12064
rect 5630 11500 5632 11520
rect 5632 11500 5684 11520
rect 5684 11500 5686 11520
rect 5630 11464 5686 11500
rect 5538 11328 5594 11384
rect 5170 10648 5226 10704
rect 5630 10240 5686 10296
rect 5538 10104 5594 10160
rect 5630 9968 5686 10024
rect 5078 9696 5134 9752
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5814 9696 5870 9752
rect 5630 9560 5686 9616
rect 4986 9424 5042 9480
rect 5262 8356 5318 8392
rect 5262 8336 5264 8356
rect 5264 8336 5316 8356
rect 5316 8336 5318 8356
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 6458 13096 6514 13152
rect 7286 14864 7342 14920
rect 6734 11328 6790 11384
rect 6918 12688 6974 12744
rect 7102 11056 7158 11112
rect 7010 10784 7066 10840
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 6274 6704 6330 6760
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 4342 3848 4398 3904
rect 3790 3304 3846 3360
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 7010 9560 7066 9616
rect 7378 12960 7434 13016
rect 7746 18964 7802 19000
rect 7746 18944 7748 18964
rect 7748 18944 7800 18964
rect 7800 18944 7802 18964
rect 7930 18128 7986 18184
rect 7562 15816 7618 15872
rect 7930 15680 7986 15736
rect 9678 18164 9680 18184
rect 9680 18164 9732 18184
rect 9732 18164 9734 18184
rect 8942 17176 8998 17232
rect 8114 15544 8170 15600
rect 8390 15700 8446 15736
rect 8390 15680 8392 15700
rect 8392 15680 8444 15700
rect 8444 15680 8446 15700
rect 8298 14728 8354 14784
rect 8298 13776 8354 13832
rect 7746 10648 7802 10704
rect 8574 12144 8630 12200
rect 9678 18128 9734 18164
rect 9310 16224 9366 16280
rect 8942 13640 8998 13696
rect 8482 11464 8538 11520
rect 8390 11192 8446 11248
rect 8850 11348 8906 11384
rect 8850 11328 8852 11348
rect 8852 11328 8904 11348
rect 8904 11328 8906 11348
rect 7378 8336 7434 8392
rect 7562 7828 7564 7848
rect 7564 7828 7616 7848
rect 7616 7828 7618 7848
rect 7010 7384 7066 7440
rect 7562 7792 7618 7828
rect 6918 6840 6974 6896
rect 7378 7284 7380 7304
rect 7380 7284 7432 7304
rect 7432 7284 7434 7304
rect 7378 7248 7434 7284
rect 6918 3984 6974 4040
rect 8390 2488 8446 2544
rect 7194 2352 7250 2408
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 9862 19352 9918 19408
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 10782 19896 10838 19952
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 12070 19352 12126 19408
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 11334 18672 11390 18728
rect 10782 18264 10838 18320
rect 9862 17584 9918 17640
rect 9862 16632 9918 16688
rect 11150 18164 11152 18184
rect 11152 18164 11204 18184
rect 11204 18164 11206 18184
rect 11150 18128 11206 18164
rect 12806 19896 12862 19952
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 10506 16632 10562 16688
rect 10414 15020 10470 15056
rect 10414 15000 10416 15020
rect 10416 15000 10468 15020
rect 10468 15000 10470 15020
rect 10322 14864 10378 14920
rect 10046 11736 10102 11792
rect 10782 16360 10838 16416
rect 11150 16360 11206 16416
rect 11518 16088 11574 16144
rect 10598 15852 10600 15872
rect 10600 15852 10652 15872
rect 10652 15852 10654 15872
rect 10598 15816 10654 15852
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10874 14476 10930 14512
rect 10874 14456 10876 14476
rect 10876 14456 10928 14476
rect 10928 14456 10930 14476
rect 10782 13504 10838 13560
rect 11334 14220 11336 14240
rect 11336 14220 11388 14240
rect 11388 14220 11390 14240
rect 11334 14184 11390 14220
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 10598 11600 10654 11656
rect 10138 10804 10194 10840
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10690 11192 10746 11248
rect 10138 10784 10140 10804
rect 10140 10784 10192 10804
rect 10192 10784 10194 10804
rect 10322 10512 10378 10568
rect 10322 10260 10378 10296
rect 10322 10240 10324 10260
rect 10324 10240 10376 10260
rect 10376 10240 10378 10260
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10782 10124 10838 10160
rect 10782 10104 10784 10124
rect 10784 10104 10836 10124
rect 10836 10104 10838 10124
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 9126 8744 9182 8800
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 11978 17720 12034 17776
rect 11610 11192 11666 11248
rect 12990 18028 12992 18048
rect 12992 18028 13044 18048
rect 13044 18028 13046 18048
rect 12990 17992 13046 18028
rect 12346 16224 12402 16280
rect 12530 15816 12586 15872
rect 12254 13524 12310 13560
rect 12254 13504 12256 13524
rect 12256 13504 12308 13524
rect 12308 13504 12310 13524
rect 12162 13096 12218 13152
rect 12162 12708 12218 12744
rect 12162 12688 12164 12708
rect 12164 12688 12216 12708
rect 12216 12688 12218 12708
rect 13542 17176 13598 17232
rect 12898 15816 12954 15872
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 14094 18708 14096 18728
rect 14096 18708 14148 18728
rect 14148 18708 14150 18728
rect 14094 18672 14150 18708
rect 13634 15136 13690 15192
rect 13542 13776 13598 13832
rect 13818 14184 13874 14240
rect 13358 13096 13414 13152
rect 12070 11600 12126 11656
rect 12990 12300 13046 12336
rect 12990 12280 12992 12300
rect 12992 12280 13044 12300
rect 13044 12280 13046 12300
rect 12990 12144 13046 12200
rect 13266 11500 13268 11520
rect 13268 11500 13320 11520
rect 13320 11500 13322 11520
rect 13266 11464 13322 11500
rect 11978 10648 12034 10704
rect 11518 7928 11574 7984
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 14094 13388 14150 13424
rect 14094 13368 14096 13388
rect 14096 13368 14148 13388
rect 14148 13368 14150 13388
rect 13634 12824 13690 12880
rect 13818 9016 13874 9072
rect 15750 19216 15806 19272
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15750 16088 15806 16144
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 15566 15952 15622 16008
rect 15382 15544 15438 15600
rect 14738 14864 14794 14920
rect 14462 14592 14518 14648
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 16026 15036 16028 15056
rect 16028 15036 16080 15056
rect 16080 15036 16082 15056
rect 16026 15000 16082 15036
rect 15014 14320 15070 14376
rect 15658 14456 15714 14512
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 14922 12552 14978 12608
rect 15106 12552 15162 12608
rect 14922 12144 14978 12200
rect 16302 13232 16358 13288
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15290 12144 15346 12200
rect 15382 11464 15438 11520
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 15842 11636 15844 11656
rect 15844 11636 15896 11656
rect 15896 11636 15898 11656
rect 15842 11600 15898 11636
rect 16210 11192 16266 11248
rect 17038 16496 17094 16552
rect 16394 11328 16450 11384
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 16486 11192 16542 11248
rect 16762 11056 16818 11112
rect 18326 17584 18382 17640
rect 17406 14592 17462 14648
rect 19982 20324 20038 20360
rect 19982 20304 19984 20324
rect 19984 20304 20036 20324
rect 20036 20304 20038 20324
rect 19430 18828 19486 18864
rect 19430 18808 19432 18828
rect 19432 18808 19484 18828
rect 19484 18808 19486 18828
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 19982 18692 20038 18728
rect 19982 18672 19984 18692
rect 19984 18672 20036 18692
rect 20036 18672 20038 18692
rect 19062 18148 19118 18184
rect 19062 18128 19064 18148
rect 19064 18128 19116 18148
rect 19116 18128 19118 18148
rect 19982 18128 20038 18184
rect 18970 16904 19026 16960
rect 18694 16632 18750 16688
rect 18510 15272 18566 15328
rect 18326 13504 18382 13560
rect 18234 13232 18290 13288
rect 18602 12960 18658 13016
rect 18602 12688 18658 12744
rect 18510 12280 18566 12336
rect 17682 11328 17738 11384
rect 16854 10240 16910 10296
rect 18142 11348 18198 11384
rect 18142 11328 18144 11348
rect 18144 11328 18196 11348
rect 18196 11328 18198 11348
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 15566 9580 15622 9616
rect 15566 9560 15568 9580
rect 15568 9560 15620 9580
rect 15620 9560 15622 9580
rect 16302 9460 16304 9480
rect 16304 9460 16356 9480
rect 16356 9460 16358 9480
rect 16302 9424 16358 9460
rect 16302 9152 16358 9208
rect 15658 8744 15714 8800
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 16946 9832 17002 9888
rect 18878 16496 18934 16552
rect 19430 16360 19486 16416
rect 19338 14048 19394 14104
rect 18970 12588 18972 12608
rect 18972 12588 19024 12608
rect 19024 12588 19026 12608
rect 18970 12552 19026 12588
rect 19338 12416 19394 12472
rect 19522 15816 19578 15872
rect 19522 15408 19578 15464
rect 19522 14048 19578 14104
rect 19522 13948 19524 13968
rect 19524 13948 19576 13968
rect 19576 13948 19578 13968
rect 19522 13912 19578 13948
rect 19982 16496 20038 16552
rect 19982 16088 20038 16144
rect 19706 14592 19762 14648
rect 19982 14456 20038 14512
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20810 16940 20812 16960
rect 20812 16940 20864 16960
rect 20864 16940 20866 16960
rect 20810 16904 20866 16940
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20902 14320 20958 14376
rect 19890 12688 19946 12744
rect 19522 12416 19578 12472
rect 19706 12144 19762 12200
rect 19890 12144 19946 12200
rect 19614 11872 19670 11928
rect 19982 11056 20038 11112
rect 19706 10920 19762 10976
rect 19706 10240 19762 10296
rect 18694 9560 18750 9616
rect 16854 9424 16910 9480
rect 16854 8880 16910 8936
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 14370 7520 14426 7576
rect 19154 9172 19210 9208
rect 19154 9152 19156 9172
rect 19156 9152 19208 9172
rect 19208 9152 19210 9172
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20626 12860 20628 12880
rect 20628 12860 20680 12880
rect 20680 12860 20682 12880
rect 20626 12824 20682 12860
rect 21362 13640 21418 13696
rect 21362 12960 21418 13016
rect 20350 10648 20406 10704
rect 18878 8336 18934 8392
rect 19614 8336 19670 8392
rect 20810 12552 20866 12608
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 21270 10920 21326 10976
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 24858 21528 24914 21584
rect 23938 20304 23994 20360
rect 22006 16768 22062 16824
rect 22834 18264 22890 18320
rect 22466 16632 22522 16688
rect 22282 16088 22338 16144
rect 22558 15544 22614 15600
rect 22006 14320 22062 14376
rect 21822 13640 21878 13696
rect 21822 13388 21878 13424
rect 21822 13368 21824 13388
rect 21824 13368 21876 13388
rect 21876 13368 21878 13388
rect 21822 12280 21878 12336
rect 20718 9968 20774 10024
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 21822 10784 21878 10840
rect 21546 8880 21602 8936
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 22006 9152 22062 9208
rect 19062 7792 19118 7848
rect 19982 7384 20038 7440
rect 24214 18128 24270 18184
rect 23202 15952 23258 16008
rect 23018 13096 23074 13152
rect 22926 11464 22982 11520
rect 22742 11076 22798 11112
rect 22742 11056 22744 11076
rect 22744 11056 22796 11076
rect 22796 11056 22798 11076
rect 23478 11872 23534 11928
rect 24030 14320 24086 14376
rect 23938 13640 23994 13696
rect 23110 9424 23166 9480
rect 23938 9460 23940 9480
rect 23940 9460 23992 9480
rect 23992 9460 23994 9480
rect 23938 9424 23994 9460
rect 25042 21256 25098 21312
rect 25778 23024 25834 23080
rect 25410 20476 25412 20496
rect 25412 20476 25464 20496
rect 25464 20476 25466 20496
rect 25870 22344 25926 22400
rect 25410 20440 25466 20476
rect 25042 19352 25098 19408
rect 24950 18128 25006 18184
rect 24582 18028 24584 18048
rect 24584 18028 24636 18048
rect 24636 18028 24638 18048
rect 24582 17992 24638 18028
rect 24398 16360 24454 16416
rect 24950 16088 25006 16144
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 26606 20596 26662 20632
rect 26606 20576 26608 20596
rect 26608 20576 26660 20596
rect 26660 20576 26662 20596
rect 28998 20576 29054 20632
rect 27158 20440 27214 20496
rect 25686 19216 25742 19272
rect 25778 19080 25834 19136
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 26514 17992 26570 18048
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25502 16224 25558 16280
rect 25870 16788 25926 16824
rect 25870 16768 25872 16788
rect 25872 16768 25924 16788
rect 25924 16768 25926 16788
rect 25778 16632 25834 16688
rect 25042 15952 25098 16008
rect 24858 15816 24914 15872
rect 24766 15408 24822 15464
rect 24582 15272 24638 15328
rect 24490 14884 24546 14920
rect 24490 14864 24492 14884
rect 24492 14864 24544 14884
rect 24544 14864 24546 14884
rect 24582 12688 24638 12744
rect 24398 11328 24454 11384
rect 24950 15408 25006 15464
rect 24858 13096 24914 13152
rect 24858 11736 24914 11792
rect 25226 14592 25282 14648
rect 25686 13368 25742 13424
rect 24950 10684 24952 10704
rect 24952 10684 25004 10704
rect 25004 10684 25006 10704
rect 24950 10648 25006 10684
rect 25134 10784 25190 10840
rect 25042 10104 25098 10160
rect 24858 9832 24914 9888
rect 24674 9696 24730 9752
rect 24030 7928 24086 7984
rect 21362 7828 21364 7848
rect 21364 7828 21416 7848
rect 21416 7828 21418 7848
rect 21362 7792 21418 7828
rect 22098 7792 22154 7848
rect 24858 7656 24914 7712
rect 19706 7112 19762 7168
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 24858 6976 24914 7032
rect 13358 5072 13414 5128
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 15474 3440 15530 3496
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 11150 2352 11206 2408
rect 9034 856 9090 912
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 19706 3984 19762 4040
rect 25318 9036 25374 9072
rect 25318 9016 25320 9036
rect 25320 9016 25372 9036
rect 25372 9016 25374 9036
rect 25318 7948 25374 7984
rect 25318 7928 25320 7948
rect 25320 7928 25372 7948
rect 25372 7928 25374 7948
rect 25502 11736 25558 11792
rect 25502 11600 25558 11656
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 26790 20032 26846 20088
rect 27342 19216 27398 19272
rect 26882 19116 26884 19136
rect 26884 19116 26936 19136
rect 26936 19116 26938 19136
rect 26882 19080 26938 19116
rect 26790 18808 26846 18864
rect 26882 17740 26938 17776
rect 26882 17720 26884 17740
rect 26884 17720 26936 17740
rect 26936 17720 26938 17740
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 25870 13776 25926 13832
rect 26514 13640 26570 13696
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25870 12144 25926 12200
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 27250 14864 27306 14920
rect 26698 14456 26754 14512
rect 26698 13932 26754 13968
rect 26698 13912 26700 13932
rect 26700 13912 26752 13932
rect 26752 13912 26754 13932
rect 26882 14320 26938 14376
rect 26790 11892 26846 11928
rect 26790 11872 26792 11892
rect 26792 11872 26844 11892
rect 26844 11872 26846 11892
rect 25594 10548 25596 10568
rect 25596 10548 25648 10568
rect 25648 10548 25650 10568
rect 25594 10512 25650 10548
rect 25594 9696 25650 9752
rect 25594 9288 25650 9344
rect 25502 8472 25558 8528
rect 25502 8084 25558 8120
rect 25502 8064 25504 8084
rect 25504 8064 25556 8084
rect 25556 8064 25558 8084
rect 25410 7384 25466 7440
rect 25042 3848 25098 3904
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 25686 3440 25742 3496
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 26514 11348 26570 11384
rect 26514 11328 26516 11348
rect 26516 11328 26568 11348
rect 26568 11328 26570 11348
rect 26514 10648 26570 10704
rect 26514 9988 26570 10024
rect 26514 9968 26516 9988
rect 26516 9968 26568 9988
rect 26568 9968 26570 9988
rect 26422 9152 26478 9208
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 26514 8336 26570 8392
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 26606 7384 26662 7440
rect 26514 6976 26570 7032
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 26882 11464 26938 11520
rect 26790 7792 26846 7848
rect 26698 6296 26754 6352
rect 26606 5480 26662 5536
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 26422 5108 26424 5128
rect 26424 5108 26476 5128
rect 26476 5108 26478 5128
rect 26422 5072 26478 5108
rect 26606 5072 26662 5128
rect 25870 4528 25926 4584
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 26422 3984 26478 4040
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 26606 2796 26608 2816
rect 26608 2796 26660 2816
rect 26660 2796 26662 2816
rect 26606 2760 26662 2796
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 26790 1400 26846 1456
rect 2686 312 2742 368
rect 29366 17176 29422 17232
rect 27710 12280 27766 12336
rect 27434 12144 27490 12200
rect 27710 10376 27766 10432
rect 27526 9560 27582 9616
rect 27710 6976 27766 7032
rect 26974 5480 27030 5536
rect 26974 2080 27030 2136
rect 29366 17040 29422 17096
rect 28170 12860 28172 12880
rect 28172 12860 28224 12880
rect 28224 12860 28226 12880
rect 28170 12824 28226 12860
rect 27802 5616 27858 5672
rect 27066 856 27122 912
rect 26882 312 26938 368
<< metal3 >>
rect 0 23626 480 23656
rect 3325 23626 3391 23629
rect 0 23624 3391 23626
rect 0 23568 3330 23624
rect 3386 23568 3391 23624
rect 0 23566 3391 23568
rect 0 23536 480 23566
rect 3325 23563 3391 23566
rect 25037 23626 25103 23629
rect 29520 23626 30000 23656
rect 25037 23624 30000 23626
rect 25037 23568 25042 23624
rect 25098 23568 30000 23624
rect 25037 23566 30000 23568
rect 25037 23563 25103 23566
rect 29520 23536 30000 23566
rect 0 23082 480 23112
rect 3509 23082 3575 23085
rect 0 23080 3575 23082
rect 0 23024 3514 23080
rect 3570 23024 3575 23080
rect 0 23022 3575 23024
rect 0 22992 480 23022
rect 3509 23019 3575 23022
rect 25773 23082 25839 23085
rect 29520 23082 30000 23112
rect 25773 23080 30000 23082
rect 25773 23024 25778 23080
rect 25834 23024 30000 23080
rect 25773 23022 30000 23024
rect 25773 23019 25839 23022
rect 29520 22992 30000 23022
rect 0 22402 480 22432
rect 2865 22402 2931 22405
rect 0 22400 2931 22402
rect 0 22344 2870 22400
rect 2926 22344 2931 22400
rect 0 22342 2931 22344
rect 0 22312 480 22342
rect 2865 22339 2931 22342
rect 25865 22402 25931 22405
rect 29520 22402 30000 22432
rect 25865 22400 30000 22402
rect 25865 22344 25870 22400
rect 25926 22344 30000 22400
rect 25865 22342 30000 22344
rect 25865 22339 25931 22342
rect 29520 22312 30000 22342
rect 0 21858 480 21888
rect 3325 21858 3391 21861
rect 29520 21858 30000 21888
rect 0 21856 3391 21858
rect 0 21800 3330 21856
rect 3386 21800 3391 21856
rect 0 21798 3391 21800
rect 0 21768 480 21798
rect 3325 21795 3391 21798
rect 26374 21798 30000 21858
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 21727 26264 21728
rect 24853 21586 24919 21589
rect 26374 21586 26434 21798
rect 29520 21768 30000 21798
rect 24853 21584 26434 21586
rect 24853 21528 24858 21584
rect 24914 21528 26434 21584
rect 24853 21526 26434 21528
rect 24853 21523 24919 21526
rect 0 21314 480 21344
rect 4061 21314 4127 21317
rect 0 21312 4127 21314
rect 0 21256 4066 21312
rect 4122 21256 4127 21312
rect 0 21254 4127 21256
rect 0 21224 480 21254
rect 4061 21251 4127 21254
rect 25037 21314 25103 21317
rect 29520 21314 30000 21344
rect 25037 21312 30000 21314
rect 25037 21256 25042 21312
rect 25098 21256 30000 21312
rect 25037 21254 30000 21256
rect 25037 21251 25103 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 29520 21224 30000 21254
rect 20944 21183 21264 21184
rect 5944 20704 6264 20705
rect 0 20634 480 20664
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 2957 20634 3023 20637
rect 0 20632 3023 20634
rect 0 20576 2962 20632
rect 3018 20576 3023 20632
rect 0 20574 3023 20576
rect 0 20544 480 20574
rect 2957 20571 3023 20574
rect 26601 20634 26667 20637
rect 28993 20634 29059 20637
rect 29520 20634 30000 20664
rect 26601 20632 29059 20634
rect 26601 20576 26606 20632
rect 26662 20576 28998 20632
rect 29054 20576 29059 20632
rect 26601 20574 29059 20576
rect 26601 20571 26667 20574
rect 28993 20571 29059 20574
rect 29134 20574 30000 20634
rect 25405 20498 25471 20501
rect 27153 20498 27219 20501
rect 25405 20496 27219 20498
rect 25405 20440 25410 20496
rect 25466 20440 27158 20496
rect 27214 20440 27219 20496
rect 25405 20438 27219 20440
rect 25405 20435 25471 20438
rect 27153 20435 27219 20438
rect 19977 20362 20043 20365
rect 23933 20362 23999 20365
rect 4294 20360 23999 20362
rect 4294 20304 19982 20360
rect 20038 20304 23938 20360
rect 23994 20304 23999 20360
rect 4294 20302 23999 20304
rect 1945 20226 2011 20229
rect 3417 20226 3483 20229
rect 1945 20224 3483 20226
rect 1945 20168 1950 20224
rect 2006 20168 3422 20224
rect 3478 20168 3483 20224
rect 1945 20166 3483 20168
rect 1945 20163 2011 20166
rect 3417 20163 3483 20166
rect 0 20090 480 20120
rect 4294 20090 4354 20302
rect 19977 20299 20043 20302
rect 23933 20299 23999 20302
rect 25262 20300 25268 20364
rect 25332 20362 25338 20364
rect 29134 20362 29194 20574
rect 29520 20544 30000 20574
rect 25332 20302 29194 20362
rect 25332 20300 25338 20302
rect 10944 20160 11264 20161
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 0 20030 4354 20090
rect 4429 20090 4495 20093
rect 6545 20090 6611 20093
rect 4429 20088 6611 20090
rect 4429 20032 4434 20088
rect 4490 20032 6550 20088
rect 6606 20032 6611 20088
rect 4429 20030 6611 20032
rect 0 20000 480 20030
rect 4429 20027 4495 20030
rect 6545 20027 6611 20030
rect 26785 20090 26851 20093
rect 29520 20090 30000 20120
rect 26785 20088 30000 20090
rect 26785 20032 26790 20088
rect 26846 20032 30000 20088
rect 26785 20030 30000 20032
rect 26785 20027 26851 20030
rect 29520 20000 30000 20030
rect 10777 19954 10843 19957
rect 12801 19954 12867 19957
rect 10777 19952 12867 19954
rect 10777 19896 10782 19952
rect 10838 19896 12806 19952
rect 12862 19896 12867 19952
rect 10777 19894 12867 19896
rect 10777 19891 10843 19894
rect 12801 19891 12867 19894
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 3918 19546 3924 19548
rect 2454 19486 3924 19546
rect 0 19410 480 19440
rect 2454 19410 2514 19486
rect 3918 19484 3924 19486
rect 3988 19484 3994 19548
rect 0 19350 2514 19410
rect 2681 19410 2747 19413
rect 4613 19410 4679 19413
rect 2681 19408 4679 19410
rect 2681 19352 2686 19408
rect 2742 19352 4618 19408
rect 4674 19352 4679 19408
rect 2681 19350 4679 19352
rect 0 19320 480 19350
rect 2681 19347 2747 19350
rect 4613 19347 4679 19350
rect 9857 19410 9923 19413
rect 12065 19410 12131 19413
rect 9857 19408 12131 19410
rect 9857 19352 9862 19408
rect 9918 19352 12070 19408
rect 12126 19352 12131 19408
rect 9857 19350 12131 19352
rect 9857 19347 9923 19350
rect 12065 19347 12131 19350
rect 25037 19410 25103 19413
rect 29520 19410 30000 19440
rect 25037 19408 30000 19410
rect 25037 19352 25042 19408
rect 25098 19352 30000 19408
rect 25037 19350 30000 19352
rect 25037 19347 25103 19350
rect 29520 19320 30000 19350
rect 3693 19274 3759 19277
rect 5349 19274 5415 19277
rect 6177 19274 6243 19277
rect 3693 19272 6243 19274
rect 3693 19216 3698 19272
rect 3754 19216 5354 19272
rect 5410 19216 6182 19272
rect 6238 19216 6243 19272
rect 3693 19214 6243 19216
rect 3693 19211 3759 19214
rect 5349 19211 5415 19214
rect 6177 19211 6243 19214
rect 15745 19274 15811 19277
rect 25681 19274 25747 19277
rect 27337 19274 27403 19277
rect 15745 19272 27403 19274
rect 15745 19216 15750 19272
rect 15806 19216 25686 19272
rect 25742 19216 27342 19272
rect 27398 19216 27403 19272
rect 15745 19214 27403 19216
rect 15745 19211 15811 19214
rect 25681 19211 25747 19214
rect 27337 19211 27403 19214
rect 3877 19138 3943 19141
rect 7281 19138 7347 19141
rect 3877 19136 7347 19138
rect 3877 19080 3882 19136
rect 3938 19080 7286 19136
rect 7342 19080 7347 19136
rect 3877 19078 7347 19080
rect 3877 19075 3943 19078
rect 7281 19075 7347 19078
rect 24894 19076 24900 19140
rect 24964 19138 24970 19140
rect 25773 19138 25839 19141
rect 26877 19138 26943 19141
rect 24964 19136 26943 19138
rect 24964 19080 25778 19136
rect 25834 19080 26882 19136
rect 26938 19080 26943 19136
rect 24964 19078 26943 19080
rect 24964 19076 24970 19078
rect 25773 19075 25839 19078
rect 26877 19075 26943 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 19007 21264 19008
rect 4981 19002 5047 19005
rect 7741 19002 7807 19005
rect 4981 19000 7807 19002
rect 4981 18944 4986 19000
rect 5042 18944 7746 19000
rect 7802 18944 7807 19000
rect 4981 18942 7807 18944
rect 4981 18939 5047 18942
rect 7741 18939 7807 18942
rect 0 18866 480 18896
rect 2037 18866 2103 18869
rect 19425 18866 19491 18869
rect 26785 18866 26851 18869
rect 29520 18866 30000 18896
rect 0 18806 1778 18866
rect 0 18776 480 18806
rect 1718 18594 1778 18806
rect 2037 18864 26851 18866
rect 2037 18808 2042 18864
rect 2098 18808 19430 18864
rect 19486 18808 26790 18864
rect 26846 18808 26851 18864
rect 2037 18806 26851 18808
rect 2037 18803 2103 18806
rect 19425 18803 19491 18806
rect 26785 18803 26851 18806
rect 26926 18806 30000 18866
rect 11329 18730 11395 18733
rect 5766 18728 11395 18730
rect 5766 18672 11334 18728
rect 11390 18672 11395 18728
rect 5766 18670 11395 18672
rect 2957 18594 3023 18597
rect 5766 18594 5826 18670
rect 11329 18667 11395 18670
rect 14089 18730 14155 18733
rect 19977 18730 20043 18733
rect 26926 18730 26986 18806
rect 29520 18776 30000 18806
rect 14089 18728 20043 18730
rect 14089 18672 14094 18728
rect 14150 18672 19982 18728
rect 20038 18672 20043 18728
rect 14089 18670 20043 18672
rect 14089 18667 14155 18670
rect 19977 18667 20043 18670
rect 24028 18670 26986 18730
rect 1718 18592 5826 18594
rect 1718 18536 2962 18592
rect 3018 18536 5826 18592
rect 1718 18534 5826 18536
rect 2957 18531 3023 18534
rect 5944 18528 6264 18529
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 0 18322 480 18352
rect 3141 18322 3207 18325
rect 0 18320 3207 18322
rect 0 18264 3146 18320
rect 3202 18264 3207 18320
rect 0 18262 3207 18264
rect 0 18232 480 18262
rect 3141 18259 3207 18262
rect 3693 18322 3759 18325
rect 6821 18322 6887 18325
rect 3693 18320 6887 18322
rect 3693 18264 3698 18320
rect 3754 18264 6826 18320
rect 6882 18264 6887 18320
rect 3693 18262 6887 18264
rect 3693 18259 3759 18262
rect 6821 18259 6887 18262
rect 10777 18322 10843 18325
rect 22829 18322 22895 18325
rect 24028 18322 24088 18670
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 10777 18320 24088 18322
rect 10777 18264 10782 18320
rect 10838 18264 22834 18320
rect 22890 18264 24088 18320
rect 10777 18262 24088 18264
rect 10777 18259 10843 18262
rect 22829 18259 22895 18262
rect 25630 18260 25636 18324
rect 25700 18322 25706 18324
rect 29520 18322 30000 18352
rect 25700 18262 30000 18322
rect 25700 18260 25706 18262
rect 29520 18232 30000 18262
rect 5717 18188 5783 18189
rect 5717 18186 5764 18188
rect 5672 18184 5764 18186
rect 5672 18128 5722 18184
rect 5672 18126 5764 18128
rect 5717 18124 5764 18126
rect 5828 18124 5834 18188
rect 7925 18186 7991 18189
rect 9673 18186 9739 18189
rect 7925 18184 9739 18186
rect 7925 18128 7930 18184
rect 7986 18128 9678 18184
rect 9734 18128 9739 18184
rect 7925 18126 9739 18128
rect 5717 18123 5783 18124
rect 7925 18123 7991 18126
rect 9673 18123 9739 18126
rect 11145 18186 11211 18189
rect 19057 18186 19123 18189
rect 11145 18184 19123 18186
rect 11145 18128 11150 18184
rect 11206 18128 19062 18184
rect 19118 18128 19123 18184
rect 11145 18126 19123 18128
rect 11145 18123 11211 18126
rect 19057 18123 19123 18126
rect 19977 18186 20043 18189
rect 24209 18186 24275 18189
rect 24945 18186 25011 18189
rect 19977 18184 25011 18186
rect 19977 18128 19982 18184
rect 20038 18128 24214 18184
rect 24270 18128 24950 18184
rect 25006 18128 25011 18184
rect 19977 18126 25011 18128
rect 19977 18123 20043 18126
rect 24209 18123 24275 18126
rect 24945 18123 25011 18126
rect 12985 18052 13051 18053
rect 12934 17988 12940 18052
rect 13004 18050 13051 18052
rect 24577 18050 24643 18053
rect 26509 18050 26575 18053
rect 13004 18048 13096 18050
rect 13046 17992 13096 18048
rect 13004 17990 13096 17992
rect 24577 18048 26575 18050
rect 24577 17992 24582 18048
rect 24638 17992 26514 18048
rect 26570 17992 26575 18048
rect 24577 17990 26575 17992
rect 13004 17988 13051 17990
rect 12985 17987 13051 17988
rect 24577 17987 24643 17990
rect 26509 17987 26575 17990
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 4981 17778 5047 17781
rect 11973 17778 12039 17781
rect 26877 17778 26943 17781
rect 4981 17776 12039 17778
rect 4981 17720 4986 17776
rect 5042 17720 11978 17776
rect 12034 17720 12039 17776
rect 4981 17718 12039 17720
rect 4981 17715 5047 17718
rect 11973 17715 12039 17718
rect 12574 17776 26943 17778
rect 12574 17720 26882 17776
rect 26938 17720 26943 17776
rect 12574 17718 26943 17720
rect 0 17642 480 17672
rect 9857 17642 9923 17645
rect 12574 17642 12634 17718
rect 26877 17715 26943 17718
rect 0 17640 9923 17642
rect 0 17584 9862 17640
rect 9918 17584 9923 17640
rect 0 17582 9923 17584
rect 0 17552 480 17582
rect 9857 17579 9923 17582
rect 12252 17582 12634 17642
rect 18321 17642 18387 17645
rect 29520 17642 30000 17672
rect 18321 17640 30000 17642
rect 18321 17584 18326 17640
rect 18382 17584 30000 17640
rect 18321 17582 30000 17584
rect 6453 17506 6519 17509
rect 12252 17506 12312 17582
rect 18321 17579 18387 17582
rect 29520 17552 30000 17582
rect 6453 17504 12312 17506
rect 6453 17448 6458 17504
rect 6514 17448 12312 17504
rect 6453 17446 12312 17448
rect 6453 17443 6519 17446
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 8937 17234 9003 17237
rect 13537 17234 13603 17237
rect 29361 17234 29427 17237
rect 8937 17232 29427 17234
rect 8937 17176 8942 17232
rect 8998 17176 13542 17232
rect 13598 17176 29366 17232
rect 29422 17176 29427 17232
rect 8937 17174 29427 17176
rect 8937 17171 9003 17174
rect 13537 17171 13603 17174
rect 29361 17171 29427 17174
rect 0 17098 480 17128
rect 6453 17098 6519 17101
rect 0 17096 6519 17098
rect 0 17040 6458 17096
rect 6514 17040 6519 17096
rect 0 17038 6519 17040
rect 0 17008 480 17038
rect 6453 17035 6519 17038
rect 29361 17098 29427 17101
rect 29520 17098 30000 17128
rect 29361 17096 30000 17098
rect 29361 17040 29366 17096
rect 29422 17040 30000 17096
rect 29361 17038 30000 17040
rect 29361 17035 29427 17038
rect 29520 17008 30000 17038
rect 18965 16962 19031 16965
rect 20805 16962 20871 16965
rect 18965 16960 20871 16962
rect 18965 16904 18970 16960
rect 19026 16904 20810 16960
rect 20866 16904 20871 16960
rect 18965 16902 20871 16904
rect 18965 16899 19031 16902
rect 20805 16899 20871 16902
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 22001 16826 22067 16829
rect 25865 16826 25931 16829
rect 22001 16824 25931 16826
rect 22001 16768 22006 16824
rect 22062 16768 25870 16824
rect 25926 16768 25931 16824
rect 22001 16766 25931 16768
rect 22001 16763 22067 16766
rect 25865 16763 25931 16766
rect 9857 16690 9923 16693
rect 10501 16690 10567 16693
rect 18689 16690 18755 16693
rect 9857 16688 18755 16690
rect 9857 16632 9862 16688
rect 9918 16632 10506 16688
rect 10562 16632 18694 16688
rect 18750 16632 18755 16688
rect 9857 16630 18755 16632
rect 9857 16627 9923 16630
rect 10501 16627 10567 16630
rect 18689 16627 18755 16630
rect 22461 16690 22527 16693
rect 25773 16690 25839 16693
rect 22461 16688 25839 16690
rect 22461 16632 22466 16688
rect 22522 16632 25778 16688
rect 25834 16632 25839 16688
rect 22461 16630 25839 16632
rect 22461 16627 22527 16630
rect 25773 16627 25839 16630
rect 17033 16554 17099 16557
rect 18873 16554 18939 16557
rect 19977 16554 20043 16557
rect 5720 16494 16866 16554
rect 0 16418 480 16448
rect 5720 16421 5780 16494
rect 5717 16418 5783 16421
rect 0 16416 5783 16418
rect 0 16360 5722 16416
rect 5778 16360 5783 16416
rect 0 16358 5783 16360
rect 0 16328 480 16358
rect 5717 16355 5783 16358
rect 7281 16418 7347 16421
rect 10777 16418 10843 16421
rect 11145 16418 11211 16421
rect 7281 16416 11211 16418
rect 7281 16360 7286 16416
rect 7342 16360 10782 16416
rect 10838 16360 11150 16416
rect 11206 16360 11211 16416
rect 7281 16358 11211 16360
rect 16806 16418 16866 16494
rect 17033 16552 20043 16554
rect 17033 16496 17038 16552
rect 17094 16496 18878 16552
rect 18934 16496 19982 16552
rect 20038 16496 20043 16552
rect 17033 16494 20043 16496
rect 17033 16491 17099 16494
rect 18873 16491 18939 16494
rect 19977 16491 20043 16494
rect 19425 16418 19491 16421
rect 24393 16418 24459 16421
rect 29520 16418 30000 16448
rect 16806 16416 24459 16418
rect 16806 16360 19430 16416
rect 19486 16360 24398 16416
rect 24454 16360 24459 16416
rect 16806 16358 24459 16360
rect 7281 16355 7347 16358
rect 10777 16355 10843 16358
rect 11145 16355 11211 16358
rect 19425 16355 19491 16358
rect 24393 16355 24459 16358
rect 26374 16358 30000 16418
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 9305 16282 9371 16285
rect 12341 16282 12407 16285
rect 25497 16282 25563 16285
rect 9305 16280 12407 16282
rect 9305 16224 9310 16280
rect 9366 16224 12346 16280
rect 12402 16224 12407 16280
rect 9305 16222 12407 16224
rect 9305 16219 9371 16222
rect 12341 16219 12407 16222
rect 24718 16280 25563 16282
rect 24718 16224 25502 16280
rect 25558 16224 25563 16280
rect 24718 16222 25563 16224
rect 11513 16146 11579 16149
rect 15745 16146 15811 16149
rect 11513 16144 15811 16146
rect 11513 16088 11518 16144
rect 11574 16088 15750 16144
rect 15806 16088 15811 16144
rect 11513 16086 15811 16088
rect 11513 16083 11579 16086
rect 15745 16083 15811 16086
rect 19977 16146 20043 16149
rect 22277 16146 22343 16149
rect 24718 16146 24778 16222
rect 25497 16219 25563 16222
rect 19977 16144 24778 16146
rect 19977 16088 19982 16144
rect 20038 16088 22282 16144
rect 22338 16088 24778 16144
rect 19977 16086 24778 16088
rect 24945 16146 25011 16149
rect 26374 16146 26434 16358
rect 29520 16328 30000 16358
rect 24945 16144 26434 16146
rect 24945 16088 24950 16144
rect 25006 16088 26434 16144
rect 24945 16086 26434 16088
rect 19977 16083 20043 16086
rect 22277 16083 22343 16086
rect 24945 16083 25011 16086
rect 15561 16010 15627 16013
rect 23197 16010 23263 16013
rect 25037 16010 25103 16013
rect 15561 16008 25103 16010
rect 15561 15952 15566 16008
rect 15622 15952 23202 16008
rect 23258 15952 25042 16008
rect 25098 15952 25103 16008
rect 15561 15950 25103 15952
rect 15561 15947 15627 15950
rect 23197 15947 23263 15950
rect 25037 15947 25103 15950
rect 0 15874 480 15904
rect 749 15874 815 15877
rect 0 15872 815 15874
rect 0 15816 754 15872
rect 810 15816 815 15872
rect 0 15814 815 15816
rect 0 15784 480 15814
rect 749 15811 815 15814
rect 2037 15874 2103 15877
rect 4521 15874 4587 15877
rect 2037 15872 4587 15874
rect 2037 15816 2042 15872
rect 2098 15816 4526 15872
rect 4582 15816 4587 15872
rect 2037 15814 4587 15816
rect 2037 15811 2103 15814
rect 4521 15811 4587 15814
rect 7557 15874 7623 15877
rect 10593 15874 10659 15877
rect 7557 15872 10659 15874
rect 7557 15816 7562 15872
rect 7618 15816 10598 15872
rect 10654 15816 10659 15872
rect 7557 15814 10659 15816
rect 7557 15811 7623 15814
rect 10593 15811 10659 15814
rect 12525 15874 12591 15877
rect 12893 15874 12959 15877
rect 19517 15874 19583 15877
rect 12525 15872 19583 15874
rect 12525 15816 12530 15872
rect 12586 15816 12898 15872
rect 12954 15816 19522 15872
rect 19578 15816 19583 15872
rect 12525 15814 19583 15816
rect 12525 15811 12591 15814
rect 12893 15811 12959 15814
rect 19517 15811 19583 15814
rect 24853 15874 24919 15877
rect 29520 15874 30000 15904
rect 24853 15872 30000 15874
rect 24853 15816 24858 15872
rect 24914 15816 30000 15872
rect 24853 15814 30000 15816
rect 24853 15811 24919 15814
rect 10944 15808 11264 15809
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 29520 15784 30000 15814
rect 20944 15743 21264 15744
rect 3141 15738 3207 15741
rect 7925 15738 7991 15741
rect 8385 15738 8451 15741
rect 3141 15736 8451 15738
rect 3141 15680 3146 15736
rect 3202 15680 7930 15736
rect 7986 15680 8390 15736
rect 8446 15680 8451 15736
rect 3141 15678 8451 15680
rect 3141 15675 3207 15678
rect 7925 15675 7991 15678
rect 8385 15675 8451 15678
rect 2037 15602 2103 15605
rect 4613 15602 4679 15605
rect 2037 15600 4679 15602
rect 2037 15544 2042 15600
rect 2098 15544 4618 15600
rect 4674 15544 4679 15600
rect 2037 15542 4679 15544
rect 2037 15539 2103 15542
rect 4613 15539 4679 15542
rect 8109 15602 8175 15605
rect 15377 15602 15443 15605
rect 22553 15602 22619 15605
rect 8109 15600 22619 15602
rect 8109 15544 8114 15600
rect 8170 15544 15382 15600
rect 15438 15544 22558 15600
rect 22614 15544 22619 15600
rect 8109 15542 22619 15544
rect 8109 15539 8175 15542
rect 15377 15539 15443 15542
rect 22553 15539 22619 15542
rect 19517 15466 19583 15469
rect 24761 15466 24827 15469
rect 19517 15464 24827 15466
rect 19517 15408 19522 15464
rect 19578 15408 24766 15464
rect 24822 15408 24827 15464
rect 19517 15406 24827 15408
rect 19517 15403 19583 15406
rect 24761 15403 24827 15406
rect 24945 15466 25011 15469
rect 24945 15464 26434 15466
rect 24945 15408 24950 15464
rect 25006 15408 26434 15464
rect 24945 15406 26434 15408
rect 24945 15403 25011 15406
rect 0 15330 480 15360
rect 3785 15330 3851 15333
rect 0 15328 3851 15330
rect 0 15272 3790 15328
rect 3846 15272 3851 15328
rect 0 15270 3851 15272
rect 0 15240 480 15270
rect 3785 15267 3851 15270
rect 18505 15330 18571 15333
rect 24577 15330 24643 15333
rect 18505 15328 24643 15330
rect 18505 15272 18510 15328
rect 18566 15272 24582 15328
rect 24638 15272 24643 15328
rect 18505 15270 24643 15272
rect 26374 15330 26434 15406
rect 29520 15330 30000 15360
rect 26374 15270 30000 15330
rect 18505 15267 18571 15270
rect 24577 15267 24643 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 29520 15240 30000 15270
rect 25944 15199 26264 15200
rect 13629 15194 13695 15197
rect 6502 15192 13695 15194
rect 6502 15136 13634 15192
rect 13690 15136 13695 15192
rect 6502 15134 13695 15136
rect 4061 15058 4127 15061
rect 6502 15058 6562 15134
rect 13629 15131 13695 15134
rect 4061 15056 6562 15058
rect 4061 15000 4066 15056
rect 4122 15000 6562 15056
rect 4061 14998 6562 15000
rect 6637 15058 6703 15061
rect 10409 15058 10475 15061
rect 16021 15058 16087 15061
rect 6637 15056 16087 15058
rect 6637 15000 6642 15056
rect 6698 15000 10414 15056
rect 10470 15000 16026 15056
rect 16082 15000 16087 15056
rect 6637 14998 16087 15000
rect 4061 14995 4127 14998
rect 6637 14995 6703 14998
rect 10409 14995 10475 14998
rect 16021 14995 16087 14998
rect 5625 14922 5691 14925
rect 7281 14922 7347 14925
rect 10317 14922 10383 14925
rect 14733 14922 14799 14925
rect 5625 14920 14799 14922
rect 5625 14864 5630 14920
rect 5686 14864 7286 14920
rect 7342 14864 10322 14920
rect 10378 14864 14738 14920
rect 14794 14864 14799 14920
rect 5625 14862 14799 14864
rect 5625 14859 5691 14862
rect 7281 14859 7347 14862
rect 10317 14859 10383 14862
rect 14733 14859 14799 14862
rect 24485 14922 24551 14925
rect 27245 14922 27311 14925
rect 24485 14920 27311 14922
rect 24485 14864 24490 14920
rect 24546 14864 27250 14920
rect 27306 14864 27311 14920
rect 24485 14862 27311 14864
rect 24485 14859 24551 14862
rect 27245 14859 27311 14862
rect 2405 14786 2471 14789
rect 2865 14786 2931 14789
rect 8293 14786 8359 14789
rect 2405 14784 8359 14786
rect 2405 14728 2410 14784
rect 2466 14728 2870 14784
rect 2926 14728 8298 14784
rect 8354 14728 8359 14784
rect 2405 14726 8359 14728
rect 2405 14723 2471 14726
rect 2865 14723 2931 14726
rect 8293 14723 8359 14726
rect 10944 14720 11264 14721
rect 0 14650 480 14680
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 6545 14650 6611 14653
rect 14457 14652 14523 14653
rect 0 14648 6611 14650
rect 0 14592 6550 14648
rect 6606 14592 6611 14648
rect 0 14590 6611 14592
rect 0 14560 480 14590
rect 6545 14587 6611 14590
rect 14406 14588 14412 14652
rect 14476 14650 14523 14652
rect 17401 14650 17467 14653
rect 19701 14650 19767 14653
rect 14476 14648 14568 14650
rect 14518 14592 14568 14648
rect 14476 14590 14568 14592
rect 17401 14648 19767 14650
rect 17401 14592 17406 14648
rect 17462 14592 19706 14648
rect 19762 14592 19767 14648
rect 17401 14590 19767 14592
rect 14476 14588 14523 14590
rect 14457 14587 14523 14588
rect 17401 14587 17467 14590
rect 19701 14587 19767 14590
rect 25221 14650 25287 14653
rect 29520 14650 30000 14680
rect 25221 14648 30000 14650
rect 25221 14592 25226 14648
rect 25282 14592 30000 14648
rect 25221 14590 30000 14592
rect 25221 14587 25287 14590
rect 29520 14560 30000 14590
rect 10869 14514 10935 14517
rect 15653 14514 15719 14517
rect 10869 14512 15719 14514
rect 10869 14456 10874 14512
rect 10930 14456 15658 14512
rect 15714 14456 15719 14512
rect 10869 14454 15719 14456
rect 10869 14451 10935 14454
rect 15653 14451 15719 14454
rect 19977 14514 20043 14517
rect 26693 14514 26759 14517
rect 19977 14512 26759 14514
rect 19977 14456 19982 14512
rect 20038 14456 26698 14512
rect 26754 14456 26759 14512
rect 19977 14454 26759 14456
rect 19977 14451 20043 14454
rect 26693 14451 26759 14454
rect 15009 14378 15075 14381
rect 20897 14378 20963 14381
rect 22001 14378 22067 14381
rect 15009 14376 22067 14378
rect 15009 14320 15014 14376
rect 15070 14320 20902 14376
rect 20958 14320 22006 14376
rect 22062 14320 22067 14376
rect 15009 14318 22067 14320
rect 15009 14315 15075 14318
rect 20897 14315 20963 14318
rect 22001 14315 22067 14318
rect 24025 14378 24091 14381
rect 26877 14378 26943 14381
rect 24025 14376 26943 14378
rect 24025 14320 24030 14376
rect 24086 14320 26882 14376
rect 26938 14320 26943 14376
rect 24025 14318 26943 14320
rect 24025 14315 24091 14318
rect 26877 14315 26943 14318
rect 11329 14242 11395 14245
rect 13813 14242 13879 14245
rect 11329 14240 13879 14242
rect 11329 14184 11334 14240
rect 11390 14184 13818 14240
rect 13874 14184 13879 14240
rect 11329 14182 13879 14184
rect 11329 14179 11395 14182
rect 13813 14179 13879 14182
rect 5944 14176 6264 14177
rect 0 14106 480 14136
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 4981 14106 5047 14109
rect 5349 14106 5415 14109
rect 0 14104 5415 14106
rect 0 14048 4986 14104
rect 5042 14048 5354 14104
rect 5410 14048 5415 14104
rect 0 14046 5415 14048
rect 0 14016 480 14046
rect 4981 14043 5047 14046
rect 5349 14043 5415 14046
rect 19333 14106 19399 14109
rect 19517 14106 19583 14109
rect 29520 14106 30000 14136
rect 19333 14104 19583 14106
rect 19333 14048 19338 14104
rect 19394 14048 19522 14104
rect 19578 14048 19583 14104
rect 19333 14046 19583 14048
rect 19333 14043 19399 14046
rect 19517 14043 19583 14046
rect 26926 14046 30000 14106
rect 19517 13970 19583 13973
rect 26693 13970 26759 13973
rect 19517 13968 26759 13970
rect 19517 13912 19522 13968
rect 19578 13912 26698 13968
rect 26754 13912 26759 13968
rect 19517 13910 26759 13912
rect 19517 13907 19583 13910
rect 26693 13907 26759 13910
rect 8293 13834 8359 13837
rect 13537 13834 13603 13837
rect 8293 13832 13603 13834
rect 8293 13776 8298 13832
rect 8354 13776 13542 13832
rect 13598 13776 13603 13832
rect 8293 13774 13603 13776
rect 8293 13771 8359 13774
rect 13537 13771 13603 13774
rect 25865 13834 25931 13837
rect 26926 13834 26986 14046
rect 29520 14016 30000 14046
rect 25865 13832 26986 13834
rect 25865 13776 25870 13832
rect 25926 13776 26986 13832
rect 25865 13774 26986 13776
rect 25865 13771 25931 13774
rect 4245 13698 4311 13701
rect 8937 13698 9003 13701
rect 4245 13696 9003 13698
rect 4245 13640 4250 13696
rect 4306 13640 8942 13696
rect 8998 13640 9003 13696
rect 4245 13638 9003 13640
rect 4245 13635 4311 13638
rect 8937 13635 9003 13638
rect 21357 13698 21423 13701
rect 21817 13698 21883 13701
rect 21357 13696 21883 13698
rect 21357 13640 21362 13696
rect 21418 13640 21822 13696
rect 21878 13640 21883 13696
rect 21357 13638 21883 13640
rect 21357 13635 21423 13638
rect 21817 13635 21883 13638
rect 23933 13698 23999 13701
rect 26509 13698 26575 13701
rect 23933 13696 26575 13698
rect 23933 13640 23938 13696
rect 23994 13640 26514 13696
rect 26570 13640 26575 13696
rect 23933 13638 26575 13640
rect 23933 13635 23999 13638
rect 26509 13635 26575 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 13567 21264 13568
rect 3969 13562 4035 13565
rect 4429 13562 4495 13565
rect 3969 13560 4495 13562
rect 3969 13504 3974 13560
rect 4030 13504 4434 13560
rect 4490 13504 4495 13560
rect 3969 13502 4495 13504
rect 3969 13499 4035 13502
rect 4429 13499 4495 13502
rect 5625 13562 5691 13565
rect 6269 13562 6335 13565
rect 10777 13562 10843 13565
rect 5625 13560 10843 13562
rect 5625 13504 5630 13560
rect 5686 13504 6274 13560
rect 6330 13504 10782 13560
rect 10838 13504 10843 13560
rect 5625 13502 10843 13504
rect 5625 13499 5691 13502
rect 6269 13499 6335 13502
rect 10777 13499 10843 13502
rect 12249 13562 12315 13565
rect 18321 13562 18387 13565
rect 12249 13560 18387 13562
rect 12249 13504 12254 13560
rect 12310 13504 18326 13560
rect 18382 13504 18387 13560
rect 12249 13502 18387 13504
rect 12249 13499 12315 13502
rect 18321 13499 18387 13502
rect 0 13426 480 13456
rect 3509 13426 3575 13429
rect 0 13424 3575 13426
rect 0 13368 3514 13424
rect 3570 13368 3575 13424
rect 0 13366 3575 13368
rect 0 13336 480 13366
rect 3509 13363 3575 13366
rect 4705 13426 4771 13429
rect 14089 13426 14155 13429
rect 21817 13426 21883 13429
rect 4705 13424 21883 13426
rect 4705 13368 4710 13424
rect 4766 13368 14094 13424
rect 14150 13368 21822 13424
rect 21878 13368 21883 13424
rect 4705 13366 21883 13368
rect 4705 13363 4771 13366
rect 14089 13363 14155 13366
rect 21817 13363 21883 13366
rect 25681 13426 25747 13429
rect 29520 13426 30000 13456
rect 25681 13424 30000 13426
rect 25681 13368 25686 13424
rect 25742 13368 30000 13424
rect 25681 13366 30000 13368
rect 25681 13363 25747 13366
rect 29520 13336 30000 13366
rect 2037 13290 2103 13293
rect 9622 13290 9628 13292
rect 2037 13288 9628 13290
rect 2037 13232 2042 13288
rect 2098 13232 9628 13288
rect 2037 13230 9628 13232
rect 2037 13227 2103 13230
rect 9622 13228 9628 13230
rect 9692 13228 9698 13292
rect 16297 13290 16363 13293
rect 18229 13290 18295 13293
rect 16297 13288 18295 13290
rect 16297 13232 16302 13288
rect 16358 13232 18234 13288
rect 18290 13232 18295 13288
rect 16297 13230 18295 13232
rect 16297 13227 16363 13230
rect 18229 13227 18295 13230
rect 6453 13154 6519 13157
rect 12157 13154 12223 13157
rect 13353 13154 13419 13157
rect 6453 13152 12223 13154
rect 6453 13096 6458 13152
rect 6514 13096 12162 13152
rect 12218 13096 12223 13152
rect 6453 13094 12223 13096
rect 6453 13091 6519 13094
rect 12157 13091 12223 13094
rect 13310 13152 13419 13154
rect 13310 13096 13358 13152
rect 13414 13096 13419 13152
rect 13310 13091 13419 13096
rect 23013 13154 23079 13157
rect 24853 13154 24919 13157
rect 23013 13152 24919 13154
rect 23013 13096 23018 13152
rect 23074 13096 24858 13152
rect 24914 13096 24919 13152
rect 23013 13094 24919 13096
rect 23013 13091 23079 13094
rect 24853 13091 24919 13094
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 7373 13018 7439 13021
rect 13310 13018 13370 13091
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 7373 13016 13370 13018
rect 7373 12960 7378 13016
rect 7434 12960 13370 13016
rect 7373 12958 13370 12960
rect 18597 13018 18663 13021
rect 21357 13018 21423 13021
rect 18597 13016 21423 13018
rect 18597 12960 18602 13016
rect 18658 12960 21362 13016
rect 21418 12960 21423 13016
rect 18597 12958 21423 12960
rect 7373 12955 7439 12958
rect 18597 12955 18663 12958
rect 21357 12955 21423 12958
rect 0 12882 480 12912
rect 0 12822 2744 12882
rect 0 12792 480 12822
rect 2684 12746 2744 12822
rect 9622 12820 9628 12884
rect 9692 12882 9698 12884
rect 13629 12882 13695 12885
rect 20621 12882 20687 12885
rect 9692 12880 20687 12882
rect 9692 12824 13634 12880
rect 13690 12824 20626 12880
rect 20682 12824 20687 12880
rect 9692 12822 20687 12824
rect 9692 12820 9698 12822
rect 13629 12819 13695 12822
rect 20621 12819 20687 12822
rect 28165 12882 28231 12885
rect 29520 12882 30000 12912
rect 28165 12880 30000 12882
rect 28165 12824 28170 12880
rect 28226 12824 30000 12880
rect 28165 12822 30000 12824
rect 28165 12819 28231 12822
rect 29520 12792 30000 12822
rect 4981 12746 5047 12749
rect 2684 12744 5047 12746
rect 2684 12688 4986 12744
rect 5042 12688 5047 12744
rect 2684 12686 5047 12688
rect 4981 12683 5047 12686
rect 5165 12746 5231 12749
rect 6913 12746 6979 12749
rect 12157 12746 12223 12749
rect 18597 12746 18663 12749
rect 5165 12744 6979 12746
rect 5165 12688 5170 12744
rect 5226 12688 6918 12744
rect 6974 12688 6979 12744
rect 5165 12686 6979 12688
rect 5165 12683 5231 12686
rect 6913 12683 6979 12686
rect 7974 12744 18663 12746
rect 7974 12688 12162 12744
rect 12218 12688 18602 12744
rect 18658 12688 18663 12744
rect 7974 12686 18663 12688
rect 4429 12610 4495 12613
rect 7974 12610 8034 12686
rect 12157 12683 12223 12686
rect 18597 12683 18663 12686
rect 19885 12746 19951 12749
rect 24577 12746 24643 12749
rect 19885 12744 24643 12746
rect 19885 12688 19890 12744
rect 19946 12688 24582 12744
rect 24638 12688 24643 12744
rect 19885 12686 24643 12688
rect 19885 12683 19951 12686
rect 24577 12683 24643 12686
rect 4429 12608 8034 12610
rect 4429 12552 4434 12608
rect 4490 12552 8034 12608
rect 4429 12550 8034 12552
rect 14917 12610 14983 12613
rect 15101 12610 15167 12613
rect 18965 12610 19031 12613
rect 20805 12610 20871 12613
rect 14917 12608 20871 12610
rect 14917 12552 14922 12608
rect 14978 12552 15106 12608
rect 15162 12552 18970 12608
rect 19026 12552 20810 12608
rect 20866 12552 20871 12608
rect 14917 12550 20871 12552
rect 4429 12547 4495 12550
rect 14917 12547 14983 12550
rect 15101 12547 15167 12550
rect 18965 12547 19031 12550
rect 20805 12547 20871 12550
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 19333 12474 19399 12477
rect 19517 12474 19583 12477
rect 19333 12472 19583 12474
rect 19333 12416 19338 12472
rect 19394 12416 19522 12472
rect 19578 12416 19583 12472
rect 19333 12414 19583 12416
rect 19333 12411 19399 12414
rect 19517 12411 19583 12414
rect 0 12338 480 12368
rect 4613 12338 4679 12341
rect 0 12336 4679 12338
rect 0 12280 4618 12336
rect 4674 12280 4679 12336
rect 0 12278 4679 12280
rect 0 12248 480 12278
rect 4613 12275 4679 12278
rect 12985 12338 13051 12341
rect 18505 12338 18571 12341
rect 12985 12336 18571 12338
rect 12985 12280 12990 12336
rect 13046 12280 18510 12336
rect 18566 12280 18571 12336
rect 12985 12278 18571 12280
rect 12985 12275 13051 12278
rect 18505 12275 18571 12278
rect 21817 12338 21883 12341
rect 27705 12338 27771 12341
rect 29520 12338 30000 12368
rect 21817 12336 30000 12338
rect 21817 12280 21822 12336
rect 21878 12280 27710 12336
rect 27766 12280 30000 12336
rect 21817 12278 30000 12280
rect 21817 12275 21883 12278
rect 27705 12275 27771 12278
rect 29520 12248 30000 12278
rect 8569 12202 8635 12205
rect 12985 12202 13051 12205
rect 14917 12202 14983 12205
rect 8569 12200 14983 12202
rect 8569 12144 8574 12200
rect 8630 12144 12990 12200
rect 13046 12144 14922 12200
rect 14978 12144 14983 12200
rect 8569 12142 14983 12144
rect 8569 12139 8635 12142
rect 12985 12139 13051 12142
rect 14917 12139 14983 12142
rect 15285 12202 15351 12205
rect 19701 12202 19767 12205
rect 19885 12202 19951 12205
rect 15285 12200 19951 12202
rect 15285 12144 15290 12200
rect 15346 12144 19706 12200
rect 19762 12144 19890 12200
rect 19946 12144 19951 12200
rect 15285 12142 19951 12144
rect 15285 12139 15351 12142
rect 19701 12139 19767 12142
rect 19885 12139 19951 12142
rect 25865 12202 25931 12205
rect 27429 12202 27495 12205
rect 25865 12200 27495 12202
rect 25865 12144 25870 12200
rect 25926 12144 27434 12200
rect 27490 12144 27495 12200
rect 25865 12142 27495 12144
rect 25865 12139 25931 12142
rect 27429 12139 27495 12142
rect 3877 12066 3943 12069
rect 5717 12066 5783 12069
rect 3877 12064 5783 12066
rect 3877 12008 3882 12064
rect 3938 12008 5722 12064
rect 5778 12008 5783 12064
rect 3877 12006 5783 12008
rect 3877 12003 3943 12006
rect 5717 12003 5783 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 19609 11930 19675 11933
rect 23473 11930 23539 11933
rect 26785 11932 26851 11933
rect 19609 11928 23539 11930
rect 19609 11872 19614 11928
rect 19670 11872 23478 11928
rect 23534 11872 23539 11928
rect 19609 11870 23539 11872
rect 19609 11867 19675 11870
rect 23473 11867 23539 11870
rect 26734 11868 26740 11932
rect 26804 11930 26851 11932
rect 26804 11928 26896 11930
rect 26846 11872 26896 11928
rect 26804 11870 26896 11872
rect 26804 11868 26851 11870
rect 26785 11867 26851 11868
rect 2129 11794 2195 11797
rect 10041 11794 10107 11797
rect 2129 11792 10107 11794
rect 2129 11736 2134 11792
rect 2190 11736 10046 11792
rect 10102 11736 10107 11792
rect 2129 11734 10107 11736
rect 2129 11731 2195 11734
rect 10041 11731 10107 11734
rect 24853 11794 24919 11797
rect 25497 11794 25563 11797
rect 24853 11792 25563 11794
rect 24853 11736 24858 11792
rect 24914 11736 25502 11792
rect 25558 11736 25563 11792
rect 24853 11734 25563 11736
rect 24853 11731 24919 11734
rect 25497 11731 25563 11734
rect 0 11658 480 11688
rect 3969 11658 4035 11661
rect 0 11656 4035 11658
rect 0 11600 3974 11656
rect 4030 11600 4035 11656
rect 0 11598 4035 11600
rect 0 11568 480 11598
rect 3969 11595 4035 11598
rect 10593 11658 10659 11661
rect 12065 11658 12131 11661
rect 15837 11658 15903 11661
rect 10593 11656 15903 11658
rect 10593 11600 10598 11656
rect 10654 11600 12070 11656
rect 12126 11600 15842 11656
rect 15898 11600 15903 11656
rect 10593 11598 15903 11600
rect 10593 11595 10659 11598
rect 12065 11595 12131 11598
rect 15837 11595 15903 11598
rect 25497 11658 25563 11661
rect 29520 11658 30000 11688
rect 25497 11656 30000 11658
rect 25497 11600 25502 11656
rect 25558 11600 30000 11656
rect 25497 11598 30000 11600
rect 25497 11595 25563 11598
rect 29520 11568 30000 11598
rect 5625 11522 5691 11525
rect 8477 11522 8543 11525
rect 5625 11520 8543 11522
rect 5625 11464 5630 11520
rect 5686 11464 8482 11520
rect 8538 11464 8543 11520
rect 5625 11462 8543 11464
rect 5625 11459 5691 11462
rect 8477 11459 8543 11462
rect 13261 11522 13327 11525
rect 15377 11522 15443 11525
rect 13261 11520 15443 11522
rect 13261 11464 13266 11520
rect 13322 11464 15382 11520
rect 15438 11464 15443 11520
rect 13261 11462 15443 11464
rect 13261 11459 13327 11462
rect 15377 11459 15443 11462
rect 22921 11522 22987 11525
rect 26877 11522 26943 11525
rect 22921 11520 26943 11522
rect 22921 11464 22926 11520
rect 22982 11464 26882 11520
rect 26938 11464 26943 11520
rect 22921 11462 26943 11464
rect 22921 11459 22987 11462
rect 26877 11459 26943 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 3417 11386 3483 11389
rect 4153 11386 4219 11389
rect 3417 11384 4219 11386
rect 3417 11328 3422 11384
rect 3478 11328 4158 11384
rect 4214 11328 4219 11384
rect 3417 11326 4219 11328
rect 3417 11323 3483 11326
rect 4153 11323 4219 11326
rect 5533 11386 5599 11389
rect 6729 11386 6795 11389
rect 8845 11386 8911 11389
rect 5533 11384 8911 11386
rect 5533 11328 5538 11384
rect 5594 11328 6734 11384
rect 6790 11328 8850 11384
rect 8906 11328 8911 11384
rect 5533 11326 8911 11328
rect 5533 11323 5599 11326
rect 6729 11323 6795 11326
rect 8845 11323 8911 11326
rect 16389 11386 16455 11389
rect 17677 11386 17743 11389
rect 18137 11386 18203 11389
rect 16389 11384 18203 11386
rect 16389 11328 16394 11384
rect 16450 11328 17682 11384
rect 17738 11328 18142 11384
rect 18198 11328 18203 11384
rect 16389 11326 18203 11328
rect 16389 11323 16455 11326
rect 17677 11323 17743 11326
rect 18137 11323 18203 11326
rect 24393 11386 24459 11389
rect 26509 11386 26575 11389
rect 24393 11384 26575 11386
rect 24393 11328 24398 11384
rect 24454 11328 26514 11384
rect 26570 11328 26575 11384
rect 24393 11326 26575 11328
rect 24393 11323 24459 11326
rect 26509 11323 26575 11326
rect 8385 11250 8451 11253
rect 8518 11250 8524 11252
rect 8385 11248 8524 11250
rect 8385 11192 8390 11248
rect 8446 11192 8524 11248
rect 8385 11190 8524 11192
rect 8385 11187 8451 11190
rect 8518 11188 8524 11190
rect 8588 11188 8594 11252
rect 10685 11250 10751 11253
rect 11605 11250 11671 11253
rect 16205 11250 16271 11253
rect 16481 11252 16547 11253
rect 10685 11248 16271 11250
rect 10685 11192 10690 11248
rect 10746 11192 11610 11248
rect 11666 11192 16210 11248
rect 16266 11192 16271 11248
rect 10685 11190 16271 11192
rect 10685 11187 10751 11190
rect 11605 11187 11671 11190
rect 16205 11187 16271 11190
rect 16430 11188 16436 11252
rect 16500 11250 16547 11252
rect 16500 11248 16592 11250
rect 16542 11192 16592 11248
rect 16500 11190 16592 11192
rect 16500 11188 16547 11190
rect 16481 11187 16547 11188
rect 0 11114 480 11144
rect 7097 11114 7163 11117
rect 0 11112 7163 11114
rect 0 11056 7102 11112
rect 7158 11056 7163 11112
rect 0 11054 7163 11056
rect 0 11024 480 11054
rect 7097 11051 7163 11054
rect 16757 11114 16823 11117
rect 19977 11114 20043 11117
rect 16757 11112 20043 11114
rect 16757 11056 16762 11112
rect 16818 11056 19982 11112
rect 20038 11056 20043 11112
rect 16757 11054 20043 11056
rect 16757 11051 16823 11054
rect 19977 11051 20043 11054
rect 22737 11114 22803 11117
rect 29520 11114 30000 11144
rect 22737 11112 30000 11114
rect 22737 11056 22742 11112
rect 22798 11056 30000 11112
rect 22737 11054 30000 11056
rect 22737 11051 22803 11054
rect 29520 11024 30000 11054
rect 19701 10978 19767 10981
rect 21265 10978 21331 10981
rect 19701 10976 21331 10978
rect 19701 10920 19706 10976
rect 19762 10920 21270 10976
rect 21326 10920 21331 10976
rect 19701 10918 21331 10920
rect 19701 10915 19767 10918
rect 21265 10915 21331 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 7005 10842 7071 10845
rect 10133 10842 10199 10845
rect 21817 10842 21883 10845
rect 25129 10842 25195 10845
rect 7005 10840 10199 10842
rect 7005 10784 7010 10840
rect 7066 10784 10138 10840
rect 10194 10784 10199 10840
rect 7005 10782 10199 10784
rect 7005 10779 7071 10782
rect 10133 10779 10199 10782
rect 19566 10840 25195 10842
rect 19566 10784 21822 10840
rect 21878 10784 25134 10840
rect 25190 10784 25195 10840
rect 19566 10782 25195 10784
rect 5165 10706 5231 10709
rect 7741 10706 7807 10709
rect 5165 10704 7807 10706
rect 5165 10648 5170 10704
rect 5226 10648 7746 10704
rect 7802 10648 7807 10704
rect 5165 10646 7807 10648
rect 5165 10643 5231 10646
rect 7741 10643 7807 10646
rect 11973 10706 12039 10709
rect 19566 10706 19626 10782
rect 21817 10779 21883 10782
rect 25129 10779 25195 10782
rect 11973 10704 19626 10706
rect 11973 10648 11978 10704
rect 12034 10648 19626 10704
rect 11973 10646 19626 10648
rect 20345 10706 20411 10709
rect 24945 10706 25011 10709
rect 20345 10704 25011 10706
rect 20345 10648 20350 10704
rect 20406 10648 24950 10704
rect 25006 10648 25011 10704
rect 20345 10646 25011 10648
rect 11973 10643 12039 10646
rect 20345 10643 20411 10646
rect 24945 10643 25011 10646
rect 25630 10644 25636 10708
rect 25700 10706 25706 10708
rect 26509 10706 26575 10709
rect 25700 10704 26575 10706
rect 25700 10648 26514 10704
rect 26570 10648 26575 10704
rect 25700 10646 26575 10648
rect 25700 10644 25706 10646
rect 26509 10643 26575 10646
rect 2497 10570 2563 10573
rect 2630 10570 2636 10572
rect 2497 10568 2636 10570
rect 2497 10512 2502 10568
rect 2558 10512 2636 10568
rect 2497 10510 2636 10512
rect 2497 10507 2563 10510
rect 2630 10508 2636 10510
rect 2700 10508 2706 10572
rect 10317 10570 10383 10573
rect 25589 10570 25655 10573
rect 10317 10568 25655 10570
rect 10317 10512 10322 10568
rect 10378 10512 25594 10568
rect 25650 10512 25655 10568
rect 10317 10510 25655 10512
rect 10317 10507 10383 10510
rect 25589 10507 25655 10510
rect 0 10434 480 10464
rect 2129 10434 2195 10437
rect 0 10432 2195 10434
rect 0 10376 2134 10432
rect 2190 10376 2195 10432
rect 0 10374 2195 10376
rect 0 10344 480 10374
rect 2129 10371 2195 10374
rect 27705 10434 27771 10437
rect 29520 10434 30000 10464
rect 27705 10432 30000 10434
rect 27705 10376 27710 10432
rect 27766 10376 30000 10432
rect 27705 10374 30000 10376
rect 27705 10371 27771 10374
rect 10944 10368 11264 10369
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 29520 10344 30000 10374
rect 20944 10303 21264 10304
rect 5625 10298 5691 10301
rect 10317 10298 10383 10301
rect 5625 10296 10383 10298
rect 5625 10240 5630 10296
rect 5686 10240 10322 10296
rect 10378 10240 10383 10296
rect 5625 10238 10383 10240
rect 5625 10235 5691 10238
rect 10317 10235 10383 10238
rect 16849 10298 16915 10301
rect 19701 10298 19767 10301
rect 16849 10296 19767 10298
rect 16849 10240 16854 10296
rect 16910 10240 19706 10296
rect 19762 10240 19767 10296
rect 16849 10238 19767 10240
rect 16849 10235 16915 10238
rect 19701 10235 19767 10238
rect 5533 10162 5599 10165
rect 10777 10162 10843 10165
rect 25037 10162 25103 10165
rect 5533 10160 25103 10162
rect 5533 10104 5538 10160
rect 5594 10104 10782 10160
rect 10838 10104 25042 10160
rect 25098 10104 25103 10160
rect 5533 10102 25103 10104
rect 5533 10099 5599 10102
rect 10777 10099 10843 10102
rect 25037 10099 25103 10102
rect 5625 10026 5691 10029
rect 5758 10026 5764 10028
rect 5625 10024 5764 10026
rect 5625 9968 5630 10024
rect 5686 9968 5764 10024
rect 5625 9966 5764 9968
rect 5625 9963 5691 9966
rect 5758 9964 5764 9966
rect 5828 10026 5834 10028
rect 20713 10026 20779 10029
rect 26509 10028 26575 10029
rect 5828 10024 20779 10026
rect 5828 9968 20718 10024
rect 20774 9968 20779 10024
rect 5828 9966 20779 9968
rect 5828 9964 5834 9966
rect 20713 9963 20779 9966
rect 24902 9966 26434 10026
rect 0 9890 480 9920
rect 24902 9893 24962 9966
rect 1485 9890 1551 9893
rect 16941 9892 17007 9893
rect 16941 9890 16988 9892
rect 0 9888 1551 9890
rect 0 9832 1490 9888
rect 1546 9832 1551 9888
rect 0 9830 1551 9832
rect 16896 9888 16988 9890
rect 16896 9832 16946 9888
rect 16896 9830 16988 9832
rect 0 9800 480 9830
rect 1485 9827 1551 9830
rect 16941 9828 16988 9830
rect 17052 9828 17058 9892
rect 24853 9888 24962 9893
rect 24853 9832 24858 9888
rect 24914 9832 24962 9888
rect 24853 9830 24962 9832
rect 26374 9890 26434 9966
rect 26509 10024 26556 10028
rect 26620 10026 26626 10028
rect 26509 9968 26514 10024
rect 26509 9964 26556 9968
rect 26620 9966 26666 10026
rect 26620 9964 26626 9966
rect 26509 9963 26575 9964
rect 29520 9890 30000 9920
rect 26374 9830 30000 9890
rect 16941 9827 17007 9828
rect 24853 9827 24919 9830
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 29520 9800 30000 9830
rect 25944 9759 26264 9760
rect 5073 9754 5139 9757
rect 5809 9754 5875 9757
rect 5073 9752 5875 9754
rect 5073 9696 5078 9752
rect 5134 9696 5814 9752
rect 5870 9696 5875 9752
rect 5073 9694 5875 9696
rect 5073 9691 5139 9694
rect 5809 9691 5875 9694
rect 24669 9754 24735 9757
rect 25589 9754 25655 9757
rect 24669 9752 25655 9754
rect 24669 9696 24674 9752
rect 24730 9696 25594 9752
rect 25650 9696 25655 9752
rect 24669 9694 25655 9696
rect 24669 9691 24735 9694
rect 25589 9691 25655 9694
rect 1393 9618 1459 9621
rect 5625 9618 5691 9621
rect 1393 9616 5691 9618
rect 1393 9560 1398 9616
rect 1454 9560 5630 9616
rect 5686 9560 5691 9616
rect 1393 9558 5691 9560
rect 1393 9555 1459 9558
rect 5625 9555 5691 9558
rect 7005 9618 7071 9621
rect 15561 9618 15627 9621
rect 7005 9616 15627 9618
rect 7005 9560 7010 9616
rect 7066 9560 15566 9616
rect 15622 9560 15627 9616
rect 7005 9558 15627 9560
rect 7005 9555 7071 9558
rect 15561 9555 15627 9558
rect 18689 9618 18755 9621
rect 27521 9618 27587 9621
rect 18689 9616 27587 9618
rect 18689 9560 18694 9616
rect 18750 9560 27526 9616
rect 27582 9560 27587 9616
rect 18689 9558 27587 9560
rect 18689 9555 18755 9558
rect 27521 9555 27587 9558
rect 2589 9482 2655 9485
rect 2957 9482 3023 9485
rect 2589 9480 3023 9482
rect 2589 9424 2594 9480
rect 2650 9424 2962 9480
rect 3018 9424 3023 9480
rect 2589 9422 3023 9424
rect 2589 9419 2655 9422
rect 2957 9419 3023 9422
rect 3141 9482 3207 9485
rect 3325 9482 3391 9485
rect 3141 9480 3391 9482
rect 3141 9424 3146 9480
rect 3202 9424 3330 9480
rect 3386 9424 3391 9480
rect 3141 9422 3391 9424
rect 3141 9419 3207 9422
rect 3325 9419 3391 9422
rect 3601 9482 3667 9485
rect 4981 9482 5047 9485
rect 16297 9482 16363 9485
rect 16849 9482 16915 9485
rect 23105 9482 23171 9485
rect 23933 9482 23999 9485
rect 3601 9480 23999 9482
rect 3601 9424 3606 9480
rect 3662 9424 4986 9480
rect 5042 9424 16302 9480
rect 16358 9424 16854 9480
rect 16910 9424 23110 9480
rect 23166 9424 23938 9480
rect 23994 9424 23999 9480
rect 3601 9422 23999 9424
rect 3601 9419 3667 9422
rect 4981 9419 5047 9422
rect 16297 9419 16363 9422
rect 16849 9419 16915 9422
rect 23105 9419 23171 9422
rect 23933 9419 23999 9422
rect 0 9346 480 9376
rect 3693 9346 3759 9349
rect 0 9344 3759 9346
rect 0 9288 3698 9344
rect 3754 9288 3759 9344
rect 0 9286 3759 9288
rect 0 9256 480 9286
rect 3693 9283 3759 9286
rect 25589 9346 25655 9349
rect 29520 9346 30000 9376
rect 25589 9344 30000 9346
rect 25589 9288 25594 9344
rect 25650 9288 30000 9344
rect 25589 9286 30000 9288
rect 25589 9283 25655 9286
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 29520 9256 30000 9286
rect 20944 9215 21264 9216
rect 16297 9210 16363 9213
rect 19149 9210 19215 9213
rect 16297 9208 19215 9210
rect 16297 9152 16302 9208
rect 16358 9152 19154 9208
rect 19210 9152 19215 9208
rect 16297 9150 19215 9152
rect 16297 9147 16363 9150
rect 19149 9147 19215 9150
rect 22001 9210 22067 9213
rect 26417 9210 26483 9213
rect 22001 9208 26483 9210
rect 22001 9152 22006 9208
rect 22062 9152 26422 9208
rect 26478 9152 26483 9208
rect 22001 9150 26483 9152
rect 22001 9147 22067 9150
rect 26417 9147 26483 9150
rect 13813 9074 13879 9077
rect 25313 9074 25379 9077
rect 13813 9072 25379 9074
rect 13813 9016 13818 9072
rect 13874 9016 25318 9072
rect 25374 9016 25379 9072
rect 13813 9014 25379 9016
rect 13813 9011 13879 9014
rect 25313 9011 25379 9014
rect 16849 8938 16915 8941
rect 21541 8938 21607 8941
rect 16849 8936 21607 8938
rect 16849 8880 16854 8936
rect 16910 8880 21546 8936
rect 21602 8880 21607 8936
rect 16849 8878 21607 8880
rect 16849 8875 16915 8878
rect 21541 8875 21607 8878
rect 9121 8802 9187 8805
rect 15653 8802 15719 8805
rect 9121 8800 15719 8802
rect 9121 8744 9126 8800
rect 9182 8744 15658 8800
rect 15714 8744 15719 8800
rect 9121 8742 15719 8744
rect 9121 8739 9187 8742
rect 15653 8739 15719 8742
rect 5944 8736 6264 8737
rect 0 8666 480 8696
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 2681 8666 2747 8669
rect 29520 8666 30000 8696
rect 0 8664 2747 8666
rect 0 8608 2686 8664
rect 2742 8608 2747 8664
rect 0 8606 2747 8608
rect 0 8576 480 8606
rect 2681 8603 2747 8606
rect 26374 8606 30000 8666
rect 25497 8530 25563 8533
rect 26374 8530 26434 8606
rect 29520 8576 30000 8606
rect 25497 8528 26434 8530
rect 25497 8472 25502 8528
rect 25558 8472 26434 8528
rect 25497 8470 26434 8472
rect 25497 8467 25563 8470
rect 5257 8394 5323 8397
rect 7373 8394 7439 8397
rect 5257 8392 7439 8394
rect 5257 8336 5262 8392
rect 5318 8336 7378 8392
rect 7434 8336 7439 8392
rect 5257 8334 7439 8336
rect 5257 8331 5323 8334
rect 7373 8331 7439 8334
rect 18873 8394 18939 8397
rect 19609 8394 19675 8397
rect 26509 8394 26575 8397
rect 18873 8392 26575 8394
rect 18873 8336 18878 8392
rect 18934 8336 19614 8392
rect 19670 8336 26514 8392
rect 26570 8336 26575 8392
rect 18873 8334 26575 8336
rect 18873 8331 18939 8334
rect 19609 8331 19675 8334
rect 26509 8331 26575 8334
rect 10944 8192 11264 8193
rect 0 8122 480 8152
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 8127 21264 8128
rect 3417 8122 3483 8125
rect 0 8120 3483 8122
rect 0 8064 3422 8120
rect 3478 8064 3483 8120
rect 0 8062 3483 8064
rect 0 8032 480 8062
rect 3417 8059 3483 8062
rect 25497 8122 25563 8125
rect 29520 8122 30000 8152
rect 25497 8120 30000 8122
rect 25497 8064 25502 8120
rect 25558 8064 30000 8120
rect 25497 8062 30000 8064
rect 25497 8059 25563 8062
rect 29520 8032 30000 8062
rect 1393 7986 1459 7989
rect 2037 7986 2103 7989
rect 11513 7986 11579 7989
rect 1393 7984 11579 7986
rect 1393 7928 1398 7984
rect 1454 7928 2042 7984
rect 2098 7928 11518 7984
rect 11574 7928 11579 7984
rect 1393 7926 11579 7928
rect 1393 7923 1459 7926
rect 2037 7923 2103 7926
rect 11513 7923 11579 7926
rect 24025 7986 24091 7989
rect 25313 7986 25379 7989
rect 24025 7984 25379 7986
rect 24025 7928 24030 7984
rect 24086 7928 25318 7984
rect 25374 7928 25379 7984
rect 24025 7926 25379 7928
rect 24025 7923 24091 7926
rect 25313 7923 25379 7926
rect 7557 7850 7623 7853
rect 19057 7850 19123 7853
rect 21357 7850 21423 7853
rect 22093 7850 22159 7853
rect 26785 7850 26851 7853
rect 7557 7848 19258 7850
rect 7557 7792 7562 7848
rect 7618 7792 19062 7848
rect 19118 7792 19258 7848
rect 7557 7790 19258 7792
rect 7557 7787 7623 7790
rect 19057 7787 19123 7790
rect 19198 7714 19258 7790
rect 21357 7848 26851 7850
rect 21357 7792 21362 7848
rect 21418 7792 22098 7848
rect 22154 7792 26790 7848
rect 26846 7792 26851 7848
rect 21357 7790 26851 7792
rect 21357 7787 21423 7790
rect 22093 7787 22159 7790
rect 26785 7787 26851 7790
rect 24853 7714 24919 7717
rect 19198 7712 24919 7714
rect 19198 7656 24858 7712
rect 24914 7656 24919 7712
rect 19198 7654 24919 7656
rect 24853 7651 24919 7654
rect 5944 7648 6264 7649
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 14365 7578 14431 7581
rect 6502 7576 14431 7578
rect 6502 7520 14370 7576
rect 14426 7520 14431 7576
rect 6502 7518 14431 7520
rect 0 7442 480 7472
rect 2681 7442 2747 7445
rect 0 7440 2747 7442
rect 0 7384 2686 7440
rect 2742 7384 2747 7440
rect 0 7382 2747 7384
rect 0 7352 480 7382
rect 2681 7379 2747 7382
rect 3141 7442 3207 7445
rect 6502 7442 6562 7518
rect 14365 7515 14431 7518
rect 3141 7440 6562 7442
rect 3141 7384 3146 7440
rect 3202 7384 6562 7440
rect 3141 7382 6562 7384
rect 7005 7442 7071 7445
rect 19977 7442 20043 7445
rect 25405 7442 25471 7445
rect 7005 7440 25471 7442
rect 7005 7384 7010 7440
rect 7066 7384 19982 7440
rect 20038 7384 25410 7440
rect 25466 7384 25471 7440
rect 7005 7382 25471 7384
rect 3141 7379 3207 7382
rect 7005 7379 7071 7382
rect 19977 7379 20043 7382
rect 25405 7379 25471 7382
rect 26601 7442 26667 7445
rect 29520 7442 30000 7472
rect 26601 7440 30000 7442
rect 26601 7384 26606 7440
rect 26662 7384 30000 7440
rect 26601 7382 30000 7384
rect 26601 7379 26667 7382
rect 29520 7352 30000 7382
rect 7373 7306 7439 7309
rect 7373 7304 11530 7306
rect 7373 7248 7378 7304
rect 7434 7248 11530 7304
rect 7373 7246 11530 7248
rect 7373 7243 7439 7246
rect 11470 7170 11530 7246
rect 19701 7170 19767 7173
rect 11470 7168 19767 7170
rect 11470 7112 19706 7168
rect 19762 7112 19767 7168
rect 11470 7110 19767 7112
rect 19701 7107 19767 7110
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 24853 7034 24919 7037
rect 26509 7034 26575 7037
rect 24853 7032 26575 7034
rect 24853 6976 24858 7032
rect 24914 6976 26514 7032
rect 26570 6976 26575 7032
rect 24853 6974 26575 6976
rect 24853 6971 24919 6974
rect 26509 6971 26575 6974
rect 27705 7034 27771 7037
rect 27705 7032 27906 7034
rect 27705 6976 27710 7032
rect 27766 6976 27906 7032
rect 27705 6974 27906 6976
rect 27705 6971 27771 6974
rect 0 6898 480 6928
rect 1577 6898 1643 6901
rect 0 6896 1643 6898
rect 0 6840 1582 6896
rect 1638 6840 1643 6896
rect 0 6838 1643 6840
rect 0 6808 480 6838
rect 1577 6835 1643 6838
rect 2405 6898 2471 6901
rect 6913 6898 6979 6901
rect 2405 6896 6979 6898
rect 2405 6840 2410 6896
rect 2466 6840 6918 6896
rect 6974 6840 6979 6896
rect 2405 6838 6979 6840
rect 27846 6898 27906 6974
rect 29520 6898 30000 6928
rect 27846 6838 30000 6898
rect 2405 6835 2471 6838
rect 6913 6835 6979 6838
rect 29520 6808 30000 6838
rect 3141 6762 3207 6765
rect 6269 6762 6335 6765
rect 3141 6760 6335 6762
rect 3141 6704 3146 6760
rect 3202 6704 6274 6760
rect 6330 6704 6335 6760
rect 3141 6702 6335 6704
rect 3141 6699 3207 6702
rect 6269 6699 6335 6702
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 0 6354 480 6384
rect 1577 6354 1643 6357
rect 0 6352 1643 6354
rect 0 6296 1582 6352
rect 1638 6296 1643 6352
rect 0 6294 1643 6296
rect 0 6264 480 6294
rect 1577 6291 1643 6294
rect 26693 6354 26759 6357
rect 29520 6354 30000 6384
rect 26693 6352 30000 6354
rect 26693 6296 26698 6352
rect 26754 6296 30000 6352
rect 26693 6294 30000 6296
rect 26693 6291 26759 6294
rect 29520 6264 30000 6294
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 0 5674 480 5704
rect 1393 5674 1459 5677
rect 0 5672 1459 5674
rect 0 5616 1398 5672
rect 1454 5616 1459 5672
rect 0 5614 1459 5616
rect 0 5584 480 5614
rect 1393 5611 1459 5614
rect 27797 5674 27863 5677
rect 29520 5674 30000 5704
rect 27797 5672 30000 5674
rect 27797 5616 27802 5672
rect 27858 5616 30000 5672
rect 27797 5614 30000 5616
rect 27797 5611 27863 5614
rect 29520 5584 30000 5614
rect 26601 5538 26667 5541
rect 26969 5538 27035 5541
rect 26601 5536 27035 5538
rect 26601 5480 26606 5536
rect 26662 5480 26974 5536
rect 27030 5480 27035 5536
rect 26601 5478 27035 5480
rect 26601 5475 26667 5478
rect 26969 5475 27035 5478
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 0 5130 480 5160
rect 3509 5130 3575 5133
rect 0 5128 3575 5130
rect 0 5072 3514 5128
rect 3570 5072 3575 5128
rect 0 5070 3575 5072
rect 0 5040 480 5070
rect 3509 5067 3575 5070
rect 13353 5130 13419 5133
rect 26417 5130 26483 5133
rect 13353 5128 26483 5130
rect 13353 5072 13358 5128
rect 13414 5072 26422 5128
rect 26478 5072 26483 5128
rect 13353 5070 26483 5072
rect 13353 5067 13419 5070
rect 26417 5067 26483 5070
rect 26601 5130 26667 5133
rect 29520 5130 30000 5160
rect 26601 5128 30000 5130
rect 26601 5072 26606 5128
rect 26662 5072 30000 5128
rect 26601 5070 30000 5072
rect 26601 5067 26667 5070
rect 29520 5040 30000 5070
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 25865 4586 25931 4589
rect 25865 4584 26434 4586
rect 25865 4528 25870 4584
rect 25926 4528 26434 4584
rect 25865 4526 26434 4528
rect 25865 4523 25931 4526
rect 0 4450 480 4480
rect 1669 4450 1735 4453
rect 0 4448 1735 4450
rect 0 4392 1674 4448
rect 1730 4392 1735 4448
rect 0 4390 1735 4392
rect 26374 4450 26434 4526
rect 29520 4450 30000 4480
rect 26374 4390 30000 4450
rect 0 4360 480 4390
rect 1669 4387 1735 4390
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 29520 4360 30000 4390
rect 25944 4319 26264 4320
rect 2037 4042 2103 4045
rect 6913 4042 6979 4045
rect 2037 4040 6979 4042
rect 2037 3984 2042 4040
rect 2098 3984 6918 4040
rect 6974 3984 6979 4040
rect 2037 3982 6979 3984
rect 2037 3979 2103 3982
rect 6913 3979 6979 3982
rect 19701 4042 19767 4045
rect 26417 4042 26483 4045
rect 19701 4040 26483 4042
rect 19701 3984 19706 4040
rect 19762 3984 26422 4040
rect 26478 3984 26483 4040
rect 19701 3982 26483 3984
rect 19701 3979 19767 3982
rect 26417 3979 26483 3982
rect 0 3906 480 3936
rect 4337 3906 4403 3909
rect 0 3904 4403 3906
rect 0 3848 4342 3904
rect 4398 3848 4403 3904
rect 0 3846 4403 3848
rect 0 3816 480 3846
rect 4337 3843 4403 3846
rect 25037 3906 25103 3909
rect 29520 3906 30000 3936
rect 25037 3904 30000 3906
rect 25037 3848 25042 3904
rect 25098 3848 30000 3904
rect 25037 3846 30000 3848
rect 25037 3843 25103 3846
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 29520 3816 30000 3846
rect 20944 3775 21264 3776
rect 3693 3498 3759 3501
rect 15469 3498 15535 3501
rect 3693 3496 15535 3498
rect 3693 3440 3698 3496
rect 3754 3440 15474 3496
rect 15530 3440 15535 3496
rect 3693 3438 15535 3440
rect 3693 3435 3759 3438
rect 15469 3435 15535 3438
rect 25681 3498 25747 3501
rect 25681 3496 26434 3498
rect 25681 3440 25686 3496
rect 25742 3440 26434 3496
rect 25681 3438 26434 3440
rect 25681 3435 25747 3438
rect 0 3362 480 3392
rect 3785 3362 3851 3365
rect 0 3360 3851 3362
rect 0 3304 3790 3360
rect 3846 3304 3851 3360
rect 0 3302 3851 3304
rect 26374 3362 26434 3438
rect 29520 3362 30000 3392
rect 26374 3302 30000 3362
rect 0 3272 480 3302
rect 3785 3299 3851 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 29520 3272 30000 3302
rect 25944 3231 26264 3232
rect 26601 2818 26667 2821
rect 26601 2816 26802 2818
rect 26601 2760 26606 2816
rect 26662 2760 26802 2816
rect 26601 2758 26802 2760
rect 26601 2755 26667 2758
rect 10944 2752 11264 2753
rect 0 2682 480 2712
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 1577 2682 1643 2685
rect 0 2680 1643 2682
rect 0 2624 1582 2680
rect 1638 2624 1643 2680
rect 0 2622 1643 2624
rect 26742 2682 26802 2758
rect 29520 2682 30000 2712
rect 26742 2622 30000 2682
rect 0 2592 480 2622
rect 1577 2619 1643 2622
rect 29520 2592 30000 2622
rect 8385 2546 8451 2549
rect 7054 2544 8451 2546
rect 7054 2488 8390 2544
rect 8446 2488 8451 2544
rect 7054 2486 8451 2488
rect 7054 2410 7114 2486
rect 8385 2483 8451 2486
rect 3190 2350 7114 2410
rect 7189 2410 7255 2413
rect 11145 2410 11211 2413
rect 7189 2408 11211 2410
rect 7189 2352 7194 2408
rect 7250 2352 11150 2408
rect 11206 2352 11211 2408
rect 7189 2350 11211 2352
rect 0 2138 480 2168
rect 3190 2138 3250 2350
rect 7189 2347 7255 2350
rect 11145 2347 11211 2350
rect 5944 2208 6264 2209
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 0 2078 3250 2138
rect 26969 2138 27035 2141
rect 29520 2138 30000 2168
rect 26969 2136 30000 2138
rect 26969 2080 26974 2136
rect 27030 2080 30000 2136
rect 26969 2078 30000 2080
rect 0 2048 480 2078
rect 26969 2075 27035 2078
rect 29520 2048 30000 2078
rect 0 1458 480 1488
rect 1393 1458 1459 1461
rect 0 1456 1459 1458
rect 0 1400 1398 1456
rect 1454 1400 1459 1456
rect 0 1398 1459 1400
rect 0 1368 480 1398
rect 1393 1395 1459 1398
rect 26785 1458 26851 1461
rect 29520 1458 30000 1488
rect 26785 1456 30000 1458
rect 26785 1400 26790 1456
rect 26846 1400 30000 1456
rect 26785 1398 30000 1400
rect 26785 1395 26851 1398
rect 29520 1368 30000 1398
rect 0 914 480 944
rect 9029 914 9095 917
rect 0 912 9095 914
rect 0 856 9034 912
rect 9090 856 9095 912
rect 0 854 9095 856
rect 0 824 480 854
rect 9029 851 9095 854
rect 27061 914 27127 917
rect 29520 914 30000 944
rect 27061 912 30000 914
rect 27061 856 27066 912
rect 27122 856 30000 912
rect 27061 854 30000 856
rect 27061 851 27127 854
rect 29520 824 30000 854
rect 0 370 480 400
rect 2681 370 2747 373
rect 0 368 2747 370
rect 0 312 2686 368
rect 2742 312 2747 368
rect 0 310 2747 312
rect 0 280 480 310
rect 2681 307 2747 310
rect 26877 370 26943 373
rect 29520 370 30000 400
rect 26877 368 30000 370
rect 26877 312 26882 368
rect 26938 312 30000 368
rect 26877 310 30000 312
rect 26877 307 26943 310
rect 29520 280 30000 310
<< via3 >>
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 25268 20300 25332 20364
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 3924 19484 3988 19548
rect 24900 19076 24964 19140
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 25636 18260 25700 18324
rect 5764 18184 5828 18188
rect 5764 18128 5778 18184
rect 5778 18128 5828 18184
rect 5764 18124 5828 18128
rect 12940 18048 13004 18052
rect 12940 17992 12990 18048
rect 12990 17992 13004 18048
rect 12940 17988 13004 17992
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 14412 14648 14476 14652
rect 14412 14592 14462 14648
rect 14462 14592 14476 14648
rect 14412 14588 14476 14592
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 9628 13228 9692 13292
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 9628 12820 9692 12884
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 26740 11928 26804 11932
rect 26740 11872 26790 11928
rect 26790 11872 26804 11928
rect 26740 11868 26804 11872
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 8524 11188 8588 11252
rect 16436 11248 16500 11252
rect 16436 11192 16486 11248
rect 16486 11192 16500 11248
rect 16436 11188 16500 11192
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 25636 10644 25700 10708
rect 2636 10508 2700 10572
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5764 9964 5828 10028
rect 16988 9888 17052 9892
rect 16988 9832 17002 9888
rect 17002 9832 17052 9888
rect 16988 9828 17052 9832
rect 26556 10024 26620 10028
rect 26556 9968 26570 10024
rect 26570 9968 26620 10024
rect 26556 9964 26620 9968
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 21792 6264 21808
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 3923 19548 3989 19549
rect 3923 19484 3924 19548
rect 3988 19484 3989 19548
rect 3923 19483 3989 19484
rect 3926 14738 3986 19483
rect 5944 18528 6264 19552
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5763 18188 5829 18189
rect 5763 18124 5764 18188
rect 5828 18124 5829 18188
rect 5763 18123 5829 18124
rect 5766 10029 5826 18123
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15264 6264 16288
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 10944 21248 11264 21808
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 19072 11264 20096
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 17984 11264 19008
rect 15944 21792 16264 21808
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 12939 18052 13005 18053
rect 12939 17988 12940 18052
rect 13004 17988 13005 18052
rect 12939 17987 13005 17988
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 9627 13292 9693 13293
rect 9627 13228 9628 13292
rect 9692 13228 9693 13292
rect 9627 13227 9693 13228
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 9630 12885 9690 13227
rect 9627 12884 9693 12885
rect 9627 12820 9628 12884
rect 9692 12820 9693 12884
rect 9627 12819 9693 12820
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 12942 12018 13002 17987
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15264 16264 16288
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5763 10028 5829 10029
rect 5763 9964 5764 10028
rect 5828 9964 5829 10028
rect 5763 9963 5829 9964
rect 5944 9824 6264 10848
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 10912 16264 11936
rect 20944 21248 21264 21808
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 25944 21792 26264 21808
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25267 20364 25333 20365
rect 25267 20300 25268 20364
rect 25332 20300 25333 20364
rect 25267 20299 25333 20300
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 24899 19140 24965 19141
rect 24899 19076 24900 19140
rect 24964 19076 24965 19140
rect 24899 19075 24965 19076
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 20944 10368 21264 11392
rect 24902 10658 24962 19075
rect 25270 11338 25330 20299
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25635 18324 25701 18325
rect 25635 18260 25636 18324
rect 25700 18260 25701 18324
rect 25635 18259 25701 18260
rect 25638 10709 25698 18259
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15264 26264 16288
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25635 10708 25701 10709
rect 25635 10644 25636 10708
rect 25700 10644 25701 10708
rect 25635 10643 25701 10644
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 25944 9824 26264 10848
rect 26555 10028 26621 10029
rect 26555 9978 26556 10028
rect 26620 9978 26621 10028
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 3838 14502 4074 14738
rect 2550 10572 2786 10658
rect 2550 10508 2636 10572
rect 2636 10508 2700 10572
rect 2700 10508 2786 10572
rect 2550 10422 2786 10508
rect 14326 14652 14562 14738
rect 14326 14588 14412 14652
rect 14412 14588 14476 14652
rect 14476 14588 14562 14652
rect 14326 14502 14562 14588
rect 12854 11782 13090 12018
rect 8438 11252 8674 11338
rect 8438 11188 8524 11252
rect 8524 11188 8588 11252
rect 8588 11188 8674 11252
rect 8438 11102 8674 11188
rect 16350 11252 16586 11338
rect 16350 11188 16436 11252
rect 16436 11188 16500 11252
rect 16500 11188 16586 11252
rect 16350 11102 16586 11188
rect 25182 11102 25418 11338
rect 26654 11932 26890 12018
rect 26654 11868 26740 11932
rect 26740 11868 26804 11932
rect 26804 11868 26890 11932
rect 26654 11782 26890 11868
rect 24814 10422 25050 10658
rect 16902 9892 17138 9978
rect 16902 9828 16988 9892
rect 16988 9828 17052 9892
rect 17052 9828 17138 9892
rect 16902 9742 17138 9828
rect 26470 9964 26556 9978
rect 26556 9964 26620 9978
rect 26620 9964 26706 9978
rect 26470 9742 26706 9964
<< metal5 >>
rect 3796 14738 14604 14780
rect 3796 14502 3838 14738
rect 4074 14502 14326 14738
rect 14562 14502 14604 14738
rect 3796 14460 14604 14502
rect 12812 12018 26932 12060
rect 12812 11782 12854 12018
rect 13090 11782 26654 12018
rect 26890 11782 26932 12018
rect 12812 11740 26932 11782
rect 8396 11338 25460 11380
rect 8396 11102 8438 11338
rect 8674 11102 16350 11338
rect 16586 11102 25182 11338
rect 25418 11102 25460 11338
rect 8396 11060 25460 11102
rect 2508 10658 25092 10700
rect 2508 10422 2550 10658
rect 2786 10422 24814 10658
rect 25050 10422 25092 10658
rect 2508 10380 25092 10422
rect 16860 9978 26748 10020
rect 16860 9742 16902 9978
rect 17138 9742 26470 9978
rect 26706 9742 26748 9978
rect 16860 9700 26748 9742
use sky130_fd_sc_hd__buf_2  _49_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1604666999
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1932 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1604666999
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 1748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_11
timestamp 1604666999
transform 1 0 2116 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1604666999
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_23
timestamp 1604666999
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_35
timestamp 1604666999
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1604666999
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 1604666999
transform 1 0 6440 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_47
timestamp 1604666999
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59
timestamp 1604666999
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 6900 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1604666999
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1604666999
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6624 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1604666999
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1604666999
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1604666999
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_82 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 8648 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_90
timestamp 1604666999
transform 1 0 9384 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1604666999
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1604666999
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1604666999
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1604666999
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_110
timestamp 1604666999
transform 1 0 11224 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1604666999
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1604666999
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1604666999
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1604666999
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1604666999
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1604666999
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1604666999
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1604666999
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1604666999
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1604666999
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1604666999
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1604666999
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1604666999
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1604666999
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1604666999
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1604666999
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1604666999
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1604666999
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1604666999
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1604666999
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1604666999
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1604666999
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1604666999
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1604666999
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1604666999
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1604666999
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1604666999
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1604666999
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1604666999
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1604666999
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1604666999
transform 1 0 24012 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1604666999
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1604666999
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1604666999
transform 1 0 26404 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1604666999
transform 1 0 25116 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1604666999
transform 1 0 26220 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_269
timestamp 1604666999
transform 1 0 25852 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1604666999
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1604666999
transform 1 0 26956 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1604666999
transform 1 0 26864 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292
timestamp 1604666999
transform 1 0 27968 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_279
timestamp 1604666999
transform 1 0 26772 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_283
timestamp 1604666999
transform 1 0 27140 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_295
timestamp 1604666999
transform 1 0 28244 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1604666999
transform -1 0 28888 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1604666999
transform -1 0 28888 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298 tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 28520 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1604666999
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1604666999
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1604666999
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1604666999
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1604666999
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1604666999
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1604666999
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1604666999
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1604666999
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1604666999
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1604666999
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1604666999
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1604666999
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1604666999
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1604666999
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1604666999
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1604666999
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1604666999
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1604666999
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1604666999
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1604666999
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1604666999
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1604666999
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1604666999
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1604666999
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1604666999
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1604666999
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1604666999
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1604666999
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1604666999
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_288
timestamp 1604666999
transform 1 0 27600 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp 1604666999
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1604666999
transform -1 0 28888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1604666999
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1604666999
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1604666999
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1604666999
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1604666999
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1604666999
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1604666999
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1604666999
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1604666999
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1604666999
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1604666999
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1604666999
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1604666999
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1604666999
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1604666999
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1604666999
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1604666999
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1604666999
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1604666999
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1604666999
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1604666999
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1604666999
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1604666999
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1604666999
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1604666999
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1604666999
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1604666999
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1604666999
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1604666999
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1604666999
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1604666999
transform 1 0 28060 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1604666999
transform -1 0 28888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1604666999
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1604666999
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1604666999
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1604666999
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1604666999
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1604666999
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1604666999
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1604666999
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1604666999
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1604666999
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1604666999
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1604666999
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1604666999
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1604666999
transform 1 0 11868 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1604666999
transform 1 0 12972 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1604666999
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1604666999
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1604666999
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1604666999
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1604666999
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1604666999
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1604666999
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1604666999
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1604666999
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1604666999
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1604666999
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1604666999
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1604666999
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1604666999
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1604666999
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_288
timestamp 1604666999
transform 1 0 27600 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_296
timestamp 1604666999
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1604666999
transform -1 0 28888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1604666999
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1604666999
transform 1 0 1564 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_3
timestamp 1604666999
transform 1 0 1380 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_7
timestamp 1604666999
transform 1 0 1748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_19
timestamp 1604666999
transform 1 0 2852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_31
timestamp 1604666999
transform 1 0 3956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_43
timestamp 1604666999
transform 1 0 5060 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_55
timestamp 1604666999
transform 1 0 6164 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1604666999
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1604666999
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1604666999
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1604666999
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1604666999
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1604666999
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1604666999
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1604666999
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1604666999
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1604666999
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1604666999
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1604666999
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1604666999
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1604666999
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1604666999
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1604666999
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1604666999
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1604666999
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1604666999
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1604666999
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1604666999
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1604666999
transform 1 0 26404 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_269
timestamp 1604666999
transform 1 0 25852 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1604666999
transform 1 0 26956 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_279
timestamp 1604666999
transform 1 0 26772 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_283
timestamp 1604666999
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_295
timestamp 1604666999
transform 1 0 28244 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1604666999
transform -1 0 28888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1604666999
transform 1 0 1748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_7
timestamp 1604666999
transform 1 0 1748 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1604666999
transform 1 0 1932 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1604666999
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1604666999
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1604666999
transform 1 0 1380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1604666999
transform 1 0 1380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp 1604666999
transform 1 0 2852 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1604666999
transform 1 0 2116 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1604666999
transform 1 0 2484 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1604666999
transform 1 0 2300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1604666999
transform 1 0 2484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_17
timestamp 1604666999
transform 1 0 2668 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1604666999
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1604666999
transform 1 0 3036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp 1604666999
transform 1 0 3772 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1604666999
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_23
timestamp 1604666999
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_35
timestamp 1604666999
transform 1 0 4324 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1604666999
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1604666999
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_43
timestamp 1604666999
transform 1 0 5060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_46
timestamp 1604666999
transform 1 0 5336 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1604666999
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1604666999
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1604666999
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1604666999
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1604666999
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1604666999
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1604666999
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1604666999
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1604666999
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1604666999
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1604666999
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1604666999
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1604666999
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1604666999
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1604666999
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1604666999
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1604666999
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1604666999
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1604666999
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1604666999
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_147
timestamp 1604666999
transform 1 0 14628 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_153
timestamp 1604666999
transform 1 0 15180 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_156
timestamp 1604666999
transform 1 0 15456 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1604666999
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1604666999
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_168
timestamp 1604666999
transform 1 0 16560 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1604666999
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1604666999
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_180
timestamp 1604666999
transform 1 0 17664 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1604666999
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1604666999
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1604666999
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1604666999
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1604666999
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1604666999
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1604666999
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1604666999
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1604666999
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1604666999
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1604666999
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1604666999
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1604666999
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1604666999
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1604666999
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1604666999
transform 1 0 26496 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1604666999
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1604666999
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_269
timestamp 1604666999
transform 1 0 25852 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_275
timestamp 1604666999
transform 1 0 26404 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_288
timestamp 1604666999
transform 1 0 27600 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_296
timestamp 1604666999
transform 1 0 28336 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_278
timestamp 1604666999
transform 1 0 26680 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_290
timestamp 1604666999
transform 1 0 27784 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1604666999
transform -1 0 28888 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1604666999
transform -1 0 28888 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_298
timestamp 1604666999
transform 1 0 28520 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1604666999
transform 1 0 2484 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1604666999
transform 1 0 1380 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1604666999
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1604666999
transform 1 0 1932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2300 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1604666999
transform 1 0 1748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1604666999
transform 1 0 2116 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_19
timestamp 1604666999
transform 1 0 2852 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1604666999
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 4600 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1604666999
transform 1 0 4048 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5152 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 5520 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_40
timestamp 1604666999
transform 1 0 4784 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1604666999
transform 1 0 5336 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_50
timestamp 1604666999
transform 1 0 5704 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_54
timestamp 1604666999
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_57
timestamp 1604666999
transform 1 0 6348 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6808 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_61
timestamp 1604666999
transform 1 0 6716 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_64
timestamp 1604666999
transform 1 0 6992 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1604666999
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1604666999
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1604666999
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1604666999
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1604666999
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1604666999
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1604666999
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 15272 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1604666999
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1604666999
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_157
timestamp 1604666999
transform 1 0 15548 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16652 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_171
timestamp 1604666999
transform 1 0 16836 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19136 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 18768 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 18400 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_183
timestamp 1604666999
transform 1 0 17940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_186
timestamp 1604666999
transform 1 0 18216 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1604666999
transform 1 0 18584 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1604666999
transform 1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_198
timestamp 1604666999
transform 1 0 19320 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1604666999
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 19964 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1604666999
transform 1 0 19780 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_207
timestamp 1604666999
transform 1 0 20148 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1604666999
transform 1 0 20700 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1604666999
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1604666999
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1604666999
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1604666999
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1604666999
transform 1 0 26496 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1604666999
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1604666999
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_280
timestamp 1604666999
transform 1 0 26864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_292
timestamp 1604666999
transform 1 0 27968 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1604666999
transform -1 0 28888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_298
timestamp 1604666999
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1604666999
transform 1 0 2484 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1604666999
transform 1 0 1380 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1604666999
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1604666999
transform 1 0 1932 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1604666999
transform 1 0 2300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1604666999
transform 1 0 1748 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_11
timestamp 1604666999
transform 1 0 2116 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_19
timestamp 1604666999
transform 1 0 2852 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1604666999
transform 1 0 3588 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 4600 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1604666999
transform 1 0 3036 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1604666999
transform 1 0 4140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_23
timestamp 1604666999
transform 1 0 3220 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1604666999
transform 1 0 3956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_35
timestamp 1604666999
transform 1 0 4324 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 5152 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6164 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4968 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1604666999
transform 1 0 4784 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_53
timestamp 1604666999
transform 1 0 5980 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1604666999
transform 1 0 6348 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1604666999
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 7820 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 8188 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1604666999
transform 1 0 7636 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_75
timestamp 1604666999
transform 1 0 8004 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_79
timestamp 1604666999
transform 1 0 8372 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 8556 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_83
timestamp 1604666999
transform 1 0 8740 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_95
timestamp 1604666999
transform 1 0 9844 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_107
timestamp 1604666999
transform 1 0 10948 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_119
timestamp 1604666999
transform 1 0 12052 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1604666999
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1604666999
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1604666999
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_147
timestamp 1604666999
transform 1 0 14628 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_155
timestamp 1604666999
transform 1 0 15364 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_158
timestamp 1604666999
transform 1 0 15640 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 16192 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17388 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 15824 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_162
timestamp 1604666999
transform 1 0 16008 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_175
timestamp 1604666999
transform 1 0 17204 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1604666999
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 1604666999
transform 1 0 17572 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 1604666999
transform 1 0 18860 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_198
timestamp 1604666999
transform 1 0 19320 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1604666999
transform 1 0 19596 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 20884 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_210
timestamp 1604666999
transform 1 0 20424 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_214
timestamp 1604666999
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1604666999
transform 1 0 21068 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 21252 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 21620 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1604666999
transform 1 0 21436 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1604666999
transform 1 0 21804 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_237
timestamp 1604666999
transform 1 0 22908 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1604666999
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_243
timestamp 1604666999
transform 1 0 23460 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1604666999
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_257
timestamp 1604666999
transform 1 0 24748 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1604666999
transform 1 0 26404 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1604666999
transform 1 0 25300 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_265
timestamp 1604666999
transform 1 0 25484 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_273
timestamp 1604666999
transform 1 0 26220 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1604666999
transform 1 0 27508 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1604666999
transform 1 0 26956 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1604666999
transform 1 0 28060 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1604666999
transform 1 0 27324 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_279
timestamp 1604666999
transform 1 0 26772 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_283
timestamp 1604666999
transform 1 0 27140 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_291
timestamp 1604666999
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_295
timestamp 1604666999
transform 1 0 28244 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1604666999
transform -1 0 28888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1604666999
transform 1 0 2484 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1604666999
transform 1 0 1380 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1604666999
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 1932 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 2300 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_7
timestamp 1604666999
transform 1 0 1748 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 1604666999
transform 1 0 2116 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 1604666999
transform 1 0 2852 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 4600 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1604666999
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 4416 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 3036 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_23
timestamp 1604666999
transform 1 0 3220 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1604666999
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_32
timestamp 1604666999
transform 1 0 4048 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6164 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5980 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 5612 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_47
timestamp 1604666999
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_51
timestamp 1604666999
transform 1 0 5796 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 7728 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1604666999
transform 1 0 6992 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1604666999
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1604666999
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_81
timestamp 1604666999
transform 1 0 8556 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_89
timestamp 1604666999
transform 1 0 9292 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1604666999
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1604666999
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1604666999
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1604666999
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1604666999
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1604666999
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_154
timestamp 1604666999
transform 1 0 15272 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16652 0 -1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 16284 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_162
timestamp 1604666999
transform 1 0 16008 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_167
timestamp 1604666999
transform 1 0 16468 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 19136 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18676 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_188
timestamp 1604666999
transform 1 0 18400 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1604666999
transform 1 0 18860 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1604666999
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20148 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1604666999
transform 1 0 19964 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_209
timestamp 1604666999
transform 1 0 20332 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_213
timestamp 1604666999
transform 1 0 20700 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_224
timestamp 1604666999
transform 1 0 21712 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_236
timestamp 1604666999
transform 1 0 22816 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_248
timestamp 1604666999
transform 1 0 23920 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1604666999
transform 1 0 25300 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1604666999
transform 1 0 26496 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1604666999
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_260
timestamp 1604666999
transform 1 0 25024 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_267
timestamp 1604666999
transform 1 0 25668 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_280
timestamp 1604666999
transform 1 0 26864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_292
timestamp 1604666999
transform 1 0 27968 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1604666999
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_298
timestamp 1604666999
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l4_in_0_
timestamp 1604666999
transform 1 0 1932 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1604666999
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 1748 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1604666999
transform 1 0 1380 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_18
timestamp 1604666999
transform 1 0 2760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1604666999
transform 1 0 3496 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1604666999
transform 1 0 4048 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4600 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 2944 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 3312 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_22
timestamp 1604666999
transform 1 0 3128 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_30
timestamp 1604666999
transform 1 0 3864 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_34
timestamp 1604666999
transform 1 0 4232 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1604666999
transform 1 0 4784 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6164 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 5796 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_49
timestamp 1604666999
transform 1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_53
timestamp 1604666999
transform 1 0 5980 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1604666999
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1604666999
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 8740 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1604666999
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1604666999
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_89
timestamp 1604666999
transform 1 0 9292 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_101
timestamp 1604666999
transform 1 0 10396 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1604666999
transform 1 0 11500 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1604666999
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1604666999
transform 1 0 12236 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1604666999
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1604666999
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 15364 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_147
timestamp 1604666999
transform 1 0 14628 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1604666999
transform 1 0 15548 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 16284 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16100 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 15732 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 17296 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1604666999
transform 1 0 15916 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_174
timestamp 1604666999
transform 1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_178
timestamp 1604666999
transform 1 0 17480 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18676 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1604666999
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 18492 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1604666999
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_188
timestamp 1604666999
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20056 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_200
timestamp 1604666999
transform 1 0 19504 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_204
timestamp 1604666999
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_208
timestamp 1604666999
transform 1 0 20240 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_212
timestamp 1604666999
transform 1 0 20608 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_224
timestamp 1604666999
transform 1 0 21712 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_236
timestamp 1604666999
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1604666999
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1604666999
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_257
timestamp 1604666999
transform 1 0 24748 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1604666999
transform 1 0 25300 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1604666999
transform 1 0 26404 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1604666999
transform 1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1604666999
transform 1 0 25116 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_267
timestamp 1604666999
transform 1 0 25668 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_271
timestamp 1604666999
transform 1 0 26036 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1604666999
transform 1 0 27508 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1604666999
transform 1 0 26956 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1604666999
transform 1 0 28060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1604666999
transform 1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_279
timestamp 1604666999
transform 1 0 26772 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_283
timestamp 1604666999
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_291
timestamp 1604666999
transform 1 0 27876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_295
timestamp 1604666999
transform 1 0 28244 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1604666999
transform -1 0 28888 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l3_in_1_
timestamp 1604666999
transform 1 0 1840 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1604666999
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1604666999
transform 1 0 1564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 2852 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1604666999
transform 1 0 1380 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1604666999
transform 1 0 1748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_17
timestamp 1604666999
transform 1 0 2668 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_21
timestamp 1604666999
transform 1 0 3036 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 3220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_25
timestamp 1604666999
transform 1 0 3404 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1604666999
transform 1 0 3772 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1604666999
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1604666999
transform 1 0 4048 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 4232 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_36
timestamp 1604666999
transform 1 0 4416 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 4692 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4876 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1604666999
transform 1 0 7360 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 6808 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7176 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1604666999
transform 1 0 6624 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1604666999
transform 1 0 6992 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_77
timestamp 1604666999
transform 1 0 8188 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1604666999
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_89
timestamp 1604666999
transform 1 0 9292 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1604666999
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1604666999
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1604666999
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1604666999
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _20_ tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1604666999
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1604666999
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1604666999
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_157
timestamp 1604666999
transform 1 0 15548 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 16284 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 16100 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 19044 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18676 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_184
timestamp 1604666999
transform 1 0 18032 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_190
timestamp 1604666999
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_193
timestamp 1604666999
transform 1 0 18860 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1604666999
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_206
timestamp 1604666999
transform 1 0 20056 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1604666999
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1604666999
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24564 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1604666999
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_251
timestamp 1604666999
transform 1 0 24196 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_257
timestamp 1604666999
transform 1 0 24748 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1604666999
transform 1 0 25300 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1604666999
transform 1 0 26496 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1604666999
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_267
timestamp 1604666999
transform 1 0 25668 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_280
timestamp 1604666999
transform 1 0 26864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_292
timestamp 1604666999
transform 1 0 27968 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1604666999
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_298
timestamp 1604666999
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1604666999
transform 1 0 1748 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1604666999
transform 1 0 1380 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_7
timestamp 1604666999
transform 1 0 1748 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 1840 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1604666999
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1604666999
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1604666999
transform 1 0 1380 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_19
timestamp 1604666999
transform 1 0 2852 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 1604666999
transform 1 0 2208 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 2392 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 2024 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l3_in_0_
timestamp 1604666999
transform 1 0 2576 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_3_
timestamp 1604666999
transform 1 0 2024 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 1604666999
transform 1 0 3772 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1604666999
transform 1 0 3220 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1604666999
transform 1 0 3772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_25
timestamp 1604666999
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3036 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3588 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 3956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1604666999
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4140 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4048 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_13_46
timestamp 1604666999
transform 1 0 5336 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_42
timestamp 1604666999
transform 1 0 4968 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 5520 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 5152 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1604666999
transform 1 0 5704 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 5980 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_53
timestamp 1604666999
transform 1 0 5980 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_51
timestamp 1604666999
transform 1 0 5796 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 6348 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1604666999
transform 1 0 6348 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_55
timestamp 1604666999
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_0_
timestamp 1604666999
transform 1 0 6532 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_68
timestamp 1604666999
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1604666999
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 6808 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1604666999
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_75
timestamp 1604666999
transform 1 0 8004 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_71
timestamp 1604666999
transform 1 0 7636 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 7912 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1604666999
transform 1 0 8096 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1604666999
transform 1 0 8096 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_78
timestamp 1604666999
transform 1 0 8280 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1604666999
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 8648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_90
timestamp 1604666999
transform 1 0 9384 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_80
timestamp 1604666999
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1604666999
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_88
timestamp 1604666999
transform 1 0 9200 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_93
timestamp 1604666999
transform 1 0 9660 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1604666999
transform 1 0 10212 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11040 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_102
timestamp 1604666999
transform 1 0 10488 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_114
timestamp 1604666999
transform 1 0 11592 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1604666999
transform 1 0 10488 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_106
timestamp 1604666999
transform 1 0 10856 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_110
timestamp 1604666999
transform 1 0 11224 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1604666999
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1604666999
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1604666999
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_122
timestamp 1604666999
transform 1 0 12328 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_134
timestamp 1604666999
transform 1 0 13432 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1604666999
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_147
timestamp 1604666999
transform 1 0 14628 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_155
timestamp 1604666999
transform 1 0 15364 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 1604666999
transform 1 0 15640 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_14_146
timestamp 1604666999
transform 1 0 14536 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1604666999
transform 1 0 15088 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1604666999
transform 1 0 15272 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_158
timestamp 1604666999
transform 1 0 15640 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_165
timestamp 1604666999
transform 1 0 16284 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1604666999
transform 1 0 15916 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1604666999
transform 1 0 16008 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 15732 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 16100 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1604666999
transform 1 0 16376 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1604666999
transform 1 0 16468 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_14_176
timestamp 1604666999
transform 1 0 17296 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_175
timestamp 1604666999
transform 1 0 17204 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 17388 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_182
timestamp 1604666999
transform 1 0 17848 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_188
timestamp 1604666999
transform 1 0 18400 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_184
timestamp 1604666999
transform 1 0 18032 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1604666999
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1604666999
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_193
timestamp 1604666999
transform 1 0 18860 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_190
timestamp 1604666999
transform 1 0 18584 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_191
timestamp 1604666999
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 19044 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_1_
timestamp 1604666999
transform 1 0 19228 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 19044 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_3_
timestamp 1604666999
transform 1 0 20884 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1604666999
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 20976 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 20240 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_214
timestamp 1604666999
transform 1 0 20792 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_218
timestamp 1604666999
transform 1 0 21160 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_206
timestamp 1604666999
transform 1 0 20056 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_210
timestamp 1604666999
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_228
timestamp 1604666999
transform 1 0 22080 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 1604666999
transform 1 0 21712 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1604666999
transform 1 0 21528 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 21712 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 21344 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 21896 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_236
timestamp 1604666999
transform 1 0 22816 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_238
timestamp 1604666999
transform 1 0 23000 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 23000 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_226
timestamp 1604666999
transform 1 0 21896 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_247
timestamp 1604666999
transform 1 0 23828 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_240
timestamp 1604666999
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_245
timestamp 1604666999
transform 1 0 23644 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 23368 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1604666999
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1604666999
transform 1 0 23552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_251
timestamp 1604666999
transform 1 0 24196 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_255
timestamp 1604666999
transform 1 0 24564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 24380 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 24012 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1604666999
transform 1 0 24012 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 24748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_1_
timestamp 1604666999
transform 1 0 24564 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1604666999
transform 1 0 24196 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_264
timestamp 1604666999
transform 1 0 25392 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_259
timestamp 1604666999
transform 1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 25116 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1604666999
transform 1 0 25300 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_274
timestamp 1604666999
transform 1 0 26312 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_271
timestamp 1604666999
transform 1 0 26036 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_267
timestamp 1604666999
transform 1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 26128 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1604666999
transform 1 0 26220 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1604666999
transform 1 0 25852 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1604666999
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1604666999
transform 1 0 26404 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1604666999
transform 1 0 26496 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_280
timestamp 1604666999
transform 1 0 26864 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_283
timestamp 1604666999
transform 1 0 27140 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_279
timestamp 1604666999
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 27048 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1604666999
transform 1 0 26956 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1604666999
transform 1 0 27508 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1604666999
transform 1 0 28336 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_295
timestamp 1604666999
transform 1 0 28244 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_291
timestamp 1604666999
transform 1 0 27876 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1604666999
transform 1 0 28060 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_284
timestamp 1604666999
transform 1 0 27232 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1604666999
transform -1 0 28888 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1604666999
transform -1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2024 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1604666999
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 1840 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1604666999
transform 1 0 1380 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_7
timestamp 1604666999
transform 1 0 1748 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_19
timestamp 1604666999
transform 1 0 2852 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 3036 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 4600 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_23
timestamp 1604666999
transform 1 0 3220 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_36
timestamp 1604666999
transform 1 0 4416 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_2_
timestamp 1604666999
transform 1 0 5152 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 4968 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 6164 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_40
timestamp 1604666999
transform 1 0 4784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_53
timestamp 1604666999
transform 1 0 5980 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1604666999
transform 1 0 6348 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7268 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1604666999
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7084 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_62
timestamp 1604666999
transform 1 0 6808 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_76
timestamp 1604666999
transform 1 0 8096 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1604666999
transform 1 0 8832 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 9752 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1604666999
transform 1 0 9384 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 8648 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_80
timestamp 1604666999
transform 1 0 8464 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1604666999
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_92
timestamp 1604666999
transform 1 0 9568 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_96
timestamp 1604666999
transform 1 0 9936 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_2_
timestamp 1604666999
transform 1 0 10304 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 11316 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_109
timestamp 1604666999
transform 1 0 11132 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1604666999
transform 1 0 11500 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_118
timestamp 1604666999
transform 1 0 11960 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1604666999
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 12144 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12604 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1604666999
transform 1 0 12420 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_127
timestamp 1604666999
transform 1 0 12788 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 15456 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1604666999
transform 1 0 13892 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_151
timestamp 1604666999
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_154
timestamp 1604666999
transform 1 0 15272 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1604666999
transform 1 0 15640 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1604666999
transform 1 0 16008 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_175
timestamp 1604666999
transform 1 0 17204 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1604666999
transform 1 0 17848 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_179
timestamp 1604666999
transform 1 0 17572 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 17664 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1604666999
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_188
timestamp 1604666999
transform 1 0 18400 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1604666999
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_192
timestamp 1604666999
transform 1 0 18768 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 18860 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_195
timestamp 1604666999
transform 1 0 19044 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 19228 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 19412 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_15_218
timestamp 1604666999
transform 1 0 21160 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_2_
timestamp 1604666999
transform 1 0 21896 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 21712 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1604666999
transform 1 0 22908 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 21344 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1604666999
transform 1 0 21528 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_235
timestamp 1604666999
transform 1 0 22724 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23644 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1604666999
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_239
timestamp 1604666999
transform 1 0 23092 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_2_
timestamp 1604666999
transform 1 0 26128 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 25944 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1604666999
transform 1 0 25576 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_264
timestamp 1604666999
transform 1 0 25392 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_268
timestamp 1604666999
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 27140 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 27508 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1604666999
transform 1 0 26956 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_285
timestamp 1604666999
transform 1 0 27324 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_289
timestamp 1604666999
transform 1 0 27692 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_297
timestamp 1604666999
transform 1 0 28428 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1604666999
transform -1 0 28888 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1604666999
transform 1 0 1380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_1_
timestamp 1604666999
transform 1 0 2392 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1604666999
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 2024 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1604666999
transform 1 0 1656 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_12
timestamp 1604666999
transform 1 0 2208 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1604666999
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 4232 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4600 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1604666999
transform 1 0 3220 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1604666999
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1604666999
transform 1 0 4048 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1604666999
transform 1 0 4416 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 4968 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_16_40
timestamp 1604666999
transform 1 0 4784 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l3_in_1_
timestamp 1604666999
transform 1 0 7452 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 6900 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7268 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_61
timestamp 1604666999
transform 1 0 6716 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_65
timestamp 1604666999
transform 1 0 7084 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1604666999
transform 1 0 8280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10212 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1604666999
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 10028 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8464 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1604666999
transform 1 0 8648 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1604666999
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_93
timestamp 1604666999
transform 1 0 9660 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_0_
timestamp 1604666999
transform 1 0 11776 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_16_108
timestamp 1604666999
transform 1 0 11040 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 13248 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_125
timestamp 1604666999
transform 1 0 12604 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_131
timestamp 1604666999
transform 1 0 13156 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_134
timestamp 1604666999
transform 1 0 13432 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1604666999
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 14812 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 15548 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_146
timestamp 1604666999
transform 1 0 14536 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1604666999
transform 1 0 14996 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1604666999
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_3_
timestamp 1604666999
transform 1 0 16100 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17112 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_159
timestamp 1604666999
transform 1 0 15732 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_172
timestamp 1604666999
transform 1 0 16928 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_176
timestamp 1604666999
transform 1 0 17296 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l2_in_0_
timestamp 1604666999
transform 1 0 17664 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19228 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18676 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 19044 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1604666999
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_193
timestamp 1604666999
transform 1 0 18860 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l3_in_1_
timestamp 1604666999
transform 1 0 20884 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1604666999
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20608 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_206
timestamp 1604666999
transform 1 0 20056 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1604666999
transform 1 0 22540 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 21896 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_224
timestamp 1604666999
transform 1 0 21712 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_228
timestamp 1604666999
transform 1 0 22080 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_232
timestamp 1604666999
transform 1 0 22448 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_237
timestamp 1604666999
transform 1 0 22908 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l3_in_1_
timestamp 1604666999
transform 1 0 23644 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 23368 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24748 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_241
timestamp 1604666999
transform 1 0 23276 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_244
timestamp 1604666999
transform 1 0 23552 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_254
timestamp 1604666999
transform 1 0 24472 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1604666999
transform 1 0 25300 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_3_
timestamp 1604666999
transform 1 0 26496 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1604666999
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 26128 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 25116 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_259
timestamp 1604666999
transform 1 0 24932 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_267
timestamp 1604666999
transform 1 0 25668 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_271
timestamp 1604666999
transform 1 0 26036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_274
timestamp 1604666999
transform 1 0 26312 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 27508 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_285
timestamp 1604666999
transform 1 0 27324 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_289
timestamp 1604666999
transform 1 0 27692 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_297
timestamp 1604666999
transform 1 0 28428 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1604666999
transform -1 0 28888 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 2300 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1604666999
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 2116 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 1564 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1604666999
transform 1 0 1380 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_7
timestamp 1604666999
transform 1 0 1748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 4600 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_32
timestamp 1604666999
transform 1 0 4048 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1604666999
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l3_in_0_
timestamp 1604666999
transform 1 0 5152 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_40
timestamp 1604666999
transform 1 0 4784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_53
timestamp 1604666999
transform 1 0 5980 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 1604666999
transform 1 0 6348 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1604666999
transform 1 0 6808 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_3_
timestamp 1604666999
transform 1 0 7912 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1604666999
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 7728 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1604666999
transform 1 0 7360 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_66
timestamp 1604666999
transform 1 0 7176 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1604666999
transform 1 0 7544 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_1_
timestamp 1604666999
transform 1 0 10212 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 10028 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 9660 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 9292 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_83
timestamp 1604666999
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_87
timestamp 1604666999
transform 1 0 9108 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_91
timestamp 1604666999
transform 1 0 9476 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1604666999
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 11776 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 11224 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_108
timestamp 1604666999
transform 1 0 11040 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_112
timestamp 1604666999
transform 1 0 11408 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_118
timestamp 1604666999
transform 1 0 11960 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_1_
timestamp 1604666999
transform 1 0 13248 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1604666999
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 12604 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 13064 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_123
timestamp 1604666999
transform 1 0 12420 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_127
timestamp 1604666999
transform 1 0 12788 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_0_
timestamp 1604666999
transform 1 0 14812 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_141
timestamp 1604666999
transform 1 0 14076 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_145
timestamp 1604666999
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_158
timestamp 1604666999
transform 1 0 15640 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_162
timestamp 1604666999
transform 1 0 16008 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1604666999
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18124 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1604666999
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1604666999
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_184
timestamp 1604666999
transform 1 0 18032 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 20884 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 20516 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 20148 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_204
timestamp 1604666999
transform 1 0 19872 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1604666999
transform 1 0 20332 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_213
timestamp 1604666999
transform 1 0 20700 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1604666999
transform 1 0 21068 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21436 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 23000 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 22448 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_230
timestamp 1604666999
transform 1 0 22264 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_234
timestamp 1604666999
transform 1 0 22632 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_2_
timestamp 1604666999
transform 1 0 23828 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1604666999
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_240
timestamp 1604666999
transform 1 0 23184 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_245
timestamp 1604666999
transform 1 0 23644 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_256
timestamp 1604666999
transform 1 0 24656 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l3_in_0_
timestamp 1604666999
transform 1 0 25392 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26404 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 24840 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 25208 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_260
timestamp 1604666999
transform 1 0 25024 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_273
timestamp 1604666999
transform 1 0 26220 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_277
timestamp 1604666999
transform 1 0 26588 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_1_
timestamp 1604666999
transform 1 0 26956 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 26772 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 27968 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_290
timestamp 1604666999
transform 1 0 27784 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_294
timestamp 1604666999
transform 1 0 28152 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1604666999
transform -1 0 28888 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_298
timestamp 1604666999
transform 1 0 28520 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l2_in_0_
timestamp 1604666999
transform 1 0 2392 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1604666999
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1564 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_3
timestamp 1604666999
transform 1 0 1380 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_7
timestamp 1604666999
transform 1 0 1748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1604666999
transform 1 0 2116 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_1.mux_l1_in_1_
timestamp 1604666999
transform 1 0 4048 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1604666999
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 3772 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_23
timestamp 1604666999
transform 1 0 3220 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1604666999
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5612 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5244 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_41
timestamp 1604666999
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_47
timestamp 1604666999
transform 1 0 5428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7544 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_68
timestamp 1604666999
transform 1 0 7360 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1604666999
transform 1 0 7728 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_76
timestamp 1604666999
transform 1 0 8096 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 10028 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1604666999
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 8740 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_81
timestamp 1604666999
transform 1 0 8556 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_85
timestamp 1604666999
transform 1 0 8924 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_91
timestamp 1604666999
transform 1 0 9476 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1604666999
transform 1 0 9660 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 11960 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_116
timestamp 1604666999
transform 1 0 11776 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l1_in_1_
timestamp 1604666999
transform 1 0 12512 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 13524 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_120
timestamp 1604666999
transform 1 0 12144 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_133
timestamp 1604666999
transform 1 0 13340 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_137
timestamp 1604666999
transform 1 0 13708 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l3_in_0_
timestamp 1604666999
transform 1 0 15548 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1604666999
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 14812 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14444 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1604666999
transform 1 0 14628 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1604666999
transform 1 0 14996 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_154
timestamp 1604666999
transform 1 0 15272 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 17112 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16928 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_166
timestamp 1604666999
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1604666999
transform 1 0 16744 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_193
timestamp 1604666999
transform 1 0 18860 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1604666999
transform 1 0 19780 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 20884 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1604666999
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 19412 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_201
timestamp 1604666999
transform 1 0 19596 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_206
timestamp 1604666999
transform 1 0 20056 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_210
timestamp 1604666999
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_234
timestamp 1604666999
transform 1 0 22632 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 23368 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1604666999
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 26128 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 25760 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 25392 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_261
timestamp 1604666999
transform 1 0 25116 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_266
timestamp 1604666999
transform 1 0 25576 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_270
timestamp 1604666999
transform 1 0 25944 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_274
timestamp 1604666999
transform 1 0 26312 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 27508 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_285
timestamp 1604666999
transform 1 0 27324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1604666999
transform 1 0 27692 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_297
timestamp 1604666999
transform 1 0 28428 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1604666999
transform -1 0 28888 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1656 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1472 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1604666999
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1604666999
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1604666999
transform 1 0 1380 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1604666999
transform 1 0 1380 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_23
timestamp 1604666999
transform 1 0 3220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1604666999
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_29
timestamp 1604666999
transform 1 0 3772 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_25
timestamp 1604666999
transform 1 0 3404 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 3772 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 3404 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_1.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3588 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_34
timestamp 1604666999
transform 1 0 4232 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1604666999
transform 1 0 4048 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1604666999
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1604666999
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_36
timestamp 1604666999
transform 1 0 4416 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_39
timestamp 1604666999
transform 1 0 4692 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4692 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_41
timestamp 1604666999
transform 1 0 4876 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 5060 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_0_
timestamp 1604666999
transform 1 0 5060 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_0_
timestamp 1604666999
transform 1 0 5244 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1604666999
transform 1 0 6440 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_54
timestamp 1604666999
transform 1 0 6072 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_56
timestamp 1604666999
transform 1 0 6256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_52
timestamp 1604666999
transform 1 0 5888 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 6072 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_64
timestamp 1604666999
transform 1 0 6992 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1604666999
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_75
timestamp 1604666999
transform 1 0 8004 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_71
timestamp 1604666999
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 8188 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 8372 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 7084 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l3_in_0_
timestamp 1604666999
transform 1 0 9936 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1604666999
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 9016 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 1604666999
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1604666999
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_88
timestamp 1604666999
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_93
timestamp 1604666999
transform 1 0 9660 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_105
timestamp 1604666999
transform 1 0 10764 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1604666999
transform 1 0 10856 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_102
timestamp 1604666999
transform 1 0 10488 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11040 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 10672 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_113
timestamp 1604666999
transform 1 0 11500 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_118
timestamp 1604666999
transform 1 0 11960 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_114
timestamp 1604666999
transform 1 0 11592 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1604666999
transform 1 0 11224 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 11776 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_2_
timestamp 1604666999
transform 1 0 11776 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_125
timestamp 1604666999
transform 1 0 12604 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 12788 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 12144 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1604666999
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l2_in_3_
timestamp 1604666999
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_20_133
timestamp 1604666999
transform 1 0 13340 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_129
timestamp 1604666999
transform 1 0 12972 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1604666999
transform 1 0 13800 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1604666999
transform 1 0 13248 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13156 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 13616 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l2_in_2_
timestamp 1604666999
transform 1 0 13616 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_145
timestamp 1604666999
transform 1 0 14444 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_146
timestamp 1604666999
transform 1 0 14536 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 1604666999
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 14352 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 13984 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_158
timestamp 1604666999
transform 1 0 15640 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_154
timestamp 1604666999
transform 1 0 15272 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1604666999
transform 1 0 15088 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_149
timestamp 1604666999
transform 1 0 14812 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1604666999
transform 1 0 15640 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 15456 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1604666999
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l3_in_1_
timestamp 1604666999
transform 1 0 14812 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1604666999
transform 1 0 16008 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1604666999
transform 1 0 16008 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 15824 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 15824 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 16192 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_10.mux_l4_in_0_
timestamp 1604666999
transform 1 0 16376 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_19_175
timestamp 1604666999
transform 1 0 17204 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 17388 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16560 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_20_187
timestamp 1604666999
transform 1 0 18308 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_188
timestamp 1604666999
transform 1 0 18400 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1604666999
transform 1 0 18032 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_179
timestamp 1604666999
transform 1 0 17572 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1604666999
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_195
timestamp 1604666999
transform 1 0 19044 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_195
timestamp 1604666999
transform 1 0 19044 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_191
timestamp 1604666999
transform 1 0 18676 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18492 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 18860 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 19228 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_1_
timestamp 1604666999
transform 1 0 19228 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1604666999
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1604666999
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_11.mux_l4_in_0_
timestamp 1604666999
transform 1 0 19412 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1604666999
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_210
timestamp 1604666999
transform 1 0 20424 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1604666999
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 20608 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 21068 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 20792 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1604666999
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_11.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 20976 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l1_in_2_
timestamp 1604666999
transform 1 0 21436 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 22908 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1604666999
transform 1 0 22724 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_219
timestamp 1604666999
transform 1 0 21252 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_230
timestamp 1604666999
transform 1 0 22264 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_238
timestamp 1604666999
transform 1 0 23000 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_242
timestamp 1604666999
transform 1 0 23368 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_245
timestamp 1604666999
transform 1 0 23644 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_239
timestamp 1604666999
transform 1 0 23092 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 23184 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 23552 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 23368 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1604666999
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l2_in_3_
timestamp 1604666999
transform 1 0 23736 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_255
timestamp 1604666999
transform 1 0 24564 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_257
timestamp 1604666999
transform 1 0 24748 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 24748 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l4_in_0_
timestamp 1604666999
transform 1 0 23920 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_267
timestamp 1604666999
transform 1 0 25668 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_259
timestamp 1604666999
transform 1 0 24932 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_265
timestamp 1604666999
transform 1 0 25484 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_261
timestamp 1604666999
transform 1 0 25116 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 25116 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 24932 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1604666999
transform 1 0 25300 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1604666999
transform 1 0 25300 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_271
timestamp 1604666999
transform 1 0 26036 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_269
timestamp 1604666999
transform 1 0 25852 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 26220 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 25852 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 25944 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1604666999
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_15.mux_l1_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26128 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 28060 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_291
timestamp 1604666999
transform 1 0 27876 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_295
timestamp 1604666999
transform 1 0 28244 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_285
timestamp 1604666999
transform 1 0 27324 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_297
timestamp 1604666999
transform 1 0 28428 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1604666999
transform -1 0 28888 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1604666999
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 2208 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1604666999
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 1840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1604666999
transform 1 0 1380 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1604666999
transform 1 0 1748 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_10
timestamp 1604666999
transform 1 0 2024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4692 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1604666999
transform 1 0 4140 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_31
timestamp 1604666999
transform 1 0 3956 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1604666999
transform 1 0 4324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 5704 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 6164 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 1604666999
transform 1 0 5520 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_52
timestamp 1604666999
transform 1 0 5888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1604666999
transform 1 0 6348 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1604666999
transform 1 0 8372 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_2_
timestamp 1604666999
transform 1 0 6808 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1604666999
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_71
timestamp 1604666999
transform 1 0 7636 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1604666999
transform 1 0 8188 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 9844 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 8832 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9660 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 9200 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp 1604666999
transform 1 0 8648 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_86
timestamp 1604666999
transform 1 0 9016 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_90
timestamp 1604666999
transform 1 0 9384 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 11776 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_114
timestamp 1604666999
transform 1 0 11592 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1604666999
transform 1 0 11960 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 12420 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1604666999
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 12144 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_1_
timestamp 1604666999
transform 1 0 14904 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 14720 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 14352 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_142
timestamp 1604666999
transform 1 0 14168 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_146
timestamp 1604666999
transform 1 0 14536 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 17112 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 17480 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 15916 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 16284 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_159
timestamp 1604666999
transform 1 0 15732 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_163
timestamp 1604666999
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_167
timestamp 1604666999
transform 1 0 16468 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1604666999
transform 1 0 17020 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1604666999
transform 1 0 17296 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1604666999
transform 1 0 18216 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1604666999
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 19320 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 18952 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1604666999
transform 1 0 17664 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1604666999
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_189
timestamp 1604666999
transform 1 0 18492 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_193
timestamp 1604666999
transform 1 0 18860 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1604666999
transform 1 0 19136 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 21068 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l3_in_0_
timestamp 1604666999
transform 1 0 19504 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 20884 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20516 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_209
timestamp 1604666999
transform 1 0 20332 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_213
timestamp 1604666999
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23000 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_236
timestamp 1604666999
transform 1 0 22816 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l3_in_1_
timestamp 1604666999
transform 1 0 24012 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1604666999
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 23828 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 23368 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_240
timestamp 1604666999
transform 1 0 23184 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_245
timestamp 1604666999
transform 1 0 23644 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 25576 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_15.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 25024 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_258
timestamp 1604666999
transform 1 0 24840 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_262
timestamp 1604666999
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 27508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 27876 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 28244 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_285
timestamp 1604666999
transform 1 0 27324 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_289
timestamp 1604666999
transform 1 0 27692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_293
timestamp 1604666999
transform 1 0 28060 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_297
timestamp 1604666999
transform 1 0 28428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1604666999
transform -1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_1_
timestamp 1604666999
transform 1 0 1840 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1604666999
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 1656 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 2852 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3
timestamp 1604666999
transform 1 0 1380 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_17
timestamp 1604666999
transform 1 0 2668 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1604666999
transform 1 0 4048 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1604666999
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 3220 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 4692 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_21
timestamp 1604666999
transform 1 0 3036 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_25
timestamp 1604666999
transform 1 0 3404 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 1604666999
transform 1 0 3772 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_36
timestamp 1604666999
transform 1 0 4416 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 5520 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 5152 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp 1604666999
transform 1 0 4876 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_46
timestamp 1604666999
transform 1 0 5336 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 7820 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_67
timestamp 1604666999
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 1604666999
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l4_in_0_
timestamp 1604666999
transform 1 0 9752 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1604666999
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 9384 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 9016 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1604666999
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_88
timestamp 1604666999
transform 1 0 9200 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp 1604666999
transform 1 0 9660 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 11316 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 10764 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 11132 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_103
timestamp 1604666999
transform 1 0 10580 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1604666999
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1604666999
transform 1 0 13800 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_5.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 13248 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 13616 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_130
timestamp 1604666999
transform 1 0 13064 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1604666999
transform 1 0 13432 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_0_
timestamp 1604666999
transform 1 0 15272 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1604666999
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 14628 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 14260 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1604666999
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_145
timestamp 1604666999
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_149
timestamp 1604666999
transform 1 0 14812 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 17112 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 16284 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_163
timestamp 1604666999
transform 1 0 16100 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_167
timestamp 1604666999
transform 1 0 16468 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_173
timestamp 1604666999
transform 1 0 17020 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 19136 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1604666999
transform 1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1604666999
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19504 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_202
timestamp 1604666999
transform 1 0 19688 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 19872 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_206
timestamp 1604666999
transform 1 0 20056 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 20240 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1604666999
transform 1 0 20424 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 20608 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1604666999
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1604666999
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 21068 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1604666999
transform 1 0 22908 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_1_
timestamp 1604666999
transform 1 0 21252 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 22724 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 22264 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_228
timestamp 1604666999
transform 1 0 22080 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_232
timestamp 1604666999
transform 1 0 22448 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 23920 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 23736 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 23368 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_240
timestamp 1604666999
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_244
timestamp 1604666999
transform 1 0 23552 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l4_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1604666999
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_267
timestamp 1604666999
transform 1 0 25668 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 27508 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_285
timestamp 1604666999
transform 1 0 27324 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_289
timestamp 1604666999
transform 1 0 27692 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_297
timestamp 1604666999
transform 1 0 28428 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1604666999
transform -1 0 28888 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_2_
timestamp 1604666999
transform 1 0 2024 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1604666999
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 1840 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1604666999
transform 1 0 1380 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1604666999
transform 1 0 1748 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_19
timestamp 1604666999
transform 1 0 2852 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_0_
timestamp 1604666999
transform 1 0 3588 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 3404 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 3036 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1604666999
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1604666999
transform 1 0 3220 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1604666999
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_4.mux_l1_in_1_
timestamp 1604666999
transform 1 0 5152 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_40
timestamp 1604666999
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_53
timestamp 1604666999
transform 1 0 5980 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1604666999
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 8096 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1604666999
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 7176 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1604666999
transform 1 0 6808 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1604666999
transform 1 0 7360 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_72
timestamp 1604666999
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_95
timestamp 1604666999
transform 1 0 9844 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_99
timestamp 1604666999
transform 1 0 10212 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_5.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 10304 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11868 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_102
timestamp 1604666999
transform 1 0 10488 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_114
timestamp 1604666999
transform 1 0 11592 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_119
timestamp 1604666999
transform 1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l3_in_0_
timestamp 1604666999
transform 1 0 13064 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1604666999
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12604 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1604666999
transform 1 0 12420 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_127
timestamp 1604666999
transform 1 0 12788 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_1_
timestamp 1604666999
transform 1 0 14628 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 14444 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 14076 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1604666999
transform 1 0 13892 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_143
timestamp 1604666999
transform 1 0 14260 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1604666999
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_0_
timestamp 1604666999
transform 1 0 16192 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 16008 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_160
timestamp 1604666999
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_173
timestamp 1604666999
transform 1 0 17020 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1604666999
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18308 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 18676 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 19320 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_181
timestamp 1604666999
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_184
timestamp 1604666999
transform 1 0 18032 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_189
timestamp 1604666999
transform 1 0 18492 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_193
timestamp 1604666999
transform 1 0 18860 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_197
timestamp 1604666999
transform 1 0 19228 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 21068 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_0_
timestamp 1604666999
transform 1 0 19504 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 20516 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_209
timestamp 1604666999
transform 1 0 20332 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_213
timestamp 1604666999
transform 1 0 20700 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 23000 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_236
timestamp 1604666999
transform 1 0 22816 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 24196 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1604666999
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 24012 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 23368 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_240
timestamp 1604666999
transform 1 0 23184 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1604666999
transform 1 0 23644 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 26496 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 26128 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_270
timestamp 1604666999
transform 1 0 25944 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_274
timestamp 1604666999
transform 1 0 26312 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26680 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 27692 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 28060 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 28428 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_287
timestamp 1604666999
transform 1 0 27508 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_291
timestamp 1604666999
transform 1 0 27876 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_295
timestamp 1604666999
transform 1 0 28244 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1604666999
transform -1 0 28888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l2_in_3_
timestamp 1604666999
transform 1 0 2024 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1604666999
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1604666999
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_7
timestamp 1604666999
transform 1 0 1748 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1604666999
transform 1 0 2852 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1604666999
transform 1 0 4048 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1604666999
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 3036 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3404 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4600 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1604666999
transform 1 0 3220 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1604666999
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_36
timestamp 1604666999
transform 1 0 4416 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 5336 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 5152 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_40
timestamp 1604666999
transform 1 0 4784 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 7820 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 1604666999
transform 1 0 7084 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1604666999
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 9016 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 10120 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 9384 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1604666999
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_88
timestamp 1604666999
transform 1 0 9200 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_93
timestamp 1604666999
transform 1 0 9660 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_97
timestamp 1604666999
transform 1 0 10028 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11868 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l1_in_0_
timestamp 1604666999
transform 1 0 10304 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_109
timestamp 1604666999
transform 1 0 11132 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 1604666999
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_136
timestamp 1604666999
transform 1 0 13616 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 15272 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1604666999
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 14628 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_140
timestamp 1604666999
transform 1 0 13984 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_146
timestamp 1604666999
transform 1 0 14536 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1604666999
transform 1 0 14812 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_173
timestamp 1604666999
transform 1 0 17020 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18308 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_181
timestamp 1604666999
transform 1 0 17756 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_186
timestamp 1604666999
transform 1 0 18216 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l3_in_0_
timestamp 1604666999
transform 1 0 21160 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1604666999
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_206
timestamp 1604666999
transform 1 0 20056 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_24_215
timestamp 1604666999
transform 1 0 20884 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_2_
timestamp 1604666999
transform 1 0 22724 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 22172 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_227
timestamp 1604666999
transform 1 0 21988 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1604666999
transform 1 0 22356 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 24656 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 24196 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 23828 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_244
timestamp 1604666999
transform 1 0 23552 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_249
timestamp 1604666999
transform 1 0 24012 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_253
timestamp 1604666999
transform 1 0 24380 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_1_
timestamp 1604666999
transform 1 0 24840 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_14.mux_l1_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1604666999
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 26128 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_267
timestamp 1604666999
transform 1 0 25668 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_271
timestamp 1604666999
transform 1 0 26036 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1604666999
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 27508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_285
timestamp 1604666999
transform 1 0 27324 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_289
timestamp 1604666999
transform 1 0 27692 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_297
timestamp 1604666999
transform 1 0 28428 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1604666999
transform -1 0 28888 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 1656 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1604666999
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1604666999
transform 1 0 1380 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4140 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 3588 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 3956 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_25
timestamp 1604666999
transform 1 0 3404 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1604666999
transform 1 0 3772 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 5520 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 5888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1604666999
transform 1 0 4968 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_46
timestamp 1604666999
transform 1 0 5336 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1604666999
transform 1 0 5704 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_54
timestamp 1604666999
transform 1 0 6072 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_62
timestamp 1604666999
transform 1 0 6808 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1604666999
transform 1 0 6624 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 7084 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1604666999
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1604666999
transform 1 0 7268 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_77
timestamp 1604666999
transform 1 0 8188 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_74
timestamp 1604666999
transform 1 0 7912 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_70
timestamp 1604666999
transform 1 0 7544 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 8280 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 10212 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1604666999
transform 1 0 10028 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_3_
timestamp 1604666999
transform 1 0 10764 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 10580 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 11776 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1604666999
transform 1 0 10396 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_114
timestamp 1604666999
transform 1 0 11592 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_118
timestamp 1604666999
transform 1 0 11960 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l1_in_2_
timestamp 1604666999
transform 1 0 13432 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1604666999
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 12144 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_123
timestamp 1604666999
transform 1 0 12420 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_127
timestamp 1604666999
transform 1 0 12788 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_130
timestamp 1604666999
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_2_
timestamp 1604666999
transform 1 0 14996 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 14812 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 14444 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 1604666999
transform 1 0 14260 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1604666999
transform 1 0 14628 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 16008 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 1604666999
transform 1 0 15824 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_164
timestamp 1604666999
transform 1 0 16192 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_176
timestamp 1604666999
transform 1 0 17296 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 18032 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1604666999
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 17756 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_179
timestamp 1604666999
transform 1 0 17572 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 19964 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 21160 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 20792 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20424 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1604666999
transform 1 0 19780 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_207
timestamp 1604666999
transform 1 0 20148 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_212
timestamp 1604666999
transform 1 0 20608 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_216
timestamp 1604666999
transform 1 0 20976 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l3_in_1_
timestamp 1604666999
transform 1 0 21436 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 22448 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 23000 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_220
timestamp 1604666999
transform 1 0 21344 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_230
timestamp 1604666999
transform 1 0 22264 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1604666999
transform 1 0 22632 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_2_
timestamp 1604666999
transform 1 0 24564 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1604666999
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 24380 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 23368 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_240
timestamp 1604666999
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_245
timestamp 1604666999
transform 1 0 23644 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_251
timestamp 1604666999
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 26128 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 25944 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 25576 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_264
timestamp 1604666999
transform 1 0 25392 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_268
timestamp 1604666999
transform 1 0 25760 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 28060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_291
timestamp 1604666999
transform 1 0 27876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_295
timestamp 1604666999
transform 1 0 28244 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1604666999
transform -1 0 28888 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 1472 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 1748 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1604666999
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1604666999
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 1564 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1604666999
transform 1 0 1380 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1604666999
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1604666999
transform 1 0 3496 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1604666999
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_23
timestamp 1604666999
transform 1 0 3220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3680 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 3772 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_2.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 3404 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_30
timestamp 1604666999
transform 1 0 3864 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_39
timestamp 1604666999
transform 1 0 4692 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_35
timestamp 1604666999
transform 1 0 4324 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 4048 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1604666999
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1604666999
transform 1 0 4048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 4232 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_4.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 5152 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 4968 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_53
timestamp 1604666999
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1604666999
transform 1 0 6348 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_67
timestamp 1604666999
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_62
timestamp 1604666999
transform 1 0 6808 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1604666999
transform 1 0 7268 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1604666999
transform 1 0 6900 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 7084 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 7452 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 7084 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 7452 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1604666999
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1604666999
transform 1 0 7636 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_6.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l4_in_0_
timestamp 1604666999
transform 1 0 7636 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_2_
timestamp 1604666999
transform 1 0 8004 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1604666999
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_80
timestamp 1604666999
transform 1 0 8464 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_84
timestamp 1604666999
transform 1 0 8832 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 9200 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 9016 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_90
timestamp 1604666999
transform 1 0 9384 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1604666999
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l2_in_0_
timestamp 1604666999
transform 1 0 9660 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 9200 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_27_107
timestamp 1604666999
transform 1 0 10948 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_107
timestamp 1604666999
transform 1 0 10948 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_102
timestamp 1604666999
transform 1 0 10488 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 11132 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 10764 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1604666999
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1604666999
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1604666999
transform 1 0 11316 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1604666999
transform 1 0 11316 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 11408 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 11408 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1604666999
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_136
timestamp 1604666999
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_132
timestamp 1604666999
transform 1 0 13248 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1604666999
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_131
timestamp 1604666999
transform 1 0 13156 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 13800 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 13432 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 13432 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1604666999
transform 1 0 14720 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1604666999
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_140
timestamp 1604666999
transform 1 0 13984 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_144
timestamp 1604666999
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_140
timestamp 1604666999
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_150
timestamp 1604666999
transform 1 0 14904 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 14996 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 14904 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1604666999
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 15088 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 15272 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 17020 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_173
timestamp 1604666999
transform 1 0 17020 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1604666999
transform 1 0 16836 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1604666999
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1604666999
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1604666999
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1604666999
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_186
timestamp 1604666999
transform 1 0 18216 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_181
timestamp 1604666999
transform 1 0 17756 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__S
timestamp 1604666999
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_10.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 18032 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1604666999
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_198
timestamp 1604666999
transform 1 0 19320 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A1
timestamp 1604666999
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_0_
timestamp 1604666999
transform 1 0 18492 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 18768 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_26_202
timestamp 1604666999
transform 1 0 19688 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_1__A0
timestamp 1604666999
transform 1 0 19504 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_218
timestamp 1604666999
transform 1 0 21160 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_215
timestamp 1604666999
transform 1 0 20884 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_211
timestamp 1604666999
transform 1 0 20516 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_215
timestamp 1604666999
transform 1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1604666999
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 20608 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 20976 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1604666999
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 21160 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l1_in_0_
timestamp 1604666999
transform 1 0 21988 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 21804 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 23000 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_237
timestamp 1604666999
transform 1 0 22908 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_223
timestamp 1604666999
transform 1 0 21620 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_236
timestamp 1604666999
transform 1 0 22816 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_1_
timestamp 1604666999
transform 1 0 23920 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_1_
timestamp 1604666999
transform 1 0 24104 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1604666999
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 23920 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 23368 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_245
timestamp 1604666999
transform 1 0 23644 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 1604666999
transform 1 0 23184 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_245
timestamp 1604666999
transform 1 0 23644 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_263
timestamp 1604666999
transform 1 0 25300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_259
timestamp 1604666999
transform 1 0 24932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1604666999
transform 1 0 25668 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 25116 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 25484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_271
timestamp 1604666999
transform 1 0 26036 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 25852 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 26220 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1604666999
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_0_
timestamp 1604666999
transform 1 0 26496 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 25668 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 27600 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 27968 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_285
timestamp 1604666999
transform 1 0 27324 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_297
timestamp 1604666999
transform 1 0 28428 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_286
timestamp 1604666999
transform 1 0 27416 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_290
timestamp 1604666999
transform 1 0 27784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_294
timestamp 1604666999
transform 1 0 28152 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1604666999
transform -1 0 28888 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1604666999
transform -1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_298
timestamp 1604666999
transform 1 0 28520 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l4_in_0_
timestamp 1604666999
transform 1 0 1656 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1604666999
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 2668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1604666999
transform 1 0 1380 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_15
timestamp 1604666999
transform 1 0 2484 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_19
timestamp 1604666999
transform 1 0 2852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1604666999
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 3312 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_1__D
timestamp 1604666999
transform 1 0 4232 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 3680 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_23
timestamp 1604666999
transform 1 0 3220 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1604666999
transform 1 0 3496 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1604666999
transform 1 0 3864 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1604666999
transform 1 0 4048 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1604666999
transform 1 0 4416 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 4968 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 4784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l3_in_1_
timestamp 1604666999
transform 1 0 8004 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_61
timestamp 1604666999
transform 1 0 6716 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_65
timestamp 1604666999
transform 1 0 7084 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_69
timestamp 1604666999
transform 1 0 7452 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_73
timestamp 1604666999
transform 1 0 7820 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1604666999
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_84
timestamp 1604666999
transform 1 0 8832 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1604666999
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_97
timestamp 1604666999
transform 1 0 10028 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1604666999
transform 1 0 10396 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l1_in_0_
timestamp 1604666999
transform 1 0 11408 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 11224 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 10856 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_104
timestamp 1604666999
transform 1 0 10672 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_108
timestamp 1604666999
transform 1 0 11040 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l4_in_0_
timestamp 1604666999
transform 1 0 13616 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 12420 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1604666999
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_125
timestamp 1604666999
transform 1 0 12604 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_129
timestamp 1604666999
transform 1 0 12972 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_133
timestamp 1604666999
transform 1 0 13340 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1604666999
transform 1 0 15272 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1604666999
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__CLK
timestamp 1604666999
transform 1 0 14628 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 1604666999
transform 1 0 14444 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_149
timestamp 1604666999
transform 1 0 14812 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_157
timestamp 1604666999
transform 1 0 15548 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 16652 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_1_
timestamp 1604666999
transform 1 0 19136 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_1__CLK
timestamp 1604666999
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_188
timestamp 1604666999
transform 1 0 18400 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1604666999
transform 1 0 18952 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l4_in_0_
timestamp 1604666999
transform 1 0 20976 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1604666999
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 20148 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1604666999
transform 1 0 19964 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_209
timestamp 1604666999
transform 1 0 20332 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_215
timestamp 1604666999
transform 1 0 20884 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 22540 0 -1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 21988 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 22356 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_225
timestamp 1604666999
transform 1 0 21804 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_229
timestamp 1604666999
transform 1 0 22172 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 24472 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_252
timestamp 1604666999
transform 1 0 24288 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_256
timestamp 1604666999
transform 1 0 24656 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_2_
timestamp 1604666999
transform 1 0 26496 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1604666999
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_14.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 25668 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 24840 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 26220 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 25208 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_260
timestamp 1604666999
transform 1 0 25024 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_264
timestamp 1604666999
transform 1 0 25392 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_269
timestamp 1604666999
transform 1 0 25852 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_285
timestamp 1604666999
transform 1 0 27324 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_297
timestamp 1604666999
transform 1 0 28428 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1604666999
transform -1 0 28888 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_2.mux_l3_in_0_
timestamp 1604666999
transform 1 0 1564 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1604666999
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 2576 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1604666999
transform 1 0 1380 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_14
timestamp 1604666999
transform 1 0 2392 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_18
timestamp 1604666999
transform 1 0 2760 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_3_
timestamp 1604666999
transform 1 0 3312 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A1
timestamp 1604666999
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 3128 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__A0
timestamp 1604666999
transform 1 0 4324 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_33
timestamp 1604666999
transform 1 0 4140 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_37
timestamp 1604666999
transform 1 0 4508 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l1_in_0_
timestamp 1604666999
transform 1 0 4876 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l1_in_0__S
timestamp 1604666999
transform 1 0 5888 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_50
timestamp 1604666999
transform 1 0 5704 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_54
timestamp 1604666999
transform 1 0 6072 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_58
timestamp 1604666999
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_1_
timestamp 1604666999
transform 1 0 6808 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1604666999
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 8372 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_71
timestamp 1604666999
transform 1 0 7636 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_75
timestamp 1604666999
transform 1 0 8004 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_6.mux_l3_in_0_
timestamp 1604666999
transform 1 0 8556 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 10212 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_90
timestamp 1604666999
transform 1 0 9384 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1604666999
transform 1 0 9844 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_2_
timestamp 1604666999
transform 1 0 10764 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 10580 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 11776 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1604666999
transform 1 0 10396 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1604666999
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1604666999
transform 1 0 11960 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_1_
timestamp 1604666999
transform 1 0 12420 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1604666999
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 12144 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1604666999
transform 1 0 13248 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_138
timestamp 1604666999
transform 1 0 13800 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0_
timestamp 1604666999
transform 1 0 13984 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 16468 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 16836 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 17388 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1604666999
transform 1 0 15732 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1604666999
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_173
timestamp 1604666999
transform 1 0 17020 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l3_in_0_
timestamp 1604666999
transform 1 0 18032 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1604666999
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 19044 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1604666999
transform 1 0 17572 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_193
timestamp 1604666999
transform 1 0 18860 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1604666999
transform 1 0 19228 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_3_
timestamp 1604666999
transform 1 0 19596 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 19412 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 21160 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1604666999
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_214
timestamp 1604666999
transform 1 0 20792 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_12.mux_l2_in_3_
timestamp 1604666999
transform 1 0 21712 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 21528 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 22724 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_220
timestamp 1604666999
transform 1 0 21344 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_233
timestamp 1604666999
transform 1 0 22540 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_237
timestamp 1604666999
transform 1 0 22908 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l3_in_0_
timestamp 1604666999
transform 1 0 24104 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1604666999
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 23092 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 23920 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_241
timestamp 1604666999
transform 1 0 23276 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_245
timestamp 1604666999
transform 1 0 23644 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 25668 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 25484 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 25116 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_259
timestamp 1604666999
transform 1 0 24932 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_263
timestamp 1604666999
transform 1 0 25300 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 27600 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 27968 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_286
timestamp 1604666999
transform 1 0 27416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_290
timestamp 1604666999
transform 1 0 27784 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_294
timestamp 1604666999
transform 1 0 28152 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1604666999
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_298
timestamp 1604666999
transform 1 0 28520 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1604666999
transform 1 0 1380 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2484 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1604666999
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1604666999
transform 1 0 1932 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 2300 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1604666999
transform 1 0 1748 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1604666999
transform 1 0 2116 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1604666999
transform 1 0 2760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1604666999
transform 1 0 3128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_26
timestamp 1604666999
transform 1 0 3496 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 3772 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1604666999
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1604666999
transform 1 0 4048 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 4232 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_36
timestamp 1604666999
transform 1 0 4416 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 4600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_3.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 4784 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_30_59
timestamp 1604666999
transform 1 0 6532 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l3_in_0_
timestamp 1604666999
transform 1 0 7268 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 6808 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_64
timestamp 1604666999
transform 1 0 6992 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_76
timestamp 1604666999
transform 1 0 8096 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9660 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1604666999
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 8556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_6.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 8924 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_80
timestamp 1604666999
transform 1 0 8464 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_83
timestamp 1604666999
transform 1 0 8740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_87
timestamp 1604666999
transform 1 0 9108 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_91
timestamp 1604666999
transform 1 0 9476 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_96
timestamp 1604666999
transform 1 0 9936 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 11132 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_104
timestamp 1604666999
transform 1 0 10672 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_107
timestamp 1604666999
transform 1 0 10948 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l2_in_3_
timestamp 1604666999
transform 1 0 13616 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 13432 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_128
timestamp 1604666999
transform 1 0 12880 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1604666999
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_8.sky130_fd_sc_hd__dfxbp_1_0__D
timestamp 1604666999
transform 1 0 14628 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 15456 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 14996 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_145
timestamp 1604666999
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_149
timestamp 1604666999
transform 1 0 14812 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1604666999
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_158
timestamp 1604666999
transform 1 0 15640 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 16468 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_166
timestamp 1604666999
transform 1 0 16376 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_2_
timestamp 1604666999
transform 1 0 18952 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 18768 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1604666999
transform 1 0 18216 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1604666999
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1604666999
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 19964 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1604666999
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_207
timestamp 1604666999
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_211
timestamp 1604666999
transform 1 0 20516 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1604666999
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_12.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 21620 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l4_in_0_
timestamp 1604666999
transform 1 0 24748 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 24564 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 24104 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1604666999
transform 1 0 23368 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_252
timestamp 1604666999
transform 1 0 24288 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l3_in_1_
timestamp 1604666999
transform 1 0 26496 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1604666999
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 25760 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 26128 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_266
timestamp 1604666999
transform 1 0 25576 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_270
timestamp 1604666999
transform 1 0 25944 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_274
timestamp 1604666999
transform 1 0 26312 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_285
timestamp 1604666999
transform 1 0 27324 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_297
timestamp 1604666999
transform 1 0 28428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1604666999
transform -1 0 28888 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1604666999
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_2.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 1932 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 2852 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1604666999
transform 1 0 1380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1604666999
transform 1 0 1748 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_11
timestamp 1604666999
transform 1 0 2116 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l4_in_0_
timestamp 1604666999
transform 1 0 3404 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A1
timestamp 1604666999
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 3220 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_21
timestamp 1604666999
transform 1 0 3036 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1604666999
transform 1 0 4232 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1604666999
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_0_
timestamp 1604666999
transform 1 0 4968 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__A0
timestamp 1604666999
transform 1 0 5980 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_2__S
timestamp 1604666999
transform 1 0 6348 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1604666999
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1604666999
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1604666999
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1604666999
transform 1 0 6808 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1604666999
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_65
timestamp 1604666999
transform 1 0 7084 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_77
timestamp 1604666999
transform 1 0 8188 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 10212 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_89
timestamp 1604666999
transform 1 0 9292 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_97
timestamp 1604666999
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l3_in_1_
timestamp 1604666999
transform 1 0 10764 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 10580 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__S
timestamp 1604666999
transform 1 0 11776 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_101
timestamp 1604666999
transform 1 0 10396 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_114
timestamp 1604666999
transform 1 0 11592 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1604666999
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 12420 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1604666999
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l3_in_1_
timestamp 1604666999
transform 1 0 14904 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1604666999
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1604666999
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1604666999
transform 1 0 16100 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_159
timestamp 1604666999
transform 1 0 15732 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1604666999
transform 1 0 16468 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_170
timestamp 1604666999
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_178
timestamp 1604666999
transform 1 0 17480 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_174
timestamp 1604666999
transform 1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 17296 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1604666999
transform 1 0 18308 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2_
timestamp 1604666999
transform 1 0 19320 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1604666999
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__CLK
timestamp 1604666999
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_9.sky130_fd_sc_hd__dfxbp_1_2__D
timestamp 1604666999
transform 1 0 18768 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_184
timestamp 1604666999
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1604666999
transform 1 0 18584 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1604666999
transform 1 0 18952 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_217
timestamp 1604666999
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1604666999
transform 1 0 21804 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 21252 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 22264 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_221
timestamp 1604666999
transform 1 0 21436 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_228
timestamp 1604666999
transform 1 0 22080 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1604666999
transform 1 0 22448 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxbp_1  mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3_
timestamp 1604666999
transform 1 0 24564 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1604666999
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_13.sky130_fd_sc_hd__dfxbp_1_3__CLK
timestamp 1604666999
transform 1 0 24380 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1604666999
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__S
timestamp 1604666999
transform 1 0 26496 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_274
timestamp 1604666999
transform 1 0 26312 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_13.mux_l2_in_3_
timestamp 1604666999
transform 1 0 27048 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A1
timestamp 1604666999
transform 1 0 26864 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1604666999
transform 1 0 26680 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_291
timestamp 1604666999
transform 1 0 27876 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1604666999
transform -1 0 28888 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1604666999
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1604666999
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_15
timestamp 1604666999
transform 1 0 2484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 4232 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1604666999
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 3404 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1604666999
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1604666999
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1604666999
transform 1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_37
timestamp 1604666999
transform 1 0 4508 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l2_in_2_
timestamp 1604666999
transform 1 0 5244 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 4968 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_41
timestamp 1604666999
transform 1 0 4876 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1604666999
transform 1 0 5152 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_54
timestamp 1604666999
transform 1 0 6072 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_66
timestamp 1604666999
transform 1 0 7176 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_78
timestamp 1604666999
transform 1 0 8280 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1604666999
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1604666999
transform 1 0 9384 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1604666999
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l3_in_0_
timestamp 1604666999
transform 1 0 11592 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A1
timestamp 1604666999
transform 1 0 11408 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 10764 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_107
timestamp 1604666999
transform 1 0 10948 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_111
timestamp 1604666999
transform 1 0 11316 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_7.sky130_fd_sc_hd__dfxbp_1_3__D
timestamp 1604666999
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_123
timestamp 1604666999
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_127
timestamp 1604666999
transform 1 0 12788 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_8.mux_l2_in_3_
timestamp 1604666999
transform 1 0 15272 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1604666999
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_139
timestamp 1604666999
transform 1 0 13892 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_147
timestamp 1604666999
transform 1 0 14628 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1604666999
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l4_in_0_
timestamp 1604666999
transform 1 0 17296 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_163
timestamp 1604666999
transform 1 0 16100 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_169
timestamp 1604666999
transform 1 0 16652 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_172
timestamp 1604666999
transform 1 0 16928 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l3_in_1_
timestamp 1604666999
transform 1 0 18860 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A0
timestamp 1604666999
transform 1 0 18584 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_185
timestamp 1604666999
transform 1 0 18124 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_189
timestamp 1604666999
transform 1 0 18492 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_192
timestamp 1604666999
transform 1 0 18768 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1604666999
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__S
timestamp 1604666999
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_202
timestamp 1604666999
transform 1 0 19688 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_206
timestamp 1604666999
transform 1 0 20056 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1604666999
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1604666999
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_218
timestamp 1604666999
transform 1 0 21160 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_229
timestamp 1604666999
transform 1 0 22172 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_241
timestamp 1604666999
transform 1 0 23276 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1604666999
transform 1 0 24380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1604666999
transform 1 0 26496 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1604666999
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_265
timestamp 1604666999
transform 1 0 25484 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_273
timestamp 1604666999
transform 1 0 26220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.mux_l2_in_3__A0
timestamp 1604666999
transform 1 0 27048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_279
timestamp 1604666999
transform 1 0 26772 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_284
timestamp 1604666999
transform 1 0 27232 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1604666999
transform 1 0 28336 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1604666999
transform -1 0 28888 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_6
timestamp 1604666999
transform 1 0 1656 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 1840 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1604666999
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1604666999
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 1380 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_17
timestamp 1604666999
transform 1 0 2668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_10
timestamp 1604666999
transform 1 0 2024 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 2852 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 2392 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1604666999
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1604666999
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1604666999
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__S
timestamp 1604666999
transform 1 0 4692 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A0
timestamp 1604666999
transform 1 0 4324 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_21
timestamp 1604666999
transform 1 0 3036 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_33
timestamp 1604666999
transform 1 0 4140 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1604666999
transform 1 0 4508 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1604666999
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_32
timestamp 1604666999
transform 1 0 4048 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_3.mux_l3_in_1_
timestamp 1604666999
transform 1 0 4876 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_3.mux_l3_in_1__A1
timestamp 1604666999
transform 1 0 4876 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_50
timestamp 1604666999
transform 1 0 5704 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_58
timestamp 1604666999
transform 1 0 6440 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 1604666999
transform 1 0 4784 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_43
timestamp 1604666999
transform 1 0 5060 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_55
timestamp 1604666999
transform 1 0 6164 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 7084 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1604666999
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_62
timestamp 1604666999
transform 1 0 6808 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_68
timestamp 1604666999
transform 1 0 7360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_72
timestamp 1604666999
transform 1 0 7728 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_67
timestamp 1604666999
transform 1 0 7268 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_79
timestamp 1604666999
transform 1 0 8372 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 9292 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1604666999
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_5.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_84
timestamp 1604666999
transform 1 0 8832 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_88
timestamp 1604666999
transform 1 0 9200 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_92
timestamp 1604666999
transform 1 0 9568 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_96
timestamp 1604666999
transform 1 0 9936 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_91
timestamp 1604666999
transform 1 0 9476 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1604666999
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l3_in_0__A0
timestamp 1604666999
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 11224 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_108
timestamp 1604666999
transform 1 0 11040 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1604666999
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_116
timestamp 1604666999
transform 1 0 11776 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1604666999
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_117
timestamp 1604666999
transform 1 0 11868 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_123
timestamp 1604666999
transform 1 0 12420 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A1
timestamp 1604666999
transform 1 0 12604 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__S
timestamp 1604666999
transform 1 0 12144 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1604666999
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 12144 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_7.mux_l4_in_0_
timestamp 1604666999
transform 1 0 12420 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_33_136
timestamp 1604666999
transform 1 0 13616 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1604666999
transform 1 0 13248 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_7.mux_l4_in_0__A0
timestamp 1604666999
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_127
timestamp 1604666999
transform 1 0 12788 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 14444 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1604666999
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_8.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 14904 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_144
timestamp 1604666999
transform 1 0 14352 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1604666999
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_152
timestamp 1604666999
transform 1 0 15088 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_139
timestamp 1604666999
transform 1 0 13892 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_151
timestamp 1604666999
transform 1 0 14996 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1604666999
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 17296 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 16744 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__S
timestamp 1604666999
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_10.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 16560 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_164
timestamp 1604666999
transform 1 0 16192 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_173
timestamp 1604666999
transform 1 0 17020 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_166
timestamp 1604666999
transform 1 0 16376 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_174
timestamp 1604666999
transform 1 0 17112 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_179
timestamp 1604666999
transform 1 0 17572 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_184
timestamp 1604666999
transform 1 0 18032 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1604666999
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A0
timestamp 1604666999
transform 1 0 18124 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__S
timestamp 1604666999
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l1_in_2__A1
timestamp 1604666999
transform 1 0 18400 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1604666999
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_0_
timestamp 1604666999
transform 1 0 18308 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_34_196
timestamp 1604666999
transform 1 0 19136 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l1_in_2_
timestamp 1604666999
transform 1 0 18584 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_34_204
timestamp 1604666999
transform 1 0 19872 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1604666999
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_199
timestamp 1604666999
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A1
timestamp 1604666999
transform 1 0 20148 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_0__A1
timestamp 1604666999
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_9.mux_l2_in_1__A0
timestamp 1604666999
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_9.mux_l2_in_1_
timestamp 1604666999
transform 1 0 20148 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1604666999
transform 1 0 20700 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1604666999
transform 1 0 20332 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1604666999
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1604666999
transform 1 0 20884 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_216
timestamp 1604666999
transform 1 0 20976 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_228
timestamp 1604666999
transform 1 0 22080 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1604666999
transform 1 0 21988 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_245
timestamp 1604666999
transform 1 0 23644 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1604666999
transform 1 0 23184 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1604666999
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_257
timestamp 1604666999
transform 1 0 24748 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_253
timestamp 1604666999
transform 1 0 24380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_249
timestamp 1604666999
transform 1 0 24012 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 24564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 24104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_251
timestamp 1604666999
transform 1 0 24196 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1604666999
transform 1 0 23092 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 25208 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1604666999
transform 1 0 26404 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1604666999
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_14.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 25668 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_261
timestamp 1604666999
transform 1 0 25116 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_265
timestamp 1604666999
transform 1 0 25484 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_33_269
timestamp 1604666999
transform 1 0 25852 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_263
timestamp 1604666999
transform 1 0 25300 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1604666999
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_15.sky130_fd_sc_hd__buf_4_0__A
timestamp 1604666999
transform 1 0 26864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1604666999
transform 1 0 26680 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_282
timestamp 1604666999
transform 1 0 27048 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_294
timestamp 1604666999
transform 1 0 28152 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1604666999
transform 1 0 27600 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1604666999
transform 1 0 28336 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1604666999
transform -1 0 28888 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1604666999
transform -1 0 28888 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_298
timestamp 1604666999
transform 1 0 28520 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1604666999
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1604666999
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1604666999
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1604666999
transform 1 0 3956 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_27
timestamp 1604666999
transform 1 0 3588 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_32
timestamp 1604666999
transform 1 0 4048 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_44
timestamp 1604666999
transform 1 0 5152 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_56
timestamp 1604666999
transform 1 0 6256 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1604666999
transform 1 0 6808 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_63
timestamp 1604666999
transform 1 0 6900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_75
timestamp 1604666999
transform 1 0 8004 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1604666999
transform 1 0 9660 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_87
timestamp 1604666999
transform 1 0 9108 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1604666999
transform 1 0 9752 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1604666999
transform 1 0 10856 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_118
timestamp 1604666999
transform 1 0 11960 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1604666999
transform 1 0 12512 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1604666999
transform 1 0 12604 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1604666999
transform 1 0 13708 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1604666999
transform 1 0 15364 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_149
timestamp 1604666999
transform 1 0 14812 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_156
timestamp 1604666999
transform 1 0 15456 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_168
timestamp 1604666999
transform 1 0 16560 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1604666999
transform 1 0 18216 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_180
timestamp 1604666999
transform 1 0 17664 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_187
timestamp 1604666999
transform 1 0 18308 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1604666999
transform 1 0 21068 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_199
timestamp 1604666999
transform 1 0 19412 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_211
timestamp 1604666999
transform 1 0 20516 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_218
timestamp 1604666999
transform 1 0 21160 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_230
timestamp 1604666999
transform 1 0 22264 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1604666999
transform 1 0 23920 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_242
timestamp 1604666999
transform 1 0 23368 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_249
timestamp 1604666999
transform 1 0 24012 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_261
timestamp 1604666999
transform 1 0 25116 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1604666999
transform 1 0 26220 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1604666999
transform 1 0 26772 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_280
timestamp 1604666999
transform 1 0 26864 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_292
timestamp 1604666999
transform 1 0 27968 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1604666999
transform -1 0 28888 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_35_298
timestamp 1604666999
transform 1 0 28520 0 1 21216
box -38 -48 130 592
<< labels >>
rlabel metal2 s 3698 0 3754 480 6 bottom_grid_pin_0_
port 0 nsew default tristate
rlabel metal2 s 11150 0 11206 480 6 ccff_head
port 1 nsew default input
rlabel metal2 s 18694 0 18750 480 6 ccff_tail
port 2 nsew default tristate
rlabel metal3 s 0 12248 480 12368 6 chanx_left_in[0]
port 3 nsew default input
rlabel metal3 s 0 18232 480 18352 6 chanx_left_in[10]
port 4 nsew default input
rlabel metal3 s 0 18776 480 18896 6 chanx_left_in[11]
port 5 nsew default input
rlabel metal3 s 0 19320 480 19440 6 chanx_left_in[12]
port 6 nsew default input
rlabel metal3 s 0 20000 480 20120 6 chanx_left_in[13]
port 7 nsew default input
rlabel metal3 s 0 20544 480 20664 6 chanx_left_in[14]
port 8 nsew default input
rlabel metal3 s 0 21224 480 21344 6 chanx_left_in[15]
port 9 nsew default input
rlabel metal3 s 0 21768 480 21888 6 chanx_left_in[16]
port 10 nsew default input
rlabel metal3 s 0 22312 480 22432 6 chanx_left_in[17]
port 11 nsew default input
rlabel metal3 s 0 22992 480 23112 6 chanx_left_in[18]
port 12 nsew default input
rlabel metal3 s 0 23536 480 23656 6 chanx_left_in[19]
port 13 nsew default input
rlabel metal3 s 0 12792 480 12912 6 chanx_left_in[1]
port 14 nsew default input
rlabel metal3 s 0 13336 480 13456 6 chanx_left_in[2]
port 15 nsew default input
rlabel metal3 s 0 14016 480 14136 6 chanx_left_in[3]
port 16 nsew default input
rlabel metal3 s 0 14560 480 14680 6 chanx_left_in[4]
port 17 nsew default input
rlabel metal3 s 0 15240 480 15360 6 chanx_left_in[5]
port 18 nsew default input
rlabel metal3 s 0 15784 480 15904 6 chanx_left_in[6]
port 19 nsew default input
rlabel metal3 s 0 16328 480 16448 6 chanx_left_in[7]
port 20 nsew default input
rlabel metal3 s 0 17008 480 17128 6 chanx_left_in[8]
port 21 nsew default input
rlabel metal3 s 0 17552 480 17672 6 chanx_left_in[9]
port 22 nsew default input
rlabel metal3 s 0 280 480 400 6 chanx_left_out[0]
port 23 nsew default tristate
rlabel metal3 s 0 6264 480 6384 6 chanx_left_out[10]
port 24 nsew default tristate
rlabel metal3 s 0 6808 480 6928 6 chanx_left_out[11]
port 25 nsew default tristate
rlabel metal3 s 0 7352 480 7472 6 chanx_left_out[12]
port 26 nsew default tristate
rlabel metal3 s 0 8032 480 8152 6 chanx_left_out[13]
port 27 nsew default tristate
rlabel metal3 s 0 8576 480 8696 6 chanx_left_out[14]
port 28 nsew default tristate
rlabel metal3 s 0 9256 480 9376 6 chanx_left_out[15]
port 29 nsew default tristate
rlabel metal3 s 0 9800 480 9920 6 chanx_left_out[16]
port 30 nsew default tristate
rlabel metal3 s 0 10344 480 10464 6 chanx_left_out[17]
port 31 nsew default tristate
rlabel metal3 s 0 11024 480 11144 6 chanx_left_out[18]
port 32 nsew default tristate
rlabel metal3 s 0 11568 480 11688 6 chanx_left_out[19]
port 33 nsew default tristate
rlabel metal3 s 0 824 480 944 6 chanx_left_out[1]
port 34 nsew default tristate
rlabel metal3 s 0 1368 480 1488 6 chanx_left_out[2]
port 35 nsew default tristate
rlabel metal3 s 0 2048 480 2168 6 chanx_left_out[3]
port 36 nsew default tristate
rlabel metal3 s 0 2592 480 2712 6 chanx_left_out[4]
port 37 nsew default tristate
rlabel metal3 s 0 3272 480 3392 6 chanx_left_out[5]
port 38 nsew default tristate
rlabel metal3 s 0 3816 480 3936 6 chanx_left_out[6]
port 39 nsew default tristate
rlabel metal3 s 0 4360 480 4480 6 chanx_left_out[7]
port 40 nsew default tristate
rlabel metal3 s 0 5040 480 5160 6 chanx_left_out[8]
port 41 nsew default tristate
rlabel metal3 s 0 5584 480 5704 6 chanx_left_out[9]
port 42 nsew default tristate
rlabel metal3 s 29520 12248 30000 12368 6 chanx_right_in[0]
port 43 nsew default input
rlabel metal3 s 29520 18232 30000 18352 6 chanx_right_in[10]
port 44 nsew default input
rlabel metal3 s 29520 18776 30000 18896 6 chanx_right_in[11]
port 45 nsew default input
rlabel metal3 s 29520 19320 30000 19440 6 chanx_right_in[12]
port 46 nsew default input
rlabel metal3 s 29520 20000 30000 20120 6 chanx_right_in[13]
port 47 nsew default input
rlabel metal3 s 29520 20544 30000 20664 6 chanx_right_in[14]
port 48 nsew default input
rlabel metal3 s 29520 21224 30000 21344 6 chanx_right_in[15]
port 49 nsew default input
rlabel metal3 s 29520 21768 30000 21888 6 chanx_right_in[16]
port 50 nsew default input
rlabel metal3 s 29520 22312 30000 22432 6 chanx_right_in[17]
port 51 nsew default input
rlabel metal3 s 29520 22992 30000 23112 6 chanx_right_in[18]
port 52 nsew default input
rlabel metal3 s 29520 23536 30000 23656 6 chanx_right_in[19]
port 53 nsew default input
rlabel metal3 s 29520 12792 30000 12912 6 chanx_right_in[1]
port 54 nsew default input
rlabel metal3 s 29520 13336 30000 13456 6 chanx_right_in[2]
port 55 nsew default input
rlabel metal3 s 29520 14016 30000 14136 6 chanx_right_in[3]
port 56 nsew default input
rlabel metal3 s 29520 14560 30000 14680 6 chanx_right_in[4]
port 57 nsew default input
rlabel metal3 s 29520 15240 30000 15360 6 chanx_right_in[5]
port 58 nsew default input
rlabel metal3 s 29520 15784 30000 15904 6 chanx_right_in[6]
port 59 nsew default input
rlabel metal3 s 29520 16328 30000 16448 6 chanx_right_in[7]
port 60 nsew default input
rlabel metal3 s 29520 17008 30000 17128 6 chanx_right_in[8]
port 61 nsew default input
rlabel metal3 s 29520 17552 30000 17672 6 chanx_right_in[9]
port 62 nsew default input
rlabel metal3 s 29520 280 30000 400 6 chanx_right_out[0]
port 63 nsew default tristate
rlabel metal3 s 29520 6264 30000 6384 6 chanx_right_out[10]
port 64 nsew default tristate
rlabel metal3 s 29520 6808 30000 6928 6 chanx_right_out[11]
port 65 nsew default tristate
rlabel metal3 s 29520 7352 30000 7472 6 chanx_right_out[12]
port 66 nsew default tristate
rlabel metal3 s 29520 8032 30000 8152 6 chanx_right_out[13]
port 67 nsew default tristate
rlabel metal3 s 29520 8576 30000 8696 6 chanx_right_out[14]
port 68 nsew default tristate
rlabel metal3 s 29520 9256 30000 9376 6 chanx_right_out[15]
port 69 nsew default tristate
rlabel metal3 s 29520 9800 30000 9920 6 chanx_right_out[16]
port 70 nsew default tristate
rlabel metal3 s 29520 10344 30000 10464 6 chanx_right_out[17]
port 71 nsew default tristate
rlabel metal3 s 29520 11024 30000 11144 6 chanx_right_out[18]
port 72 nsew default tristate
rlabel metal3 s 29520 11568 30000 11688 6 chanx_right_out[19]
port 73 nsew default tristate
rlabel metal3 s 29520 824 30000 944 6 chanx_right_out[1]
port 74 nsew default tristate
rlabel metal3 s 29520 1368 30000 1488 6 chanx_right_out[2]
port 75 nsew default tristate
rlabel metal3 s 29520 2048 30000 2168 6 chanx_right_out[3]
port 76 nsew default tristate
rlabel metal3 s 29520 2592 30000 2712 6 chanx_right_out[4]
port 77 nsew default tristate
rlabel metal3 s 29520 3272 30000 3392 6 chanx_right_out[5]
port 78 nsew default tristate
rlabel metal3 s 29520 3816 30000 3936 6 chanx_right_out[6]
port 79 nsew default tristate
rlabel metal3 s 29520 4360 30000 4480 6 chanx_right_out[7]
port 80 nsew default tristate
rlabel metal3 s 29520 5040 30000 5160 6 chanx_right_out[8]
port 81 nsew default tristate
rlabel metal3 s 29520 5584 30000 5704 6 chanx_right_out[9]
port 82 nsew default tristate
rlabel metal2 s 26146 0 26202 480 6 prog_clk
port 83 nsew default input
rlabel metal2 s 938 23520 994 24000 6 top_grid_pin_16_
port 84 nsew default tristate
rlabel metal2 s 2778 23520 2834 24000 6 top_grid_pin_17_
port 85 nsew default tristate
rlabel metal2 s 4618 23520 4674 24000 6 top_grid_pin_18_
port 86 nsew default tristate
rlabel metal2 s 6550 23520 6606 24000 6 top_grid_pin_19_
port 87 nsew default tristate
rlabel metal2 s 8390 23520 8446 24000 6 top_grid_pin_20_
port 88 nsew default tristate
rlabel metal2 s 10230 23520 10286 24000 6 top_grid_pin_21_
port 89 nsew default tristate
rlabel metal2 s 12162 23520 12218 24000 6 top_grid_pin_22_
port 90 nsew default tristate
rlabel metal2 s 14002 23520 14058 24000 6 top_grid_pin_23_
port 91 nsew default tristate
rlabel metal2 s 15934 23520 15990 24000 6 top_grid_pin_24_
port 92 nsew default tristate
rlabel metal2 s 17774 23520 17830 24000 6 top_grid_pin_25_
port 93 nsew default tristate
rlabel metal2 s 19614 23520 19670 24000 6 top_grid_pin_26_
port 94 nsew default tristate
rlabel metal2 s 21546 23520 21602 24000 6 top_grid_pin_27_
port 95 nsew default tristate
rlabel metal2 s 23386 23520 23442 24000 6 top_grid_pin_28_
port 96 nsew default tristate
rlabel metal2 s 25226 23520 25282 24000 6 top_grid_pin_29_
port 97 nsew default tristate
rlabel metal2 s 27158 23520 27214 24000 6 top_grid_pin_30_
port 98 nsew default tristate
rlabel metal2 s 28998 23520 29054 24000 6 top_grid_pin_31_
port 99 nsew default tristate
rlabel metal4 s 5944 2128 6264 21808 6 VPWR
port 100 nsew default input
rlabel metal4 s 10944 2128 11264 21808 6 VGND
port 101 nsew default input
<< properties >>
string FIXED_BBOX 0 0 30000 24000
<< end >>
